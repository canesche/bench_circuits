// Benchmark "testing" written by ABC on Thu Oct  8 22:16:41 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A139  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A139;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2254]_ , \new_[2255]_ , \new_[2256]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2260]_ ,
    \new_[2261]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2271]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2274]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2277]_ , \new_[2278]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2290]_ , \new_[2291]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2310]_ , \new_[2311]_ , \new_[2312]_ ,
    \new_[2313]_ , \new_[2314]_ , \new_[2315]_ , \new_[2316]_ ,
    \new_[2317]_ , \new_[2318]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2326]_ , \new_[2327]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2333]_ , \new_[2334]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2337]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2342]_ , \new_[2343]_ , \new_[2344]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2350]_ , \new_[2351]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2382]_ , \new_[2383]_ , \new_[2384]_ ,
    \new_[2385]_ , \new_[2386]_ , \new_[2387]_ , \new_[2388]_ ,
    \new_[2389]_ , \new_[2390]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2394]_ , \new_[2395]_ , \new_[2396]_ ,
    \new_[2397]_ , \new_[2398]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2407]_ , \new_[2408]_ ,
    \new_[2409]_ , \new_[2410]_ , \new_[2411]_ , \new_[2412]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2445]_ , \new_[2446]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2470]_ , \new_[2471]_ , \new_[2472]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2477]_ , \new_[2478]_ , \new_[2479]_ , \new_[2480]_ ,
    \new_[2481]_ , \new_[2482]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2489]_ , \new_[2490]_ , \new_[2491]_ , \new_[2492]_ ,
    \new_[2493]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2512]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2518]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2525]_ , \new_[2526]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2552]_ ,
    \new_[2553]_ , \new_[2554]_ , \new_[2555]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2559]_ , \new_[2560]_ ,
    \new_[2561]_ , \new_[2562]_ , \new_[2563]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2567]_ , \new_[2568]_ ,
    \new_[2569]_ , \new_[2570]_ , \new_[2571]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2574]_ , \new_[2575]_ , \new_[2576]_ ,
    \new_[2577]_ , \new_[2578]_ , \new_[2579]_ , \new_[2580]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2584]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2587]_ , \new_[2588]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2599]_ , \new_[2600]_ ,
    \new_[2601]_ , \new_[2602]_ , \new_[2603]_ , \new_[2604]_ ,
    \new_[2605]_ , \new_[2606]_ , \new_[2607]_ , \new_[2608]_ ,
    \new_[2609]_ , \new_[2610]_ , \new_[2611]_ , \new_[2612]_ ,
    \new_[2613]_ , \new_[2614]_ , \new_[2615]_ , \new_[2616]_ ,
    \new_[2617]_ , \new_[2618]_ , \new_[2619]_ , \new_[2620]_ ,
    \new_[2621]_ , \new_[2622]_ , \new_[2623]_ , \new_[2624]_ ,
    \new_[2625]_ , \new_[2626]_ , \new_[2627]_ , \new_[2628]_ ,
    \new_[2629]_ , \new_[2630]_ , \new_[2631]_ , \new_[2632]_ ,
    \new_[2633]_ , \new_[2634]_ , \new_[2635]_ , \new_[2636]_ ,
    \new_[2637]_ , \new_[2638]_ , \new_[2639]_ , \new_[2640]_ ,
    \new_[2641]_ , \new_[2642]_ , \new_[2643]_ , \new_[2644]_ ,
    \new_[2645]_ , \new_[2646]_ , \new_[2647]_ , \new_[2648]_ ,
    \new_[2649]_ , \new_[2650]_ , \new_[2651]_ , \new_[2652]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2655]_ , \new_[2656]_ ,
    \new_[2657]_ , \new_[2658]_ , \new_[2659]_ , \new_[2660]_ ,
    \new_[2661]_ , \new_[2662]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2669]_ , \new_[2670]_ , \new_[2671]_ , \new_[2672]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2724]_ ,
    \new_[2725]_ , \new_[2726]_ , \new_[2727]_ , \new_[2728]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2731]_ , \new_[2732]_ ,
    \new_[2733]_ , \new_[2734]_ , \new_[2735]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2743]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2746]_ , \new_[2747]_ , \new_[2748]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2758]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2778]_ , \new_[2779]_ , \new_[2780]_ ,
    \new_[2781]_ , \new_[2782]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2785]_ , \new_[2786]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2796]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2803]_ , \new_[2804]_ ,
    \new_[2805]_ , \new_[2806]_ , \new_[2807]_ , \new_[2808]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2812]_ ,
    \new_[2813]_ , \new_[2814]_ , \new_[2815]_ , \new_[2816]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2819]_ , \new_[2820]_ ,
    \new_[2821]_ , \new_[2822]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2829]_ , \new_[2830]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2836]_ ,
    \new_[2837]_ , \new_[2838]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2843]_ , \new_[2844]_ ,
    \new_[2845]_ , \new_[2846]_ , \new_[2847]_ , \new_[2848]_ ,
    \new_[2849]_ , \new_[2850]_ , \new_[2851]_ , \new_[2852]_ ,
    \new_[2853]_ , \new_[2854]_ , \new_[2855]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2858]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2861]_ , \new_[2862]_ , \new_[2863]_ , \new_[2864]_ ,
    \new_[2865]_ , \new_[2866]_ , \new_[2867]_ , \new_[2868]_ ,
    \new_[2869]_ , \new_[2870]_ , \new_[2871]_ , \new_[2872]_ ,
    \new_[2873]_ , \new_[2874]_ , \new_[2875]_ , \new_[2876]_ ,
    \new_[2877]_ , \new_[2878]_ , \new_[2879]_ , \new_[2880]_ ,
    \new_[2881]_ , \new_[2882]_ , \new_[2883]_ , \new_[2884]_ ,
    \new_[2885]_ , \new_[2886]_ , \new_[2887]_ , \new_[2888]_ ,
    \new_[2889]_ , \new_[2890]_ , \new_[2891]_ , \new_[2892]_ ,
    \new_[2893]_ , \new_[2894]_ , \new_[2895]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2898]_ , \new_[2899]_ , \new_[2900]_ ,
    \new_[2901]_ , \new_[2902]_ , \new_[2903]_ , \new_[2904]_ ,
    \new_[2905]_ , \new_[2906]_ , \new_[2907]_ , \new_[2908]_ ,
    \new_[2909]_ , \new_[2910]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2915]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2934]_ , \new_[2935]_ , \new_[2936]_ ,
    \new_[2937]_ , \new_[2938]_ , \new_[2939]_ , \new_[2940]_ ,
    \new_[2941]_ , \new_[2942]_ , \new_[2943]_ , \new_[2944]_ ,
    \new_[2945]_ , \new_[2946]_ , \new_[2947]_ , \new_[2948]_ ,
    \new_[2949]_ , \new_[2950]_ , \new_[2951]_ , \new_[2952]_ ,
    \new_[2953]_ , \new_[2954]_ , \new_[2955]_ , \new_[2956]_ ,
    \new_[2957]_ , \new_[2958]_ , \new_[2959]_ , \new_[2960]_ ,
    \new_[2961]_ , \new_[2962]_ , \new_[2963]_ , \new_[2964]_ ,
    \new_[2965]_ , \new_[2966]_ , \new_[2967]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2970]_ , \new_[2971]_ , \new_[2972]_ ,
    \new_[2973]_ , \new_[2974]_ , \new_[2975]_ , \new_[2976]_ ,
    \new_[2977]_ , \new_[2978]_ , \new_[2979]_ , \new_[2980]_ ,
    \new_[2981]_ , \new_[2982]_ , \new_[2983]_ , \new_[2984]_ ,
    \new_[2985]_ , \new_[2986]_ , \new_[2987]_ , \new_[2988]_ ,
    \new_[2989]_ , \new_[2990]_ , \new_[2991]_ , \new_[2992]_ ,
    \new_[2993]_ , \new_[2994]_ , \new_[2995]_ , \new_[2996]_ ,
    \new_[2997]_ , \new_[2998]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3003]_ , \new_[3004]_ ,
    \new_[3005]_ , \new_[3006]_ , \new_[3007]_ , \new_[3008]_ ,
    \new_[3009]_ , \new_[3010]_ , \new_[3011]_ , \new_[3012]_ ,
    \new_[3013]_ , \new_[3014]_ , \new_[3015]_ , \new_[3016]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3019]_ , \new_[3020]_ ,
    \new_[3021]_ , \new_[3022]_ , \new_[3023]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3026]_ , \new_[3027]_ , \new_[3028]_ ,
    \new_[3029]_ , \new_[3030]_ , \new_[3031]_ , \new_[3032]_ ,
    \new_[3033]_ , \new_[3034]_ , \new_[3035]_ , \new_[3036]_ ,
    \new_[3037]_ , \new_[3038]_ , \new_[3039]_ , \new_[3040]_ ,
    \new_[3041]_ , \new_[3042]_ , \new_[3043]_ , \new_[3044]_ ,
    \new_[3045]_ , \new_[3046]_ , \new_[3047]_ , \new_[3048]_ ,
    \new_[3049]_ , \new_[3050]_ , \new_[3051]_ , \new_[3052]_ ,
    \new_[3053]_ , \new_[3054]_ , \new_[3055]_ , \new_[3056]_ ,
    \new_[3057]_ , \new_[3058]_ , \new_[3059]_ , \new_[3060]_ ,
    \new_[3061]_ , \new_[3062]_ , \new_[3063]_ , \new_[3064]_ ,
    \new_[3065]_ , \new_[3066]_ , \new_[3067]_ , \new_[3068]_ ,
    \new_[3069]_ , \new_[3070]_ , \new_[3071]_ , \new_[3072]_ ,
    \new_[3073]_ , \new_[3074]_ , \new_[3075]_ , \new_[3076]_ ,
    \new_[3077]_ , \new_[3078]_ , \new_[3079]_ , \new_[3080]_ ,
    \new_[3081]_ , \new_[3082]_ , \new_[3083]_ , \new_[3084]_ ,
    \new_[3085]_ , \new_[3086]_ , \new_[3087]_ , \new_[3088]_ ,
    \new_[3089]_ , \new_[3090]_ , \new_[3091]_ , \new_[3092]_ ,
    \new_[3093]_ , \new_[3094]_ , \new_[3095]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ , \new_[3100]_ ,
    \new_[3101]_ , \new_[3102]_ , \new_[3103]_ , \new_[3104]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3107]_ , \new_[3108]_ ,
    \new_[3109]_ , \new_[3110]_ , \new_[3111]_ , \new_[3112]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3115]_ , \new_[3116]_ ,
    \new_[3117]_ , \new_[3118]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3124]_ ,
    \new_[3125]_ , \new_[3126]_ , \new_[3127]_ , \new_[3128]_ ,
    \new_[3129]_ , \new_[3130]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3135]_ , \new_[3136]_ ,
    \new_[3137]_ , \new_[3138]_ , \new_[3139]_ , \new_[3140]_ ,
    \new_[3141]_ , \new_[3142]_ , \new_[3143]_ , \new_[3144]_ ,
    \new_[3145]_ , \new_[3146]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3150]_ , \new_[3151]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3156]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3162]_ , \new_[3163]_ , \new_[3164]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3173]_ , \new_[3174]_ , \new_[3175]_ , \new_[3176]_ ,
    \new_[3177]_ , \new_[3178]_ , \new_[3179]_ , \new_[3180]_ ,
    \new_[3181]_ , \new_[3182]_ , \new_[3183]_ , \new_[3184]_ ,
    \new_[3185]_ , \new_[3186]_ , \new_[3187]_ , \new_[3188]_ ,
    \new_[3189]_ , \new_[3190]_ , \new_[3191]_ , \new_[3192]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3197]_ , \new_[3198]_ , \new_[3199]_ , \new_[3200]_ ,
    \new_[3201]_ , \new_[3202]_ , \new_[3203]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3222]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3226]_ , \new_[3227]_ , \new_[3228]_ ,
    \new_[3229]_ , \new_[3230]_ , \new_[3231]_ , \new_[3232]_ ,
    \new_[3233]_ , \new_[3234]_ , \new_[3235]_ , \new_[3236]_ ,
    \new_[3237]_ , \new_[3238]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3246]_ , \new_[3247]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3251]_ , \new_[3252]_ ,
    \new_[3253]_ , \new_[3254]_ , \new_[3255]_ , \new_[3256]_ ,
    \new_[3257]_ , \new_[3258]_ , \new_[3259]_ , \new_[3260]_ ,
    \new_[3261]_ , \new_[3262]_ , \new_[3263]_ , \new_[3264]_ ,
    \new_[3265]_ , \new_[3266]_ , \new_[3267]_ , \new_[3268]_ ,
    \new_[3269]_ , \new_[3270]_ , \new_[3271]_ , \new_[3272]_ ,
    \new_[3273]_ , \new_[3274]_ , \new_[3275]_ , \new_[3276]_ ,
    \new_[3277]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3281]_ , \new_[3282]_ , \new_[3283]_ , \new_[3284]_ ,
    \new_[3285]_ , \new_[3286]_ , \new_[3287]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3294]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3299]_ , \new_[3300]_ ,
    \new_[3301]_ , \new_[3302]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3305]_ , \new_[3306]_ , \new_[3307]_ , \new_[3308]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3319]_ , \new_[3320]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3323]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3332]_ ,
    \new_[3333]_ , \new_[3334]_ , \new_[3335]_ , \new_[3336]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3341]_ , \new_[3342]_ , \new_[3343]_ , \new_[3344]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3398]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3402]_ , \new_[3403]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3416]_ ,
    \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3426]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3429]_ , \new_[3430]_ , \new_[3431]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3438]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3444]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3492]_ ,
    \new_[3493]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3504]_ ,
    \new_[3505]_ , \new_[3506]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3516]_ ,
    \new_[3517]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3523]_ , \new_[3524]_ ,
    \new_[3525]_ , \new_[3526]_ , \new_[3527]_ , \new_[3528]_ ,
    \new_[3529]_ , \new_[3530]_ , \new_[3531]_ , \new_[3532]_ ,
    \new_[3533]_ , \new_[3534]_ , \new_[3535]_ , \new_[3536]_ ,
    \new_[3537]_ , \new_[3538]_ , \new_[3539]_ , \new_[3540]_ ,
    \new_[3541]_ , \new_[3542]_ , \new_[3543]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3546]_ , \new_[3547]_ , \new_[3548]_ ,
    \new_[3549]_ , \new_[3550]_ , \new_[3551]_ , \new_[3552]_ ,
    \new_[3553]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3557]_ , \new_[3558]_ , \new_[3559]_ , \new_[3560]_ ,
    \new_[3561]_ , \new_[3562]_ , \new_[3563]_ , \new_[3564]_ ,
    \new_[3565]_ , \new_[3566]_ , \new_[3567]_ , \new_[3568]_ ,
    \new_[3569]_ , \new_[3570]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3573]_ , \new_[3574]_ , \new_[3575]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3582]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3587]_ , \new_[3588]_ ,
    \new_[3589]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3593]_ , \new_[3594]_ , \new_[3595]_ , \new_[3596]_ ,
    \new_[3597]_ , \new_[3598]_ , \new_[3599]_ , \new_[3600]_ ,
    \new_[3601]_ , \new_[3602]_ , \new_[3603]_ , \new_[3604]_ ,
    \new_[3605]_ , \new_[3606]_ , \new_[3607]_ , \new_[3608]_ ,
    \new_[3609]_ , \new_[3610]_ , \new_[3611]_ , \new_[3612]_ ,
    \new_[3613]_ , \new_[3614]_ , \new_[3615]_ , \new_[3616]_ ,
    \new_[3617]_ , \new_[3618]_ , \new_[3619]_ , \new_[3620]_ ,
    \new_[3621]_ , \new_[3622]_ , \new_[3623]_ , \new_[3624]_ ,
    \new_[3625]_ , \new_[3626]_ , \new_[3627]_ , \new_[3628]_ ,
    \new_[3629]_ , \new_[3630]_ , \new_[3631]_ , \new_[3632]_ ,
    \new_[3633]_ , \new_[3634]_ , \new_[3635]_ , \new_[3636]_ ,
    \new_[3637]_ , \new_[3638]_ , \new_[3639]_ , \new_[3640]_ ,
    \new_[3641]_ , \new_[3642]_ , \new_[3643]_ , \new_[3644]_ ,
    \new_[3645]_ , \new_[3646]_ , \new_[3647]_ , \new_[3648]_ ,
    \new_[3649]_ , \new_[3650]_ , \new_[3651]_ , \new_[3652]_ ,
    \new_[3653]_ , \new_[3654]_ , \new_[3655]_ , \new_[3656]_ ,
    \new_[3657]_ , \new_[3658]_ , \new_[3659]_ , \new_[3660]_ ,
    \new_[3661]_ , \new_[3662]_ , \new_[3663]_ , \new_[3664]_ ,
    \new_[3665]_ , \new_[3666]_ , \new_[3667]_ , \new_[3668]_ ,
    \new_[3669]_ , \new_[3670]_ , \new_[3671]_ , \new_[3672]_ ,
    \new_[3673]_ , \new_[3674]_ , \new_[3675]_ , \new_[3676]_ ,
    \new_[3677]_ , \new_[3678]_ , \new_[3679]_ , \new_[3680]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3683]_ , \new_[3684]_ ,
    \new_[3685]_ , \new_[3686]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3690]_ , \new_[3691]_ , \new_[3692]_ ,
    \new_[3693]_ , \new_[3694]_ , \new_[3695]_ , \new_[3696]_ ,
    \new_[3697]_ , \new_[3698]_ , \new_[3699]_ , \new_[3700]_ ,
    \new_[3701]_ , \new_[3702]_ , \new_[3706]_ , \new_[3707]_ ,
    \new_[3710]_ , \new_[3713]_ , \new_[3714]_ , \new_[3715]_ ,
    \new_[3719]_ , \new_[3720]_ , \new_[3723]_ , \new_[3726]_ ,
    \new_[3727]_ , \new_[3728]_ , \new_[3729]_ , \new_[3733]_ ,
    \new_[3734]_ , \new_[3737]_ , \new_[3740]_ , \new_[3741]_ ,
    \new_[3742]_ , \new_[3746]_ , \new_[3747]_ , \new_[3750]_ ,
    \new_[3753]_ , \new_[3754]_ , \new_[3755]_ , \new_[3756]_ ,
    \new_[3757]_ , \new_[3761]_ , \new_[3762]_ , \new_[3765]_ ,
    \new_[3768]_ , \new_[3769]_ , \new_[3770]_ , \new_[3774]_ ,
    \new_[3775]_ , \new_[3778]_ , \new_[3781]_ , \new_[3782]_ ,
    \new_[3783]_ , \new_[3784]_ , \new_[3788]_ , \new_[3789]_ ,
    \new_[3792]_ , \new_[3795]_ , \new_[3796]_ , \new_[3797]_ ,
    \new_[3800]_ , \new_[3803]_ , \new_[3804]_ , \new_[3807]_ ,
    \new_[3810]_ , \new_[3811]_ , \new_[3812]_ , \new_[3813]_ ,
    \new_[3814]_ , \new_[3815]_ , \new_[3819]_ , \new_[3820]_ ,
    \new_[3823]_ , \new_[3826]_ , \new_[3827]_ , \new_[3828]_ ,
    \new_[3832]_ , \new_[3833]_ , \new_[3836]_ , \new_[3839]_ ,
    \new_[3840]_ , \new_[3841]_ , \new_[3842]_ , \new_[3846]_ ,
    \new_[3847]_ , \new_[3850]_ , \new_[3853]_ , \new_[3854]_ ,
    \new_[3855]_ , \new_[3858]_ , \new_[3861]_ , \new_[3862]_ ,
    \new_[3865]_ , \new_[3868]_ , \new_[3869]_ , \new_[3870]_ ,
    \new_[3871]_ , \new_[3872]_ , \new_[3876]_ , \new_[3877]_ ,
    \new_[3880]_ , \new_[3883]_ , \new_[3884]_ , \new_[3885]_ ,
    \new_[3889]_ , \new_[3890]_ , \new_[3893]_ , \new_[3896]_ ,
    \new_[3897]_ , \new_[3898]_ , \new_[3899]_ , \new_[3903]_ ,
    \new_[3904]_ , \new_[3907]_ , \new_[3910]_ , \new_[3911]_ ,
    \new_[3912]_ , \new_[3915]_ , \new_[3918]_ , \new_[3919]_ ,
    \new_[3922]_ , \new_[3925]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3928]_ , \new_[3929]_ , \new_[3930]_ , \new_[3931]_ ,
    \new_[3935]_ , \new_[3936]_ , \new_[3939]_ , \new_[3942]_ ,
    \new_[3943]_ , \new_[3944]_ , \new_[3948]_ , \new_[3949]_ ,
    \new_[3952]_ , \new_[3955]_ , \new_[3956]_ , \new_[3957]_ ,
    \new_[3958]_ , \new_[3962]_ , \new_[3963]_ , \new_[3966]_ ,
    \new_[3969]_ , \new_[3970]_ , \new_[3971]_ , \new_[3974]_ ,
    \new_[3977]_ , \new_[3978]_ , \new_[3981]_ , \new_[3984]_ ,
    \new_[3985]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3992]_ , \new_[3993]_ , \new_[3996]_ , \new_[3999]_ ,
    \new_[4000]_ , \new_[4001]_ , \new_[4005]_ , \new_[4006]_ ,
    \new_[4009]_ , \new_[4012]_ , \new_[4013]_ , \new_[4014]_ ,
    \new_[4015]_ , \new_[4019]_ , \new_[4020]_ , \new_[4023]_ ,
    \new_[4026]_ , \new_[4027]_ , \new_[4028]_ , \new_[4031]_ ,
    \new_[4034]_ , \new_[4035]_ , \new_[4038]_ , \new_[4041]_ ,
    \new_[4042]_ , \new_[4043]_ , \new_[4044]_ , \new_[4045]_ ,
    \new_[4046]_ , \new_[4050]_ , \new_[4051]_ , \new_[4054]_ ,
    \new_[4057]_ , \new_[4058]_ , \new_[4059]_ , \new_[4063]_ ,
    \new_[4064]_ , \new_[4067]_ , \new_[4070]_ , \new_[4071]_ ,
    \new_[4072]_ , \new_[4073]_ , \new_[4077]_ , \new_[4078]_ ,
    \new_[4081]_ , \new_[4084]_ , \new_[4085]_ , \new_[4086]_ ,
    \new_[4089]_ , \new_[4092]_ , \new_[4093]_ , \new_[4096]_ ,
    \new_[4099]_ , \new_[4100]_ , \new_[4101]_ , \new_[4102]_ ,
    \new_[4103]_ , \new_[4107]_ , \new_[4108]_ , \new_[4111]_ ,
    \new_[4114]_ , \new_[4115]_ , \new_[4116]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4124]_ , \new_[4127]_ , \new_[4128]_ ,
    \new_[4129]_ , \new_[4130]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4138]_ , \new_[4141]_ , \new_[4142]_ , \new_[4143]_ ,
    \new_[4146]_ , \new_[4149]_ , \new_[4150]_ , \new_[4153]_ ,
    \new_[4156]_ , \new_[4157]_ , \new_[4158]_ , \new_[4159]_ ,
    \new_[4160]_ , \new_[4161]_ , \new_[4162]_ , \new_[4163]_ ,
    \new_[4167]_ , \new_[4168]_ , \new_[4171]_ , \new_[4174]_ ,
    \new_[4175]_ , \new_[4176]_ , \new_[4180]_ , \new_[4181]_ ,
    \new_[4184]_ , \new_[4187]_ , \new_[4188]_ , \new_[4189]_ ,
    \new_[4190]_ , \new_[4194]_ , \new_[4195]_ , \new_[4198]_ ,
    \new_[4201]_ , \new_[4202]_ , \new_[4203]_ , \new_[4207]_ ,
    \new_[4208]_ , \new_[4211]_ , \new_[4214]_ , \new_[4215]_ ,
    \new_[4216]_ , \new_[4217]_ , \new_[4218]_ , \new_[4222]_ ,
    \new_[4223]_ , \new_[4226]_ , \new_[4229]_ , \new_[4230]_ ,
    \new_[4231]_ , \new_[4235]_ , \new_[4236]_ , \new_[4239]_ ,
    \new_[4242]_ , \new_[4243]_ , \new_[4244]_ , \new_[4245]_ ,
    \new_[4249]_ , \new_[4250]_ , \new_[4253]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4261]_ , \new_[4264]_ ,
    \new_[4265]_ , \new_[4268]_ , \new_[4271]_ , \new_[4272]_ ,
    \new_[4273]_ , \new_[4274]_ , \new_[4275]_ , \new_[4276]_ ,
    \new_[4280]_ , \new_[4281]_ , \new_[4284]_ , \new_[4287]_ ,
    \new_[4288]_ , \new_[4289]_ , \new_[4293]_ , \new_[4294]_ ,
    \new_[4297]_ , \new_[4300]_ , \new_[4301]_ , \new_[4302]_ ,
    \new_[4303]_ , \new_[4307]_ , \new_[4308]_ , \new_[4311]_ ,
    \new_[4314]_ , \new_[4315]_ , \new_[4316]_ , \new_[4319]_ ,
    \new_[4322]_ , \new_[4323]_ , \new_[4326]_ , \new_[4329]_ ,
    \new_[4330]_ , \new_[4331]_ , \new_[4332]_ , \new_[4333]_ ,
    \new_[4337]_ , \new_[4338]_ , \new_[4341]_ , \new_[4344]_ ,
    \new_[4345]_ , \new_[4346]_ , \new_[4350]_ , \new_[4351]_ ,
    \new_[4354]_ , \new_[4357]_ , \new_[4358]_ , \new_[4359]_ ,
    \new_[4360]_ , \new_[4364]_ , \new_[4365]_ , \new_[4368]_ ,
    \new_[4371]_ , \new_[4372]_ , \new_[4373]_ , \new_[4376]_ ,
    \new_[4379]_ , \new_[4380]_ , \new_[4383]_ , \new_[4386]_ ,
    \new_[4387]_ , \new_[4388]_ , \new_[4389]_ , \new_[4390]_ ,
    \new_[4391]_ , \new_[4392]_ , \new_[4396]_ , \new_[4397]_ ,
    \new_[4400]_ , \new_[4403]_ , \new_[4404]_ , \new_[4405]_ ,
    \new_[4409]_ , \new_[4410]_ , \new_[4413]_ , \new_[4416]_ ,
    \new_[4417]_ , \new_[4418]_ , \new_[4419]_ , \new_[4423]_ ,
    \new_[4424]_ , \new_[4427]_ , \new_[4430]_ , \new_[4431]_ ,
    \new_[4432]_ , \new_[4435]_ , \new_[4438]_ , \new_[4439]_ ,
    \new_[4442]_ , \new_[4445]_ , \new_[4446]_ , \new_[4447]_ ,
    \new_[4448]_ , \new_[4449]_ , \new_[4453]_ , \new_[4454]_ ,
    \new_[4457]_ , \new_[4460]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4466]_ , \new_[4467]_ , \new_[4470]_ , \new_[4473]_ ,
    \new_[4474]_ , \new_[4475]_ , \new_[4476]_ , \new_[4480]_ ,
    \new_[4481]_ , \new_[4484]_ , \new_[4487]_ , \new_[4488]_ ,
    \new_[4489]_ , \new_[4492]_ , \new_[4495]_ , \new_[4496]_ ,
    \new_[4499]_ , \new_[4502]_ , \new_[4503]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4507]_ , \new_[4511]_ ,
    \new_[4512]_ , \new_[4515]_ , \new_[4518]_ , \new_[4519]_ ,
    \new_[4520]_ , \new_[4524]_ , \new_[4525]_ , \new_[4528]_ ,
    \new_[4531]_ , \new_[4532]_ , \new_[4533]_ , \new_[4534]_ ,
    \new_[4538]_ , \new_[4539]_ , \new_[4542]_ , \new_[4545]_ ,
    \new_[4546]_ , \new_[4547]_ , \new_[4550]_ , \new_[4553]_ ,
    \new_[4554]_ , \new_[4557]_ , \new_[4560]_ , \new_[4561]_ ,
    \new_[4562]_ , \new_[4563]_ , \new_[4564]_ , \new_[4568]_ ,
    \new_[4569]_ , \new_[4572]_ , \new_[4575]_ , \new_[4576]_ ,
    \new_[4577]_ , \new_[4581]_ , \new_[4582]_ , \new_[4585]_ ,
    \new_[4588]_ , \new_[4589]_ , \new_[4590]_ , \new_[4591]_ ,
    \new_[4595]_ , \new_[4596]_ , \new_[4599]_ , \new_[4602]_ ,
    \new_[4603]_ , \new_[4604]_ , \new_[4607]_ , \new_[4610]_ ,
    \new_[4611]_ , \new_[4614]_ , \new_[4617]_ , \new_[4618]_ ,
    \new_[4619]_ , \new_[4620]_ , \new_[4621]_ , \new_[4622]_ ,
    \new_[4623]_ , \new_[4624]_ , \new_[4625]_ , \new_[4629]_ ,
    \new_[4630]_ , \new_[4633]_ , \new_[4636]_ , \new_[4637]_ ,
    \new_[4638]_ , \new_[4642]_ , \new_[4643]_ , \new_[4646]_ ,
    \new_[4649]_ , \new_[4650]_ , \new_[4651]_ , \new_[4652]_ ,
    \new_[4656]_ , \new_[4657]_ , \new_[4660]_ , \new_[4663]_ ,
    \new_[4664]_ , \new_[4665]_ , \new_[4669]_ , \new_[4670]_ ,
    \new_[4673]_ , \new_[4676]_ , \new_[4677]_ , \new_[4678]_ ,
    \new_[4679]_ , \new_[4680]_ , \new_[4684]_ , \new_[4685]_ ,
    \new_[4688]_ , \new_[4691]_ , \new_[4692]_ , \new_[4693]_ ,
    \new_[4697]_ , \new_[4698]_ , \new_[4701]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4706]_ , \new_[4707]_ , \new_[4711]_ ,
    \new_[4712]_ , \new_[4715]_ , \new_[4718]_ , \new_[4719]_ ,
    \new_[4720]_ , \new_[4723]_ , \new_[4726]_ , \new_[4727]_ ,
    \new_[4730]_ , \new_[4733]_ , \new_[4734]_ , \new_[4735]_ ,
    \new_[4736]_ , \new_[4737]_ , \new_[4738]_ , \new_[4742]_ ,
    \new_[4743]_ , \new_[4746]_ , \new_[4749]_ , \new_[4750]_ ,
    \new_[4751]_ , \new_[4755]_ , \new_[4756]_ , \new_[4759]_ ,
    \new_[4762]_ , \new_[4763]_ , \new_[4764]_ , \new_[4765]_ ,
    \new_[4769]_ , \new_[4770]_ , \new_[4773]_ , \new_[4776]_ ,
    \new_[4777]_ , \new_[4778]_ , \new_[4781]_ , \new_[4784]_ ,
    \new_[4785]_ , \new_[4788]_ , \new_[4791]_ , \new_[4792]_ ,
    \new_[4793]_ , \new_[4794]_ , \new_[4795]_ , \new_[4799]_ ,
    \new_[4800]_ , \new_[4803]_ , \new_[4806]_ , \new_[4807]_ ,
    \new_[4808]_ , \new_[4812]_ , \new_[4813]_ , \new_[4816]_ ,
    \new_[4819]_ , \new_[4820]_ , \new_[4821]_ , \new_[4822]_ ,
    \new_[4826]_ , \new_[4827]_ , \new_[4830]_ , \new_[4833]_ ,
    \new_[4834]_ , \new_[4835]_ , \new_[4838]_ , \new_[4841]_ ,
    \new_[4842]_ , \new_[4845]_ , \new_[4848]_ , \new_[4849]_ ,
    \new_[4850]_ , \new_[4851]_ , \new_[4852]_ , \new_[4853]_ ,
    \new_[4854]_ , \new_[4858]_ , \new_[4859]_ , \new_[4862]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4871]_ ,
    \new_[4872]_ , \new_[4875]_ , \new_[4878]_ , \new_[4879]_ ,
    \new_[4880]_ , \new_[4881]_ , \new_[4885]_ , \new_[4886]_ ,
    \new_[4889]_ , \new_[4892]_ , \new_[4893]_ , \new_[4894]_ ,
    \new_[4897]_ , \new_[4900]_ , \new_[4901]_ , \new_[4904]_ ,
    \new_[4907]_ , \new_[4908]_ , \new_[4909]_ , \new_[4910]_ ,
    \new_[4911]_ , \new_[4915]_ , \new_[4916]_ , \new_[4919]_ ,
    \new_[4922]_ , \new_[4923]_ , \new_[4924]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4932]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4942]_ , \new_[4943]_ ,
    \new_[4946]_ , \new_[4949]_ , \new_[4950]_ , \new_[4951]_ ,
    \new_[4954]_ , \new_[4957]_ , \new_[4958]_ , \new_[4961]_ ,
    \new_[4964]_ , \new_[4965]_ , \new_[4966]_ , \new_[4967]_ ,
    \new_[4968]_ , \new_[4969]_ , \new_[4973]_ , \new_[4974]_ ,
    \new_[4977]_ , \new_[4980]_ , \new_[4981]_ , \new_[4982]_ ,
    \new_[4986]_ , \new_[4987]_ , \new_[4990]_ , \new_[4993]_ ,
    \new_[4994]_ , \new_[4995]_ , \new_[4996]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5004]_ , \new_[5007]_ , \new_[5008]_ ,
    \new_[5009]_ , \new_[5012]_ , \new_[5015]_ , \new_[5016]_ ,
    \new_[5019]_ , \new_[5022]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5025]_ , \new_[5026]_ , \new_[5030]_ , \new_[5031]_ ,
    \new_[5034]_ , \new_[5037]_ , \new_[5038]_ , \new_[5039]_ ,
    \new_[5043]_ , \new_[5044]_ , \new_[5047]_ , \new_[5050]_ ,
    \new_[5051]_ , \new_[5052]_ , \new_[5053]_ , \new_[5057]_ ,
    \new_[5058]_ , \new_[5061]_ , \new_[5064]_ , \new_[5065]_ ,
    \new_[5066]_ , \new_[5069]_ , \new_[5072]_ , \new_[5073]_ ,
    \new_[5076]_ , \new_[5079]_ , \new_[5080]_ , \new_[5081]_ ,
    \new_[5082]_ , \new_[5083]_ , \new_[5084]_ , \new_[5085]_ ,
    \new_[5086]_ , \new_[5090]_ , \new_[5091]_ , \new_[5094]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5099]_ , \new_[5103]_ ,
    \new_[5104]_ , \new_[5107]_ , \new_[5110]_ , \new_[5111]_ ,
    \new_[5112]_ , \new_[5113]_ , \new_[5117]_ , \new_[5118]_ ,
    \new_[5121]_ , \new_[5124]_ , \new_[5125]_ , \new_[5126]_ ,
    \new_[5129]_ , \new_[5132]_ , \new_[5133]_ , \new_[5136]_ ,
    \new_[5139]_ , \new_[5140]_ , \new_[5141]_ , \new_[5142]_ ,
    \new_[5143]_ , \new_[5147]_ , \new_[5148]_ , \new_[5151]_ ,
    \new_[5154]_ , \new_[5155]_ , \new_[5156]_ , \new_[5160]_ ,
    \new_[5161]_ , \new_[5164]_ , \new_[5167]_ , \new_[5168]_ ,
    \new_[5169]_ , \new_[5170]_ , \new_[5174]_ , \new_[5175]_ ,
    \new_[5178]_ , \new_[5181]_ , \new_[5182]_ , \new_[5183]_ ,
    \new_[5186]_ , \new_[5189]_ , \new_[5190]_ , \new_[5193]_ ,
    \new_[5196]_ , \new_[5197]_ , \new_[5198]_ , \new_[5199]_ ,
    \new_[5200]_ , \new_[5201]_ , \new_[5205]_ , \new_[5206]_ ,
    \new_[5209]_ , \new_[5212]_ , \new_[5213]_ , \new_[5214]_ ,
    \new_[5218]_ , \new_[5219]_ , \new_[5222]_ , \new_[5225]_ ,
    \new_[5226]_ , \new_[5227]_ , \new_[5228]_ , \new_[5232]_ ,
    \new_[5233]_ , \new_[5236]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5241]_ , \new_[5244]_ , \new_[5247]_ , \new_[5248]_ ,
    \new_[5251]_ , \new_[5254]_ , \new_[5255]_ , \new_[5256]_ ,
    \new_[5257]_ , \new_[5258]_ , \new_[5262]_ , \new_[5263]_ ,
    \new_[5266]_ , \new_[5269]_ , \new_[5270]_ , \new_[5271]_ ,
    \new_[5275]_ , \new_[5276]_ , \new_[5279]_ , \new_[5282]_ ,
    \new_[5283]_ , \new_[5284]_ , \new_[5285]_ , \new_[5289]_ ,
    \new_[5290]_ , \new_[5293]_ , \new_[5296]_ , \new_[5297]_ ,
    \new_[5298]_ , \new_[5301]_ , \new_[5304]_ , \new_[5305]_ ,
    \new_[5308]_ , \new_[5311]_ , \new_[5312]_ , \new_[5313]_ ,
    \new_[5314]_ , \new_[5315]_ , \new_[5316]_ , \new_[5317]_ ,
    \new_[5321]_ , \new_[5322]_ , \new_[5325]_ , \new_[5328]_ ,
    \new_[5329]_ , \new_[5330]_ , \new_[5334]_ , \new_[5335]_ ,
    \new_[5338]_ , \new_[5341]_ , \new_[5342]_ , \new_[5343]_ ,
    \new_[5344]_ , \new_[5348]_ , \new_[5349]_ , \new_[5352]_ ,
    \new_[5355]_ , \new_[5356]_ , \new_[5357]_ , \new_[5360]_ ,
    \new_[5363]_ , \new_[5364]_ , \new_[5367]_ , \new_[5370]_ ,
    \new_[5371]_ , \new_[5372]_ , \new_[5373]_ , \new_[5374]_ ,
    \new_[5378]_ , \new_[5379]_ , \new_[5382]_ , \new_[5385]_ ,
    \new_[5386]_ , \new_[5387]_ , \new_[5391]_ , \new_[5392]_ ,
    \new_[5395]_ , \new_[5398]_ , \new_[5399]_ , \new_[5400]_ ,
    \new_[5401]_ , \new_[5405]_ , \new_[5406]_ , \new_[5409]_ ,
    \new_[5412]_ , \new_[5413]_ , \new_[5414]_ , \new_[5417]_ ,
    \new_[5420]_ , \new_[5421]_ , \new_[5424]_ , \new_[5427]_ ,
    \new_[5428]_ , \new_[5429]_ , \new_[5430]_ , \new_[5431]_ ,
    \new_[5432]_ , \new_[5436]_ , \new_[5437]_ , \new_[5440]_ ,
    \new_[5443]_ , \new_[5444]_ , \new_[5445]_ , \new_[5449]_ ,
    \new_[5450]_ , \new_[5453]_ , \new_[5456]_ , \new_[5457]_ ,
    \new_[5458]_ , \new_[5459]_ , \new_[5463]_ , \new_[5464]_ ,
    \new_[5467]_ , \new_[5470]_ , \new_[5471]_ , \new_[5472]_ ,
    \new_[5475]_ , \new_[5478]_ , \new_[5479]_ , \new_[5482]_ ,
    \new_[5485]_ , \new_[5486]_ , \new_[5487]_ , \new_[5488]_ ,
    \new_[5489]_ , \new_[5493]_ , \new_[5494]_ , \new_[5497]_ ,
    \new_[5500]_ , \new_[5501]_ , \new_[5502]_ , \new_[5506]_ ,
    \new_[5507]_ , \new_[5510]_ , \new_[5513]_ , \new_[5514]_ ,
    \new_[5515]_ , \new_[5516]_ , \new_[5520]_ , \new_[5521]_ ,
    \new_[5524]_ , \new_[5527]_ , \new_[5528]_ , \new_[5529]_ ,
    \new_[5532]_ , \new_[5535]_ , \new_[5536]_ , \new_[5539]_ ,
    \new_[5542]_ , \new_[5543]_ , \new_[5544]_ , \new_[5545]_ ,
    \new_[5546]_ , \new_[5547]_ , \new_[5548]_ , \new_[5549]_ ,
    \new_[5550]_ , \new_[5551]_ , \new_[5555]_ , \new_[5556]_ ,
    \new_[5559]_ , \new_[5562]_ , \new_[5563]_ , \new_[5564]_ ,
    \new_[5568]_ , \new_[5569]_ , \new_[5572]_ , \new_[5575]_ ,
    \new_[5576]_ , \new_[5577]_ , \new_[5578]_ , \new_[5582]_ ,
    \new_[5583]_ , \new_[5586]_ , \new_[5589]_ , \new_[5590]_ ,
    \new_[5591]_ , \new_[5595]_ , \new_[5596]_ , \new_[5599]_ ,
    \new_[5602]_ , \new_[5603]_ , \new_[5604]_ , \new_[5605]_ ,
    \new_[5606]_ , \new_[5610]_ , \new_[5611]_ , \new_[5614]_ ,
    \new_[5617]_ , \new_[5618]_ , \new_[5619]_ , \new_[5623]_ ,
    \new_[5624]_ , \new_[5627]_ , \new_[5630]_ , \new_[5631]_ ,
    \new_[5632]_ , \new_[5633]_ , \new_[5637]_ , \new_[5638]_ ,
    \new_[5641]_ , \new_[5644]_ , \new_[5645]_ , \new_[5646]_ ,
    \new_[5649]_ , \new_[5652]_ , \new_[5653]_ , \new_[5656]_ ,
    \new_[5659]_ , \new_[5660]_ , \new_[5661]_ , \new_[5662]_ ,
    \new_[5663]_ , \new_[5664]_ , \new_[5668]_ , \new_[5669]_ ,
    \new_[5672]_ , \new_[5675]_ , \new_[5676]_ , \new_[5677]_ ,
    \new_[5681]_ , \new_[5682]_ , \new_[5685]_ , \new_[5688]_ ,
    \new_[5689]_ , \new_[5690]_ , \new_[5691]_ , \new_[5695]_ ,
    \new_[5696]_ , \new_[5699]_ , \new_[5702]_ , \new_[5703]_ ,
    \new_[5704]_ , \new_[5707]_ , \new_[5710]_ , \new_[5711]_ ,
    \new_[5714]_ , \new_[5717]_ , \new_[5718]_ , \new_[5719]_ ,
    \new_[5720]_ , \new_[5721]_ , \new_[5725]_ , \new_[5726]_ ,
    \new_[5729]_ , \new_[5732]_ , \new_[5733]_ , \new_[5734]_ ,
    \new_[5738]_ , \new_[5739]_ , \new_[5742]_ , \new_[5745]_ ,
    \new_[5746]_ , \new_[5747]_ , \new_[5748]_ , \new_[5752]_ ,
    \new_[5753]_ , \new_[5756]_ , \new_[5759]_ , \new_[5760]_ ,
    \new_[5761]_ , \new_[5764]_ , \new_[5767]_ , \new_[5768]_ ,
    \new_[5771]_ , \new_[5774]_ , \new_[5775]_ , \new_[5776]_ ,
    \new_[5777]_ , \new_[5778]_ , \new_[5779]_ , \new_[5780]_ ,
    \new_[5784]_ , \new_[5785]_ , \new_[5788]_ , \new_[5791]_ ,
    \new_[5792]_ , \new_[5793]_ , \new_[5797]_ , \new_[5798]_ ,
    \new_[5801]_ , \new_[5804]_ , \new_[5805]_ , \new_[5806]_ ,
    \new_[5807]_ , \new_[5811]_ , \new_[5812]_ , \new_[5815]_ ,
    \new_[5818]_ , \new_[5819]_ , \new_[5820]_ , \new_[5823]_ ,
    \new_[5826]_ , \new_[5827]_ , \new_[5830]_ , \new_[5833]_ ,
    \new_[5834]_ , \new_[5835]_ , \new_[5836]_ , \new_[5837]_ ,
    \new_[5841]_ , \new_[5842]_ , \new_[5845]_ , \new_[5848]_ ,
    \new_[5849]_ , \new_[5850]_ , \new_[5854]_ , \new_[5855]_ ,
    \new_[5858]_ , \new_[5861]_ , \new_[5862]_ , \new_[5863]_ ,
    \new_[5864]_ , \new_[5868]_ , \new_[5869]_ , \new_[5872]_ ,
    \new_[5875]_ , \new_[5876]_ , \new_[5877]_ , \new_[5880]_ ,
    \new_[5883]_ , \new_[5884]_ , \new_[5887]_ , \new_[5890]_ ,
    \new_[5891]_ , \new_[5892]_ , \new_[5893]_ , \new_[5894]_ ,
    \new_[5895]_ , \new_[5899]_ , \new_[5900]_ , \new_[5903]_ ,
    \new_[5906]_ , \new_[5907]_ , \new_[5908]_ , \new_[5912]_ ,
    \new_[5913]_ , \new_[5916]_ , \new_[5919]_ , \new_[5920]_ ,
    \new_[5921]_ , \new_[5922]_ , \new_[5926]_ , \new_[5927]_ ,
    \new_[5930]_ , \new_[5933]_ , \new_[5934]_ , \new_[5935]_ ,
    \new_[5938]_ , \new_[5941]_ , \new_[5942]_ , \new_[5945]_ ,
    \new_[5948]_ , \new_[5949]_ , \new_[5950]_ , \new_[5951]_ ,
    \new_[5952]_ , \new_[5956]_ , \new_[5957]_ , \new_[5960]_ ,
    \new_[5963]_ , \new_[5964]_ , \new_[5965]_ , \new_[5969]_ ,
    \new_[5970]_ , \new_[5973]_ , \new_[5976]_ , \new_[5977]_ ,
    \new_[5978]_ , \new_[5979]_ , \new_[5983]_ , \new_[5984]_ ,
    \new_[5987]_ , \new_[5990]_ , \new_[5991]_ , \new_[5992]_ ,
    \new_[5995]_ , \new_[5998]_ , \new_[5999]_ , \new_[6002]_ ,
    \new_[6005]_ , \new_[6006]_ , \new_[6007]_ , \new_[6008]_ ,
    \new_[6009]_ , \new_[6010]_ , \new_[6011]_ , \new_[6012]_ ,
    \new_[6016]_ , \new_[6017]_ , \new_[6020]_ , \new_[6023]_ ,
    \new_[6024]_ , \new_[6025]_ , \new_[6029]_ , \new_[6030]_ ,
    \new_[6033]_ , \new_[6036]_ , \new_[6037]_ , \new_[6038]_ ,
    \new_[6039]_ , \new_[6043]_ , \new_[6044]_ , \new_[6047]_ ,
    \new_[6050]_ , \new_[6051]_ , \new_[6052]_ , \new_[6055]_ ,
    \new_[6058]_ , \new_[6059]_ , \new_[6062]_ , \new_[6065]_ ,
    \new_[6066]_ , \new_[6067]_ , \new_[6068]_ , \new_[6069]_ ,
    \new_[6073]_ , \new_[6074]_ , \new_[6077]_ , \new_[6080]_ ,
    \new_[6081]_ , \new_[6082]_ , \new_[6086]_ , \new_[6087]_ ,
    \new_[6090]_ , \new_[6093]_ , \new_[6094]_ , \new_[6095]_ ,
    \new_[6096]_ , \new_[6100]_ , \new_[6101]_ , \new_[6104]_ ,
    \new_[6107]_ , \new_[6108]_ , \new_[6109]_ , \new_[6112]_ ,
    \new_[6115]_ , \new_[6116]_ , \new_[6119]_ , \new_[6122]_ ,
    \new_[6123]_ , \new_[6124]_ , \new_[6125]_ , \new_[6126]_ ,
    \new_[6127]_ , \new_[6131]_ , \new_[6132]_ , \new_[6135]_ ,
    \new_[6138]_ , \new_[6139]_ , \new_[6140]_ , \new_[6144]_ ,
    \new_[6145]_ , \new_[6148]_ , \new_[6151]_ , \new_[6152]_ ,
    \new_[6153]_ , \new_[6154]_ , \new_[6158]_ , \new_[6159]_ ,
    \new_[6162]_ , \new_[6165]_ , \new_[6166]_ , \new_[6167]_ ,
    \new_[6170]_ , \new_[6173]_ , \new_[6174]_ , \new_[6177]_ ,
    \new_[6180]_ , \new_[6181]_ , \new_[6182]_ , \new_[6183]_ ,
    \new_[6184]_ , \new_[6188]_ , \new_[6189]_ , \new_[6192]_ ,
    \new_[6195]_ , \new_[6196]_ , \new_[6197]_ , \new_[6201]_ ,
    \new_[6202]_ , \new_[6205]_ , \new_[6208]_ , \new_[6209]_ ,
    \new_[6210]_ , \new_[6211]_ , \new_[6215]_ , \new_[6216]_ ,
    \new_[6219]_ , \new_[6222]_ , \new_[6223]_ , \new_[6224]_ ,
    \new_[6227]_ , \new_[6230]_ , \new_[6231]_ , \new_[6234]_ ,
    \new_[6237]_ , \new_[6238]_ , \new_[6239]_ , \new_[6240]_ ,
    \new_[6241]_ , \new_[6242]_ , \new_[6243]_ , \new_[6247]_ ,
    \new_[6248]_ , \new_[6251]_ , \new_[6254]_ , \new_[6255]_ ,
    \new_[6256]_ , \new_[6260]_ , \new_[6261]_ , \new_[6264]_ ,
    \new_[6267]_ , \new_[6268]_ , \new_[6269]_ , \new_[6270]_ ,
    \new_[6274]_ , \new_[6275]_ , \new_[6278]_ , \new_[6281]_ ,
    \new_[6282]_ , \new_[6283]_ , \new_[6286]_ , \new_[6289]_ ,
    \new_[6290]_ , \new_[6293]_ , \new_[6296]_ , \new_[6297]_ ,
    \new_[6298]_ , \new_[6299]_ , \new_[6300]_ , \new_[6304]_ ,
    \new_[6305]_ , \new_[6308]_ , \new_[6311]_ , \new_[6312]_ ,
    \new_[6313]_ , \new_[6317]_ , \new_[6318]_ , \new_[6321]_ ,
    \new_[6324]_ , \new_[6325]_ , \new_[6326]_ , \new_[6327]_ ,
    \new_[6331]_ , \new_[6332]_ , \new_[6335]_ , \new_[6338]_ ,
    \new_[6339]_ , \new_[6340]_ , \new_[6343]_ , \new_[6346]_ ,
    \new_[6347]_ , \new_[6350]_ , \new_[6353]_ , \new_[6354]_ ,
    \new_[6355]_ , \new_[6356]_ , \new_[6357]_ , \new_[6358]_ ,
    \new_[6362]_ , \new_[6363]_ , \new_[6366]_ , \new_[6369]_ ,
    \new_[6370]_ , \new_[6371]_ , \new_[6375]_ , \new_[6376]_ ,
    \new_[6379]_ , \new_[6382]_ , \new_[6383]_ , \new_[6384]_ ,
    \new_[6385]_ , \new_[6389]_ , \new_[6390]_ , \new_[6393]_ ,
    \new_[6396]_ , \new_[6397]_ , \new_[6398]_ , \new_[6401]_ ,
    \new_[6404]_ , \new_[6405]_ , \new_[6408]_ , \new_[6411]_ ,
    \new_[6412]_ , \new_[6413]_ , \new_[6414]_ , \new_[6415]_ ,
    \new_[6419]_ , \new_[6420]_ , \new_[6423]_ , \new_[6426]_ ,
    \new_[6427]_ , \new_[6428]_ , \new_[6432]_ , \new_[6433]_ ,
    \new_[6436]_ , \new_[6439]_ , \new_[6440]_ , \new_[6441]_ ,
    \new_[6442]_ , \new_[6446]_ , \new_[6447]_ , \new_[6450]_ ,
    \new_[6453]_ , \new_[6454]_ , \new_[6455]_ , \new_[6458]_ ,
    \new_[6461]_ , \new_[6462]_ , \new_[6465]_ , \new_[6468]_ ,
    \new_[6469]_ , \new_[6470]_ , \new_[6471]_ , \new_[6472]_ ,
    \new_[6473]_ , \new_[6474]_ , \new_[6475]_ , \new_[6476]_ ,
    \new_[6480]_ , \new_[6481]_ , \new_[6484]_ , \new_[6487]_ ,
    \new_[6488]_ , \new_[6489]_ , \new_[6493]_ , \new_[6494]_ ,
    \new_[6497]_ , \new_[6500]_ , \new_[6501]_ , \new_[6502]_ ,
    \new_[6503]_ , \new_[6507]_ , \new_[6508]_ , \new_[6511]_ ,
    \new_[6514]_ , \new_[6515]_ , \new_[6516]_ , \new_[6520]_ ,
    \new_[6521]_ , \new_[6524]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6529]_ , \new_[6530]_ , \new_[6531]_ , \new_[6535]_ ,
    \new_[6536]_ , \new_[6539]_ , \new_[6542]_ , \new_[6543]_ ,
    \new_[6544]_ , \new_[6548]_ , \new_[6549]_ , \new_[6552]_ ,
    \new_[6555]_ , \new_[6556]_ , \new_[6557]_ , \new_[6558]_ ,
    \new_[6562]_ , \new_[6563]_ , \new_[6566]_ , \new_[6569]_ ,
    \new_[6570]_ , \new_[6571]_ , \new_[6574]_ , \new_[6577]_ ,
    \new_[6578]_ , \new_[6581]_ , \new_[6584]_ , \new_[6585]_ ,
    \new_[6586]_ , \new_[6587]_ , \new_[6588]_ , \new_[6589]_ ,
    \new_[6593]_ , \new_[6594]_ , \new_[6597]_ , \new_[6600]_ ,
    \new_[6601]_ , \new_[6602]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6610]_ , \new_[6613]_ , \new_[6614]_ , \new_[6615]_ ,
    \new_[6616]_ , \new_[6620]_ , \new_[6621]_ , \new_[6624]_ ,
    \new_[6627]_ , \new_[6628]_ , \new_[6629]_ , \new_[6632]_ ,
    \new_[6635]_ , \new_[6636]_ , \new_[6639]_ , \new_[6642]_ ,
    \new_[6643]_ , \new_[6644]_ , \new_[6645]_ , \new_[6646]_ ,
    \new_[6650]_ , \new_[6651]_ , \new_[6654]_ , \new_[6657]_ ,
    \new_[6658]_ , \new_[6659]_ , \new_[6663]_ , \new_[6664]_ ,
    \new_[6667]_ , \new_[6670]_ , \new_[6671]_ , \new_[6672]_ ,
    \new_[6673]_ , \new_[6677]_ , \new_[6678]_ , \new_[6681]_ ,
    \new_[6684]_ , \new_[6685]_ , \new_[6686]_ , \new_[6689]_ ,
    \new_[6692]_ , \new_[6693]_ , \new_[6696]_ , \new_[6699]_ ,
    \new_[6700]_ , \new_[6701]_ , \new_[6702]_ , \new_[6703]_ ,
    \new_[6704]_ , \new_[6705]_ , \new_[6709]_ , \new_[6710]_ ,
    \new_[6713]_ , \new_[6716]_ , \new_[6717]_ , \new_[6718]_ ,
    \new_[6722]_ , \new_[6723]_ , \new_[6726]_ , \new_[6729]_ ,
    \new_[6730]_ , \new_[6731]_ , \new_[6732]_ , \new_[6736]_ ,
    \new_[6737]_ , \new_[6740]_ , \new_[6743]_ , \new_[6744]_ ,
    \new_[6745]_ , \new_[6748]_ , \new_[6751]_ , \new_[6752]_ ,
    \new_[6755]_ , \new_[6758]_ , \new_[6759]_ , \new_[6760]_ ,
    \new_[6761]_ , \new_[6762]_ , \new_[6766]_ , \new_[6767]_ ,
    \new_[6770]_ , \new_[6773]_ , \new_[6774]_ , \new_[6775]_ ,
    \new_[6779]_ , \new_[6780]_ , \new_[6783]_ , \new_[6786]_ ,
    \new_[6787]_ , \new_[6788]_ , \new_[6789]_ , \new_[6793]_ ,
    \new_[6794]_ , \new_[6797]_ , \new_[6800]_ , \new_[6801]_ ,
    \new_[6802]_ , \new_[6805]_ , \new_[6808]_ , \new_[6809]_ ,
    \new_[6812]_ , \new_[6815]_ , \new_[6816]_ , \new_[6817]_ ,
    \new_[6818]_ , \new_[6819]_ , \new_[6820]_ , \new_[6824]_ ,
    \new_[6825]_ , \new_[6828]_ , \new_[6831]_ , \new_[6832]_ ,
    \new_[6833]_ , \new_[6837]_ , \new_[6838]_ , \new_[6841]_ ,
    \new_[6844]_ , \new_[6845]_ , \new_[6846]_ , \new_[6847]_ ,
    \new_[6851]_ , \new_[6852]_ , \new_[6855]_ , \new_[6858]_ ,
    \new_[6859]_ , \new_[6860]_ , \new_[6863]_ , \new_[6866]_ ,
    \new_[6867]_ , \new_[6870]_ , \new_[6873]_ , \new_[6874]_ ,
    \new_[6875]_ , \new_[6876]_ , \new_[6877]_ , \new_[6881]_ ,
    \new_[6882]_ , \new_[6885]_ , \new_[6888]_ , \new_[6889]_ ,
    \new_[6890]_ , \new_[6894]_ , \new_[6895]_ , \new_[6898]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6908]_ , \new_[6909]_ , \new_[6912]_ , \new_[6915]_ ,
    \new_[6916]_ , \new_[6917]_ , \new_[6920]_ , \new_[6923]_ ,
    \new_[6924]_ , \new_[6927]_ , \new_[6930]_ , \new_[6931]_ ,
    \new_[6932]_ , \new_[6933]_ , \new_[6934]_ , \new_[6935]_ ,
    \new_[6936]_ , \new_[6937]_ , \new_[6941]_ , \new_[6942]_ ,
    \new_[6945]_ , \new_[6948]_ , \new_[6949]_ , \new_[6950]_ ,
    \new_[6954]_ , \new_[6955]_ , \new_[6958]_ , \new_[6961]_ ,
    \new_[6962]_ , \new_[6963]_ , \new_[6964]_ , \new_[6968]_ ,
    \new_[6969]_ , \new_[6972]_ , \new_[6975]_ , \new_[6976]_ ,
    \new_[6977]_ , \new_[6980]_ , \new_[6983]_ , \new_[6984]_ ,
    \new_[6987]_ , \new_[6990]_ , \new_[6991]_ , \new_[6992]_ ,
    \new_[6993]_ , \new_[6994]_ , \new_[6998]_ , \new_[6999]_ ,
    \new_[7002]_ , \new_[7005]_ , \new_[7006]_ , \new_[7007]_ ,
    \new_[7011]_ , \new_[7012]_ , \new_[7015]_ , \new_[7018]_ ,
    \new_[7019]_ , \new_[7020]_ , \new_[7021]_ , \new_[7025]_ ,
    \new_[7026]_ , \new_[7029]_ , \new_[7032]_ , \new_[7033]_ ,
    \new_[7034]_ , \new_[7037]_ , \new_[7040]_ , \new_[7041]_ ,
    \new_[7044]_ , \new_[7047]_ , \new_[7048]_ , \new_[7049]_ ,
    \new_[7050]_ , \new_[7051]_ , \new_[7052]_ , \new_[7056]_ ,
    \new_[7057]_ , \new_[7060]_ , \new_[7063]_ , \new_[7064]_ ,
    \new_[7065]_ , \new_[7069]_ , \new_[7070]_ , \new_[7073]_ ,
    \new_[7076]_ , \new_[7077]_ , \new_[7078]_ , \new_[7079]_ ,
    \new_[7083]_ , \new_[7084]_ , \new_[7087]_ , \new_[7090]_ ,
    \new_[7091]_ , \new_[7092]_ , \new_[7095]_ , \new_[7098]_ ,
    \new_[7099]_ , \new_[7102]_ , \new_[7105]_ , \new_[7106]_ ,
    \new_[7107]_ , \new_[7108]_ , \new_[7109]_ , \new_[7113]_ ,
    \new_[7114]_ , \new_[7117]_ , \new_[7120]_ , \new_[7121]_ ,
    \new_[7122]_ , \new_[7126]_ , \new_[7127]_ , \new_[7130]_ ,
    \new_[7133]_ , \new_[7134]_ , \new_[7135]_ , \new_[7136]_ ,
    \new_[7140]_ , \new_[7141]_ , \new_[7144]_ , \new_[7147]_ ,
    \new_[7148]_ , \new_[7149]_ , \new_[7152]_ , \new_[7155]_ ,
    \new_[7156]_ , \new_[7159]_ , \new_[7162]_ , \new_[7163]_ ,
    \new_[7164]_ , \new_[7165]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7168]_ , \new_[7172]_ , \new_[7173]_ , \new_[7176]_ ,
    \new_[7179]_ , \new_[7180]_ , \new_[7181]_ , \new_[7185]_ ,
    \new_[7186]_ , \new_[7189]_ , \new_[7192]_ , \new_[7193]_ ,
    \new_[7194]_ , \new_[7195]_ , \new_[7199]_ , \new_[7200]_ ,
    \new_[7203]_ , \new_[7206]_ , \new_[7207]_ , \new_[7208]_ ,
    \new_[7211]_ , \new_[7214]_ , \new_[7215]_ , \new_[7218]_ ,
    \new_[7221]_ , \new_[7222]_ , \new_[7223]_ , \new_[7224]_ ,
    \new_[7225]_ , \new_[7229]_ , \new_[7230]_ , \new_[7233]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7242]_ ,
    \new_[7243]_ , \new_[7246]_ , \new_[7249]_ , \new_[7250]_ ,
    \new_[7251]_ , \new_[7252]_ , \new_[7256]_ , \new_[7257]_ ,
    \new_[7260]_ , \new_[7263]_ , \new_[7264]_ , \new_[7265]_ ,
    \new_[7268]_ , \new_[7271]_ , \new_[7272]_ , \new_[7275]_ ,
    \new_[7278]_ , \new_[7279]_ , \new_[7280]_ , \new_[7281]_ ,
    \new_[7282]_ , \new_[7283]_ , \new_[7287]_ , \new_[7288]_ ,
    \new_[7291]_ , \new_[7294]_ , \new_[7295]_ , \new_[7296]_ ,
    \new_[7300]_ , \new_[7301]_ , \new_[7304]_ , \new_[7307]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7310]_ , \new_[7314]_ ,
    \new_[7315]_ , \new_[7318]_ , \new_[7321]_ , \new_[7322]_ ,
    \new_[7323]_ , \new_[7326]_ , \new_[7329]_ , \new_[7330]_ ,
    \new_[7333]_ , \new_[7336]_ , \new_[7337]_ , \new_[7338]_ ,
    \new_[7339]_ , \new_[7340]_ , \new_[7344]_ , \new_[7345]_ ,
    \new_[7348]_ , \new_[7351]_ , \new_[7352]_ , \new_[7353]_ ,
    \new_[7357]_ , \new_[7358]_ , \new_[7361]_ , \new_[7364]_ ,
    \new_[7365]_ , \new_[7366]_ , \new_[7367]_ , \new_[7371]_ ,
    \new_[7372]_ , \new_[7375]_ , \new_[7378]_ , \new_[7379]_ ,
    \new_[7380]_ , \new_[7383]_ , \new_[7386]_ , \new_[7387]_ ,
    \new_[7390]_ , \new_[7393]_ , \new_[7394]_ , \new_[7395]_ ,
    \new_[7396]_ , \new_[7397]_ , \new_[7398]_ , \new_[7399]_ ,
    \new_[7400]_ , \new_[7401]_ , \new_[7402]_ , \new_[7403]_ ,
    \new_[7407]_ , \new_[7408]_ , \new_[7411]_ , \new_[7414]_ ,
    \new_[7415]_ , \new_[7416]_ , \new_[7420]_ , \new_[7421]_ ,
    \new_[7424]_ , \new_[7427]_ , \new_[7428]_ , \new_[7429]_ ,
    \new_[7430]_ , \new_[7434]_ , \new_[7435]_ , \new_[7438]_ ,
    \new_[7441]_ , \new_[7442]_ , \new_[7443]_ , \new_[7447]_ ,
    \new_[7448]_ , \new_[7451]_ , \new_[7454]_ , \new_[7455]_ ,
    \new_[7456]_ , \new_[7457]_ , \new_[7458]_ , \new_[7462]_ ,
    \new_[7463]_ , \new_[7466]_ , \new_[7469]_ , \new_[7470]_ ,
    \new_[7471]_ , \new_[7475]_ , \new_[7476]_ , \new_[7479]_ ,
    \new_[7482]_ , \new_[7483]_ , \new_[7484]_ , \new_[7485]_ ,
    \new_[7489]_ , \new_[7490]_ , \new_[7493]_ , \new_[7496]_ ,
    \new_[7497]_ , \new_[7498]_ , \new_[7501]_ , \new_[7504]_ ,
    \new_[7505]_ , \new_[7508]_ , \new_[7511]_ , \new_[7512]_ ,
    \new_[7513]_ , \new_[7514]_ , \new_[7515]_ , \new_[7516]_ ,
    \new_[7520]_ , \new_[7521]_ , \new_[7524]_ , \new_[7527]_ ,
    \new_[7528]_ , \new_[7529]_ , \new_[7533]_ , \new_[7534]_ ,
    \new_[7537]_ , \new_[7540]_ , \new_[7541]_ , \new_[7542]_ ,
    \new_[7543]_ , \new_[7547]_ , \new_[7548]_ , \new_[7551]_ ,
    \new_[7554]_ , \new_[7555]_ , \new_[7556]_ , \new_[7559]_ ,
    \new_[7562]_ , \new_[7563]_ , \new_[7566]_ , \new_[7569]_ ,
    \new_[7570]_ , \new_[7571]_ , \new_[7572]_ , \new_[7573]_ ,
    \new_[7577]_ , \new_[7578]_ , \new_[7581]_ , \new_[7584]_ ,
    \new_[7585]_ , \new_[7586]_ , \new_[7590]_ , \new_[7591]_ ,
    \new_[7594]_ , \new_[7597]_ , \new_[7598]_ , \new_[7599]_ ,
    \new_[7600]_ , \new_[7604]_ , \new_[7605]_ , \new_[7608]_ ,
    \new_[7611]_ , \new_[7612]_ , \new_[7613]_ , \new_[7616]_ ,
    \new_[7619]_ , \new_[7620]_ , \new_[7623]_ , \new_[7626]_ ,
    \new_[7627]_ , \new_[7628]_ , \new_[7629]_ , \new_[7630]_ ,
    \new_[7631]_ , \new_[7632]_ , \new_[7636]_ , \new_[7637]_ ,
    \new_[7640]_ , \new_[7643]_ , \new_[7644]_ , \new_[7645]_ ,
    \new_[7649]_ , \new_[7650]_ , \new_[7653]_ , \new_[7656]_ ,
    \new_[7657]_ , \new_[7658]_ , \new_[7659]_ , \new_[7663]_ ,
    \new_[7664]_ , \new_[7667]_ , \new_[7670]_ , \new_[7671]_ ,
    \new_[7672]_ , \new_[7675]_ , \new_[7678]_ , \new_[7679]_ ,
    \new_[7682]_ , \new_[7685]_ , \new_[7686]_ , \new_[7687]_ ,
    \new_[7688]_ , \new_[7689]_ , \new_[7693]_ , \new_[7694]_ ,
    \new_[7697]_ , \new_[7700]_ , \new_[7701]_ , \new_[7702]_ ,
    \new_[7706]_ , \new_[7707]_ , \new_[7710]_ , \new_[7713]_ ,
    \new_[7714]_ , \new_[7715]_ , \new_[7716]_ , \new_[7720]_ ,
    \new_[7721]_ , \new_[7724]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7732]_ , \new_[7735]_ , \new_[7736]_ ,
    \new_[7739]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7745]_ , \new_[7746]_ , \new_[7747]_ , \new_[7751]_ ,
    \new_[7752]_ , \new_[7755]_ , \new_[7758]_ , \new_[7759]_ ,
    \new_[7760]_ , \new_[7764]_ , \new_[7765]_ , \new_[7768]_ ,
    \new_[7771]_ , \new_[7772]_ , \new_[7773]_ , \new_[7774]_ ,
    \new_[7778]_ , \new_[7779]_ , \new_[7782]_ , \new_[7785]_ ,
    \new_[7786]_ , \new_[7787]_ , \new_[7790]_ , \new_[7793]_ ,
    \new_[7794]_ , \new_[7797]_ , \new_[7800]_ , \new_[7801]_ ,
    \new_[7802]_ , \new_[7803]_ , \new_[7804]_ , \new_[7808]_ ,
    \new_[7809]_ , \new_[7812]_ , \new_[7815]_ , \new_[7816]_ ,
    \new_[7817]_ , \new_[7821]_ , \new_[7822]_ , \new_[7825]_ ,
    \new_[7828]_ , \new_[7829]_ , \new_[7830]_ , \new_[7831]_ ,
    \new_[7835]_ , \new_[7836]_ , \new_[7839]_ , \new_[7842]_ ,
    \new_[7843]_ , \new_[7844]_ , \new_[7847]_ , \new_[7850]_ ,
    \new_[7851]_ , \new_[7854]_ , \new_[7857]_ , \new_[7858]_ ,
    \new_[7859]_ , \new_[7860]_ , \new_[7861]_ , \new_[7862]_ ,
    \new_[7863]_ , \new_[7864]_ , \new_[7868]_ , \new_[7869]_ ,
    \new_[7872]_ , \new_[7875]_ , \new_[7876]_ , \new_[7877]_ ,
    \new_[7881]_ , \new_[7882]_ , \new_[7885]_ , \new_[7888]_ ,
    \new_[7889]_ , \new_[7890]_ , \new_[7891]_ , \new_[7895]_ ,
    \new_[7896]_ , \new_[7899]_ , \new_[7902]_ , \new_[7903]_ ,
    \new_[7904]_ , \new_[7908]_ , \new_[7909]_ , \new_[7912]_ ,
    \new_[7915]_ , \new_[7916]_ , \new_[7917]_ , \new_[7918]_ ,
    \new_[7919]_ , \new_[7923]_ , \new_[7924]_ , \new_[7927]_ ,
    \new_[7930]_ , \new_[7931]_ , \new_[7932]_ , \new_[7936]_ ,
    \new_[7937]_ , \new_[7940]_ , \new_[7943]_ , \new_[7944]_ ,
    \new_[7945]_ , \new_[7946]_ , \new_[7950]_ , \new_[7951]_ ,
    \new_[7954]_ , \new_[7957]_ , \new_[7958]_ , \new_[7959]_ ,
    \new_[7962]_ , \new_[7965]_ , \new_[7966]_ , \new_[7969]_ ,
    \new_[7972]_ , \new_[7973]_ , \new_[7974]_ , \new_[7975]_ ,
    \new_[7976]_ , \new_[7977]_ , \new_[7981]_ , \new_[7982]_ ,
    \new_[7985]_ , \new_[7988]_ , \new_[7989]_ , \new_[7990]_ ,
    \new_[7994]_ , \new_[7995]_ , \new_[7998]_ , \new_[8001]_ ,
    \new_[8002]_ , \new_[8003]_ , \new_[8004]_ , \new_[8008]_ ,
    \new_[8009]_ , \new_[8012]_ , \new_[8015]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8020]_ , \new_[8023]_ , \new_[8024]_ ,
    \new_[8027]_ , \new_[8030]_ , \new_[8031]_ , \new_[8032]_ ,
    \new_[8033]_ , \new_[8034]_ , \new_[8038]_ , \new_[8039]_ ,
    \new_[8042]_ , \new_[8045]_ , \new_[8046]_ , \new_[8047]_ ,
    \new_[8051]_ , \new_[8052]_ , \new_[8055]_ , \new_[8058]_ ,
    \new_[8059]_ , \new_[8060]_ , \new_[8061]_ , \new_[8065]_ ,
    \new_[8066]_ , \new_[8069]_ , \new_[8072]_ , \new_[8073]_ ,
    \new_[8074]_ , \new_[8077]_ , \new_[8080]_ , \new_[8081]_ ,
    \new_[8084]_ , \new_[8087]_ , \new_[8088]_ , \new_[8089]_ ,
    \new_[8090]_ , \new_[8091]_ , \new_[8092]_ , \new_[8093]_ ,
    \new_[8097]_ , \new_[8098]_ , \new_[8101]_ , \new_[8104]_ ,
    \new_[8105]_ , \new_[8106]_ , \new_[8110]_ , \new_[8111]_ ,
    \new_[8114]_ , \new_[8117]_ , \new_[8118]_ , \new_[8119]_ ,
    \new_[8120]_ , \new_[8124]_ , \new_[8125]_ , \new_[8128]_ ,
    \new_[8131]_ , \new_[8132]_ , \new_[8133]_ , \new_[8136]_ ,
    \new_[8139]_ , \new_[8140]_ , \new_[8143]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8148]_ , \new_[8149]_ , \new_[8150]_ ,
    \new_[8154]_ , \new_[8155]_ , \new_[8158]_ , \new_[8161]_ ,
    \new_[8162]_ , \new_[8163]_ , \new_[8167]_ , \new_[8168]_ ,
    \new_[8171]_ , \new_[8174]_ , \new_[8175]_ , \new_[8176]_ ,
    \new_[8177]_ , \new_[8181]_ , \new_[8182]_ , \new_[8185]_ ,
    \new_[8188]_ , \new_[8189]_ , \new_[8190]_ , \new_[8193]_ ,
    \new_[8196]_ , \new_[8197]_ , \new_[8200]_ , \new_[8203]_ ,
    \new_[8204]_ , \new_[8205]_ , \new_[8206]_ , \new_[8207]_ ,
    \new_[8208]_ , \new_[8212]_ , \new_[8213]_ , \new_[8216]_ ,
    \new_[8219]_ , \new_[8220]_ , \new_[8221]_ , \new_[8225]_ ,
    \new_[8226]_ , \new_[8229]_ , \new_[8232]_ , \new_[8233]_ ,
    \new_[8234]_ , \new_[8235]_ , \new_[8239]_ , \new_[8240]_ ,
    \new_[8243]_ , \new_[8246]_ , \new_[8247]_ , \new_[8248]_ ,
    \new_[8251]_ , \new_[8254]_ , \new_[8255]_ , \new_[8258]_ ,
    \new_[8261]_ , \new_[8262]_ , \new_[8263]_ , \new_[8264]_ ,
    \new_[8265]_ , \new_[8269]_ , \new_[8270]_ , \new_[8273]_ ,
    \new_[8276]_ , \new_[8277]_ , \new_[8278]_ , \new_[8282]_ ,
    \new_[8283]_ , \new_[8286]_ , \new_[8289]_ , \new_[8290]_ ,
    \new_[8291]_ , \new_[8292]_ , \new_[8296]_ , \new_[8297]_ ,
    \new_[8300]_ , \new_[8303]_ , \new_[8304]_ , \new_[8305]_ ,
    \new_[8308]_ , \new_[8311]_ , \new_[8312]_ , \new_[8315]_ ,
    \new_[8318]_ , \new_[8319]_ , \new_[8320]_ , \new_[8321]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8324]_ , \new_[8325]_ ,
    \new_[8326]_ , \new_[8330]_ , \new_[8331]_ , \new_[8334]_ ,
    \new_[8337]_ , \new_[8338]_ , \new_[8339]_ , \new_[8343]_ ,
    \new_[8344]_ , \new_[8347]_ , \new_[8350]_ , \new_[8351]_ ,
    \new_[8352]_ , \new_[8353]_ , \new_[8357]_ , \new_[8358]_ ,
    \new_[8361]_ , \new_[8364]_ , \new_[8365]_ , \new_[8366]_ ,
    \new_[8370]_ , \new_[8371]_ , \new_[8374]_ , \new_[8377]_ ,
    \new_[8378]_ , \new_[8379]_ , \new_[8380]_ , \new_[8381]_ ,
    \new_[8385]_ , \new_[8386]_ , \new_[8389]_ , \new_[8392]_ ,
    \new_[8393]_ , \new_[8394]_ , \new_[8398]_ , \new_[8399]_ ,
    \new_[8402]_ , \new_[8405]_ , \new_[8406]_ , \new_[8407]_ ,
    \new_[8408]_ , \new_[8412]_ , \new_[8413]_ , \new_[8416]_ ,
    \new_[8419]_ , \new_[8420]_ , \new_[8421]_ , \new_[8424]_ ,
    \new_[8427]_ , \new_[8428]_ , \new_[8431]_ , \new_[8434]_ ,
    \new_[8435]_ , \new_[8436]_ , \new_[8437]_ , \new_[8438]_ ,
    \new_[8439]_ , \new_[8443]_ , \new_[8444]_ , \new_[8447]_ ,
    \new_[8450]_ , \new_[8451]_ , \new_[8452]_ , \new_[8456]_ ,
    \new_[8457]_ , \new_[8460]_ , \new_[8463]_ , \new_[8464]_ ,
    \new_[8465]_ , \new_[8466]_ , \new_[8470]_ , \new_[8471]_ ,
    \new_[8474]_ , \new_[8477]_ , \new_[8478]_ , \new_[8479]_ ,
    \new_[8482]_ , \new_[8485]_ , \new_[8486]_ , \new_[8489]_ ,
    \new_[8492]_ , \new_[8493]_ , \new_[8494]_ , \new_[8495]_ ,
    \new_[8496]_ , \new_[8500]_ , \new_[8501]_ , \new_[8504]_ ,
    \new_[8507]_ , \new_[8508]_ , \new_[8509]_ , \new_[8513]_ ,
    \new_[8514]_ , \new_[8517]_ , \new_[8520]_ , \new_[8521]_ ,
    \new_[8522]_ , \new_[8523]_ , \new_[8527]_ , \new_[8528]_ ,
    \new_[8531]_ , \new_[8534]_ , \new_[8535]_ , \new_[8536]_ ,
    \new_[8539]_ , \new_[8542]_ , \new_[8543]_ , \new_[8546]_ ,
    \new_[8549]_ , \new_[8550]_ , \new_[8551]_ , \new_[8552]_ ,
    \new_[8553]_ , \new_[8554]_ , \new_[8555]_ , \new_[8559]_ ,
    \new_[8560]_ , \new_[8563]_ , \new_[8566]_ , \new_[8567]_ ,
    \new_[8568]_ , \new_[8572]_ , \new_[8573]_ , \new_[8576]_ ,
    \new_[8579]_ , \new_[8580]_ , \new_[8581]_ , \new_[8582]_ ,
    \new_[8586]_ , \new_[8587]_ , \new_[8590]_ , \new_[8593]_ ,
    \new_[8594]_ , \new_[8595]_ , \new_[8598]_ , \new_[8601]_ ,
    \new_[8602]_ , \new_[8605]_ , \new_[8608]_ , \new_[8609]_ ,
    \new_[8610]_ , \new_[8611]_ , \new_[8612]_ , \new_[8616]_ ,
    \new_[8617]_ , \new_[8620]_ , \new_[8623]_ , \new_[8624]_ ,
    \new_[8625]_ , \new_[8629]_ , \new_[8630]_ , \new_[8633]_ ,
    \new_[8636]_ , \new_[8637]_ , \new_[8638]_ , \new_[8639]_ ,
    \new_[8643]_ , \new_[8644]_ , \new_[8647]_ , \new_[8650]_ ,
    \new_[8651]_ , \new_[8652]_ , \new_[8655]_ , \new_[8658]_ ,
    \new_[8659]_ , \new_[8662]_ , \new_[8665]_ , \new_[8666]_ ,
    \new_[8667]_ , \new_[8668]_ , \new_[8669]_ , \new_[8670]_ ,
    \new_[8674]_ , \new_[8675]_ , \new_[8678]_ , \new_[8681]_ ,
    \new_[8682]_ , \new_[8683]_ , \new_[8687]_ , \new_[8688]_ ,
    \new_[8691]_ , \new_[8694]_ , \new_[8695]_ , \new_[8696]_ ,
    \new_[8697]_ , \new_[8701]_ , \new_[8702]_ , \new_[8705]_ ,
    \new_[8708]_ , \new_[8709]_ , \new_[8710]_ , \new_[8713]_ ,
    \new_[8716]_ , \new_[8717]_ , \new_[8720]_ , \new_[8723]_ ,
    \new_[8724]_ , \new_[8725]_ , \new_[8726]_ , \new_[8727]_ ,
    \new_[8731]_ , \new_[8732]_ , \new_[8735]_ , \new_[8738]_ ,
    \new_[8739]_ , \new_[8740]_ , \new_[8744]_ , \new_[8745]_ ,
    \new_[8748]_ , \new_[8751]_ , \new_[8752]_ , \new_[8753]_ ,
    \new_[8754]_ , \new_[8758]_ , \new_[8759]_ , \new_[8762]_ ,
    \new_[8765]_ , \new_[8766]_ , \new_[8767]_ , \new_[8770]_ ,
    \new_[8773]_ , \new_[8774]_ , \new_[8777]_ , \new_[8780]_ ,
    \new_[8781]_ , \new_[8782]_ , \new_[8783]_ , \new_[8784]_ ,
    \new_[8785]_ , \new_[8786]_ , \new_[8787]_ , \new_[8791]_ ,
    \new_[8792]_ , \new_[8795]_ , \new_[8798]_ , \new_[8799]_ ,
    \new_[8800]_ , \new_[8804]_ , \new_[8805]_ , \new_[8808]_ ,
    \new_[8811]_ , \new_[8812]_ , \new_[8813]_ , \new_[8814]_ ,
    \new_[8818]_ , \new_[8819]_ , \new_[8822]_ , \new_[8825]_ ,
    \new_[8826]_ , \new_[8827]_ , \new_[8830]_ , \new_[8833]_ ,
    \new_[8834]_ , \new_[8837]_ , \new_[8840]_ , \new_[8841]_ ,
    \new_[8842]_ , \new_[8843]_ , \new_[8844]_ , \new_[8848]_ ,
    \new_[8849]_ , \new_[8852]_ , \new_[8855]_ , \new_[8856]_ ,
    \new_[8857]_ , \new_[8861]_ , \new_[8862]_ , \new_[8865]_ ,
    \new_[8868]_ , \new_[8869]_ , \new_[8870]_ , \new_[8871]_ ,
    \new_[8875]_ , \new_[8876]_ , \new_[8879]_ , \new_[8882]_ ,
    \new_[8883]_ , \new_[8884]_ , \new_[8887]_ , \new_[8890]_ ,
    \new_[8891]_ , \new_[8894]_ , \new_[8897]_ , \new_[8898]_ ,
    \new_[8899]_ , \new_[8900]_ , \new_[8901]_ , \new_[8902]_ ,
    \new_[8906]_ , \new_[8907]_ , \new_[8910]_ , \new_[8913]_ ,
    \new_[8914]_ , \new_[8915]_ , \new_[8919]_ , \new_[8920]_ ,
    \new_[8923]_ , \new_[8926]_ , \new_[8927]_ , \new_[8928]_ ,
    \new_[8929]_ , \new_[8933]_ , \new_[8934]_ , \new_[8937]_ ,
    \new_[8940]_ , \new_[8941]_ , \new_[8942]_ , \new_[8945]_ ,
    \new_[8948]_ , \new_[8949]_ , \new_[8952]_ , \new_[8955]_ ,
    \new_[8956]_ , \new_[8957]_ , \new_[8958]_ , \new_[8959]_ ,
    \new_[8963]_ , \new_[8964]_ , \new_[8967]_ , \new_[8970]_ ,
    \new_[8971]_ , \new_[8972]_ , \new_[8976]_ , \new_[8977]_ ,
    \new_[8980]_ , \new_[8983]_ , \new_[8984]_ , \new_[8985]_ ,
    \new_[8986]_ , \new_[8990]_ , \new_[8991]_ , \new_[8994]_ ,
    \new_[8997]_ , \new_[8998]_ , \new_[8999]_ , \new_[9002]_ ,
    \new_[9005]_ , \new_[9006]_ , \new_[9009]_ , \new_[9012]_ ,
    \new_[9013]_ , \new_[9014]_ , \new_[9015]_ , \new_[9016]_ ,
    \new_[9017]_ , \new_[9018]_ , \new_[9022]_ , \new_[9023]_ ,
    \new_[9026]_ , \new_[9029]_ , \new_[9030]_ , \new_[9031]_ ,
    \new_[9035]_ , \new_[9036]_ , \new_[9039]_ , \new_[9042]_ ,
    \new_[9043]_ , \new_[9044]_ , \new_[9045]_ , \new_[9049]_ ,
    \new_[9050]_ , \new_[9053]_ , \new_[9056]_ , \new_[9057]_ ,
    \new_[9058]_ , \new_[9061]_ , \new_[9064]_ , \new_[9065]_ ,
    \new_[9068]_ , \new_[9071]_ , \new_[9072]_ , \new_[9073]_ ,
    \new_[9074]_ , \new_[9075]_ , \new_[9079]_ , \new_[9080]_ ,
    \new_[9083]_ , \new_[9086]_ , \new_[9087]_ , \new_[9088]_ ,
    \new_[9092]_ , \new_[9093]_ , \new_[9096]_ , \new_[9099]_ ,
    \new_[9100]_ , \new_[9101]_ , \new_[9102]_ , \new_[9106]_ ,
    \new_[9107]_ , \new_[9110]_ , \new_[9113]_ , \new_[9114]_ ,
    \new_[9115]_ , \new_[9118]_ , \new_[9121]_ , \new_[9122]_ ,
    \new_[9125]_ , \new_[9128]_ , \new_[9129]_ , \new_[9130]_ ,
    \new_[9131]_ , \new_[9132]_ , \new_[9133]_ , \new_[9137]_ ,
    \new_[9138]_ , \new_[9141]_ , \new_[9144]_ , \new_[9145]_ ,
    \new_[9146]_ , \new_[9150]_ , \new_[9151]_ , \new_[9154]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9164]_ , \new_[9165]_ , \new_[9168]_ , \new_[9171]_ ,
    \new_[9172]_ , \new_[9173]_ , \new_[9176]_ , \new_[9179]_ ,
    \new_[9180]_ , \new_[9183]_ , \new_[9186]_ , \new_[9187]_ ,
    \new_[9188]_ , \new_[9189]_ , \new_[9190]_ , \new_[9194]_ ,
    \new_[9195]_ , \new_[9198]_ , \new_[9201]_ , \new_[9202]_ ,
    \new_[9203]_ , \new_[9207]_ , \new_[9208]_ , \new_[9211]_ ,
    \new_[9214]_ , \new_[9215]_ , \new_[9216]_ , \new_[9217]_ ,
    \new_[9221]_ , \new_[9222]_ , \new_[9225]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9230]_ , \new_[9233]_ , \new_[9236]_ ,
    \new_[9237]_ , \new_[9240]_ , \new_[9243]_ , \new_[9244]_ ,
    \new_[9245]_ , \new_[9246]_ , \new_[9247]_ , \new_[9248]_ ,
    \new_[9249]_ , \new_[9250]_ , \new_[9251]_ , \new_[9252]_ ,
    \new_[9256]_ , \new_[9257]_ , \new_[9260]_ , \new_[9263]_ ,
    \new_[9264]_ , \new_[9265]_ , \new_[9269]_ , \new_[9270]_ ,
    \new_[9273]_ , \new_[9276]_ , \new_[9277]_ , \new_[9278]_ ,
    \new_[9279]_ , \new_[9283]_ , \new_[9284]_ , \new_[9287]_ ,
    \new_[9290]_ , \new_[9291]_ , \new_[9292]_ , \new_[9296]_ ,
    \new_[9297]_ , \new_[9300]_ , \new_[9303]_ , \new_[9304]_ ,
    \new_[9305]_ , \new_[9306]_ , \new_[9307]_ , \new_[9311]_ ,
    \new_[9312]_ , \new_[9315]_ , \new_[9318]_ , \new_[9319]_ ,
    \new_[9320]_ , \new_[9324]_ , \new_[9325]_ , \new_[9328]_ ,
    \new_[9331]_ , \new_[9332]_ , \new_[9333]_ , \new_[9334]_ ,
    \new_[9338]_ , \new_[9339]_ , \new_[9342]_ , \new_[9345]_ ,
    \new_[9346]_ , \new_[9347]_ , \new_[9350]_ , \new_[9353]_ ,
    \new_[9354]_ , \new_[9357]_ , \new_[9360]_ , \new_[9361]_ ,
    \new_[9362]_ , \new_[9363]_ , \new_[9364]_ , \new_[9365]_ ,
    \new_[9369]_ , \new_[9370]_ , \new_[9373]_ , \new_[9376]_ ,
    \new_[9377]_ , \new_[9378]_ , \new_[9382]_ , \new_[9383]_ ,
    \new_[9386]_ , \new_[9389]_ , \new_[9390]_ , \new_[9391]_ ,
    \new_[9392]_ , \new_[9396]_ , \new_[9397]_ , \new_[9400]_ ,
    \new_[9403]_ , \new_[9404]_ , \new_[9405]_ , \new_[9408]_ ,
    \new_[9411]_ , \new_[9412]_ , \new_[9415]_ , \new_[9418]_ ,
    \new_[9419]_ , \new_[9420]_ , \new_[9421]_ , \new_[9422]_ ,
    \new_[9426]_ , \new_[9427]_ , \new_[9430]_ , \new_[9433]_ ,
    \new_[9434]_ , \new_[9435]_ , \new_[9439]_ , \new_[9440]_ ,
    \new_[9443]_ , \new_[9446]_ , \new_[9447]_ , \new_[9448]_ ,
    \new_[9449]_ , \new_[9453]_ , \new_[9454]_ , \new_[9457]_ ,
    \new_[9460]_ , \new_[9461]_ , \new_[9462]_ , \new_[9465]_ ,
    \new_[9468]_ , \new_[9469]_ , \new_[9472]_ , \new_[9475]_ ,
    \new_[9476]_ , \new_[9477]_ , \new_[9478]_ , \new_[9479]_ ,
    \new_[9480]_ , \new_[9481]_ , \new_[9485]_ , \new_[9486]_ ,
    \new_[9489]_ , \new_[9492]_ , \new_[9493]_ , \new_[9494]_ ,
    \new_[9498]_ , \new_[9499]_ , \new_[9502]_ , \new_[9505]_ ,
    \new_[9506]_ , \new_[9507]_ , \new_[9508]_ , \new_[9512]_ ,
    \new_[9513]_ , \new_[9516]_ , \new_[9519]_ , \new_[9520]_ ,
    \new_[9521]_ , \new_[9524]_ , \new_[9527]_ , \new_[9528]_ ,
    \new_[9531]_ , \new_[9534]_ , \new_[9535]_ , \new_[9536]_ ,
    \new_[9537]_ , \new_[9538]_ , \new_[9542]_ , \new_[9543]_ ,
    \new_[9546]_ , \new_[9549]_ , \new_[9550]_ , \new_[9551]_ ,
    \new_[9555]_ , \new_[9556]_ , \new_[9559]_ , \new_[9562]_ ,
    \new_[9563]_ , \new_[9564]_ , \new_[9565]_ , \new_[9569]_ ,
    \new_[9570]_ , \new_[9573]_ , \new_[9576]_ , \new_[9577]_ ,
    \new_[9578]_ , \new_[9581]_ , \new_[9584]_ , \new_[9585]_ ,
    \new_[9588]_ , \new_[9591]_ , \new_[9592]_ , \new_[9593]_ ,
    \new_[9594]_ , \new_[9595]_ , \new_[9596]_ , \new_[9600]_ ,
    \new_[9601]_ , \new_[9604]_ , \new_[9607]_ , \new_[9608]_ ,
    \new_[9609]_ , \new_[9613]_ , \new_[9614]_ , \new_[9617]_ ,
    \new_[9620]_ , \new_[9621]_ , \new_[9622]_ , \new_[9623]_ ,
    \new_[9627]_ , \new_[9628]_ , \new_[9631]_ , \new_[9634]_ ,
    \new_[9635]_ , \new_[9636]_ , \new_[9639]_ , \new_[9642]_ ,
    \new_[9643]_ , \new_[9646]_ , \new_[9649]_ , \new_[9650]_ ,
    \new_[9651]_ , \new_[9652]_ , \new_[9653]_ , \new_[9657]_ ,
    \new_[9658]_ , \new_[9661]_ , \new_[9664]_ , \new_[9665]_ ,
    \new_[9666]_ , \new_[9670]_ , \new_[9671]_ , \new_[9674]_ ,
    \new_[9677]_ , \new_[9678]_ , \new_[9679]_ , \new_[9680]_ ,
    \new_[9684]_ , \new_[9685]_ , \new_[9688]_ , \new_[9691]_ ,
    \new_[9692]_ , \new_[9693]_ , \new_[9696]_ , \new_[9699]_ ,
    \new_[9700]_ , \new_[9703]_ , \new_[9706]_ , \new_[9707]_ ,
    \new_[9708]_ , \new_[9709]_ , \new_[9710]_ , \new_[9711]_ ,
    \new_[9712]_ , \new_[9713]_ , \new_[9717]_ , \new_[9718]_ ,
    \new_[9721]_ , \new_[9724]_ , \new_[9725]_ , \new_[9726]_ ,
    \new_[9730]_ , \new_[9731]_ , \new_[9734]_ , \new_[9737]_ ,
    \new_[9738]_ , \new_[9739]_ , \new_[9740]_ , \new_[9744]_ ,
    \new_[9745]_ , \new_[9748]_ , \new_[9751]_ , \new_[9752]_ ,
    \new_[9753]_ , \new_[9756]_ , \new_[9759]_ , \new_[9760]_ ,
    \new_[9763]_ , \new_[9766]_ , \new_[9767]_ , \new_[9768]_ ,
    \new_[9769]_ , \new_[9770]_ , \new_[9774]_ , \new_[9775]_ ,
    \new_[9778]_ , \new_[9781]_ , \new_[9782]_ , \new_[9783]_ ,
    \new_[9787]_ , \new_[9788]_ , \new_[9791]_ , \new_[9794]_ ,
    \new_[9795]_ , \new_[9796]_ , \new_[9797]_ , \new_[9801]_ ,
    \new_[9802]_ , \new_[9805]_ , \new_[9808]_ , \new_[9809]_ ,
    \new_[9810]_ , \new_[9813]_ , \new_[9816]_ , \new_[9817]_ ,
    \new_[9820]_ , \new_[9823]_ , \new_[9824]_ , \new_[9825]_ ,
    \new_[9826]_ , \new_[9827]_ , \new_[9828]_ , \new_[9832]_ ,
    \new_[9833]_ , \new_[9836]_ , \new_[9839]_ , \new_[9840]_ ,
    \new_[9841]_ , \new_[9845]_ , \new_[9846]_ , \new_[9849]_ ,
    \new_[9852]_ , \new_[9853]_ , \new_[9854]_ , \new_[9855]_ ,
    \new_[9859]_ , \new_[9860]_ , \new_[9863]_ , \new_[9866]_ ,
    \new_[9867]_ , \new_[9868]_ , \new_[9871]_ , \new_[9874]_ ,
    \new_[9875]_ , \new_[9878]_ , \new_[9881]_ , \new_[9882]_ ,
    \new_[9883]_ , \new_[9884]_ , \new_[9885]_ , \new_[9889]_ ,
    \new_[9890]_ , \new_[9893]_ , \new_[9896]_ , \new_[9897]_ ,
    \new_[9898]_ , \new_[9902]_ , \new_[9903]_ , \new_[9906]_ ,
    \new_[9909]_ , \new_[9910]_ , \new_[9911]_ , \new_[9912]_ ,
    \new_[9916]_ , \new_[9917]_ , \new_[9920]_ , \new_[9923]_ ,
    \new_[9924]_ , \new_[9925]_ , \new_[9928]_ , \new_[9931]_ ,
    \new_[9932]_ , \new_[9935]_ , \new_[9938]_ , \new_[9939]_ ,
    \new_[9940]_ , \new_[9941]_ , \new_[9942]_ , \new_[9943]_ ,
    \new_[9944]_ , \new_[9948]_ , \new_[9949]_ , \new_[9952]_ ,
    \new_[9955]_ , \new_[9956]_ , \new_[9957]_ , \new_[9961]_ ,
    \new_[9962]_ , \new_[9965]_ , \new_[9968]_ , \new_[9969]_ ,
    \new_[9970]_ , \new_[9971]_ , \new_[9975]_ , \new_[9976]_ ,
    \new_[9979]_ , \new_[9982]_ , \new_[9983]_ , \new_[9984]_ ,
    \new_[9987]_ , \new_[9990]_ , \new_[9991]_ , \new_[9994]_ ,
    \new_[9997]_ , \new_[9998]_ , \new_[9999]_ , \new_[10000]_ ,
    \new_[10001]_ , \new_[10005]_ , \new_[10006]_ , \new_[10009]_ ,
    \new_[10012]_ , \new_[10013]_ , \new_[10014]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10022]_ , \new_[10025]_ , \new_[10026]_ ,
    \new_[10027]_ , \new_[10028]_ , \new_[10032]_ , \new_[10033]_ ,
    \new_[10036]_ , \new_[10039]_ , \new_[10040]_ , \new_[10041]_ ,
    \new_[10044]_ , \new_[10047]_ , \new_[10048]_ , \new_[10051]_ ,
    \new_[10054]_ , \new_[10055]_ , \new_[10056]_ , \new_[10057]_ ,
    \new_[10058]_ , \new_[10059]_ , \new_[10063]_ , \new_[10064]_ ,
    \new_[10067]_ , \new_[10070]_ , \new_[10071]_ , \new_[10072]_ ,
    \new_[10076]_ , \new_[10077]_ , \new_[10080]_ , \new_[10083]_ ,
    \new_[10084]_ , \new_[10085]_ , \new_[10086]_ , \new_[10090]_ ,
    \new_[10091]_ , \new_[10094]_ , \new_[10097]_ , \new_[10098]_ ,
    \new_[10099]_ , \new_[10102]_ , \new_[10105]_ , \new_[10106]_ ,
    \new_[10109]_ , \new_[10112]_ , \new_[10113]_ , \new_[10114]_ ,
    \new_[10115]_ , \new_[10116]_ , \new_[10120]_ , \new_[10121]_ ,
    \new_[10124]_ , \new_[10127]_ , \new_[10128]_ , \new_[10129]_ ,
    \new_[10133]_ , \new_[10134]_ , \new_[10137]_ , \new_[10140]_ ,
    \new_[10141]_ , \new_[10142]_ , \new_[10143]_ , \new_[10147]_ ,
    \new_[10148]_ , \new_[10151]_ , \new_[10154]_ , \new_[10155]_ ,
    \new_[10156]_ , \new_[10159]_ , \new_[10162]_ , \new_[10163]_ ,
    \new_[10166]_ , \new_[10169]_ , \new_[10170]_ , \new_[10171]_ ,
    \new_[10172]_ , \new_[10173]_ , \new_[10174]_ , \new_[10175]_ ,
    \new_[10176]_ , \new_[10177]_ , \new_[10181]_ , \new_[10182]_ ,
    \new_[10185]_ , \new_[10188]_ , \new_[10189]_ , \new_[10190]_ ,
    \new_[10194]_ , \new_[10195]_ , \new_[10198]_ , \new_[10201]_ ,
    \new_[10202]_ , \new_[10203]_ , \new_[10204]_ , \new_[10208]_ ,
    \new_[10209]_ , \new_[10212]_ , \new_[10215]_ , \new_[10216]_ ,
    \new_[10217]_ , \new_[10221]_ , \new_[10222]_ , \new_[10225]_ ,
    \new_[10228]_ , \new_[10229]_ , \new_[10230]_ , \new_[10231]_ ,
    \new_[10232]_ , \new_[10236]_ , \new_[10237]_ , \new_[10240]_ ,
    \new_[10243]_ , \new_[10244]_ , \new_[10245]_ , \new_[10249]_ ,
    \new_[10250]_ , \new_[10253]_ , \new_[10256]_ , \new_[10257]_ ,
    \new_[10258]_ , \new_[10259]_ , \new_[10263]_ , \new_[10264]_ ,
    \new_[10267]_ , \new_[10270]_ , \new_[10271]_ , \new_[10272]_ ,
    \new_[10275]_ , \new_[10278]_ , \new_[10279]_ , \new_[10282]_ ,
    \new_[10285]_ , \new_[10286]_ , \new_[10287]_ , \new_[10288]_ ,
    \new_[10289]_ , \new_[10290]_ , \new_[10294]_ , \new_[10295]_ ,
    \new_[10298]_ , \new_[10301]_ , \new_[10302]_ , \new_[10303]_ ,
    \new_[10307]_ , \new_[10308]_ , \new_[10311]_ , \new_[10314]_ ,
    \new_[10315]_ , \new_[10316]_ , \new_[10317]_ , \new_[10321]_ ,
    \new_[10322]_ , \new_[10325]_ , \new_[10328]_ , \new_[10329]_ ,
    \new_[10330]_ , \new_[10333]_ , \new_[10336]_ , \new_[10337]_ ,
    \new_[10340]_ , \new_[10343]_ , \new_[10344]_ , \new_[10345]_ ,
    \new_[10346]_ , \new_[10347]_ , \new_[10351]_ , \new_[10352]_ ,
    \new_[10355]_ , \new_[10358]_ , \new_[10359]_ , \new_[10360]_ ,
    \new_[10364]_ , \new_[10365]_ , \new_[10368]_ , \new_[10371]_ ,
    \new_[10372]_ , \new_[10373]_ , \new_[10374]_ , \new_[10378]_ ,
    \new_[10379]_ , \new_[10382]_ , \new_[10385]_ , \new_[10386]_ ,
    \new_[10387]_ , \new_[10390]_ , \new_[10393]_ , \new_[10394]_ ,
    \new_[10397]_ , \new_[10400]_ , \new_[10401]_ , \new_[10402]_ ,
    \new_[10403]_ , \new_[10404]_ , \new_[10405]_ , \new_[10406]_ ,
    \new_[10410]_ , \new_[10411]_ , \new_[10414]_ , \new_[10417]_ ,
    \new_[10418]_ , \new_[10419]_ , \new_[10423]_ , \new_[10424]_ ,
    \new_[10427]_ , \new_[10430]_ , \new_[10431]_ , \new_[10432]_ ,
    \new_[10433]_ , \new_[10437]_ , \new_[10438]_ , \new_[10441]_ ,
    \new_[10444]_ , \new_[10445]_ , \new_[10446]_ , \new_[10449]_ ,
    \new_[10452]_ , \new_[10453]_ , \new_[10456]_ , \new_[10459]_ ,
    \new_[10460]_ , \new_[10461]_ , \new_[10462]_ , \new_[10463]_ ,
    \new_[10467]_ , \new_[10468]_ , \new_[10471]_ , \new_[10474]_ ,
    \new_[10475]_ , \new_[10476]_ , \new_[10480]_ , \new_[10481]_ ,
    \new_[10484]_ , \new_[10487]_ , \new_[10488]_ , \new_[10489]_ ,
    \new_[10490]_ , \new_[10494]_ , \new_[10495]_ , \new_[10498]_ ,
    \new_[10501]_ , \new_[10502]_ , \new_[10503]_ , \new_[10506]_ ,
    \new_[10509]_ , \new_[10510]_ , \new_[10513]_ , \new_[10516]_ ,
    \new_[10517]_ , \new_[10518]_ , \new_[10519]_ , \new_[10520]_ ,
    \new_[10521]_ , \new_[10525]_ , \new_[10526]_ , \new_[10529]_ ,
    \new_[10532]_ , \new_[10533]_ , \new_[10534]_ , \new_[10538]_ ,
    \new_[10539]_ , \new_[10542]_ , \new_[10545]_ , \new_[10546]_ ,
    \new_[10547]_ , \new_[10548]_ , \new_[10552]_ , \new_[10553]_ ,
    \new_[10556]_ , \new_[10559]_ , \new_[10560]_ , \new_[10561]_ ,
    \new_[10564]_ , \new_[10567]_ , \new_[10568]_ , \new_[10571]_ ,
    \new_[10574]_ , \new_[10575]_ , \new_[10576]_ , \new_[10577]_ ,
    \new_[10578]_ , \new_[10582]_ , \new_[10583]_ , \new_[10586]_ ,
    \new_[10589]_ , \new_[10590]_ , \new_[10591]_ , \new_[10595]_ ,
    \new_[10596]_ , \new_[10599]_ , \new_[10602]_ , \new_[10603]_ ,
    \new_[10604]_ , \new_[10605]_ , \new_[10609]_ , \new_[10610]_ ,
    \new_[10613]_ , \new_[10616]_ , \new_[10617]_ , \new_[10618]_ ,
    \new_[10621]_ , \new_[10624]_ , \new_[10625]_ , \new_[10628]_ ,
    \new_[10631]_ , \new_[10632]_ , \new_[10633]_ , \new_[10634]_ ,
    \new_[10635]_ , \new_[10636]_ , \new_[10637]_ , \new_[10638]_ ,
    \new_[10642]_ , \new_[10643]_ , \new_[10646]_ , \new_[10649]_ ,
    \new_[10650]_ , \new_[10651]_ , \new_[10655]_ , \new_[10656]_ ,
    \new_[10659]_ , \new_[10662]_ , \new_[10663]_ , \new_[10664]_ ,
    \new_[10665]_ , \new_[10669]_ , \new_[10670]_ , \new_[10673]_ ,
    \new_[10676]_ , \new_[10677]_ , \new_[10678]_ , \new_[10681]_ ,
    \new_[10684]_ , \new_[10685]_ , \new_[10688]_ , \new_[10691]_ ,
    \new_[10692]_ , \new_[10693]_ , \new_[10694]_ , \new_[10695]_ ,
    \new_[10699]_ , \new_[10700]_ , \new_[10703]_ , \new_[10706]_ ,
    \new_[10707]_ , \new_[10708]_ , \new_[10712]_ , \new_[10713]_ ,
    \new_[10716]_ , \new_[10719]_ , \new_[10720]_ , \new_[10721]_ ,
    \new_[10722]_ , \new_[10726]_ , \new_[10727]_ , \new_[10730]_ ,
    \new_[10733]_ , \new_[10734]_ , \new_[10735]_ , \new_[10738]_ ,
    \new_[10741]_ , \new_[10742]_ , \new_[10745]_ , \new_[10748]_ ,
    \new_[10749]_ , \new_[10750]_ , \new_[10751]_ , \new_[10752]_ ,
    \new_[10753]_ , \new_[10757]_ , \new_[10758]_ , \new_[10761]_ ,
    \new_[10764]_ , \new_[10765]_ , \new_[10766]_ , \new_[10770]_ ,
    \new_[10771]_ , \new_[10774]_ , \new_[10777]_ , \new_[10778]_ ,
    \new_[10779]_ , \new_[10780]_ , \new_[10784]_ , \new_[10785]_ ,
    \new_[10788]_ , \new_[10791]_ , \new_[10792]_ , \new_[10793]_ ,
    \new_[10796]_ , \new_[10799]_ , \new_[10800]_ , \new_[10803]_ ,
    \new_[10806]_ , \new_[10807]_ , \new_[10808]_ , \new_[10809]_ ,
    \new_[10810]_ , \new_[10814]_ , \new_[10815]_ , \new_[10818]_ ,
    \new_[10821]_ , \new_[10822]_ , \new_[10823]_ , \new_[10827]_ ,
    \new_[10828]_ , \new_[10831]_ , \new_[10834]_ , \new_[10835]_ ,
    \new_[10836]_ , \new_[10837]_ , \new_[10841]_ , \new_[10842]_ ,
    \new_[10845]_ , \new_[10848]_ , \new_[10849]_ , \new_[10850]_ ,
    \new_[10853]_ , \new_[10856]_ , \new_[10857]_ , \new_[10860]_ ,
    \new_[10863]_ , \new_[10864]_ , \new_[10865]_ , \new_[10866]_ ,
    \new_[10867]_ , \new_[10868]_ , \new_[10869]_ , \new_[10873]_ ,
    \new_[10874]_ , \new_[10877]_ , \new_[10880]_ , \new_[10881]_ ,
    \new_[10882]_ , \new_[10886]_ , \new_[10887]_ , \new_[10890]_ ,
    \new_[10893]_ , \new_[10894]_ , \new_[10895]_ , \new_[10896]_ ,
    \new_[10900]_ , \new_[10901]_ , \new_[10904]_ , \new_[10907]_ ,
    \new_[10908]_ , \new_[10909]_ , \new_[10912]_ , \new_[10915]_ ,
    \new_[10916]_ , \new_[10919]_ , \new_[10922]_ , \new_[10923]_ ,
    \new_[10924]_ , \new_[10925]_ , \new_[10926]_ , \new_[10930]_ ,
    \new_[10931]_ , \new_[10934]_ , \new_[10937]_ , \new_[10938]_ ,
    \new_[10939]_ , \new_[10943]_ , \new_[10944]_ , \new_[10947]_ ,
    \new_[10950]_ , \new_[10951]_ , \new_[10952]_ , \new_[10953]_ ,
    \new_[10957]_ , \new_[10958]_ , \new_[10961]_ , \new_[10964]_ ,
    \new_[10965]_ , \new_[10966]_ , \new_[10969]_ , \new_[10972]_ ,
    \new_[10973]_ , \new_[10976]_ , \new_[10979]_ , \new_[10980]_ ,
    \new_[10981]_ , \new_[10982]_ , \new_[10983]_ , \new_[10984]_ ,
    \new_[10988]_ , \new_[10989]_ , \new_[10992]_ , \new_[10995]_ ,
    \new_[10996]_ , \new_[10997]_ , \new_[11001]_ , \new_[11002]_ ,
    \new_[11005]_ , \new_[11008]_ , \new_[11009]_ , \new_[11010]_ ,
    \new_[11011]_ , \new_[11015]_ , \new_[11016]_ , \new_[11019]_ ,
    \new_[11022]_ , \new_[11023]_ , \new_[11024]_ , \new_[11027]_ ,
    \new_[11030]_ , \new_[11031]_ , \new_[11034]_ , \new_[11037]_ ,
    \new_[11038]_ , \new_[11039]_ , \new_[11040]_ , \new_[11041]_ ,
    \new_[11045]_ , \new_[11046]_ , \new_[11049]_ , \new_[11052]_ ,
    \new_[11053]_ , \new_[11054]_ , \new_[11058]_ , \new_[11059]_ ,
    \new_[11062]_ , \new_[11065]_ , \new_[11066]_ , \new_[11067]_ ,
    \new_[11068]_ , \new_[11072]_ , \new_[11073]_ , \new_[11076]_ ,
    \new_[11079]_ , \new_[11080]_ , \new_[11081]_ , \new_[11084]_ ,
    \new_[11087]_ , \new_[11088]_ , \new_[11091]_ , \new_[11094]_ ,
    \new_[11095]_ , \new_[11096]_ , \new_[11097]_ , \new_[11098]_ ,
    \new_[11099]_ , \new_[11100]_ , \new_[11101]_ , \new_[11102]_ ,
    \new_[11103]_ , \new_[11104]_ , \new_[11107]_ , \new_[11110]_ ,
    \new_[11111]_ , \new_[11114]_ , \new_[11117]_ , \new_[11118]_ ,
    \new_[11121]_ , \new_[11124]_ , \new_[11125]_ , \new_[11128]_ ,
    \new_[11131]_ , \new_[11132]_ , \new_[11135]_ , \new_[11138]_ ,
    \new_[11139]_ , \new_[11142]_ , \new_[11145]_ , \new_[11146]_ ,
    \new_[11149]_ , \new_[11152]_ , \new_[11153]_ , \new_[11156]_ ,
    \new_[11159]_ , \new_[11160]_ , \new_[11163]_ , \new_[11166]_ ,
    \new_[11167]_ , \new_[11170]_ , \new_[11173]_ , \new_[11174]_ ,
    \new_[11177]_ , \new_[11180]_ , \new_[11181]_ , \new_[11184]_ ,
    \new_[11187]_ , \new_[11188]_ , \new_[11191]_ , \new_[11194]_ ,
    \new_[11195]_ , \new_[11198]_ , \new_[11201]_ , \new_[11202]_ ,
    \new_[11205]_ , \new_[11208]_ , \new_[11209]_ , \new_[11212]_ ,
    \new_[11215]_ , \new_[11216]_ , \new_[11219]_ , \new_[11222]_ ,
    \new_[11223]_ , \new_[11226]_ , \new_[11229]_ , \new_[11230]_ ,
    \new_[11233]_ , \new_[11236]_ , \new_[11237]_ , \new_[11240]_ ,
    \new_[11243]_ , \new_[11244]_ , \new_[11247]_ , \new_[11250]_ ,
    \new_[11251]_ , \new_[11254]_ , \new_[11257]_ , \new_[11258]_ ,
    \new_[11261]_ , \new_[11264]_ , \new_[11265]_ , \new_[11268]_ ,
    \new_[11271]_ , \new_[11272]_ , \new_[11275]_ , \new_[11278]_ ,
    \new_[11279]_ , \new_[11282]_ , \new_[11285]_ , \new_[11286]_ ,
    \new_[11289]_ , \new_[11292]_ , \new_[11293]_ , \new_[11296]_ ,
    \new_[11299]_ , \new_[11300]_ , \new_[11303]_ , \new_[11306]_ ,
    \new_[11307]_ , \new_[11310]_ , \new_[11313]_ , \new_[11314]_ ,
    \new_[11317]_ , \new_[11320]_ , \new_[11321]_ , \new_[11324]_ ,
    \new_[11327]_ , \new_[11328]_ , \new_[11331]_ , \new_[11334]_ ,
    \new_[11335]_ , \new_[11338]_ , \new_[11341]_ , \new_[11342]_ ,
    \new_[11345]_ , \new_[11348]_ , \new_[11349]_ , \new_[11352]_ ,
    \new_[11355]_ , \new_[11356]_ , \new_[11359]_ , \new_[11362]_ ,
    \new_[11363]_ , \new_[11366]_ , \new_[11369]_ , \new_[11370]_ ,
    \new_[11373]_ , \new_[11376]_ , \new_[11377]_ , \new_[11380]_ ,
    \new_[11383]_ , \new_[11384]_ , \new_[11387]_ , \new_[11390]_ ,
    \new_[11391]_ , \new_[11394]_ , \new_[11397]_ , \new_[11398]_ ,
    \new_[11401]_ , \new_[11404]_ , \new_[11405]_ , \new_[11408]_ ,
    \new_[11411]_ , \new_[11412]_ , \new_[11415]_ , \new_[11418]_ ,
    \new_[11419]_ , \new_[11422]_ , \new_[11425]_ , \new_[11426]_ ,
    \new_[11429]_ , \new_[11432]_ , \new_[11433]_ , \new_[11436]_ ,
    \new_[11439]_ , \new_[11440]_ , \new_[11443]_ , \new_[11446]_ ,
    \new_[11447]_ , \new_[11450]_ , \new_[11453]_ , \new_[11454]_ ,
    \new_[11457]_ , \new_[11460]_ , \new_[11461]_ , \new_[11464]_ ,
    \new_[11467]_ , \new_[11468]_ , \new_[11471]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11478]_ , \new_[11481]_ , \new_[11482]_ ,
    \new_[11485]_ , \new_[11488]_ , \new_[11489]_ , \new_[11492]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11499]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11506]_ , \new_[11509]_ , \new_[11510]_ ,
    \new_[11513]_ , \new_[11516]_ , \new_[11517]_ , \new_[11520]_ ,
    \new_[11523]_ , \new_[11524]_ , \new_[11527]_ , \new_[11530]_ ,
    \new_[11531]_ , \new_[11534]_ , \new_[11537]_ , \new_[11538]_ ,
    \new_[11541]_ , \new_[11544]_ , \new_[11545]_ , \new_[11548]_ ,
    \new_[11551]_ , \new_[11552]_ , \new_[11555]_ , \new_[11558]_ ,
    \new_[11559]_ , \new_[11562]_ , \new_[11566]_ , \new_[11567]_ ,
    \new_[11568]_ , \new_[11571]_ , \new_[11574]_ , \new_[11575]_ ,
    \new_[11578]_ , \new_[11582]_ , \new_[11583]_ , \new_[11584]_ ,
    \new_[11587]_ , \new_[11590]_ , \new_[11591]_ , \new_[11594]_ ,
    \new_[11598]_ , \new_[11599]_ , \new_[11600]_ , \new_[11603]_ ,
    \new_[11606]_ , \new_[11607]_ , \new_[11610]_ , \new_[11614]_ ,
    \new_[11615]_ , \new_[11616]_ , \new_[11619]_ , \new_[11622]_ ,
    \new_[11623]_ , \new_[11626]_ , \new_[11630]_ , \new_[11631]_ ,
    \new_[11632]_ , \new_[11635]_ , \new_[11638]_ , \new_[11639]_ ,
    \new_[11642]_ , \new_[11646]_ , \new_[11647]_ , \new_[11648]_ ,
    \new_[11651]_ , \new_[11654]_ , \new_[11655]_ , \new_[11658]_ ,
    \new_[11662]_ , \new_[11663]_ , \new_[11664]_ , \new_[11667]_ ,
    \new_[11670]_ , \new_[11671]_ , \new_[11674]_ , \new_[11678]_ ,
    \new_[11679]_ , \new_[11680]_ , \new_[11683]_ , \new_[11686]_ ,
    \new_[11687]_ , \new_[11690]_ , \new_[11694]_ , \new_[11695]_ ,
    \new_[11696]_ , \new_[11699]_ , \new_[11702]_ , \new_[11703]_ ,
    \new_[11706]_ , \new_[11710]_ , \new_[11711]_ , \new_[11712]_ ,
    \new_[11715]_ , \new_[11718]_ , \new_[11719]_ , \new_[11722]_ ,
    \new_[11726]_ , \new_[11727]_ , \new_[11728]_ , \new_[11731]_ ,
    \new_[11734]_ , \new_[11735]_ , \new_[11738]_ , \new_[11742]_ ,
    \new_[11743]_ , \new_[11744]_ , \new_[11747]_ , \new_[11750]_ ,
    \new_[11751]_ , \new_[11754]_ , \new_[11758]_ , \new_[11759]_ ,
    \new_[11760]_ , \new_[11763]_ , \new_[11766]_ , \new_[11767]_ ,
    \new_[11770]_ , \new_[11774]_ , \new_[11775]_ , \new_[11776]_ ,
    \new_[11779]_ , \new_[11782]_ , \new_[11783]_ , \new_[11786]_ ,
    \new_[11790]_ , \new_[11791]_ , \new_[11792]_ , \new_[11795]_ ,
    \new_[11798]_ , \new_[11799]_ , \new_[11802]_ , \new_[11806]_ ,
    \new_[11807]_ , \new_[11808]_ , \new_[11811]_ , \new_[11814]_ ,
    \new_[11815]_ , \new_[11818]_ , \new_[11822]_ , \new_[11823]_ ,
    \new_[11824]_ , \new_[11827]_ , \new_[11830]_ , \new_[11831]_ ,
    \new_[11834]_ , \new_[11838]_ , \new_[11839]_ , \new_[11840]_ ,
    \new_[11843]_ , \new_[11846]_ , \new_[11847]_ , \new_[11850]_ ,
    \new_[11854]_ , \new_[11855]_ , \new_[11856]_ , \new_[11859]_ ,
    \new_[11862]_ , \new_[11863]_ , \new_[11866]_ , \new_[11870]_ ,
    \new_[11871]_ , \new_[11872]_ , \new_[11875]_ , \new_[11878]_ ,
    \new_[11879]_ , \new_[11882]_ , \new_[11886]_ , \new_[11887]_ ,
    \new_[11888]_ , \new_[11891]_ , \new_[11894]_ , \new_[11895]_ ,
    \new_[11898]_ , \new_[11902]_ , \new_[11903]_ , \new_[11904]_ ,
    \new_[11907]_ , \new_[11910]_ , \new_[11911]_ , \new_[11914]_ ,
    \new_[11918]_ , \new_[11919]_ , \new_[11920]_ , \new_[11923]_ ,
    \new_[11926]_ , \new_[11927]_ , \new_[11930]_ , \new_[11934]_ ,
    \new_[11935]_ , \new_[11936]_ , \new_[11939]_ , \new_[11942]_ ,
    \new_[11943]_ , \new_[11946]_ , \new_[11950]_ , \new_[11951]_ ,
    \new_[11952]_ , \new_[11955]_ , \new_[11958]_ , \new_[11959]_ ,
    \new_[11962]_ , \new_[11966]_ , \new_[11967]_ , \new_[11968]_ ,
    \new_[11971]_ , \new_[11974]_ , \new_[11975]_ , \new_[11978]_ ,
    \new_[11982]_ , \new_[11983]_ , \new_[11984]_ , \new_[11987]_ ,
    \new_[11990]_ , \new_[11991]_ , \new_[11994]_ , \new_[11998]_ ,
    \new_[11999]_ , \new_[12000]_ , \new_[12003]_ , \new_[12006]_ ,
    \new_[12007]_ , \new_[12010]_ , \new_[12014]_ , \new_[12015]_ ,
    \new_[12016]_ , \new_[12019]_ , \new_[12022]_ , \new_[12023]_ ,
    \new_[12026]_ , \new_[12030]_ , \new_[12031]_ , \new_[12032]_ ,
    \new_[12035]_ , \new_[12038]_ , \new_[12039]_ , \new_[12042]_ ,
    \new_[12046]_ , \new_[12047]_ , \new_[12048]_ , \new_[12051]_ ,
    \new_[12054]_ , \new_[12055]_ , \new_[12058]_ , \new_[12062]_ ,
    \new_[12063]_ , \new_[12064]_ , \new_[12067]_ , \new_[12071]_ ,
    \new_[12072]_ , \new_[12073]_ , \new_[12076]_ , \new_[12080]_ ,
    \new_[12081]_ , \new_[12082]_ , \new_[12085]_ , \new_[12089]_ ,
    \new_[12090]_ , \new_[12091]_ , \new_[12094]_ , \new_[12098]_ ,
    \new_[12099]_ , \new_[12100]_ , \new_[12103]_ , \new_[12107]_ ,
    \new_[12108]_ , \new_[12109]_ , \new_[12112]_ , \new_[12116]_ ,
    \new_[12117]_ , \new_[12118]_ , \new_[12121]_ , \new_[12125]_ ,
    \new_[12126]_ , \new_[12127]_ , \new_[12130]_ , \new_[12134]_ ,
    \new_[12135]_ , \new_[12136]_ , \new_[12139]_ , \new_[12143]_ ,
    \new_[12144]_ , \new_[12145]_ , \new_[12148]_ , \new_[12152]_ ,
    \new_[12153]_ , \new_[12154]_ , \new_[12157]_ , \new_[12161]_ ,
    \new_[12162]_ , \new_[12163]_ , \new_[12166]_ , \new_[12170]_ ,
    \new_[12171]_ , \new_[12172]_ , \new_[12175]_ , \new_[12179]_ ,
    \new_[12180]_ , \new_[12181]_ , \new_[12184]_ , \new_[12188]_ ,
    \new_[12189]_ , \new_[12190]_ , \new_[12193]_ , \new_[12197]_ ,
    \new_[12198]_ , \new_[12199]_ , \new_[12202]_ , \new_[12206]_ ,
    \new_[12207]_ , \new_[12208]_ , \new_[12211]_ , \new_[12215]_ ,
    \new_[12216]_ , \new_[12217]_ , \new_[12220]_ , \new_[12224]_ ,
    \new_[12225]_ , \new_[12226]_ , \new_[12229]_ , \new_[12233]_ ,
    \new_[12234]_ , \new_[12235]_ , \new_[12238]_ , \new_[12242]_ ,
    \new_[12243]_ , \new_[12244]_ , \new_[12247]_ , \new_[12251]_ ,
    \new_[12252]_ , \new_[12253]_ , \new_[12256]_ , \new_[12260]_ ,
    \new_[12261]_ , \new_[12262]_ , \new_[12265]_ , \new_[12269]_ ,
    \new_[12270]_ , \new_[12271]_ , \new_[12274]_ , \new_[12278]_ ,
    \new_[12279]_ , \new_[12280]_ , \new_[12283]_ , \new_[12287]_ ,
    \new_[12288]_ , \new_[12289]_ , \new_[12292]_ , \new_[12296]_ ,
    \new_[12297]_ , \new_[12298]_ , \new_[12301]_ , \new_[12305]_ ,
    \new_[12306]_ , \new_[12307]_ , \new_[12310]_ , \new_[12314]_ ,
    \new_[12315]_ , \new_[12316]_ , \new_[12319]_ , \new_[12323]_ ,
    \new_[12324]_ , \new_[12325]_ , \new_[12328]_ , \new_[12332]_ ,
    \new_[12333]_ , \new_[12334]_ , \new_[12337]_ , \new_[12341]_ ,
    \new_[12342]_ , \new_[12343]_ , \new_[12346]_ , \new_[12350]_ ,
    \new_[12351]_ , \new_[12352]_ , \new_[12355]_ , \new_[12359]_ ,
    \new_[12360]_ , \new_[12361]_ , \new_[12364]_ , \new_[12368]_ ,
    \new_[12369]_ , \new_[12370]_ , \new_[12373]_ , \new_[12377]_ ,
    \new_[12378]_ , \new_[12379]_ , \new_[12382]_ , \new_[12386]_ ,
    \new_[12387]_ , \new_[12388]_ , \new_[12391]_ , \new_[12395]_ ,
    \new_[12396]_ , \new_[12397]_ , \new_[12400]_ , \new_[12404]_ ,
    \new_[12405]_ , \new_[12406]_ , \new_[12409]_ , \new_[12413]_ ,
    \new_[12414]_ , \new_[12415]_ , \new_[12418]_ , \new_[12422]_ ,
    \new_[12423]_ , \new_[12424]_ , \new_[12427]_ , \new_[12431]_ ,
    \new_[12432]_ , \new_[12433]_ , \new_[12436]_ , \new_[12440]_ ,
    \new_[12441]_ , \new_[12442]_ , \new_[12445]_ , \new_[12449]_ ,
    \new_[12450]_ , \new_[12451]_ , \new_[12454]_ , \new_[12458]_ ,
    \new_[12459]_ , \new_[12460]_ , \new_[12463]_ , \new_[12467]_ ,
    \new_[12468]_ , \new_[12469]_ , \new_[12472]_ , \new_[12476]_ ,
    \new_[12477]_ , \new_[12478]_ , \new_[12481]_ , \new_[12485]_ ,
    \new_[12486]_ , \new_[12487]_ , \new_[12490]_ , \new_[12494]_ ,
    \new_[12495]_ , \new_[12496]_ , \new_[12499]_ , \new_[12503]_ ,
    \new_[12504]_ , \new_[12505]_ , \new_[12508]_ , \new_[12512]_ ,
    \new_[12513]_ , \new_[12514]_ , \new_[12517]_ , \new_[12521]_ ,
    \new_[12522]_ , \new_[12523]_ , \new_[12526]_ , \new_[12530]_ ,
    \new_[12531]_ , \new_[12532]_ , \new_[12535]_ , \new_[12539]_ ,
    \new_[12540]_ , \new_[12541]_ , \new_[12544]_ , \new_[12548]_ ,
    \new_[12549]_ , \new_[12550]_ , \new_[12553]_ , \new_[12557]_ ,
    \new_[12558]_ , \new_[12559]_ , \new_[12562]_ , \new_[12566]_ ,
    \new_[12567]_ , \new_[12568]_ , \new_[12571]_ , \new_[12575]_ ,
    \new_[12576]_ , \new_[12577]_ , \new_[12580]_ , \new_[12584]_ ,
    \new_[12585]_ , \new_[12586]_ , \new_[12589]_ , \new_[12593]_ ,
    \new_[12594]_ , \new_[12595]_ , \new_[12598]_ , \new_[12602]_ ,
    \new_[12603]_ , \new_[12604]_ , \new_[12607]_ , \new_[12611]_ ,
    \new_[12612]_ , \new_[12613]_ , \new_[12616]_ , \new_[12620]_ ,
    \new_[12621]_ , \new_[12622]_ , \new_[12625]_ , \new_[12629]_ ,
    \new_[12630]_ , \new_[12631]_ , \new_[12634]_ , \new_[12638]_ ,
    \new_[12639]_ , \new_[12640]_ , \new_[12643]_ , \new_[12647]_ ,
    \new_[12648]_ , \new_[12649]_ , \new_[12652]_ , \new_[12656]_ ,
    \new_[12657]_ , \new_[12658]_ , \new_[12661]_ , \new_[12665]_ ,
    \new_[12666]_ , \new_[12667]_ , \new_[12670]_ , \new_[12674]_ ,
    \new_[12675]_ , \new_[12676]_ , \new_[12679]_ , \new_[12683]_ ,
    \new_[12684]_ , \new_[12685]_ , \new_[12688]_ , \new_[12692]_ ,
    \new_[12693]_ , \new_[12694]_ , \new_[12697]_ , \new_[12701]_ ,
    \new_[12702]_ , \new_[12703]_ , \new_[12706]_ , \new_[12710]_ ,
    \new_[12711]_ , \new_[12712]_ , \new_[12715]_ , \new_[12719]_ ,
    \new_[12720]_ , \new_[12721]_ , \new_[12724]_ , \new_[12728]_ ,
    \new_[12729]_ , \new_[12730]_ , \new_[12733]_ , \new_[12737]_ ,
    \new_[12738]_ , \new_[12739]_ , \new_[12742]_ , \new_[12746]_ ,
    \new_[12747]_ , \new_[12748]_ , \new_[12751]_ , \new_[12755]_ ,
    \new_[12756]_ , \new_[12757]_ , \new_[12760]_ , \new_[12764]_ ,
    \new_[12765]_ , \new_[12766]_ , \new_[12769]_ , \new_[12773]_ ,
    \new_[12774]_ , \new_[12775]_ , \new_[12778]_ , \new_[12782]_ ,
    \new_[12783]_ , \new_[12784]_ , \new_[12787]_ , \new_[12791]_ ,
    \new_[12792]_ , \new_[12793]_ , \new_[12796]_ , \new_[12800]_ ,
    \new_[12801]_ , \new_[12802]_ , \new_[12805]_ , \new_[12809]_ ,
    \new_[12810]_ , \new_[12811]_ , \new_[12814]_ , \new_[12818]_ ,
    \new_[12819]_ , \new_[12820]_ , \new_[12823]_ , \new_[12827]_ ,
    \new_[12828]_ , \new_[12829]_ , \new_[12832]_ , \new_[12836]_ ,
    \new_[12837]_ , \new_[12838]_ , \new_[12841]_ , \new_[12845]_ ,
    \new_[12846]_ , \new_[12847]_ , \new_[12850]_ , \new_[12854]_ ,
    \new_[12855]_ , \new_[12856]_ , \new_[12859]_ , \new_[12863]_ ,
    \new_[12864]_ , \new_[12865]_ , \new_[12868]_ , \new_[12872]_ ,
    \new_[12873]_ , \new_[12874]_ , \new_[12877]_ , \new_[12881]_ ,
    \new_[12882]_ , \new_[12883]_ , \new_[12886]_ , \new_[12890]_ ,
    \new_[12891]_ , \new_[12892]_ , \new_[12895]_ , \new_[12899]_ ,
    \new_[12900]_ , \new_[12901]_ , \new_[12904]_ , \new_[12908]_ ,
    \new_[12909]_ , \new_[12910]_ , \new_[12913]_ , \new_[12917]_ ,
    \new_[12918]_ , \new_[12919]_ , \new_[12922]_ , \new_[12926]_ ,
    \new_[12927]_ , \new_[12928]_ , \new_[12931]_ , \new_[12935]_ ,
    \new_[12936]_ , \new_[12937]_ , \new_[12940]_ , \new_[12944]_ ,
    \new_[12945]_ , \new_[12946]_ , \new_[12949]_ , \new_[12953]_ ,
    \new_[12954]_ , \new_[12955]_ , \new_[12958]_ , \new_[12962]_ ,
    \new_[12963]_ , \new_[12964]_ , \new_[12967]_ , \new_[12971]_ ,
    \new_[12972]_ , \new_[12973]_ , \new_[12976]_ , \new_[12980]_ ,
    \new_[12981]_ , \new_[12982]_ , \new_[12985]_ , \new_[12989]_ ,
    \new_[12990]_ , \new_[12991]_ , \new_[12994]_ , \new_[12998]_ ,
    \new_[12999]_ , \new_[13000]_ , \new_[13003]_ , \new_[13007]_ ,
    \new_[13008]_ , \new_[13009]_ , \new_[13012]_ , \new_[13016]_ ,
    \new_[13017]_ , \new_[13018]_ , \new_[13021]_ , \new_[13025]_ ,
    \new_[13026]_ , \new_[13027]_ , \new_[13030]_ , \new_[13034]_ ,
    \new_[13035]_ , \new_[13036]_ , \new_[13039]_ , \new_[13043]_ ,
    \new_[13044]_ , \new_[13045]_ , \new_[13048]_ , \new_[13052]_ ,
    \new_[13053]_ , \new_[13054]_ , \new_[13057]_ , \new_[13061]_ ,
    \new_[13062]_ , \new_[13063]_ , \new_[13066]_ , \new_[13070]_ ,
    \new_[13071]_ , \new_[13072]_ , \new_[13075]_ , \new_[13079]_ ,
    \new_[13080]_ , \new_[13081]_ , \new_[13084]_ , \new_[13088]_ ,
    \new_[13089]_ , \new_[13090]_ , \new_[13093]_ , \new_[13097]_ ,
    \new_[13098]_ , \new_[13099]_ , \new_[13102]_ , \new_[13106]_ ,
    \new_[13107]_ , \new_[13108]_ , \new_[13111]_ , \new_[13115]_ ,
    \new_[13116]_ , \new_[13117]_ , \new_[13120]_ , \new_[13124]_ ,
    \new_[13125]_ , \new_[13126]_ , \new_[13129]_ , \new_[13133]_ ,
    \new_[13134]_ , \new_[13135]_ , \new_[13138]_ , \new_[13142]_ ,
    \new_[13143]_ , \new_[13144]_ , \new_[13147]_ , \new_[13151]_ ,
    \new_[13152]_ , \new_[13153]_ , \new_[13156]_ , \new_[13160]_ ,
    \new_[13161]_ , \new_[13162]_ , \new_[13165]_ , \new_[13169]_ ,
    \new_[13170]_ , \new_[13171]_ , \new_[13174]_ , \new_[13178]_ ,
    \new_[13179]_ , \new_[13180]_ , \new_[13183]_ , \new_[13187]_ ,
    \new_[13188]_ , \new_[13189]_ , \new_[13192]_ , \new_[13196]_ ,
    \new_[13197]_ , \new_[13198]_ , \new_[13201]_ , \new_[13205]_ ,
    \new_[13206]_ , \new_[13207]_ , \new_[13210]_ , \new_[13214]_ ,
    \new_[13215]_ , \new_[13216]_ , \new_[13219]_ , \new_[13223]_ ,
    \new_[13224]_ , \new_[13225]_ , \new_[13228]_ , \new_[13232]_ ,
    \new_[13233]_ , \new_[13234]_ , \new_[13237]_ , \new_[13241]_ ,
    \new_[13242]_ , \new_[13243]_ , \new_[13246]_ , \new_[13250]_ ,
    \new_[13251]_ , \new_[13252]_ , \new_[13255]_ , \new_[13259]_ ,
    \new_[13260]_ , \new_[13261]_ , \new_[13264]_ , \new_[13268]_ ,
    \new_[13269]_ , \new_[13270]_ , \new_[13273]_ , \new_[13277]_ ,
    \new_[13278]_ , \new_[13279]_ , \new_[13282]_ , \new_[13286]_ ,
    \new_[13287]_ , \new_[13288]_ , \new_[13291]_ , \new_[13295]_ ,
    \new_[13296]_ , \new_[13297]_ , \new_[13300]_ , \new_[13304]_ ,
    \new_[13305]_ , \new_[13306]_ , \new_[13309]_ , \new_[13313]_ ,
    \new_[13314]_ , \new_[13315]_ , \new_[13318]_ , \new_[13322]_ ,
    \new_[13323]_ , \new_[13324]_ , \new_[13327]_ , \new_[13331]_ ,
    \new_[13332]_ , \new_[13333]_ , \new_[13336]_ , \new_[13340]_ ,
    \new_[13341]_ , \new_[13342]_ , \new_[13345]_ , \new_[13349]_ ,
    \new_[13350]_ , \new_[13351]_ , \new_[13354]_ , \new_[13358]_ ,
    \new_[13359]_ , \new_[13360]_ , \new_[13363]_ , \new_[13367]_ ,
    \new_[13368]_ , \new_[13369]_ , \new_[13372]_ , \new_[13376]_ ,
    \new_[13377]_ , \new_[13378]_ , \new_[13381]_ , \new_[13385]_ ,
    \new_[13386]_ , \new_[13387]_ , \new_[13390]_ , \new_[13394]_ ,
    \new_[13395]_ , \new_[13396]_ , \new_[13399]_ , \new_[13403]_ ,
    \new_[13404]_ , \new_[13405]_ , \new_[13408]_ , \new_[13412]_ ,
    \new_[13413]_ , \new_[13414]_ , \new_[13417]_ , \new_[13421]_ ,
    \new_[13422]_ , \new_[13423]_ , \new_[13426]_ , \new_[13430]_ ,
    \new_[13431]_ , \new_[13432]_ , \new_[13435]_ , \new_[13439]_ ,
    \new_[13440]_ , \new_[13441]_ , \new_[13444]_ , \new_[13448]_ ,
    \new_[13449]_ , \new_[13450]_ , \new_[13453]_ , \new_[13457]_ ,
    \new_[13458]_ , \new_[13459]_ , \new_[13462]_ , \new_[13466]_ ,
    \new_[13467]_ , \new_[13468]_ , \new_[13471]_ , \new_[13475]_ ,
    \new_[13476]_ , \new_[13477]_ , \new_[13480]_ , \new_[13484]_ ,
    \new_[13485]_ , \new_[13486]_ , \new_[13489]_ , \new_[13493]_ ,
    \new_[13494]_ , \new_[13495]_ , \new_[13498]_ , \new_[13502]_ ,
    \new_[13503]_ , \new_[13504]_ , \new_[13507]_ , \new_[13511]_ ,
    \new_[13512]_ , \new_[13513]_ , \new_[13516]_ , \new_[13520]_ ,
    \new_[13521]_ , \new_[13522]_ , \new_[13525]_ , \new_[13529]_ ,
    \new_[13530]_ , \new_[13531]_ , \new_[13534]_ , \new_[13538]_ ,
    \new_[13539]_ , \new_[13540]_ , \new_[13543]_ , \new_[13547]_ ,
    \new_[13548]_ , \new_[13549]_ , \new_[13552]_ , \new_[13556]_ ,
    \new_[13557]_ , \new_[13558]_ , \new_[13561]_ , \new_[13565]_ ,
    \new_[13566]_ , \new_[13567]_ , \new_[13570]_ , \new_[13574]_ ,
    \new_[13575]_ , \new_[13576]_ , \new_[13579]_ , \new_[13583]_ ,
    \new_[13584]_ , \new_[13585]_ , \new_[13588]_ , \new_[13592]_ ,
    \new_[13593]_ , \new_[13594]_ , \new_[13597]_ , \new_[13601]_ ,
    \new_[13602]_ , \new_[13603]_ , \new_[13606]_ , \new_[13610]_ ,
    \new_[13611]_ , \new_[13612]_ , \new_[13615]_ , \new_[13619]_ ,
    \new_[13620]_ , \new_[13621]_ , \new_[13624]_ , \new_[13628]_ ,
    \new_[13629]_ , \new_[13630]_ , \new_[13633]_ , \new_[13637]_ ,
    \new_[13638]_ , \new_[13639]_ , \new_[13642]_ , \new_[13646]_ ,
    \new_[13647]_ , \new_[13648]_ , \new_[13651]_ , \new_[13655]_ ,
    \new_[13656]_ , \new_[13657]_ , \new_[13660]_ , \new_[13664]_ ,
    \new_[13665]_ , \new_[13666]_ , \new_[13669]_ , \new_[13673]_ ,
    \new_[13674]_ , \new_[13675]_ , \new_[13678]_ , \new_[13682]_ ,
    \new_[13683]_ , \new_[13684]_ , \new_[13687]_ , \new_[13691]_ ,
    \new_[13692]_ , \new_[13693]_ , \new_[13696]_ , \new_[13700]_ ,
    \new_[13701]_ , \new_[13702]_ , \new_[13705]_ , \new_[13709]_ ,
    \new_[13710]_ , \new_[13711]_ , \new_[13714]_ , \new_[13718]_ ,
    \new_[13719]_ , \new_[13720]_ , \new_[13723]_ , \new_[13727]_ ,
    \new_[13728]_ , \new_[13729]_ , \new_[13732]_ , \new_[13736]_ ,
    \new_[13737]_ , \new_[13738]_ , \new_[13741]_ , \new_[13745]_ ,
    \new_[13746]_ , \new_[13747]_ , \new_[13750]_ , \new_[13754]_ ,
    \new_[13755]_ , \new_[13756]_ , \new_[13759]_ , \new_[13763]_ ,
    \new_[13764]_ , \new_[13765]_ , \new_[13768]_ , \new_[13772]_ ,
    \new_[13773]_ , \new_[13774]_ , \new_[13777]_ , \new_[13781]_ ,
    \new_[13782]_ , \new_[13783]_ , \new_[13786]_ , \new_[13790]_ ,
    \new_[13791]_ , \new_[13792]_ , \new_[13795]_ , \new_[13799]_ ,
    \new_[13800]_ , \new_[13801]_ , \new_[13804]_ , \new_[13808]_ ,
    \new_[13809]_ , \new_[13810]_ , \new_[13813]_ , \new_[13817]_ ,
    \new_[13818]_ , \new_[13819]_ , \new_[13822]_ , \new_[13826]_ ,
    \new_[13827]_ , \new_[13828]_ , \new_[13831]_ , \new_[13835]_ ,
    \new_[13836]_ , \new_[13837]_ , \new_[13840]_ , \new_[13844]_ ,
    \new_[13845]_ , \new_[13846]_ , \new_[13849]_ , \new_[13853]_ ,
    \new_[13854]_ , \new_[13855]_ , \new_[13858]_ , \new_[13862]_ ,
    \new_[13863]_ , \new_[13864]_ , \new_[13867]_ , \new_[13871]_ ,
    \new_[13872]_ , \new_[13873]_ , \new_[13876]_ , \new_[13880]_ ,
    \new_[13881]_ , \new_[13882]_ , \new_[13885]_ , \new_[13889]_ ,
    \new_[13890]_ , \new_[13891]_ , \new_[13894]_ , \new_[13898]_ ,
    \new_[13899]_ , \new_[13900]_ , \new_[13903]_ , \new_[13907]_ ,
    \new_[13908]_ , \new_[13909]_ , \new_[13912]_ , \new_[13916]_ ,
    \new_[13917]_ , \new_[13918]_ , \new_[13921]_ , \new_[13925]_ ,
    \new_[13926]_ , \new_[13927]_ , \new_[13930]_ , \new_[13934]_ ,
    \new_[13935]_ , \new_[13936]_ , \new_[13939]_ , \new_[13943]_ ,
    \new_[13944]_ , \new_[13945]_ , \new_[13948]_ , \new_[13952]_ ,
    \new_[13953]_ , \new_[13954]_ , \new_[13957]_ , \new_[13961]_ ,
    \new_[13962]_ , \new_[13963]_ , \new_[13966]_ , \new_[13970]_ ,
    \new_[13971]_ , \new_[13972]_ , \new_[13975]_ , \new_[13979]_ ,
    \new_[13980]_ , \new_[13981]_ , \new_[13984]_ , \new_[13988]_ ,
    \new_[13989]_ , \new_[13990]_ , \new_[13993]_ , \new_[13997]_ ,
    \new_[13998]_ , \new_[13999]_ , \new_[14002]_ , \new_[14006]_ ,
    \new_[14007]_ , \new_[14008]_ , \new_[14011]_ , \new_[14015]_ ,
    \new_[14016]_ , \new_[14017]_ , \new_[14020]_ , \new_[14024]_ ,
    \new_[14025]_ , \new_[14026]_ , \new_[14029]_ , \new_[14033]_ ,
    \new_[14034]_ , \new_[14035]_ , \new_[14038]_ , \new_[14042]_ ,
    \new_[14043]_ , \new_[14044]_ , \new_[14047]_ , \new_[14051]_ ,
    \new_[14052]_ , \new_[14053]_ , \new_[14056]_ , \new_[14060]_ ,
    \new_[14061]_ , \new_[14062]_ , \new_[14065]_ , \new_[14069]_ ,
    \new_[14070]_ , \new_[14071]_ , \new_[14074]_ , \new_[14078]_ ,
    \new_[14079]_ , \new_[14080]_ , \new_[14083]_ , \new_[14087]_ ,
    \new_[14088]_ , \new_[14089]_ , \new_[14092]_ , \new_[14096]_ ,
    \new_[14097]_ , \new_[14098]_ , \new_[14101]_ , \new_[14105]_ ,
    \new_[14106]_ , \new_[14107]_ , \new_[14110]_ , \new_[14114]_ ,
    \new_[14115]_ , \new_[14116]_ , \new_[14119]_ , \new_[14123]_ ,
    \new_[14124]_ , \new_[14125]_ , \new_[14128]_ , \new_[14132]_ ,
    \new_[14133]_ , \new_[14134]_ , \new_[14137]_ , \new_[14141]_ ,
    \new_[14142]_ , \new_[14143]_ , \new_[14146]_ , \new_[14150]_ ,
    \new_[14151]_ , \new_[14152]_ , \new_[14155]_ , \new_[14159]_ ,
    \new_[14160]_ , \new_[14161]_ , \new_[14164]_ , \new_[14168]_ ,
    \new_[14169]_ , \new_[14170]_ , \new_[14173]_ , \new_[14177]_ ,
    \new_[14178]_ , \new_[14179]_ , \new_[14182]_ , \new_[14186]_ ,
    \new_[14187]_ , \new_[14188]_ , \new_[14191]_ , \new_[14195]_ ,
    \new_[14196]_ , \new_[14197]_ , \new_[14200]_ , \new_[14204]_ ,
    \new_[14205]_ , \new_[14206]_ , \new_[14209]_ , \new_[14213]_ ,
    \new_[14214]_ , \new_[14215]_ , \new_[14218]_ , \new_[14222]_ ,
    \new_[14223]_ , \new_[14224]_ , \new_[14227]_ , \new_[14231]_ ,
    \new_[14232]_ , \new_[14233]_ , \new_[14236]_ , \new_[14240]_ ,
    \new_[14241]_ , \new_[14242]_ , \new_[14245]_ , \new_[14249]_ ,
    \new_[14250]_ , \new_[14251]_ , \new_[14254]_ , \new_[14258]_ ,
    \new_[14259]_ , \new_[14260]_ , \new_[14263]_ , \new_[14267]_ ,
    \new_[14268]_ , \new_[14269]_ , \new_[14272]_ , \new_[14276]_ ,
    \new_[14277]_ , \new_[14278]_ , \new_[14281]_ , \new_[14285]_ ,
    \new_[14286]_ , \new_[14287]_ , \new_[14290]_ , \new_[14294]_ ,
    \new_[14295]_ , \new_[14296]_ , \new_[14299]_ , \new_[14303]_ ,
    \new_[14304]_ , \new_[14305]_ , \new_[14308]_ , \new_[14312]_ ,
    \new_[14313]_ , \new_[14314]_ , \new_[14317]_ , \new_[14321]_ ,
    \new_[14322]_ , \new_[14323]_ , \new_[14326]_ , \new_[14330]_ ,
    \new_[14331]_ , \new_[14332]_ , \new_[14335]_ , \new_[14339]_ ,
    \new_[14340]_ , \new_[14341]_ , \new_[14344]_ , \new_[14348]_ ,
    \new_[14349]_ , \new_[14350]_ , \new_[14353]_ , \new_[14357]_ ,
    \new_[14358]_ , \new_[14359]_ , \new_[14362]_ , \new_[14366]_ ,
    \new_[14367]_ , \new_[14368]_ , \new_[14371]_ , \new_[14375]_ ,
    \new_[14376]_ , \new_[14377]_ , \new_[14380]_ , \new_[14384]_ ,
    \new_[14385]_ , \new_[14386]_ , \new_[14389]_ , \new_[14393]_ ,
    \new_[14394]_ , \new_[14395]_ , \new_[14398]_ , \new_[14402]_ ,
    \new_[14403]_ , \new_[14404]_ , \new_[14407]_ , \new_[14411]_ ,
    \new_[14412]_ , \new_[14413]_ , \new_[14416]_ , \new_[14420]_ ,
    \new_[14421]_ , \new_[14422]_ , \new_[14425]_ , \new_[14429]_ ,
    \new_[14430]_ , \new_[14431]_ , \new_[14434]_ , \new_[14438]_ ,
    \new_[14439]_ , \new_[14440]_ , \new_[14443]_ , \new_[14447]_ ,
    \new_[14448]_ , \new_[14449]_ , \new_[14452]_ , \new_[14456]_ ,
    \new_[14457]_ , \new_[14458]_ , \new_[14461]_ , \new_[14465]_ ,
    \new_[14466]_ , \new_[14467]_ , \new_[14470]_ , \new_[14474]_ ,
    \new_[14475]_ , \new_[14476]_ , \new_[14479]_ , \new_[14483]_ ,
    \new_[14484]_ , \new_[14485]_ , \new_[14488]_ , \new_[14492]_ ,
    \new_[14493]_ , \new_[14494]_ , \new_[14497]_ , \new_[14501]_ ,
    \new_[14502]_ , \new_[14503]_ , \new_[14506]_ , \new_[14510]_ ,
    \new_[14511]_ , \new_[14512]_ , \new_[14515]_ , \new_[14519]_ ,
    \new_[14520]_ , \new_[14521]_ , \new_[14524]_ , \new_[14528]_ ,
    \new_[14529]_ , \new_[14530]_ , \new_[14533]_ , \new_[14537]_ ,
    \new_[14538]_ , \new_[14539]_ , \new_[14542]_ , \new_[14546]_ ,
    \new_[14547]_ , \new_[14548]_ , \new_[14551]_ , \new_[14555]_ ,
    \new_[14556]_ , \new_[14557]_ , \new_[14560]_ , \new_[14564]_ ,
    \new_[14565]_ , \new_[14566]_ , \new_[14569]_ , \new_[14573]_ ,
    \new_[14574]_ , \new_[14575]_ , \new_[14578]_ , \new_[14582]_ ,
    \new_[14583]_ , \new_[14584]_ , \new_[14587]_ , \new_[14591]_ ,
    \new_[14592]_ , \new_[14593]_ , \new_[14596]_ , \new_[14600]_ ,
    \new_[14601]_ , \new_[14602]_ , \new_[14605]_ , \new_[14609]_ ,
    \new_[14610]_ , \new_[14611]_ , \new_[14614]_ , \new_[14618]_ ,
    \new_[14619]_ , \new_[14620]_ , \new_[14623]_ , \new_[14627]_ ,
    \new_[14628]_ , \new_[14629]_ , \new_[14632]_ , \new_[14636]_ ,
    \new_[14637]_ , \new_[14638]_ , \new_[14641]_ , \new_[14645]_ ,
    \new_[14646]_ , \new_[14647]_ , \new_[14650]_ , \new_[14654]_ ,
    \new_[14655]_ , \new_[14656]_ , \new_[14659]_ , \new_[14663]_ ,
    \new_[14664]_ , \new_[14665]_ , \new_[14668]_ , \new_[14672]_ ,
    \new_[14673]_ , \new_[14674]_ , \new_[14677]_ , \new_[14681]_ ,
    \new_[14682]_ , \new_[14683]_ , \new_[14686]_ , \new_[14690]_ ,
    \new_[14691]_ , \new_[14692]_ , \new_[14695]_ , \new_[14699]_ ,
    \new_[14700]_ , \new_[14701]_ , \new_[14704]_ , \new_[14708]_ ,
    \new_[14709]_ , \new_[14710]_ , \new_[14713]_ , \new_[14717]_ ,
    \new_[14718]_ , \new_[14719]_ , \new_[14722]_ , \new_[14726]_ ,
    \new_[14727]_ , \new_[14728]_ , \new_[14731]_ , \new_[14735]_ ,
    \new_[14736]_ , \new_[14737]_ , \new_[14740]_ , \new_[14744]_ ,
    \new_[14745]_ , \new_[14746]_ , \new_[14749]_ , \new_[14753]_ ,
    \new_[14754]_ , \new_[14755]_ , \new_[14758]_ , \new_[14762]_ ,
    \new_[14763]_ , \new_[14764]_ , \new_[14767]_ , \new_[14771]_ ,
    \new_[14772]_ , \new_[14773]_ , \new_[14776]_ , \new_[14780]_ ,
    \new_[14781]_ , \new_[14782]_ , \new_[14785]_ , \new_[14789]_ ,
    \new_[14790]_ , \new_[14791]_ , \new_[14794]_ , \new_[14798]_ ,
    \new_[14799]_ , \new_[14800]_ , \new_[14803]_ , \new_[14807]_ ,
    \new_[14808]_ , \new_[14809]_ , \new_[14812]_ , \new_[14816]_ ,
    \new_[14817]_ , \new_[14818]_ , \new_[14821]_ , \new_[14825]_ ,
    \new_[14826]_ , \new_[14827]_ , \new_[14830]_ , \new_[14834]_ ,
    \new_[14835]_ , \new_[14836]_ , \new_[14839]_ , \new_[14843]_ ,
    \new_[14844]_ , \new_[14845]_ , \new_[14848]_ , \new_[14852]_ ,
    \new_[14853]_ , \new_[14854]_ , \new_[14857]_ , \new_[14861]_ ,
    \new_[14862]_ , \new_[14863]_ , \new_[14866]_ , \new_[14870]_ ,
    \new_[14871]_ , \new_[14872]_ , \new_[14875]_ , \new_[14879]_ ,
    \new_[14880]_ , \new_[14881]_ , \new_[14884]_ , \new_[14888]_ ,
    \new_[14889]_ , \new_[14890]_ , \new_[14893]_ , \new_[14897]_ ,
    \new_[14898]_ , \new_[14899]_ , \new_[14902]_ , \new_[14906]_ ,
    \new_[14907]_ , \new_[14908]_ , \new_[14911]_ , \new_[14915]_ ,
    \new_[14916]_ , \new_[14917]_ , \new_[14920]_ , \new_[14924]_ ,
    \new_[14925]_ , \new_[14926]_ , \new_[14929]_ , \new_[14933]_ ,
    \new_[14934]_ , \new_[14935]_ , \new_[14938]_ , \new_[14942]_ ,
    \new_[14943]_ , \new_[14944]_ , \new_[14947]_ , \new_[14951]_ ,
    \new_[14952]_ , \new_[14953]_ , \new_[14956]_ , \new_[14960]_ ,
    \new_[14961]_ , \new_[14962]_ , \new_[14965]_ , \new_[14969]_ ,
    \new_[14970]_ , \new_[14971]_ , \new_[14974]_ , \new_[14978]_ ,
    \new_[14979]_ , \new_[14980]_ , \new_[14983]_ , \new_[14987]_ ,
    \new_[14988]_ , \new_[14989]_ , \new_[14992]_ , \new_[14996]_ ,
    \new_[14997]_ , \new_[14998]_ , \new_[15001]_ , \new_[15005]_ ,
    \new_[15006]_ , \new_[15007]_ , \new_[15010]_ , \new_[15014]_ ,
    \new_[15015]_ , \new_[15016]_ , \new_[15019]_ , \new_[15023]_ ,
    \new_[15024]_ , \new_[15025]_ , \new_[15028]_ , \new_[15032]_ ,
    \new_[15033]_ , \new_[15034]_ , \new_[15037]_ , \new_[15041]_ ,
    \new_[15042]_ , \new_[15043]_ , \new_[15046]_ , \new_[15050]_ ,
    \new_[15051]_ , \new_[15052]_ , \new_[15055]_ , \new_[15059]_ ,
    \new_[15060]_ , \new_[15061]_ , \new_[15064]_ , \new_[15068]_ ,
    \new_[15069]_ , \new_[15070]_ , \new_[15073]_ , \new_[15077]_ ,
    \new_[15078]_ , \new_[15079]_ , \new_[15082]_ , \new_[15086]_ ,
    \new_[15087]_ , \new_[15088]_ , \new_[15091]_ , \new_[15095]_ ,
    \new_[15096]_ , \new_[15097]_ , \new_[15100]_ , \new_[15104]_ ,
    \new_[15105]_ , \new_[15106]_ , \new_[15109]_ , \new_[15113]_ ,
    \new_[15114]_ , \new_[15115]_ , \new_[15118]_ , \new_[15122]_ ,
    \new_[15123]_ , \new_[15124]_ , \new_[15127]_ , \new_[15131]_ ,
    \new_[15132]_ , \new_[15133]_ , \new_[15136]_ , \new_[15140]_ ,
    \new_[15141]_ , \new_[15142]_ , \new_[15145]_ , \new_[15149]_ ,
    \new_[15150]_ , \new_[15151]_ , \new_[15154]_ , \new_[15158]_ ,
    \new_[15159]_ , \new_[15160]_ , \new_[15163]_ , \new_[15167]_ ,
    \new_[15168]_ , \new_[15169]_ , \new_[15172]_ , \new_[15176]_ ,
    \new_[15177]_ , \new_[15178]_ , \new_[15181]_ , \new_[15185]_ ,
    \new_[15186]_ , \new_[15187]_ , \new_[15190]_ , \new_[15194]_ ,
    \new_[15195]_ , \new_[15196]_ , \new_[15199]_ , \new_[15203]_ ,
    \new_[15204]_ , \new_[15205]_ , \new_[15208]_ , \new_[15212]_ ,
    \new_[15213]_ , \new_[15214]_ , \new_[15217]_ , \new_[15221]_ ,
    \new_[15222]_ , \new_[15223]_ , \new_[15226]_ , \new_[15230]_ ,
    \new_[15231]_ , \new_[15232]_ , \new_[15235]_ , \new_[15239]_ ,
    \new_[15240]_ , \new_[15241]_ , \new_[15244]_ , \new_[15248]_ ,
    \new_[15249]_ , \new_[15250]_ , \new_[15253]_ , \new_[15257]_ ,
    \new_[15258]_ , \new_[15259]_ , \new_[15262]_ , \new_[15266]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15271]_ , \new_[15275]_ ,
    \new_[15276]_ , \new_[15277]_ , \new_[15280]_ , \new_[15284]_ ,
    \new_[15285]_ , \new_[15286]_ , \new_[15289]_ , \new_[15293]_ ,
    \new_[15294]_ , \new_[15295]_ , \new_[15298]_ , \new_[15302]_ ,
    \new_[15303]_ , \new_[15304]_ , \new_[15307]_ , \new_[15311]_ ,
    \new_[15312]_ , \new_[15313]_ , \new_[15316]_ , \new_[15320]_ ,
    \new_[15321]_ , \new_[15322]_ , \new_[15325]_ , \new_[15329]_ ,
    \new_[15330]_ , \new_[15331]_ , \new_[15334]_ , \new_[15338]_ ,
    \new_[15339]_ , \new_[15340]_ , \new_[15343]_ , \new_[15347]_ ,
    \new_[15348]_ , \new_[15349]_ , \new_[15352]_ , \new_[15356]_ ,
    \new_[15357]_ , \new_[15358]_ , \new_[15361]_ , \new_[15365]_ ,
    \new_[15366]_ , \new_[15367]_ , \new_[15370]_ , \new_[15374]_ ,
    \new_[15375]_ , \new_[15376]_ , \new_[15379]_ , \new_[15383]_ ,
    \new_[15384]_ , \new_[15385]_ , \new_[15388]_ , \new_[15392]_ ,
    \new_[15393]_ , \new_[15394]_ , \new_[15397]_ , \new_[15401]_ ,
    \new_[15402]_ , \new_[15403]_ , \new_[15406]_ , \new_[15410]_ ,
    \new_[15411]_ , \new_[15412]_ , \new_[15415]_ , \new_[15419]_ ,
    \new_[15420]_ , \new_[15421]_ , \new_[15424]_ , \new_[15428]_ ,
    \new_[15429]_ , \new_[15430]_ , \new_[15433]_ , \new_[15437]_ ,
    \new_[15438]_ , \new_[15439]_ , \new_[15442]_ , \new_[15446]_ ,
    \new_[15447]_ , \new_[15448]_ , \new_[15451]_ , \new_[15455]_ ,
    \new_[15456]_ , \new_[15457]_ , \new_[15460]_ , \new_[15464]_ ,
    \new_[15465]_ , \new_[15466]_ , \new_[15469]_ , \new_[15473]_ ,
    \new_[15474]_ , \new_[15475]_ , \new_[15478]_ , \new_[15482]_ ,
    \new_[15483]_ , \new_[15484]_ , \new_[15487]_ , \new_[15491]_ ,
    \new_[15492]_ , \new_[15493]_ , \new_[15496]_ , \new_[15500]_ ,
    \new_[15501]_ , \new_[15502]_ , \new_[15505]_ , \new_[15509]_ ,
    \new_[15510]_ , \new_[15511]_ , \new_[15514]_ , \new_[15518]_ ,
    \new_[15519]_ , \new_[15520]_ , \new_[15523]_ , \new_[15527]_ ,
    \new_[15528]_ , \new_[15529]_ , \new_[15532]_ , \new_[15536]_ ,
    \new_[15537]_ , \new_[15538]_ , \new_[15541]_ , \new_[15545]_ ,
    \new_[15546]_ , \new_[15547]_ , \new_[15550]_ , \new_[15554]_ ,
    \new_[15555]_ , \new_[15556]_ , \new_[15559]_ , \new_[15563]_ ,
    \new_[15564]_ , \new_[15565]_ , \new_[15568]_ , \new_[15572]_ ,
    \new_[15573]_ , \new_[15574]_ , \new_[15577]_ , \new_[15581]_ ,
    \new_[15582]_ , \new_[15583]_ , \new_[15586]_ , \new_[15590]_ ,
    \new_[15591]_ , \new_[15592]_ , \new_[15595]_ , \new_[15599]_ ,
    \new_[15600]_ , \new_[15601]_ , \new_[15604]_ , \new_[15608]_ ,
    \new_[15609]_ , \new_[15610]_ , \new_[15613]_ , \new_[15617]_ ,
    \new_[15618]_ , \new_[15619]_ , \new_[15622]_ , \new_[15626]_ ,
    \new_[15627]_ , \new_[15628]_ , \new_[15631]_ , \new_[15635]_ ,
    \new_[15636]_ , \new_[15637]_ , \new_[15640]_ , \new_[15644]_ ,
    \new_[15645]_ , \new_[15646]_ , \new_[15649]_ , \new_[15653]_ ,
    \new_[15654]_ , \new_[15655]_ , \new_[15658]_ , \new_[15662]_ ,
    \new_[15663]_ , \new_[15664]_ , \new_[15667]_ , \new_[15671]_ ,
    \new_[15672]_ , \new_[15673]_ , \new_[15676]_ , \new_[15680]_ ,
    \new_[15681]_ , \new_[15682]_ , \new_[15685]_ , \new_[15689]_ ,
    \new_[15690]_ , \new_[15691]_ , \new_[15694]_ , \new_[15698]_ ,
    \new_[15699]_ , \new_[15700]_ , \new_[15703]_ , \new_[15707]_ ,
    \new_[15708]_ , \new_[15709]_ , \new_[15712]_ , \new_[15716]_ ,
    \new_[15717]_ , \new_[15718]_ , \new_[15721]_ , \new_[15725]_ ,
    \new_[15726]_ , \new_[15727]_ , \new_[15730]_ , \new_[15734]_ ,
    \new_[15735]_ , \new_[15736]_ , \new_[15739]_ , \new_[15743]_ ,
    \new_[15744]_ , \new_[15745]_ , \new_[15748]_ , \new_[15752]_ ,
    \new_[15753]_ , \new_[15754]_ , \new_[15757]_ , \new_[15761]_ ,
    \new_[15762]_ , \new_[15763]_ , \new_[15766]_ , \new_[15770]_ ,
    \new_[15771]_ , \new_[15772]_ , \new_[15775]_ , \new_[15779]_ ,
    \new_[15780]_ , \new_[15781]_ , \new_[15784]_ , \new_[15788]_ ,
    \new_[15789]_ , \new_[15790]_ , \new_[15793]_ , \new_[15797]_ ,
    \new_[15798]_ , \new_[15799]_ , \new_[15802]_ , \new_[15806]_ ,
    \new_[15807]_ , \new_[15808]_ , \new_[15811]_ , \new_[15815]_ ,
    \new_[15816]_ , \new_[15817]_ , \new_[15820]_ , \new_[15824]_ ,
    \new_[15825]_ , \new_[15826]_ , \new_[15829]_ , \new_[15833]_ ,
    \new_[15834]_ , \new_[15835]_ , \new_[15838]_ , \new_[15842]_ ,
    \new_[15843]_ , \new_[15844]_ , \new_[15847]_ , \new_[15851]_ ,
    \new_[15852]_ , \new_[15853]_ , \new_[15856]_ , \new_[15860]_ ,
    \new_[15861]_ , \new_[15862]_ , \new_[15865]_ , \new_[15869]_ ,
    \new_[15870]_ , \new_[15871]_ , \new_[15874]_ , \new_[15878]_ ,
    \new_[15879]_ , \new_[15880]_ , \new_[15883]_ , \new_[15887]_ ,
    \new_[15888]_ , \new_[15889]_ , \new_[15892]_ , \new_[15896]_ ,
    \new_[15897]_ , \new_[15898]_ , \new_[15901]_ , \new_[15905]_ ,
    \new_[15906]_ , \new_[15907]_ , \new_[15910]_ , \new_[15914]_ ,
    \new_[15915]_ , \new_[15916]_ , \new_[15919]_ , \new_[15923]_ ,
    \new_[15924]_ , \new_[15925]_ , \new_[15928]_ , \new_[15932]_ ,
    \new_[15933]_ , \new_[15934]_ , \new_[15937]_ , \new_[15941]_ ,
    \new_[15942]_ , \new_[15943]_ , \new_[15946]_ , \new_[15950]_ ,
    \new_[15951]_ , \new_[15952]_ , \new_[15955]_ , \new_[15959]_ ,
    \new_[15960]_ , \new_[15961]_ , \new_[15964]_ , \new_[15968]_ ,
    \new_[15969]_ , \new_[15970]_ , \new_[15973]_ , \new_[15977]_ ,
    \new_[15978]_ , \new_[15979]_ , \new_[15982]_ , \new_[15986]_ ,
    \new_[15987]_ , \new_[15988]_ , \new_[15991]_ , \new_[15995]_ ,
    \new_[15996]_ , \new_[15997]_ , \new_[16000]_ , \new_[16004]_ ,
    \new_[16005]_ , \new_[16006]_ , \new_[16009]_ , \new_[16013]_ ,
    \new_[16014]_ , \new_[16015]_ , \new_[16018]_ , \new_[16022]_ ,
    \new_[16023]_ , \new_[16024]_ , \new_[16027]_ , \new_[16031]_ ,
    \new_[16032]_ , \new_[16033]_ , \new_[16036]_ , \new_[16040]_ ,
    \new_[16041]_ , \new_[16042]_ , \new_[16045]_ , \new_[16049]_ ,
    \new_[16050]_ , \new_[16051]_ , \new_[16054]_ , \new_[16058]_ ,
    \new_[16059]_ , \new_[16060]_ , \new_[16063]_ , \new_[16067]_ ,
    \new_[16068]_ , \new_[16069]_ , \new_[16072]_ , \new_[16076]_ ,
    \new_[16077]_ , \new_[16078]_ , \new_[16081]_ , \new_[16085]_ ,
    \new_[16086]_ , \new_[16087]_ , \new_[16090]_ , \new_[16094]_ ,
    \new_[16095]_ , \new_[16096]_ , \new_[16099]_ , \new_[16103]_ ,
    \new_[16104]_ , \new_[16105]_ , \new_[16108]_ , \new_[16112]_ ,
    \new_[16113]_ , \new_[16114]_ , \new_[16117]_ , \new_[16121]_ ,
    \new_[16122]_ , \new_[16123]_ , \new_[16126]_ , \new_[16130]_ ,
    \new_[16131]_ , \new_[16132]_ , \new_[16135]_ , \new_[16139]_ ,
    \new_[16140]_ , \new_[16141]_ , \new_[16144]_ , \new_[16148]_ ,
    \new_[16149]_ , \new_[16150]_ , \new_[16153]_ , \new_[16157]_ ,
    \new_[16158]_ , \new_[16159]_ , \new_[16162]_ , \new_[16166]_ ,
    \new_[16167]_ , \new_[16168]_ , \new_[16171]_ , \new_[16175]_ ,
    \new_[16176]_ , \new_[16177]_ , \new_[16180]_ , \new_[16184]_ ,
    \new_[16185]_ , \new_[16186]_ , \new_[16189]_ , \new_[16193]_ ,
    \new_[16194]_ , \new_[16195]_ , \new_[16198]_ , \new_[16202]_ ,
    \new_[16203]_ , \new_[16204]_ , \new_[16207]_ , \new_[16211]_ ,
    \new_[16212]_ , \new_[16213]_ , \new_[16216]_ , \new_[16220]_ ,
    \new_[16221]_ , \new_[16222]_ , \new_[16225]_ , \new_[16229]_ ,
    \new_[16230]_ , \new_[16231]_ , \new_[16234]_ , \new_[16238]_ ,
    \new_[16239]_ , \new_[16240]_ , \new_[16243]_ , \new_[16247]_ ,
    \new_[16248]_ , \new_[16249]_ , \new_[16252]_ , \new_[16256]_ ,
    \new_[16257]_ , \new_[16258]_ , \new_[16261]_ , \new_[16265]_ ,
    \new_[16266]_ , \new_[16267]_ , \new_[16270]_ , \new_[16274]_ ,
    \new_[16275]_ , \new_[16276]_ , \new_[16279]_ , \new_[16283]_ ,
    \new_[16284]_ , \new_[16285]_ , \new_[16288]_ , \new_[16292]_ ,
    \new_[16293]_ , \new_[16294]_ , \new_[16297]_ , \new_[16301]_ ,
    \new_[16302]_ , \new_[16303]_ , \new_[16306]_ , \new_[16310]_ ,
    \new_[16311]_ , \new_[16312]_ , \new_[16315]_ , \new_[16319]_ ,
    \new_[16320]_ , \new_[16321]_ , \new_[16324]_ , \new_[16328]_ ,
    \new_[16329]_ , \new_[16330]_ , \new_[16333]_ , \new_[16337]_ ,
    \new_[16338]_ , \new_[16339]_ , \new_[16342]_ , \new_[16346]_ ,
    \new_[16347]_ , \new_[16348]_ , \new_[16351]_ , \new_[16355]_ ,
    \new_[16356]_ , \new_[16357]_ , \new_[16360]_ , \new_[16364]_ ,
    \new_[16365]_ , \new_[16366]_ , \new_[16369]_ , \new_[16373]_ ,
    \new_[16374]_ , \new_[16375]_ , \new_[16378]_ , \new_[16382]_ ,
    \new_[16383]_ , \new_[16384]_ , \new_[16387]_ , \new_[16391]_ ,
    \new_[16392]_ , \new_[16393]_ , \new_[16396]_ , \new_[16400]_ ,
    \new_[16401]_ , \new_[16402]_ , \new_[16405]_ , \new_[16409]_ ,
    \new_[16410]_ , \new_[16411]_ , \new_[16414]_ , \new_[16418]_ ,
    \new_[16419]_ , \new_[16420]_ , \new_[16423]_ , \new_[16427]_ ,
    \new_[16428]_ , \new_[16429]_ , \new_[16432]_ , \new_[16436]_ ,
    \new_[16437]_ , \new_[16438]_ , \new_[16441]_ , \new_[16445]_ ,
    \new_[16446]_ , \new_[16447]_ , \new_[16450]_ , \new_[16454]_ ,
    \new_[16455]_ , \new_[16456]_ , \new_[16459]_ , \new_[16463]_ ,
    \new_[16464]_ , \new_[16465]_ , \new_[16468]_ , \new_[16472]_ ,
    \new_[16473]_ , \new_[16474]_ , \new_[16477]_ , \new_[16481]_ ,
    \new_[16482]_ , \new_[16483]_ , \new_[16486]_ , \new_[16490]_ ,
    \new_[16491]_ , \new_[16492]_ , \new_[16495]_ , \new_[16499]_ ,
    \new_[16500]_ , \new_[16501]_ , \new_[16504]_ , \new_[16508]_ ,
    \new_[16509]_ , \new_[16510]_ , \new_[16513]_ , \new_[16517]_ ,
    \new_[16518]_ , \new_[16519]_ , \new_[16522]_ , \new_[16526]_ ,
    \new_[16527]_ , \new_[16528]_ , \new_[16531]_ , \new_[16535]_ ,
    \new_[16536]_ , \new_[16537]_ , \new_[16540]_ , \new_[16544]_ ,
    \new_[16545]_ , \new_[16546]_ , \new_[16549]_ , \new_[16553]_ ,
    \new_[16554]_ , \new_[16555]_ , \new_[16558]_ , \new_[16562]_ ,
    \new_[16563]_ , \new_[16564]_ , \new_[16567]_ , \new_[16571]_ ,
    \new_[16572]_ , \new_[16573]_ , \new_[16576]_ , \new_[16580]_ ,
    \new_[16581]_ , \new_[16582]_ , \new_[16585]_ , \new_[16589]_ ,
    \new_[16590]_ , \new_[16591]_ , \new_[16594]_ , \new_[16598]_ ,
    \new_[16599]_ , \new_[16600]_ , \new_[16603]_ , \new_[16607]_ ,
    \new_[16608]_ , \new_[16609]_ , \new_[16612]_ , \new_[16616]_ ,
    \new_[16617]_ , \new_[16618]_ , \new_[16621]_ , \new_[16625]_ ,
    \new_[16626]_ , \new_[16627]_ , \new_[16630]_ , \new_[16634]_ ,
    \new_[16635]_ , \new_[16636]_ , \new_[16639]_ , \new_[16643]_ ,
    \new_[16644]_ , \new_[16645]_ , \new_[16648]_ , \new_[16652]_ ,
    \new_[16653]_ , \new_[16654]_ , \new_[16657]_ , \new_[16661]_ ,
    \new_[16662]_ , \new_[16663]_ , \new_[16666]_ , \new_[16670]_ ,
    \new_[16671]_ , \new_[16672]_ , \new_[16675]_ , \new_[16679]_ ,
    \new_[16680]_ , \new_[16681]_ , \new_[16684]_ , \new_[16688]_ ,
    \new_[16689]_ , \new_[16690]_ , \new_[16693]_ , \new_[16697]_ ,
    \new_[16698]_ , \new_[16699]_ , \new_[16702]_ , \new_[16706]_ ,
    \new_[16707]_ , \new_[16708]_ , \new_[16711]_ , \new_[16715]_ ,
    \new_[16716]_ , \new_[16717]_ , \new_[16720]_ , \new_[16724]_ ,
    \new_[16725]_ , \new_[16726]_ , \new_[16729]_ , \new_[16733]_ ,
    \new_[16734]_ , \new_[16735]_ , \new_[16738]_ , \new_[16742]_ ,
    \new_[16743]_ , \new_[16744]_ , \new_[16747]_ , \new_[16751]_ ,
    \new_[16752]_ , \new_[16753]_ , \new_[16756]_ , \new_[16760]_ ,
    \new_[16761]_ , \new_[16762]_ , \new_[16765]_ , \new_[16769]_ ,
    \new_[16770]_ , \new_[16771]_ , \new_[16774]_ , \new_[16778]_ ,
    \new_[16779]_ , \new_[16780]_ , \new_[16783]_ , \new_[16787]_ ,
    \new_[16788]_ , \new_[16789]_ , \new_[16792]_ , \new_[16796]_ ,
    \new_[16797]_ , \new_[16798]_ , \new_[16801]_ , \new_[16805]_ ,
    \new_[16806]_ , \new_[16807]_ , \new_[16810]_ , \new_[16814]_ ,
    \new_[16815]_ , \new_[16816]_ , \new_[16819]_ , \new_[16823]_ ,
    \new_[16824]_ , \new_[16825]_ , \new_[16829]_ , \new_[16830]_ ,
    \new_[16834]_ , \new_[16835]_ , \new_[16836]_ , \new_[16839]_ ,
    \new_[16843]_ , \new_[16844]_ , \new_[16845]_ , \new_[16849]_ ,
    \new_[16850]_ , \new_[16854]_ , \new_[16855]_ , \new_[16856]_ ,
    \new_[16859]_ , \new_[16863]_ , \new_[16864]_ , \new_[16865]_ ,
    \new_[16869]_ , \new_[16870]_ , \new_[16874]_ , \new_[16875]_ ,
    \new_[16876]_ , \new_[16879]_ , \new_[16883]_ , \new_[16884]_ ,
    \new_[16885]_ , \new_[16889]_ , \new_[16890]_ , \new_[16894]_ ,
    \new_[16895]_ , \new_[16896]_ , \new_[16899]_ , \new_[16903]_ ,
    \new_[16904]_ , \new_[16905]_ , \new_[16909]_ , \new_[16910]_ ,
    \new_[16914]_ , \new_[16915]_ , \new_[16916]_ , \new_[16919]_ ,
    \new_[16923]_ , \new_[16924]_ , \new_[16925]_ , \new_[16929]_ ,
    \new_[16930]_ , \new_[16934]_ , \new_[16935]_ , \new_[16936]_ ,
    \new_[16939]_ , \new_[16943]_ , \new_[16944]_ , \new_[16945]_ ,
    \new_[16949]_ , \new_[16950]_ , \new_[16954]_ , \new_[16955]_ ,
    \new_[16956]_ , \new_[16959]_ , \new_[16963]_ , \new_[16964]_ ,
    \new_[16965]_ , \new_[16969]_ , \new_[16970]_ , \new_[16974]_ ,
    \new_[16975]_ , \new_[16976]_ , \new_[16979]_ , \new_[16983]_ ,
    \new_[16984]_ , \new_[16985]_ , \new_[16989]_ , \new_[16990]_ ,
    \new_[16994]_ , \new_[16995]_ , \new_[16996]_ , \new_[16999]_ ,
    \new_[17003]_ , \new_[17004]_ , \new_[17005]_ , \new_[17009]_ ,
    \new_[17010]_ , \new_[17014]_ , \new_[17015]_ , \new_[17016]_ ,
    \new_[17019]_ , \new_[17023]_ , \new_[17024]_ , \new_[17025]_ ,
    \new_[17029]_ , \new_[17030]_ , \new_[17034]_ , \new_[17035]_ ,
    \new_[17036]_ , \new_[17039]_ , \new_[17043]_ , \new_[17044]_ ,
    \new_[17045]_ , \new_[17049]_ , \new_[17050]_ , \new_[17054]_ ,
    \new_[17055]_ , \new_[17056]_ , \new_[17059]_ , \new_[17063]_ ,
    \new_[17064]_ , \new_[17065]_ , \new_[17069]_ , \new_[17070]_ ,
    \new_[17074]_ , \new_[17075]_ , \new_[17076]_ , \new_[17079]_ ,
    \new_[17083]_ , \new_[17084]_ , \new_[17085]_ , \new_[17089]_ ,
    \new_[17090]_ , \new_[17094]_ , \new_[17095]_ , \new_[17096]_ ,
    \new_[17099]_ , \new_[17103]_ , \new_[17104]_ , \new_[17105]_ ,
    \new_[17109]_ , \new_[17110]_ , \new_[17114]_ , \new_[17115]_ ,
    \new_[17116]_ , \new_[17119]_ , \new_[17123]_ , \new_[17124]_ ,
    \new_[17125]_ , \new_[17129]_ , \new_[17130]_ , \new_[17134]_ ,
    \new_[17135]_ , \new_[17136]_ , \new_[17139]_ , \new_[17143]_ ,
    \new_[17144]_ , \new_[17145]_ , \new_[17149]_ , \new_[17150]_ ,
    \new_[17154]_ , \new_[17155]_ , \new_[17156]_ , \new_[17159]_ ,
    \new_[17163]_ , \new_[17164]_ , \new_[17165]_ , \new_[17169]_ ,
    \new_[17170]_ , \new_[17174]_ , \new_[17175]_ , \new_[17176]_ ,
    \new_[17179]_ , \new_[17183]_ , \new_[17184]_ , \new_[17185]_ ,
    \new_[17189]_ , \new_[17190]_ , \new_[17194]_ , \new_[17195]_ ,
    \new_[17196]_ , \new_[17199]_ , \new_[17203]_ , \new_[17204]_ ,
    \new_[17205]_ , \new_[17209]_ , \new_[17210]_ , \new_[17214]_ ,
    \new_[17215]_ , \new_[17216]_ , \new_[17219]_ , \new_[17223]_ ,
    \new_[17224]_ , \new_[17225]_ , \new_[17229]_ , \new_[17230]_ ,
    \new_[17234]_ , \new_[17235]_ , \new_[17236]_ , \new_[17239]_ ,
    \new_[17243]_ , \new_[17244]_ , \new_[17245]_ , \new_[17249]_ ,
    \new_[17250]_ , \new_[17254]_ , \new_[17255]_ , \new_[17256]_ ,
    \new_[17259]_ , \new_[17263]_ , \new_[17264]_ , \new_[17265]_ ,
    \new_[17269]_ , \new_[17270]_ , \new_[17274]_ , \new_[17275]_ ,
    \new_[17276]_ , \new_[17279]_ , \new_[17283]_ , \new_[17284]_ ,
    \new_[17285]_ , \new_[17289]_ , \new_[17290]_ , \new_[17294]_ ,
    \new_[17295]_ , \new_[17296]_ , \new_[17299]_ , \new_[17303]_ ,
    \new_[17304]_ , \new_[17305]_ , \new_[17309]_ , \new_[17310]_ ,
    \new_[17314]_ , \new_[17315]_ , \new_[17316]_ , \new_[17319]_ ,
    \new_[17323]_ , \new_[17324]_ , \new_[17325]_ , \new_[17329]_ ,
    \new_[17330]_ , \new_[17334]_ , \new_[17335]_ , \new_[17336]_ ,
    \new_[17339]_ , \new_[17343]_ , \new_[17344]_ , \new_[17345]_ ,
    \new_[17349]_ , \new_[17350]_ , \new_[17354]_ , \new_[17355]_ ,
    \new_[17356]_ , \new_[17359]_ , \new_[17363]_ , \new_[17364]_ ,
    \new_[17365]_ , \new_[17369]_ , \new_[17370]_ , \new_[17374]_ ,
    \new_[17375]_ , \new_[17376]_ , \new_[17379]_ , \new_[17383]_ ,
    \new_[17384]_ , \new_[17385]_ , \new_[17389]_ , \new_[17390]_ ,
    \new_[17394]_ , \new_[17395]_ , \new_[17396]_ , \new_[17399]_ ,
    \new_[17403]_ , \new_[17404]_ , \new_[17405]_ , \new_[17409]_ ,
    \new_[17410]_ , \new_[17414]_ , \new_[17415]_ , \new_[17416]_ ,
    \new_[17419]_ , \new_[17423]_ , \new_[17424]_ , \new_[17425]_ ,
    \new_[17429]_ , \new_[17430]_ , \new_[17434]_ , \new_[17435]_ ,
    \new_[17436]_ , \new_[17439]_ , \new_[17443]_ , \new_[17444]_ ,
    \new_[17445]_ , \new_[17449]_ , \new_[17450]_ , \new_[17454]_ ,
    \new_[17455]_ , \new_[17456]_ , \new_[17459]_ , \new_[17463]_ ,
    \new_[17464]_ , \new_[17465]_ , \new_[17469]_ , \new_[17470]_ ,
    \new_[17474]_ , \new_[17475]_ , \new_[17476]_ , \new_[17479]_ ,
    \new_[17483]_ , \new_[17484]_ , \new_[17485]_ , \new_[17489]_ ,
    \new_[17490]_ , \new_[17494]_ , \new_[17495]_ , \new_[17496]_ ,
    \new_[17499]_ , \new_[17503]_ , \new_[17504]_ , \new_[17505]_ ,
    \new_[17509]_ , \new_[17510]_ , \new_[17514]_ , \new_[17515]_ ,
    \new_[17516]_ , \new_[17519]_ , \new_[17523]_ , \new_[17524]_ ,
    \new_[17525]_ , \new_[17529]_ , \new_[17530]_ , \new_[17534]_ ,
    \new_[17535]_ , \new_[17536]_ , \new_[17539]_ , \new_[17543]_ ,
    \new_[17544]_ , \new_[17545]_ , \new_[17549]_ , \new_[17550]_ ,
    \new_[17554]_ , \new_[17555]_ , \new_[17556]_ , \new_[17559]_ ,
    \new_[17563]_ , \new_[17564]_ , \new_[17565]_ , \new_[17569]_ ,
    \new_[17570]_ , \new_[17574]_ , \new_[17575]_ , \new_[17576]_ ,
    \new_[17579]_ , \new_[17583]_ , \new_[17584]_ , \new_[17585]_ ,
    \new_[17589]_ , \new_[17590]_ , \new_[17594]_ , \new_[17595]_ ,
    \new_[17596]_ , \new_[17599]_ , \new_[17603]_ , \new_[17604]_ ,
    \new_[17605]_ , \new_[17609]_ , \new_[17610]_ , \new_[17614]_ ,
    \new_[17615]_ , \new_[17616]_ , \new_[17619]_ , \new_[17623]_ ,
    \new_[17624]_ , \new_[17625]_ , \new_[17629]_ , \new_[17630]_ ,
    \new_[17634]_ , \new_[17635]_ , \new_[17636]_ , \new_[17639]_ ,
    \new_[17643]_ , \new_[17644]_ , \new_[17645]_ , \new_[17649]_ ,
    \new_[17650]_ , \new_[17654]_ , \new_[17655]_ , \new_[17656]_ ,
    \new_[17659]_ , \new_[17663]_ , \new_[17664]_ , \new_[17665]_ ,
    \new_[17669]_ , \new_[17670]_ , \new_[17674]_ , \new_[17675]_ ,
    \new_[17676]_ , \new_[17679]_ , \new_[17683]_ , \new_[17684]_ ,
    \new_[17685]_ , \new_[17689]_ , \new_[17690]_ , \new_[17694]_ ,
    \new_[17695]_ , \new_[17696]_ , \new_[17699]_ , \new_[17703]_ ,
    \new_[17704]_ , \new_[17705]_ , \new_[17709]_ , \new_[17710]_ ,
    \new_[17714]_ , \new_[17715]_ , \new_[17716]_ , \new_[17719]_ ,
    \new_[17723]_ , \new_[17724]_ , \new_[17725]_ , \new_[17729]_ ,
    \new_[17730]_ , \new_[17734]_ , \new_[17735]_ , \new_[17736]_ ,
    \new_[17739]_ , \new_[17743]_ , \new_[17744]_ , \new_[17745]_ ,
    \new_[17749]_ , \new_[17750]_ , \new_[17754]_ , \new_[17755]_ ,
    \new_[17756]_ , \new_[17759]_ , \new_[17763]_ , \new_[17764]_ ,
    \new_[17765]_ , \new_[17769]_ , \new_[17770]_ , \new_[17774]_ ,
    \new_[17775]_ , \new_[17776]_ , \new_[17779]_ , \new_[17783]_ ,
    \new_[17784]_ , \new_[17785]_ , \new_[17789]_ , \new_[17790]_ ,
    \new_[17794]_ , \new_[17795]_ , \new_[17796]_ , \new_[17799]_ ,
    \new_[17803]_ , \new_[17804]_ , \new_[17805]_ , \new_[17809]_ ,
    \new_[17810]_ , \new_[17814]_ , \new_[17815]_ , \new_[17816]_ ,
    \new_[17819]_ , \new_[17823]_ , \new_[17824]_ , \new_[17825]_ ,
    \new_[17829]_ , \new_[17830]_ , \new_[17834]_ , \new_[17835]_ ,
    \new_[17836]_ , \new_[17839]_ , \new_[17843]_ , \new_[17844]_ ,
    \new_[17845]_ , \new_[17849]_ , \new_[17850]_ , \new_[17854]_ ,
    \new_[17855]_ , \new_[17856]_ , \new_[17859]_ , \new_[17863]_ ,
    \new_[17864]_ , \new_[17865]_ , \new_[17869]_ , \new_[17870]_ ,
    \new_[17874]_ , \new_[17875]_ , \new_[17876]_ , \new_[17879]_ ,
    \new_[17883]_ , \new_[17884]_ , \new_[17885]_ , \new_[17889]_ ,
    \new_[17890]_ , \new_[17894]_ , \new_[17895]_ , \new_[17896]_ ,
    \new_[17899]_ , \new_[17903]_ , \new_[17904]_ , \new_[17905]_ ,
    \new_[17909]_ , \new_[17910]_ , \new_[17914]_ , \new_[17915]_ ,
    \new_[17916]_ , \new_[17919]_ , \new_[17923]_ , \new_[17924]_ ,
    \new_[17925]_ , \new_[17929]_ , \new_[17930]_ , \new_[17934]_ ,
    \new_[17935]_ , \new_[17936]_ , \new_[17939]_ , \new_[17943]_ ,
    \new_[17944]_ , \new_[17945]_ , \new_[17949]_ , \new_[17950]_ ,
    \new_[17954]_ , \new_[17955]_ , \new_[17956]_ , \new_[17959]_ ,
    \new_[17963]_ , \new_[17964]_ , \new_[17965]_ , \new_[17969]_ ,
    \new_[17970]_ , \new_[17974]_ , \new_[17975]_ , \new_[17976]_ ,
    \new_[17979]_ , \new_[17983]_ , \new_[17984]_ , \new_[17985]_ ,
    \new_[17989]_ , \new_[17990]_ , \new_[17994]_ , \new_[17995]_ ,
    \new_[17996]_ , \new_[17999]_ , \new_[18003]_ , \new_[18004]_ ,
    \new_[18005]_ , \new_[18009]_ , \new_[18010]_ , \new_[18014]_ ,
    \new_[18015]_ , \new_[18016]_ , \new_[18019]_ , \new_[18023]_ ,
    \new_[18024]_ , \new_[18025]_ , \new_[18029]_ , \new_[18030]_ ,
    \new_[18034]_ , \new_[18035]_ , \new_[18036]_ , \new_[18039]_ ,
    \new_[18043]_ , \new_[18044]_ , \new_[18045]_ , \new_[18049]_ ,
    \new_[18050]_ , \new_[18054]_ , \new_[18055]_ , \new_[18056]_ ,
    \new_[18059]_ , \new_[18063]_ , \new_[18064]_ , \new_[18065]_ ,
    \new_[18069]_ , \new_[18070]_ , \new_[18074]_ , \new_[18075]_ ,
    \new_[18076]_ , \new_[18079]_ , \new_[18083]_ , \new_[18084]_ ,
    \new_[18085]_ , \new_[18089]_ , \new_[18090]_ , \new_[18094]_ ,
    \new_[18095]_ , \new_[18096]_ , \new_[18099]_ , \new_[18103]_ ,
    \new_[18104]_ , \new_[18105]_ , \new_[18109]_ , \new_[18110]_ ,
    \new_[18114]_ , \new_[18115]_ , \new_[18116]_ , \new_[18119]_ ,
    \new_[18123]_ , \new_[18124]_ , \new_[18125]_ , \new_[18129]_ ,
    \new_[18130]_ , \new_[18134]_ , \new_[18135]_ , \new_[18136]_ ,
    \new_[18139]_ , \new_[18143]_ , \new_[18144]_ , \new_[18145]_ ,
    \new_[18149]_ , \new_[18150]_ , \new_[18154]_ , \new_[18155]_ ,
    \new_[18156]_ , \new_[18159]_ , \new_[18163]_ , \new_[18164]_ ,
    \new_[18165]_ , \new_[18169]_ , \new_[18170]_ , \new_[18174]_ ,
    \new_[18175]_ , \new_[18176]_ , \new_[18179]_ , \new_[18183]_ ,
    \new_[18184]_ , \new_[18185]_ , \new_[18189]_ , \new_[18190]_ ,
    \new_[18194]_ , \new_[18195]_ , \new_[18196]_ , \new_[18199]_ ,
    \new_[18203]_ , \new_[18204]_ , \new_[18205]_ , \new_[18209]_ ,
    \new_[18210]_ , \new_[18214]_ , \new_[18215]_ , \new_[18216]_ ,
    \new_[18219]_ , \new_[18223]_ , \new_[18224]_ , \new_[18225]_ ,
    \new_[18229]_ , \new_[18230]_ , \new_[18234]_ , \new_[18235]_ ,
    \new_[18236]_ , \new_[18239]_ , \new_[18243]_ , \new_[18244]_ ,
    \new_[18245]_ , \new_[18249]_ , \new_[18250]_ , \new_[18254]_ ,
    \new_[18255]_ , \new_[18256]_ , \new_[18259]_ , \new_[18263]_ ,
    \new_[18264]_ , \new_[18265]_ , \new_[18269]_ , \new_[18270]_ ,
    \new_[18274]_ , \new_[18275]_ , \new_[18276]_ , \new_[18279]_ ,
    \new_[18283]_ , \new_[18284]_ , \new_[18285]_ , \new_[18289]_ ,
    \new_[18290]_ , \new_[18294]_ , \new_[18295]_ , \new_[18296]_ ,
    \new_[18299]_ , \new_[18303]_ , \new_[18304]_ , \new_[18305]_ ,
    \new_[18309]_ , \new_[18310]_ , \new_[18314]_ , \new_[18315]_ ,
    \new_[18316]_ , \new_[18319]_ , \new_[18323]_ , \new_[18324]_ ,
    \new_[18325]_ , \new_[18329]_ , \new_[18330]_ , \new_[18334]_ ,
    \new_[18335]_ , \new_[18336]_ , \new_[18339]_ , \new_[18343]_ ,
    \new_[18344]_ , \new_[18345]_ , \new_[18349]_ , \new_[18350]_ ,
    \new_[18354]_ , \new_[18355]_ , \new_[18356]_ , \new_[18359]_ ,
    \new_[18363]_ , \new_[18364]_ , \new_[18365]_ , \new_[18369]_ ,
    \new_[18370]_ , \new_[18374]_ , \new_[18375]_ , \new_[18376]_ ,
    \new_[18379]_ , \new_[18383]_ , \new_[18384]_ , \new_[18385]_ ,
    \new_[18389]_ , \new_[18390]_ , \new_[18394]_ , \new_[18395]_ ,
    \new_[18396]_ , \new_[18399]_ , \new_[18403]_ , \new_[18404]_ ,
    \new_[18405]_ , \new_[18409]_ , \new_[18410]_ , \new_[18414]_ ,
    \new_[18415]_ , \new_[18416]_ , \new_[18419]_ , \new_[18423]_ ,
    \new_[18424]_ , \new_[18425]_ , \new_[18429]_ , \new_[18430]_ ,
    \new_[18434]_ , \new_[18435]_ , \new_[18436]_ , \new_[18439]_ ,
    \new_[18443]_ , \new_[18444]_ , \new_[18445]_ , \new_[18449]_ ,
    \new_[18450]_ , \new_[18454]_ , \new_[18455]_ , \new_[18456]_ ,
    \new_[18459]_ , \new_[18463]_ , \new_[18464]_ , \new_[18465]_ ,
    \new_[18469]_ , \new_[18470]_ , \new_[18474]_ , \new_[18475]_ ,
    \new_[18476]_ , \new_[18479]_ , \new_[18483]_ , \new_[18484]_ ,
    \new_[18485]_ , \new_[18489]_ , \new_[18490]_ , \new_[18494]_ ,
    \new_[18495]_ , \new_[18496]_ , \new_[18499]_ , \new_[18503]_ ,
    \new_[18504]_ , \new_[18505]_ , \new_[18509]_ , \new_[18510]_ ,
    \new_[18514]_ , \new_[18515]_ , \new_[18516]_ , \new_[18519]_ ,
    \new_[18523]_ , \new_[18524]_ , \new_[18525]_ , \new_[18529]_ ,
    \new_[18530]_ , \new_[18534]_ , \new_[18535]_ , \new_[18536]_ ,
    \new_[18539]_ , \new_[18543]_ , \new_[18544]_ , \new_[18545]_ ,
    \new_[18549]_ , \new_[18550]_ , \new_[18554]_ , \new_[18555]_ ,
    \new_[18556]_ , \new_[18559]_ , \new_[18563]_ , \new_[18564]_ ,
    \new_[18565]_ , \new_[18569]_ , \new_[18570]_ , \new_[18574]_ ,
    \new_[18575]_ , \new_[18576]_ , \new_[18579]_ , \new_[18583]_ ,
    \new_[18584]_ , \new_[18585]_ , \new_[18589]_ , \new_[18590]_ ,
    \new_[18594]_ , \new_[18595]_ , \new_[18596]_ , \new_[18599]_ ,
    \new_[18603]_ , \new_[18604]_ , \new_[18605]_ , \new_[18609]_ ,
    \new_[18610]_ , \new_[18614]_ , \new_[18615]_ , \new_[18616]_ ,
    \new_[18619]_ , \new_[18623]_ , \new_[18624]_ , \new_[18625]_ ,
    \new_[18629]_ , \new_[18630]_ , \new_[18634]_ , \new_[18635]_ ,
    \new_[18636]_ , \new_[18639]_ , \new_[18643]_ , \new_[18644]_ ,
    \new_[18645]_ , \new_[18649]_ , \new_[18650]_ , \new_[18654]_ ,
    \new_[18655]_ , \new_[18656]_ , \new_[18659]_ , \new_[18663]_ ,
    \new_[18664]_ , \new_[18665]_ , \new_[18669]_ , \new_[18670]_ ,
    \new_[18674]_ , \new_[18675]_ , \new_[18676]_ , \new_[18679]_ ,
    \new_[18683]_ , \new_[18684]_ , \new_[18685]_ , \new_[18689]_ ,
    \new_[18690]_ , \new_[18694]_ , \new_[18695]_ , \new_[18696]_ ,
    \new_[18699]_ , \new_[18703]_ , \new_[18704]_ , \new_[18705]_ ,
    \new_[18709]_ , \new_[18710]_ , \new_[18714]_ , \new_[18715]_ ,
    \new_[18716]_ , \new_[18719]_ , \new_[18723]_ , \new_[18724]_ ,
    \new_[18725]_ , \new_[18729]_ , \new_[18730]_ , \new_[18734]_ ,
    \new_[18735]_ , \new_[18736]_ , \new_[18739]_ , \new_[18743]_ ,
    \new_[18744]_ , \new_[18745]_ , \new_[18749]_ , \new_[18750]_ ,
    \new_[18754]_ , \new_[18755]_ , \new_[18756]_ , \new_[18759]_ ,
    \new_[18763]_ , \new_[18764]_ , \new_[18765]_ , \new_[18769]_ ,
    \new_[18770]_ , \new_[18774]_ , \new_[18775]_ , \new_[18776]_ ,
    \new_[18779]_ , \new_[18783]_ , \new_[18784]_ , \new_[18785]_ ,
    \new_[18789]_ , \new_[18790]_ , \new_[18794]_ , \new_[18795]_ ,
    \new_[18796]_ , \new_[18799]_ , \new_[18803]_ , \new_[18804]_ ,
    \new_[18805]_ , \new_[18809]_ , \new_[18810]_ , \new_[18814]_ ,
    \new_[18815]_ , \new_[18816]_ , \new_[18819]_ , \new_[18823]_ ,
    \new_[18824]_ , \new_[18825]_ , \new_[18829]_ , \new_[18830]_ ,
    \new_[18834]_ , \new_[18835]_ , \new_[18836]_ , \new_[18839]_ ,
    \new_[18843]_ , \new_[18844]_ , \new_[18845]_ , \new_[18849]_ ,
    \new_[18850]_ , \new_[18854]_ , \new_[18855]_ , \new_[18856]_ ,
    \new_[18859]_ , \new_[18863]_ , \new_[18864]_ , \new_[18865]_ ,
    \new_[18869]_ , \new_[18870]_ , \new_[18874]_ , \new_[18875]_ ,
    \new_[18876]_ , \new_[18879]_ , \new_[18883]_ , \new_[18884]_ ,
    \new_[18885]_ , \new_[18889]_ , \new_[18890]_ , \new_[18894]_ ,
    \new_[18895]_ , \new_[18896]_ , \new_[18899]_ , \new_[18903]_ ,
    \new_[18904]_ , \new_[18905]_ , \new_[18909]_ , \new_[18910]_ ,
    \new_[18914]_ , \new_[18915]_ , \new_[18916]_ , \new_[18919]_ ,
    \new_[18923]_ , \new_[18924]_ , \new_[18925]_ , \new_[18929]_ ,
    \new_[18930]_ , \new_[18934]_ , \new_[18935]_ , \new_[18936]_ ,
    \new_[18939]_ , \new_[18943]_ , \new_[18944]_ , \new_[18945]_ ,
    \new_[18949]_ , \new_[18950]_ , \new_[18954]_ , \new_[18955]_ ,
    \new_[18956]_ , \new_[18959]_ , \new_[18963]_ , \new_[18964]_ ,
    \new_[18965]_ , \new_[18969]_ , \new_[18970]_ , \new_[18974]_ ,
    \new_[18975]_ , \new_[18976]_ , \new_[18979]_ , \new_[18983]_ ,
    \new_[18984]_ , \new_[18985]_ , \new_[18989]_ , \new_[18990]_ ,
    \new_[18994]_ , \new_[18995]_ , \new_[18996]_ , \new_[18999]_ ,
    \new_[19003]_ , \new_[19004]_ , \new_[19005]_ , \new_[19009]_ ,
    \new_[19010]_ , \new_[19014]_ , \new_[19015]_ , \new_[19016]_ ,
    \new_[19019]_ , \new_[19023]_ , \new_[19024]_ , \new_[19025]_ ,
    \new_[19029]_ , \new_[19030]_ , \new_[19034]_ , \new_[19035]_ ,
    \new_[19036]_ , \new_[19039]_ , \new_[19043]_ , \new_[19044]_ ,
    \new_[19045]_ , \new_[19049]_ , \new_[19050]_ , \new_[19054]_ ,
    \new_[19055]_ , \new_[19056]_ , \new_[19059]_ , \new_[19063]_ ,
    \new_[19064]_ , \new_[19065]_ , \new_[19069]_ , \new_[19070]_ ,
    \new_[19074]_ , \new_[19075]_ , \new_[19076]_ , \new_[19079]_ ,
    \new_[19083]_ , \new_[19084]_ , \new_[19085]_ , \new_[19089]_ ,
    \new_[19090]_ , \new_[19094]_ , \new_[19095]_ , \new_[19096]_ ,
    \new_[19099]_ , \new_[19103]_ , \new_[19104]_ , \new_[19105]_ ,
    \new_[19109]_ , \new_[19110]_ , \new_[19114]_ , \new_[19115]_ ,
    \new_[19116]_ , \new_[19119]_ , \new_[19123]_ , \new_[19124]_ ,
    \new_[19125]_ , \new_[19129]_ , \new_[19130]_ , \new_[19134]_ ,
    \new_[19135]_ , \new_[19136]_ , \new_[19139]_ , \new_[19143]_ ,
    \new_[19144]_ , \new_[19145]_ , \new_[19149]_ , \new_[19150]_ ,
    \new_[19154]_ , \new_[19155]_ , \new_[19156]_ , \new_[19159]_ ,
    \new_[19163]_ , \new_[19164]_ , \new_[19165]_ , \new_[19169]_ ,
    \new_[19170]_ , \new_[19174]_ , \new_[19175]_ , \new_[19176]_ ,
    \new_[19179]_ , \new_[19183]_ , \new_[19184]_ , \new_[19185]_ ,
    \new_[19189]_ , \new_[19190]_ , \new_[19194]_ , \new_[19195]_ ,
    \new_[19196]_ , \new_[19199]_ , \new_[19203]_ , \new_[19204]_ ,
    \new_[19205]_ , \new_[19209]_ , \new_[19210]_ , \new_[19214]_ ,
    \new_[19215]_ , \new_[19216]_ , \new_[19219]_ , \new_[19223]_ ,
    \new_[19224]_ , \new_[19225]_ , \new_[19229]_ , \new_[19230]_ ,
    \new_[19234]_ , \new_[19235]_ , \new_[19236]_ , \new_[19239]_ ,
    \new_[19243]_ , \new_[19244]_ , \new_[19245]_ , \new_[19249]_ ,
    \new_[19250]_ , \new_[19254]_ , \new_[19255]_ , \new_[19256]_ ,
    \new_[19259]_ , \new_[19263]_ , \new_[19264]_ , \new_[19265]_ ,
    \new_[19269]_ , \new_[19270]_ , \new_[19274]_ , \new_[19275]_ ,
    \new_[19276]_ , \new_[19279]_ , \new_[19283]_ , \new_[19284]_ ,
    \new_[19285]_ , \new_[19289]_ , \new_[19290]_ , \new_[19294]_ ,
    \new_[19295]_ , \new_[19296]_ , \new_[19299]_ , \new_[19303]_ ,
    \new_[19304]_ , \new_[19305]_ , \new_[19309]_ , \new_[19310]_ ,
    \new_[19314]_ , \new_[19315]_ , \new_[19316]_ , \new_[19319]_ ,
    \new_[19323]_ , \new_[19324]_ , \new_[19325]_ , \new_[19329]_ ,
    \new_[19330]_ , \new_[19334]_ , \new_[19335]_ , \new_[19336]_ ,
    \new_[19339]_ , \new_[19343]_ , \new_[19344]_ , \new_[19345]_ ,
    \new_[19349]_ , \new_[19350]_ , \new_[19354]_ , \new_[19355]_ ,
    \new_[19356]_ , \new_[19359]_ , \new_[19363]_ , \new_[19364]_ ,
    \new_[19365]_ , \new_[19369]_ , \new_[19370]_ , \new_[19374]_ ,
    \new_[19375]_ , \new_[19376]_ , \new_[19379]_ , \new_[19383]_ ,
    \new_[19384]_ , \new_[19385]_ , \new_[19389]_ , \new_[19390]_ ,
    \new_[19394]_ , \new_[19395]_ , \new_[19396]_ , \new_[19399]_ ,
    \new_[19403]_ , \new_[19404]_ , \new_[19405]_ , \new_[19409]_ ,
    \new_[19410]_ , \new_[19414]_ , \new_[19415]_ , \new_[19416]_ ,
    \new_[19419]_ , \new_[19423]_ , \new_[19424]_ , \new_[19425]_ ,
    \new_[19429]_ , \new_[19430]_ , \new_[19434]_ , \new_[19435]_ ,
    \new_[19436]_ , \new_[19439]_ , \new_[19443]_ , \new_[19444]_ ,
    \new_[19445]_ , \new_[19449]_ , \new_[19450]_ , \new_[19454]_ ,
    \new_[19455]_ , \new_[19456]_ , \new_[19459]_ , \new_[19463]_ ,
    \new_[19464]_ , \new_[19465]_ , \new_[19469]_ , \new_[19470]_ ,
    \new_[19474]_ , \new_[19475]_ , \new_[19476]_ , \new_[19479]_ ,
    \new_[19483]_ , \new_[19484]_ , \new_[19485]_ , \new_[19489]_ ,
    \new_[19490]_ , \new_[19494]_ , \new_[19495]_ , \new_[19496]_ ,
    \new_[19499]_ , \new_[19503]_ , \new_[19504]_ , \new_[19505]_ ,
    \new_[19509]_ , \new_[19510]_ , \new_[19514]_ , \new_[19515]_ ,
    \new_[19516]_ , \new_[19519]_ , \new_[19523]_ , \new_[19524]_ ,
    \new_[19525]_ , \new_[19529]_ , \new_[19530]_ , \new_[19534]_ ,
    \new_[19535]_ , \new_[19536]_ , \new_[19539]_ , \new_[19543]_ ,
    \new_[19544]_ , \new_[19545]_ , \new_[19549]_ , \new_[19550]_ ,
    \new_[19554]_ , \new_[19555]_ , \new_[19556]_ , \new_[19559]_ ,
    \new_[19563]_ , \new_[19564]_ , \new_[19565]_ , \new_[19569]_ ,
    \new_[19570]_ , \new_[19574]_ , \new_[19575]_ , \new_[19576]_ ,
    \new_[19579]_ , \new_[19583]_ , \new_[19584]_ , \new_[19585]_ ,
    \new_[19589]_ , \new_[19590]_ , \new_[19594]_ , \new_[19595]_ ,
    \new_[19596]_ , \new_[19599]_ , \new_[19603]_ , \new_[19604]_ ,
    \new_[19605]_ , \new_[19609]_ , \new_[19610]_ , \new_[19614]_ ,
    \new_[19615]_ , \new_[19616]_ , \new_[19619]_ , \new_[19623]_ ,
    \new_[19624]_ , \new_[19625]_ , \new_[19629]_ , \new_[19630]_ ,
    \new_[19634]_ , \new_[19635]_ , \new_[19636]_ , \new_[19639]_ ,
    \new_[19643]_ , \new_[19644]_ , \new_[19645]_ , \new_[19649]_ ,
    \new_[19650]_ , \new_[19654]_ , \new_[19655]_ , \new_[19656]_ ,
    \new_[19659]_ , \new_[19663]_ , \new_[19664]_ , \new_[19665]_ ,
    \new_[19669]_ , \new_[19670]_ , \new_[19674]_ , \new_[19675]_ ,
    \new_[19676]_ , \new_[19679]_ , \new_[19683]_ , \new_[19684]_ ,
    \new_[19685]_ , \new_[19689]_ , \new_[19690]_ , \new_[19694]_ ,
    \new_[19695]_ , \new_[19696]_ , \new_[19699]_ , \new_[19703]_ ,
    \new_[19704]_ , \new_[19705]_ , \new_[19709]_ , \new_[19710]_ ,
    \new_[19714]_ , \new_[19715]_ , \new_[19716]_ , \new_[19719]_ ,
    \new_[19723]_ , \new_[19724]_ , \new_[19725]_ , \new_[19729]_ ,
    \new_[19730]_ , \new_[19734]_ , \new_[19735]_ , \new_[19736]_ ,
    \new_[19739]_ , \new_[19743]_ , \new_[19744]_ , \new_[19745]_ ,
    \new_[19749]_ , \new_[19750]_ , \new_[19754]_ , \new_[19755]_ ,
    \new_[19756]_ , \new_[19759]_ , \new_[19763]_ , \new_[19764]_ ,
    \new_[19765]_ , \new_[19769]_ , \new_[19770]_ , \new_[19774]_ ,
    \new_[19775]_ , \new_[19776]_ , \new_[19779]_ , \new_[19783]_ ,
    \new_[19784]_ , \new_[19785]_ , \new_[19789]_ , \new_[19790]_ ,
    \new_[19794]_ , \new_[19795]_ , \new_[19796]_ , \new_[19799]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19805]_ , \new_[19809]_ ,
    \new_[19810]_ , \new_[19814]_ , \new_[19815]_ , \new_[19816]_ ,
    \new_[19819]_ , \new_[19823]_ , \new_[19824]_ , \new_[19825]_ ,
    \new_[19829]_ , \new_[19830]_ , \new_[19834]_ , \new_[19835]_ ,
    \new_[19836]_ , \new_[19839]_ , \new_[19843]_ , \new_[19844]_ ,
    \new_[19845]_ , \new_[19849]_ , \new_[19850]_ , \new_[19854]_ ,
    \new_[19855]_ , \new_[19856]_ , \new_[19859]_ , \new_[19863]_ ,
    \new_[19864]_ , \new_[19865]_ , \new_[19869]_ , \new_[19870]_ ,
    \new_[19874]_ , \new_[19875]_ , \new_[19876]_ , \new_[19879]_ ,
    \new_[19883]_ , \new_[19884]_ , \new_[19885]_ , \new_[19889]_ ,
    \new_[19890]_ , \new_[19894]_ , \new_[19895]_ , \new_[19896]_ ,
    \new_[19899]_ , \new_[19903]_ , \new_[19904]_ , \new_[19905]_ ,
    \new_[19909]_ , \new_[19910]_ , \new_[19914]_ , \new_[19915]_ ,
    \new_[19916]_ , \new_[19919]_ , \new_[19923]_ , \new_[19924]_ ,
    \new_[19925]_ , \new_[19929]_ , \new_[19930]_ , \new_[19934]_ ,
    \new_[19935]_ , \new_[19936]_ , \new_[19939]_ , \new_[19943]_ ,
    \new_[19944]_ , \new_[19945]_ , \new_[19949]_ , \new_[19950]_ ,
    \new_[19954]_ , \new_[19955]_ , \new_[19956]_ , \new_[19959]_ ,
    \new_[19963]_ , \new_[19964]_ , \new_[19965]_ , \new_[19969]_ ,
    \new_[19970]_ , \new_[19974]_ , \new_[19975]_ , \new_[19976]_ ,
    \new_[19979]_ , \new_[19983]_ , \new_[19984]_ , \new_[19985]_ ,
    \new_[19989]_ , \new_[19990]_ , \new_[19994]_ , \new_[19995]_ ,
    \new_[19996]_ , \new_[19999]_ , \new_[20003]_ , \new_[20004]_ ,
    \new_[20005]_ , \new_[20009]_ , \new_[20010]_ , \new_[20014]_ ,
    \new_[20015]_ , \new_[20016]_ , \new_[20019]_ , \new_[20023]_ ,
    \new_[20024]_ , \new_[20025]_ , \new_[20029]_ , \new_[20030]_ ,
    \new_[20034]_ , \new_[20035]_ , \new_[20036]_ , \new_[20039]_ ,
    \new_[20043]_ , \new_[20044]_ , \new_[20045]_ , \new_[20049]_ ,
    \new_[20050]_ , \new_[20054]_ , \new_[20055]_ , \new_[20056]_ ,
    \new_[20059]_ , \new_[20063]_ , \new_[20064]_ , \new_[20065]_ ,
    \new_[20069]_ , \new_[20070]_ , \new_[20074]_ , \new_[20075]_ ,
    \new_[20076]_ , \new_[20079]_ , \new_[20083]_ , \new_[20084]_ ,
    \new_[20085]_ , \new_[20089]_ , \new_[20090]_ , \new_[20094]_ ,
    \new_[20095]_ , \new_[20096]_ , \new_[20099]_ , \new_[20103]_ ,
    \new_[20104]_ , \new_[20105]_ , \new_[20109]_ , \new_[20110]_ ,
    \new_[20114]_ , \new_[20115]_ , \new_[20116]_ , \new_[20119]_ ,
    \new_[20123]_ , \new_[20124]_ , \new_[20125]_ , \new_[20129]_ ,
    \new_[20130]_ , \new_[20134]_ , \new_[20135]_ , \new_[20136]_ ,
    \new_[20139]_ , \new_[20143]_ , \new_[20144]_ , \new_[20145]_ ,
    \new_[20149]_ , \new_[20150]_ , \new_[20154]_ , \new_[20155]_ ,
    \new_[20156]_ , \new_[20159]_ , \new_[20163]_ , \new_[20164]_ ,
    \new_[20165]_ , \new_[20169]_ , \new_[20170]_ , \new_[20174]_ ,
    \new_[20175]_ , \new_[20176]_ , \new_[20179]_ , \new_[20183]_ ,
    \new_[20184]_ , \new_[20185]_ , \new_[20189]_ , \new_[20190]_ ,
    \new_[20194]_ , \new_[20195]_ , \new_[20196]_ , \new_[20199]_ ,
    \new_[20203]_ , \new_[20204]_ , \new_[20205]_ , \new_[20209]_ ,
    \new_[20210]_ , \new_[20214]_ , \new_[20215]_ , \new_[20216]_ ,
    \new_[20219]_ , \new_[20223]_ , \new_[20224]_ , \new_[20225]_ ,
    \new_[20229]_ , \new_[20230]_ , \new_[20234]_ , \new_[20235]_ ,
    \new_[20236]_ , \new_[20239]_ , \new_[20243]_ , \new_[20244]_ ,
    \new_[20245]_ , \new_[20249]_ , \new_[20250]_ , \new_[20254]_ ,
    \new_[20255]_ , \new_[20256]_ , \new_[20259]_ , \new_[20263]_ ,
    \new_[20264]_ , \new_[20265]_ , \new_[20269]_ , \new_[20270]_ ,
    \new_[20274]_ , \new_[20275]_ , \new_[20276]_ , \new_[20279]_ ,
    \new_[20283]_ , \new_[20284]_ , \new_[20285]_ , \new_[20289]_ ,
    \new_[20290]_ , \new_[20294]_ , \new_[20295]_ , \new_[20296]_ ,
    \new_[20299]_ , \new_[20303]_ , \new_[20304]_ , \new_[20305]_ ,
    \new_[20309]_ , \new_[20310]_ , \new_[20314]_ , \new_[20315]_ ,
    \new_[20316]_ , \new_[20319]_ , \new_[20323]_ , \new_[20324]_ ,
    \new_[20325]_ , \new_[20329]_ , \new_[20330]_ , \new_[20334]_ ,
    \new_[20335]_ , \new_[20336]_ , \new_[20339]_ , \new_[20343]_ ,
    \new_[20344]_ , \new_[20345]_ , \new_[20349]_ , \new_[20350]_ ,
    \new_[20354]_ , \new_[20355]_ , \new_[20356]_ , \new_[20359]_ ,
    \new_[20363]_ , \new_[20364]_ , \new_[20365]_ , \new_[20369]_ ,
    \new_[20370]_ , \new_[20374]_ , \new_[20375]_ , \new_[20376]_ ,
    \new_[20379]_ , \new_[20383]_ , \new_[20384]_ , \new_[20385]_ ,
    \new_[20389]_ , \new_[20390]_ , \new_[20394]_ , \new_[20395]_ ,
    \new_[20396]_ , \new_[20399]_ , \new_[20403]_ , \new_[20404]_ ,
    \new_[20405]_ , \new_[20409]_ , \new_[20410]_ , \new_[20414]_ ,
    \new_[20415]_ , \new_[20416]_ , \new_[20419]_ , \new_[20423]_ ,
    \new_[20424]_ , \new_[20425]_ , \new_[20429]_ , \new_[20430]_ ,
    \new_[20434]_ , \new_[20435]_ , \new_[20436]_ , \new_[20439]_ ,
    \new_[20443]_ , \new_[20444]_ , \new_[20445]_ , \new_[20449]_ ,
    \new_[20450]_ , \new_[20454]_ , \new_[20455]_ , \new_[20456]_ ,
    \new_[20459]_ , \new_[20463]_ , \new_[20464]_ , \new_[20465]_ ,
    \new_[20469]_ , \new_[20470]_ , \new_[20474]_ , \new_[20475]_ ,
    \new_[20476]_ , \new_[20479]_ , \new_[20483]_ , \new_[20484]_ ,
    \new_[20485]_ , \new_[20489]_ , \new_[20490]_ , \new_[20494]_ ,
    \new_[20495]_ , \new_[20496]_ , \new_[20499]_ , \new_[20503]_ ,
    \new_[20504]_ , \new_[20505]_ , \new_[20509]_ , \new_[20510]_ ,
    \new_[20514]_ , \new_[20515]_ , \new_[20516]_ , \new_[20519]_ ,
    \new_[20523]_ , \new_[20524]_ , \new_[20525]_ , \new_[20529]_ ,
    \new_[20530]_ , \new_[20534]_ , \new_[20535]_ , \new_[20536]_ ,
    \new_[20539]_ , \new_[20543]_ , \new_[20544]_ , \new_[20545]_ ,
    \new_[20549]_ , \new_[20550]_ , \new_[20554]_ , \new_[20555]_ ,
    \new_[20556]_ , \new_[20559]_ , \new_[20563]_ , \new_[20564]_ ,
    \new_[20565]_ , \new_[20569]_ , \new_[20570]_ , \new_[20574]_ ,
    \new_[20575]_ , \new_[20576]_ , \new_[20579]_ , \new_[20583]_ ,
    \new_[20584]_ , \new_[20585]_ , \new_[20589]_ , \new_[20590]_ ,
    \new_[20594]_ , \new_[20595]_ , \new_[20596]_ , \new_[20599]_ ,
    \new_[20603]_ , \new_[20604]_ , \new_[20605]_ , \new_[20609]_ ,
    \new_[20610]_ , \new_[20614]_ , \new_[20615]_ , \new_[20616]_ ,
    \new_[20619]_ , \new_[20623]_ , \new_[20624]_ , \new_[20625]_ ,
    \new_[20629]_ , \new_[20630]_ , \new_[20634]_ , \new_[20635]_ ,
    \new_[20636]_ , \new_[20639]_ , \new_[20643]_ , \new_[20644]_ ,
    \new_[20645]_ , \new_[20649]_ , \new_[20650]_ , \new_[20654]_ ,
    \new_[20655]_ , \new_[20656]_ , \new_[20659]_ , \new_[20663]_ ,
    \new_[20664]_ , \new_[20665]_ , \new_[20669]_ , \new_[20670]_ ,
    \new_[20674]_ , \new_[20675]_ , \new_[20676]_ , \new_[20679]_ ,
    \new_[20683]_ , \new_[20684]_ , \new_[20685]_ , \new_[20689]_ ,
    \new_[20690]_ , \new_[20694]_ , \new_[20695]_ , \new_[20696]_ ,
    \new_[20699]_ , \new_[20703]_ , \new_[20704]_ , \new_[20705]_ ,
    \new_[20709]_ , \new_[20710]_ , \new_[20714]_ , \new_[20715]_ ,
    \new_[20716]_ , \new_[20719]_ , \new_[20723]_ , \new_[20724]_ ,
    \new_[20725]_ , \new_[20729]_ , \new_[20730]_ , \new_[20734]_ ,
    \new_[20735]_ , \new_[20736]_ , \new_[20739]_ , \new_[20743]_ ,
    \new_[20744]_ , \new_[20745]_ , \new_[20749]_ , \new_[20750]_ ,
    \new_[20754]_ , \new_[20755]_ , \new_[20756]_ , \new_[20759]_ ,
    \new_[20763]_ , \new_[20764]_ , \new_[20765]_ , \new_[20769]_ ,
    \new_[20770]_ , \new_[20774]_ , \new_[20775]_ , \new_[20776]_ ,
    \new_[20779]_ , \new_[20783]_ , \new_[20784]_ , \new_[20785]_ ,
    \new_[20789]_ , \new_[20790]_ , \new_[20794]_ , \new_[20795]_ ,
    \new_[20796]_ , \new_[20799]_ , \new_[20803]_ , \new_[20804]_ ,
    \new_[20805]_ , \new_[20809]_ , \new_[20810]_ , \new_[20814]_ ,
    \new_[20815]_ , \new_[20816]_ , \new_[20819]_ , \new_[20823]_ ,
    \new_[20824]_ , \new_[20825]_ , \new_[20829]_ , \new_[20830]_ ,
    \new_[20834]_ , \new_[20835]_ , \new_[20836]_ , \new_[20839]_ ,
    \new_[20843]_ , \new_[20844]_ , \new_[20845]_ , \new_[20849]_ ,
    \new_[20850]_ , \new_[20854]_ , \new_[20855]_ , \new_[20856]_ ,
    \new_[20859]_ , \new_[20863]_ , \new_[20864]_ , \new_[20865]_ ,
    \new_[20869]_ , \new_[20870]_ , \new_[20874]_ , \new_[20875]_ ,
    \new_[20876]_ , \new_[20879]_ , \new_[20883]_ , \new_[20884]_ ,
    \new_[20885]_ , \new_[20889]_ , \new_[20890]_ , \new_[20894]_ ,
    \new_[20895]_ , \new_[20896]_ , \new_[20899]_ , \new_[20903]_ ,
    \new_[20904]_ , \new_[20905]_ , \new_[20909]_ , \new_[20910]_ ,
    \new_[20914]_ , \new_[20915]_ , \new_[20916]_ , \new_[20919]_ ,
    \new_[20923]_ , \new_[20924]_ , \new_[20925]_ , \new_[20929]_ ,
    \new_[20930]_ , \new_[20934]_ , \new_[20935]_ , \new_[20936]_ ,
    \new_[20939]_ , \new_[20943]_ , \new_[20944]_ , \new_[20945]_ ,
    \new_[20949]_ , \new_[20950]_ , \new_[20954]_ , \new_[20955]_ ,
    \new_[20956]_ , \new_[20959]_ , \new_[20963]_ , \new_[20964]_ ,
    \new_[20965]_ , \new_[20969]_ , \new_[20970]_ , \new_[20974]_ ,
    \new_[20975]_ , \new_[20976]_ , \new_[20979]_ , \new_[20983]_ ,
    \new_[20984]_ , \new_[20985]_ , \new_[20989]_ , \new_[20990]_ ,
    \new_[20994]_ , \new_[20995]_ , \new_[20996]_ , \new_[20999]_ ,
    \new_[21003]_ , \new_[21004]_ , \new_[21005]_ , \new_[21009]_ ,
    \new_[21010]_ , \new_[21014]_ , \new_[21015]_ , \new_[21016]_ ,
    \new_[21019]_ , \new_[21023]_ , \new_[21024]_ , \new_[21025]_ ,
    \new_[21029]_ , \new_[21030]_ , \new_[21034]_ , \new_[21035]_ ,
    \new_[21036]_ , \new_[21039]_ , \new_[21043]_ , \new_[21044]_ ,
    \new_[21045]_ , \new_[21049]_ , \new_[21050]_ , \new_[21054]_ ,
    \new_[21055]_ , \new_[21056]_ , \new_[21059]_ , \new_[21063]_ ,
    \new_[21064]_ , \new_[21065]_ , \new_[21069]_ , \new_[21070]_ ,
    \new_[21074]_ , \new_[21075]_ , \new_[21076]_ , \new_[21079]_ ,
    \new_[21083]_ , \new_[21084]_ , \new_[21085]_ , \new_[21089]_ ,
    \new_[21090]_ , \new_[21094]_ , \new_[21095]_ , \new_[21096]_ ,
    \new_[21099]_ , \new_[21103]_ , \new_[21104]_ , \new_[21105]_ ,
    \new_[21109]_ , \new_[21110]_ , \new_[21114]_ , \new_[21115]_ ,
    \new_[21116]_ , \new_[21119]_ , \new_[21123]_ , \new_[21124]_ ,
    \new_[21125]_ , \new_[21129]_ , \new_[21130]_ , \new_[21134]_ ,
    \new_[21135]_ , \new_[21136]_ , \new_[21139]_ , \new_[21143]_ ,
    \new_[21144]_ , \new_[21145]_ , \new_[21149]_ , \new_[21150]_ ,
    \new_[21154]_ , \new_[21155]_ , \new_[21156]_ , \new_[21159]_ ,
    \new_[21163]_ , \new_[21164]_ , \new_[21165]_ , \new_[21169]_ ,
    \new_[21170]_ , \new_[21174]_ , \new_[21175]_ , \new_[21176]_ ,
    \new_[21179]_ , \new_[21183]_ , \new_[21184]_ , \new_[21185]_ ,
    \new_[21189]_ , \new_[21190]_ , \new_[21194]_ , \new_[21195]_ ,
    \new_[21196]_ , \new_[21199]_ , \new_[21203]_ , \new_[21204]_ ,
    \new_[21205]_ , \new_[21209]_ , \new_[21210]_ , \new_[21214]_ ,
    \new_[21215]_ , \new_[21216]_ , \new_[21219]_ , \new_[21223]_ ,
    \new_[21224]_ , \new_[21225]_ , \new_[21229]_ , \new_[21230]_ ,
    \new_[21234]_ , \new_[21235]_ , \new_[21236]_ , \new_[21239]_ ,
    \new_[21243]_ , \new_[21244]_ , \new_[21245]_ , \new_[21249]_ ,
    \new_[21250]_ , \new_[21254]_ , \new_[21255]_ , \new_[21256]_ ,
    \new_[21259]_ , \new_[21263]_ , \new_[21264]_ , \new_[21265]_ ,
    \new_[21269]_ , \new_[21270]_ , \new_[21274]_ , \new_[21275]_ ,
    \new_[21276]_ , \new_[21279]_ , \new_[21283]_ , \new_[21284]_ ,
    \new_[21285]_ , \new_[21289]_ , \new_[21290]_ , \new_[21294]_ ,
    \new_[21295]_ , \new_[21296]_ , \new_[21299]_ , \new_[21303]_ ,
    \new_[21304]_ , \new_[21305]_ , \new_[21309]_ , \new_[21310]_ ,
    \new_[21314]_ , \new_[21315]_ , \new_[21316]_ , \new_[21319]_ ,
    \new_[21323]_ , \new_[21324]_ , \new_[21325]_ , \new_[21329]_ ,
    \new_[21330]_ , \new_[21334]_ , \new_[21335]_ , \new_[21336]_ ,
    \new_[21339]_ , \new_[21343]_ , \new_[21344]_ , \new_[21345]_ ,
    \new_[21349]_ , \new_[21350]_ , \new_[21354]_ , \new_[21355]_ ,
    \new_[21356]_ , \new_[21359]_ , \new_[21363]_ , \new_[21364]_ ,
    \new_[21365]_ , \new_[21369]_ , \new_[21370]_ , \new_[21374]_ ,
    \new_[21375]_ , \new_[21376]_ , \new_[21379]_ , \new_[21383]_ ,
    \new_[21384]_ , \new_[21385]_ , \new_[21389]_ , \new_[21390]_ ,
    \new_[21394]_ , \new_[21395]_ , \new_[21396]_ , \new_[21399]_ ,
    \new_[21403]_ , \new_[21404]_ , \new_[21405]_ , \new_[21409]_ ,
    \new_[21410]_ , \new_[21414]_ , \new_[21415]_ , \new_[21416]_ ,
    \new_[21419]_ , \new_[21423]_ , \new_[21424]_ , \new_[21425]_ ,
    \new_[21429]_ , \new_[21430]_ , \new_[21434]_ , \new_[21435]_ ,
    \new_[21436]_ , \new_[21439]_ , \new_[21443]_ , \new_[21444]_ ,
    \new_[21445]_ , \new_[21449]_ , \new_[21450]_ , \new_[21454]_ ,
    \new_[21455]_ , \new_[21456]_ , \new_[21459]_ , \new_[21463]_ ,
    \new_[21464]_ , \new_[21465]_ , \new_[21469]_ , \new_[21470]_ ,
    \new_[21474]_ , \new_[21475]_ , \new_[21476]_ , \new_[21479]_ ,
    \new_[21483]_ , \new_[21484]_ , \new_[21485]_ , \new_[21489]_ ,
    \new_[21490]_ , \new_[21494]_ , \new_[21495]_ , \new_[21496]_ ,
    \new_[21499]_ , \new_[21503]_ , \new_[21504]_ , \new_[21505]_ ,
    \new_[21509]_ , \new_[21510]_ , \new_[21514]_ , \new_[21515]_ ,
    \new_[21516]_ , \new_[21519]_ , \new_[21523]_ , \new_[21524]_ ,
    \new_[21525]_ , \new_[21529]_ , \new_[21530]_ , \new_[21534]_ ,
    \new_[21535]_ , \new_[21536]_ , \new_[21539]_ , \new_[21543]_ ,
    \new_[21544]_ , \new_[21545]_ , \new_[21549]_ , \new_[21550]_ ,
    \new_[21554]_ , \new_[21555]_ , \new_[21556]_ , \new_[21559]_ ,
    \new_[21563]_ , \new_[21564]_ , \new_[21565]_ , \new_[21569]_ ,
    \new_[21570]_ , \new_[21574]_ , \new_[21575]_ , \new_[21576]_ ,
    \new_[21579]_ , \new_[21583]_ , \new_[21584]_ , \new_[21585]_ ,
    \new_[21589]_ , \new_[21590]_ , \new_[21594]_ , \new_[21595]_ ,
    \new_[21596]_ , \new_[21599]_ , \new_[21603]_ , \new_[21604]_ ,
    \new_[21605]_ , \new_[21609]_ , \new_[21610]_ , \new_[21614]_ ,
    \new_[21615]_ , \new_[21616]_ , \new_[21619]_ , \new_[21623]_ ,
    \new_[21624]_ , \new_[21625]_ , \new_[21629]_ , \new_[21630]_ ,
    \new_[21634]_ , \new_[21635]_ , \new_[21636]_ , \new_[21639]_ ,
    \new_[21643]_ , \new_[21644]_ , \new_[21645]_ , \new_[21649]_ ,
    \new_[21650]_ , \new_[21654]_ , \new_[21655]_ , \new_[21656]_ ,
    \new_[21659]_ , \new_[21663]_ , \new_[21664]_ , \new_[21665]_ ,
    \new_[21669]_ , \new_[21670]_ , \new_[21674]_ , \new_[21675]_ ,
    \new_[21676]_ , \new_[21679]_ , \new_[21683]_ , \new_[21684]_ ,
    \new_[21685]_ , \new_[21689]_ , \new_[21690]_ , \new_[21694]_ ,
    \new_[21695]_ , \new_[21696]_ , \new_[21699]_ , \new_[21703]_ ,
    \new_[21704]_ , \new_[21705]_ , \new_[21709]_ , \new_[21710]_ ,
    \new_[21714]_ , \new_[21715]_ , \new_[21716]_ , \new_[21719]_ ,
    \new_[21723]_ , \new_[21724]_ , \new_[21725]_ , \new_[21729]_ ,
    \new_[21730]_ , \new_[21734]_ , \new_[21735]_ , \new_[21736]_ ,
    \new_[21739]_ , \new_[21743]_ , \new_[21744]_ , \new_[21745]_ ,
    \new_[21749]_ , \new_[21750]_ , \new_[21754]_ , \new_[21755]_ ,
    \new_[21756]_ , \new_[21759]_ , \new_[21763]_ , \new_[21764]_ ,
    \new_[21765]_ , \new_[21769]_ , \new_[21770]_ , \new_[21774]_ ,
    \new_[21775]_ , \new_[21776]_ , \new_[21779]_ , \new_[21783]_ ,
    \new_[21784]_ , \new_[21785]_ , \new_[21789]_ , \new_[21790]_ ,
    \new_[21794]_ , \new_[21795]_ , \new_[21796]_ , \new_[21799]_ ,
    \new_[21803]_ , \new_[21804]_ , \new_[21805]_ , \new_[21809]_ ,
    \new_[21810]_ , \new_[21814]_ , \new_[21815]_ , \new_[21816]_ ,
    \new_[21819]_ , \new_[21823]_ , \new_[21824]_ , \new_[21825]_ ,
    \new_[21829]_ , \new_[21830]_ , \new_[21834]_ , \new_[21835]_ ,
    \new_[21836]_ , \new_[21839]_ , \new_[21843]_ , \new_[21844]_ ,
    \new_[21845]_ , \new_[21849]_ , \new_[21850]_ , \new_[21854]_ ,
    \new_[21855]_ , \new_[21856]_ , \new_[21859]_ , \new_[21863]_ ,
    \new_[21864]_ , \new_[21865]_ , \new_[21869]_ , \new_[21870]_ ,
    \new_[21874]_ , \new_[21875]_ , \new_[21876]_ , \new_[21879]_ ,
    \new_[21883]_ , \new_[21884]_ , \new_[21885]_ , \new_[21889]_ ,
    \new_[21890]_ , \new_[21894]_ , \new_[21895]_ , \new_[21896]_ ,
    \new_[21899]_ , \new_[21903]_ , \new_[21904]_ , \new_[21905]_ ,
    \new_[21909]_ , \new_[21910]_ , \new_[21914]_ , \new_[21915]_ ,
    \new_[21916]_ , \new_[21919]_ , \new_[21923]_ , \new_[21924]_ ,
    \new_[21925]_ , \new_[21929]_ , \new_[21930]_ , \new_[21934]_ ,
    \new_[21935]_ , \new_[21936]_ , \new_[21939]_ , \new_[21943]_ ,
    \new_[21944]_ , \new_[21945]_ , \new_[21949]_ , \new_[21950]_ ,
    \new_[21954]_ , \new_[21955]_ , \new_[21956]_ , \new_[21959]_ ,
    \new_[21963]_ , \new_[21964]_ , \new_[21965]_ , \new_[21969]_ ,
    \new_[21970]_ , \new_[21974]_ , \new_[21975]_ , \new_[21976]_ ,
    \new_[21979]_ , \new_[21983]_ , \new_[21984]_ , \new_[21985]_ ,
    \new_[21989]_ , \new_[21990]_ , \new_[21994]_ , \new_[21995]_ ,
    \new_[21996]_ , \new_[21999]_ , \new_[22003]_ , \new_[22004]_ ,
    \new_[22005]_ , \new_[22009]_ , \new_[22010]_ , \new_[22014]_ ,
    \new_[22015]_ , \new_[22016]_ , \new_[22019]_ , \new_[22023]_ ,
    \new_[22024]_ , \new_[22025]_ , \new_[22029]_ , \new_[22030]_ ,
    \new_[22034]_ , \new_[22035]_ , \new_[22036]_ , \new_[22039]_ ,
    \new_[22043]_ , \new_[22044]_ , \new_[22045]_ , \new_[22049]_ ,
    \new_[22050]_ , \new_[22054]_ , \new_[22055]_ , \new_[22056]_ ,
    \new_[22059]_ , \new_[22063]_ , \new_[22064]_ , \new_[22065]_ ,
    \new_[22069]_ , \new_[22070]_ , \new_[22074]_ , \new_[22075]_ ,
    \new_[22076]_ , \new_[22079]_ , \new_[22083]_ , \new_[22084]_ ,
    \new_[22085]_ , \new_[22089]_ , \new_[22090]_ , \new_[22094]_ ,
    \new_[22095]_ , \new_[22096]_ , \new_[22099]_ , \new_[22103]_ ,
    \new_[22104]_ , \new_[22105]_ , \new_[22109]_ , \new_[22110]_ ,
    \new_[22114]_ , \new_[22115]_ , \new_[22116]_ , \new_[22119]_ ,
    \new_[22123]_ , \new_[22124]_ , \new_[22125]_ , \new_[22129]_ ,
    \new_[22130]_ , \new_[22134]_ , \new_[22135]_ , \new_[22136]_ ,
    \new_[22139]_ , \new_[22143]_ , \new_[22144]_ , \new_[22145]_ ,
    \new_[22149]_ , \new_[22150]_ , \new_[22154]_ , \new_[22155]_ ,
    \new_[22156]_ , \new_[22159]_ , \new_[22163]_ , \new_[22164]_ ,
    \new_[22165]_ , \new_[22169]_ , \new_[22170]_ , \new_[22174]_ ,
    \new_[22175]_ , \new_[22176]_ , \new_[22179]_ , \new_[22183]_ ,
    \new_[22184]_ , \new_[22185]_ , \new_[22189]_ , \new_[22190]_ ,
    \new_[22194]_ , \new_[22195]_ , \new_[22196]_ , \new_[22199]_ ,
    \new_[22203]_ , \new_[22204]_ , \new_[22205]_ , \new_[22209]_ ,
    \new_[22210]_ , \new_[22214]_ , \new_[22215]_ , \new_[22216]_ ,
    \new_[22219]_ , \new_[22223]_ , \new_[22224]_ , \new_[22225]_ ,
    \new_[22229]_ , \new_[22230]_ , \new_[22234]_ , \new_[22235]_ ,
    \new_[22236]_ , \new_[22239]_ , \new_[22243]_ , \new_[22244]_ ,
    \new_[22245]_ , \new_[22249]_ , \new_[22250]_ , \new_[22254]_ ,
    \new_[22255]_ , \new_[22256]_ , \new_[22259]_ , \new_[22263]_ ,
    \new_[22264]_ , \new_[22265]_ , \new_[22269]_ , \new_[22270]_ ,
    \new_[22274]_ , \new_[22275]_ , \new_[22276]_ , \new_[22279]_ ,
    \new_[22283]_ , \new_[22284]_ , \new_[22285]_ , \new_[22289]_ ,
    \new_[22290]_ , \new_[22294]_ , \new_[22295]_ , \new_[22296]_ ,
    \new_[22299]_ , \new_[22303]_ , \new_[22304]_ , \new_[22305]_ ,
    \new_[22309]_ , \new_[22310]_ , \new_[22314]_ , \new_[22315]_ ,
    \new_[22316]_ , \new_[22319]_ , \new_[22323]_ , \new_[22324]_ ,
    \new_[22325]_ , \new_[22329]_ , \new_[22330]_ , \new_[22334]_ ,
    \new_[22335]_ , \new_[22336]_ , \new_[22339]_ , \new_[22343]_ ,
    \new_[22344]_ , \new_[22345]_ , \new_[22349]_ , \new_[22350]_ ,
    \new_[22354]_ , \new_[22355]_ , \new_[22356]_ , \new_[22359]_ ,
    \new_[22363]_ , \new_[22364]_ , \new_[22365]_ , \new_[22369]_ ,
    \new_[22370]_ , \new_[22374]_ , \new_[22375]_ , \new_[22376]_ ,
    \new_[22379]_ , \new_[22383]_ , \new_[22384]_ , \new_[22385]_ ,
    \new_[22389]_ , \new_[22390]_ , \new_[22394]_ , \new_[22395]_ ,
    \new_[22396]_ , \new_[22399]_ , \new_[22403]_ , \new_[22404]_ ,
    \new_[22405]_ , \new_[22409]_ , \new_[22410]_ , \new_[22414]_ ,
    \new_[22415]_ , \new_[22416]_ , \new_[22419]_ , \new_[22423]_ ,
    \new_[22424]_ , \new_[22425]_ , \new_[22429]_ , \new_[22430]_ ,
    \new_[22434]_ , \new_[22435]_ , \new_[22436]_ , \new_[22439]_ ,
    \new_[22443]_ , \new_[22444]_ , \new_[22445]_ , \new_[22449]_ ,
    \new_[22450]_ , \new_[22454]_ , \new_[22455]_ , \new_[22456]_ ,
    \new_[22459]_ , \new_[22463]_ , \new_[22464]_ , \new_[22465]_ ,
    \new_[22469]_ , \new_[22470]_ , \new_[22474]_ , \new_[22475]_ ,
    \new_[22476]_ , \new_[22479]_ , \new_[22483]_ , \new_[22484]_ ,
    \new_[22485]_ , \new_[22489]_ , \new_[22490]_ , \new_[22494]_ ,
    \new_[22495]_ , \new_[22496]_ , \new_[22499]_ , \new_[22503]_ ,
    \new_[22504]_ , \new_[22505]_ , \new_[22509]_ , \new_[22510]_ ,
    \new_[22514]_ , \new_[22515]_ , \new_[22516]_ , \new_[22519]_ ,
    \new_[22523]_ , \new_[22524]_ , \new_[22525]_ , \new_[22529]_ ,
    \new_[22530]_ , \new_[22534]_ , \new_[22535]_ , \new_[22536]_ ,
    \new_[22539]_ , \new_[22543]_ , \new_[22544]_ , \new_[22545]_ ,
    \new_[22549]_ , \new_[22550]_ , \new_[22554]_ , \new_[22555]_ ,
    \new_[22556]_ , \new_[22559]_ , \new_[22563]_ , \new_[22564]_ ,
    \new_[22565]_ , \new_[22569]_ , \new_[22570]_ , \new_[22574]_ ,
    \new_[22575]_ , \new_[22576]_ , \new_[22579]_ , \new_[22583]_ ,
    \new_[22584]_ , \new_[22585]_ , \new_[22589]_ , \new_[22590]_ ,
    \new_[22594]_ , \new_[22595]_ , \new_[22596]_ , \new_[22599]_ ,
    \new_[22603]_ , \new_[22604]_ , \new_[22605]_ , \new_[22609]_ ,
    \new_[22610]_ , \new_[22614]_ , \new_[22615]_ , \new_[22616]_ ,
    \new_[22619]_ , \new_[22623]_ , \new_[22624]_ , \new_[22625]_ ,
    \new_[22629]_ , \new_[22630]_ , \new_[22634]_ , \new_[22635]_ ,
    \new_[22636]_ , \new_[22639]_ , \new_[22643]_ , \new_[22644]_ ,
    \new_[22645]_ , \new_[22649]_ , \new_[22650]_ , \new_[22654]_ ,
    \new_[22655]_ , \new_[22656]_ , \new_[22659]_ , \new_[22663]_ ,
    \new_[22664]_ , \new_[22665]_ , \new_[22669]_ , \new_[22670]_ ,
    \new_[22674]_ , \new_[22675]_ , \new_[22676]_ , \new_[22679]_ ,
    \new_[22683]_ , \new_[22684]_ , \new_[22685]_ , \new_[22689]_ ,
    \new_[22690]_ , \new_[22694]_ , \new_[22695]_ , \new_[22696]_ ,
    \new_[22699]_ , \new_[22703]_ , \new_[22704]_ , \new_[22705]_ ,
    \new_[22709]_ , \new_[22710]_ , \new_[22714]_ , \new_[22715]_ ,
    \new_[22716]_ , \new_[22719]_ , \new_[22723]_ , \new_[22724]_ ,
    \new_[22725]_ , \new_[22729]_ , \new_[22730]_ , \new_[22734]_ ,
    \new_[22735]_ , \new_[22736]_ , \new_[22739]_ , \new_[22743]_ ,
    \new_[22744]_ , \new_[22745]_ , \new_[22749]_ , \new_[22750]_ ,
    \new_[22754]_ , \new_[22755]_ , \new_[22756]_ , \new_[22759]_ ,
    \new_[22763]_ , \new_[22764]_ , \new_[22765]_ , \new_[22769]_ ,
    \new_[22770]_ , \new_[22774]_ , \new_[22775]_ , \new_[22776]_ ,
    \new_[22779]_ , \new_[22783]_ , \new_[22784]_ , \new_[22785]_ ,
    \new_[22789]_ , \new_[22790]_ , \new_[22794]_ , \new_[22795]_ ,
    \new_[22796]_ , \new_[22799]_ , \new_[22803]_ , \new_[22804]_ ,
    \new_[22805]_ , \new_[22809]_ , \new_[22810]_ , \new_[22814]_ ,
    \new_[22815]_ , \new_[22816]_ , \new_[22819]_ , \new_[22823]_ ,
    \new_[22824]_ , \new_[22825]_ , \new_[22829]_ , \new_[22830]_ ,
    \new_[22834]_ , \new_[22835]_ , \new_[22836]_ , \new_[22839]_ ,
    \new_[22843]_ , \new_[22844]_ , \new_[22845]_ , \new_[22849]_ ,
    \new_[22850]_ , \new_[22854]_ , \new_[22855]_ , \new_[22856]_ ,
    \new_[22859]_ , \new_[22863]_ , \new_[22864]_ , \new_[22865]_ ,
    \new_[22869]_ , \new_[22870]_ , \new_[22874]_ , \new_[22875]_ ,
    \new_[22876]_ , \new_[22879]_ , \new_[22883]_ , \new_[22884]_ ,
    \new_[22885]_ , \new_[22889]_ , \new_[22890]_ , \new_[22894]_ ,
    \new_[22895]_ , \new_[22896]_ , \new_[22899]_ , \new_[22903]_ ,
    \new_[22904]_ , \new_[22905]_ , \new_[22909]_ , \new_[22910]_ ,
    \new_[22914]_ , \new_[22915]_ , \new_[22916]_ , \new_[22919]_ ,
    \new_[22923]_ , \new_[22924]_ , \new_[22925]_ , \new_[22929]_ ,
    \new_[22930]_ , \new_[22934]_ , \new_[22935]_ , \new_[22936]_ ,
    \new_[22939]_ , \new_[22943]_ , \new_[22944]_ , \new_[22945]_ ,
    \new_[22949]_ , \new_[22950]_ , \new_[22954]_ , \new_[22955]_ ,
    \new_[22956]_ , \new_[22959]_ , \new_[22963]_ , \new_[22964]_ ,
    \new_[22965]_ , \new_[22969]_ , \new_[22970]_ , \new_[22974]_ ,
    \new_[22975]_ , \new_[22976]_ , \new_[22979]_ , \new_[22983]_ ,
    \new_[22984]_ , \new_[22985]_ , \new_[22989]_ , \new_[22990]_ ,
    \new_[22994]_ , \new_[22995]_ , \new_[22996]_ , \new_[22999]_ ,
    \new_[23003]_ , \new_[23004]_ , \new_[23005]_ , \new_[23009]_ ,
    \new_[23010]_ , \new_[23014]_ , \new_[23015]_ , \new_[23016]_ ,
    \new_[23019]_ , \new_[23023]_ , \new_[23024]_ , \new_[23025]_ ,
    \new_[23029]_ , \new_[23030]_ , \new_[23034]_ , \new_[23035]_ ,
    \new_[23036]_ , \new_[23039]_ , \new_[23043]_ , \new_[23044]_ ,
    \new_[23045]_ , \new_[23049]_ , \new_[23050]_ , \new_[23054]_ ,
    \new_[23055]_ , \new_[23056]_ , \new_[23059]_ , \new_[23063]_ ,
    \new_[23064]_ , \new_[23065]_ , \new_[23069]_ , \new_[23070]_ ,
    \new_[23074]_ , \new_[23075]_ , \new_[23076]_ , \new_[23079]_ ,
    \new_[23083]_ , \new_[23084]_ , \new_[23085]_ , \new_[23089]_ ,
    \new_[23090]_ , \new_[23094]_ , \new_[23095]_ , \new_[23096]_ ,
    \new_[23099]_ , \new_[23103]_ , \new_[23104]_ , \new_[23105]_ ,
    \new_[23109]_ , \new_[23110]_ , \new_[23114]_ , \new_[23115]_ ,
    \new_[23116]_ , \new_[23119]_ , \new_[23123]_ , \new_[23124]_ ,
    \new_[23125]_ , \new_[23129]_ , \new_[23130]_ , \new_[23134]_ ,
    \new_[23135]_ , \new_[23136]_ , \new_[23139]_ , \new_[23143]_ ,
    \new_[23144]_ , \new_[23145]_ , \new_[23149]_ , \new_[23150]_ ,
    \new_[23154]_ , \new_[23155]_ , \new_[23156]_ , \new_[23159]_ ,
    \new_[23163]_ , \new_[23164]_ , \new_[23165]_ , \new_[23169]_ ,
    \new_[23170]_ , \new_[23174]_ , \new_[23175]_ , \new_[23176]_ ,
    \new_[23179]_ , \new_[23183]_ , \new_[23184]_ , \new_[23185]_ ,
    \new_[23189]_ , \new_[23190]_ , \new_[23194]_ , \new_[23195]_ ,
    \new_[23196]_ , \new_[23199]_ , \new_[23203]_ , \new_[23204]_ ,
    \new_[23205]_ , \new_[23209]_ , \new_[23210]_ , \new_[23214]_ ,
    \new_[23215]_ , \new_[23216]_ , \new_[23220]_ , \new_[23221]_ ,
    \new_[23225]_ , \new_[23226]_ , \new_[23227]_ , \new_[23231]_ ,
    \new_[23232]_ , \new_[23236]_ , \new_[23237]_ , \new_[23238]_ ,
    \new_[23242]_ , \new_[23243]_ , \new_[23247]_ , \new_[23248]_ ,
    \new_[23249]_ , \new_[23253]_ , \new_[23254]_ , \new_[23258]_ ,
    \new_[23259]_ , \new_[23260]_ , \new_[23264]_ , \new_[23265]_ ,
    \new_[23269]_ , \new_[23270]_ , \new_[23271]_ , \new_[23275]_ ,
    \new_[23276]_ , \new_[23280]_ , \new_[23281]_ , \new_[23282]_ ,
    \new_[23286]_ , \new_[23287]_ , \new_[23291]_ , \new_[23292]_ ,
    \new_[23293]_ , \new_[23297]_ , \new_[23298]_ , \new_[23302]_ ,
    \new_[23303]_ , \new_[23304]_ , \new_[23308]_ , \new_[23309]_ ,
    \new_[23313]_ , \new_[23314]_ , \new_[23315]_ , \new_[23319]_ ,
    \new_[23320]_ , \new_[23324]_ , \new_[23325]_ , \new_[23326]_ ,
    \new_[23330]_ , \new_[23331]_ , \new_[23335]_ , \new_[23336]_ ,
    \new_[23337]_ , \new_[23341]_ , \new_[23342]_ , \new_[23346]_ ,
    \new_[23347]_ , \new_[23348]_ , \new_[23352]_ , \new_[23353]_ ,
    \new_[23357]_ , \new_[23358]_ , \new_[23359]_ , \new_[23363]_ ,
    \new_[23364]_ , \new_[23368]_ , \new_[23369]_ , \new_[23370]_ ,
    \new_[23374]_ , \new_[23375]_ , \new_[23379]_ , \new_[23380]_ ,
    \new_[23381]_ , \new_[23385]_ , \new_[23386]_ , \new_[23390]_ ,
    \new_[23391]_ , \new_[23392]_ , \new_[23396]_ , \new_[23397]_ ,
    \new_[23401]_ , \new_[23402]_ , \new_[23403]_ , \new_[23407]_ ,
    \new_[23408]_ , \new_[23412]_ , \new_[23413]_ , \new_[23414]_ ,
    \new_[23418]_ , \new_[23419]_ , \new_[23423]_ , \new_[23424]_ ,
    \new_[23425]_ , \new_[23429]_ , \new_[23430]_ , \new_[23434]_ ,
    \new_[23435]_ , \new_[23436]_ , \new_[23440]_ , \new_[23441]_ ,
    \new_[23445]_ , \new_[23446]_ , \new_[23447]_ , \new_[23451]_ ,
    \new_[23452]_ , \new_[23456]_ , \new_[23457]_ , \new_[23458]_ ,
    \new_[23462]_ , \new_[23463]_ , \new_[23467]_ , \new_[23468]_ ,
    \new_[23469]_ , \new_[23473]_ , \new_[23474]_ , \new_[23478]_ ,
    \new_[23479]_ , \new_[23480]_ , \new_[23484]_ , \new_[23485]_ ,
    \new_[23489]_ , \new_[23490]_ , \new_[23491]_ , \new_[23495]_ ,
    \new_[23496]_ , \new_[23500]_ , \new_[23501]_ , \new_[23502]_ ,
    \new_[23506]_ , \new_[23507]_ , \new_[23511]_ , \new_[23512]_ ,
    \new_[23513]_ , \new_[23517]_ , \new_[23518]_ , \new_[23522]_ ,
    \new_[23523]_ , \new_[23524]_ , \new_[23528]_ , \new_[23529]_ ,
    \new_[23533]_ , \new_[23534]_ , \new_[23535]_ , \new_[23539]_ ,
    \new_[23540]_ , \new_[23544]_ , \new_[23545]_ , \new_[23546]_ ,
    \new_[23550]_ , \new_[23551]_ , \new_[23555]_ , \new_[23556]_ ,
    \new_[23557]_ , \new_[23561]_ , \new_[23562]_ , \new_[23566]_ ,
    \new_[23567]_ , \new_[23568]_ , \new_[23572]_ , \new_[23573]_ ,
    \new_[23577]_ , \new_[23578]_ , \new_[23579]_ , \new_[23583]_ ,
    \new_[23584]_ , \new_[23588]_ , \new_[23589]_ , \new_[23590]_ ,
    \new_[23594]_ , \new_[23595]_ , \new_[23599]_ , \new_[23600]_ ,
    \new_[23601]_ , \new_[23605]_ , \new_[23606]_ , \new_[23610]_ ,
    \new_[23611]_ , \new_[23612]_ , \new_[23616]_ , \new_[23617]_ ,
    \new_[23621]_ , \new_[23622]_ , \new_[23623]_ , \new_[23627]_ ,
    \new_[23628]_ , \new_[23632]_ , \new_[23633]_ , \new_[23634]_ ,
    \new_[23638]_ , \new_[23639]_ , \new_[23643]_ , \new_[23644]_ ,
    \new_[23645]_ , \new_[23649]_ , \new_[23650]_ , \new_[23654]_ ,
    \new_[23655]_ , \new_[23656]_ , \new_[23660]_ , \new_[23661]_ ,
    \new_[23665]_ , \new_[23666]_ , \new_[23667]_ , \new_[23671]_ ,
    \new_[23672]_ , \new_[23676]_ , \new_[23677]_ , \new_[23678]_ ,
    \new_[23682]_ , \new_[23683]_ , \new_[23687]_ , \new_[23688]_ ,
    \new_[23689]_ , \new_[23693]_ , \new_[23694]_ , \new_[23698]_ ,
    \new_[23699]_ , \new_[23700]_ , \new_[23704]_ , \new_[23705]_ ,
    \new_[23709]_ , \new_[23710]_ , \new_[23711]_ , \new_[23715]_ ,
    \new_[23716]_ , \new_[23720]_ , \new_[23721]_ , \new_[23722]_ ,
    \new_[23726]_ , \new_[23727]_ , \new_[23731]_ , \new_[23732]_ ,
    \new_[23733]_ , \new_[23737]_ , \new_[23738]_ , \new_[23742]_ ,
    \new_[23743]_ , \new_[23744]_ , \new_[23748]_ , \new_[23749]_ ,
    \new_[23753]_ , \new_[23754]_ , \new_[23755]_ , \new_[23759]_ ,
    \new_[23760]_ , \new_[23764]_ , \new_[23765]_ , \new_[23766]_ ,
    \new_[23770]_ , \new_[23771]_ , \new_[23775]_ , \new_[23776]_ ,
    \new_[23777]_ , \new_[23781]_ , \new_[23782]_ , \new_[23786]_ ,
    \new_[23787]_ , \new_[23788]_ , \new_[23792]_ , \new_[23793]_ ,
    \new_[23797]_ , \new_[23798]_ , \new_[23799]_ , \new_[23803]_ ,
    \new_[23804]_ , \new_[23808]_ , \new_[23809]_ , \new_[23810]_ ,
    \new_[23814]_ , \new_[23815]_ , \new_[23819]_ , \new_[23820]_ ,
    \new_[23821]_ , \new_[23825]_ , \new_[23826]_ , \new_[23830]_ ,
    \new_[23831]_ , \new_[23832]_ , \new_[23836]_ , \new_[23837]_ ,
    \new_[23841]_ , \new_[23842]_ , \new_[23843]_ , \new_[23847]_ ,
    \new_[23848]_ , \new_[23852]_ , \new_[23853]_ , \new_[23854]_ ,
    \new_[23858]_ , \new_[23859]_ , \new_[23863]_ , \new_[23864]_ ,
    \new_[23865]_ , \new_[23869]_ , \new_[23870]_ , \new_[23874]_ ,
    \new_[23875]_ , \new_[23876]_ , \new_[23880]_ , \new_[23881]_ ,
    \new_[23885]_ , \new_[23886]_ , \new_[23887]_ , \new_[23891]_ ,
    \new_[23892]_ , \new_[23896]_ , \new_[23897]_ , \new_[23898]_ ,
    \new_[23902]_ , \new_[23903]_ , \new_[23907]_ , \new_[23908]_ ,
    \new_[23909]_ , \new_[23913]_ , \new_[23914]_ , \new_[23918]_ ,
    \new_[23919]_ , \new_[23920]_ , \new_[23924]_ , \new_[23925]_ ,
    \new_[23929]_ , \new_[23930]_ , \new_[23931]_ , \new_[23935]_ ,
    \new_[23936]_ , \new_[23940]_ , \new_[23941]_ , \new_[23942]_ ,
    \new_[23946]_ , \new_[23947]_ , \new_[23951]_ , \new_[23952]_ ,
    \new_[23953]_ , \new_[23957]_ , \new_[23958]_ , \new_[23962]_ ,
    \new_[23963]_ , \new_[23964]_ , \new_[23968]_ , \new_[23969]_ ,
    \new_[23973]_ , \new_[23974]_ , \new_[23975]_ , \new_[23979]_ ,
    \new_[23980]_ , \new_[23984]_ , \new_[23985]_ , \new_[23986]_ ,
    \new_[23990]_ , \new_[23991]_ , \new_[23995]_ , \new_[23996]_ ,
    \new_[23997]_ , \new_[24001]_ , \new_[24002]_ , \new_[24006]_ ,
    \new_[24007]_ , \new_[24008]_ , \new_[24012]_ , \new_[24013]_ ,
    \new_[24017]_ , \new_[24018]_ , \new_[24019]_ , \new_[24023]_ ,
    \new_[24024]_ , \new_[24028]_ , \new_[24029]_ , \new_[24030]_ ,
    \new_[24034]_ , \new_[24035]_ , \new_[24039]_ , \new_[24040]_ ,
    \new_[24041]_ , \new_[24045]_ , \new_[24046]_ , \new_[24050]_ ,
    \new_[24051]_ , \new_[24052]_ , \new_[24056]_ , \new_[24057]_ ,
    \new_[24061]_ , \new_[24062]_ , \new_[24063]_ , \new_[24067]_ ,
    \new_[24068]_ , \new_[24072]_ , \new_[24073]_ , \new_[24074]_ ,
    \new_[24078]_ , \new_[24079]_ , \new_[24083]_ , \new_[24084]_ ,
    \new_[24085]_ , \new_[24089]_ , \new_[24090]_ , \new_[24094]_ ,
    \new_[24095]_ , \new_[24096]_ , \new_[24100]_ , \new_[24101]_ ,
    \new_[24105]_ , \new_[24106]_ , \new_[24107]_ , \new_[24111]_ ,
    \new_[24112]_ , \new_[24116]_ , \new_[24117]_ , \new_[24118]_ ,
    \new_[24122]_ , \new_[24123]_ , \new_[24127]_ , \new_[24128]_ ,
    \new_[24129]_ , \new_[24133]_ , \new_[24134]_ , \new_[24138]_ ,
    \new_[24139]_ , \new_[24140]_ , \new_[24144]_ , \new_[24145]_ ,
    \new_[24149]_ , \new_[24150]_ , \new_[24151]_ , \new_[24155]_ ,
    \new_[24156]_ , \new_[24160]_ , \new_[24161]_ , \new_[24162]_ ,
    \new_[24166]_ , \new_[24167]_ , \new_[24171]_ , \new_[24172]_ ,
    \new_[24173]_ , \new_[24177]_ , \new_[24178]_ , \new_[24182]_ ,
    \new_[24183]_ , \new_[24184]_ , \new_[24188]_ , \new_[24189]_ ,
    \new_[24193]_ , \new_[24194]_ , \new_[24195]_ , \new_[24199]_ ,
    \new_[24200]_ , \new_[24204]_ , \new_[24205]_ , \new_[24206]_ ,
    \new_[24210]_ , \new_[24211]_ , \new_[24215]_ , \new_[24216]_ ,
    \new_[24217]_ , \new_[24221]_ , \new_[24222]_ , \new_[24226]_ ,
    \new_[24227]_ , \new_[24228]_ , \new_[24232]_ , \new_[24233]_ ,
    \new_[24237]_ , \new_[24238]_ , \new_[24239]_ , \new_[24243]_ ,
    \new_[24244]_ , \new_[24248]_ , \new_[24249]_ , \new_[24250]_ ,
    \new_[24254]_ , \new_[24255]_ , \new_[24259]_ , \new_[24260]_ ,
    \new_[24261]_ , \new_[24265]_ , \new_[24266]_ , \new_[24270]_ ,
    \new_[24271]_ , \new_[24272]_ , \new_[24276]_ , \new_[24277]_ ,
    \new_[24281]_ , \new_[24282]_ , \new_[24283]_ , \new_[24287]_ ,
    \new_[24288]_ , \new_[24292]_ , \new_[24293]_ , \new_[24294]_ ,
    \new_[24298]_ , \new_[24299]_ , \new_[24303]_ , \new_[24304]_ ,
    \new_[24305]_ , \new_[24309]_ , \new_[24310]_ , \new_[24314]_ ,
    \new_[24315]_ , \new_[24316]_ , \new_[24320]_ , \new_[24321]_ ,
    \new_[24325]_ , \new_[24326]_ , \new_[24327]_ , \new_[24331]_ ,
    \new_[24332]_ , \new_[24336]_ , \new_[24337]_ , \new_[24338]_ ,
    \new_[24342]_ , \new_[24343]_ , \new_[24347]_ , \new_[24348]_ ,
    \new_[24349]_ , \new_[24353]_ , \new_[24354]_ , \new_[24358]_ ,
    \new_[24359]_ , \new_[24360]_ , \new_[24364]_ , \new_[24365]_ ,
    \new_[24369]_ , \new_[24370]_ , \new_[24371]_ , \new_[24375]_ ,
    \new_[24376]_ , \new_[24380]_ , \new_[24381]_ , \new_[24382]_ ,
    \new_[24386]_ , \new_[24387]_ , \new_[24391]_ , \new_[24392]_ ,
    \new_[24393]_ , \new_[24397]_ , \new_[24398]_ , \new_[24402]_ ,
    \new_[24403]_ , \new_[24404]_ , \new_[24408]_ , \new_[24409]_ ,
    \new_[24413]_ , \new_[24414]_ , \new_[24415]_ , \new_[24419]_ ,
    \new_[24420]_ , \new_[24424]_ , \new_[24425]_ , \new_[24426]_ ,
    \new_[24430]_ , \new_[24431]_ , \new_[24435]_ , \new_[24436]_ ,
    \new_[24437]_ , \new_[24441]_ , \new_[24442]_ , \new_[24446]_ ,
    \new_[24447]_ , \new_[24448]_ , \new_[24452]_ , \new_[24453]_ ,
    \new_[24457]_ , \new_[24458]_ , \new_[24459]_ , \new_[24463]_ ,
    \new_[24464]_ , \new_[24468]_ , \new_[24469]_ , \new_[24470]_ ,
    \new_[24474]_ , \new_[24475]_ , \new_[24479]_ , \new_[24480]_ ,
    \new_[24481]_ , \new_[24485]_ , \new_[24486]_ , \new_[24490]_ ,
    \new_[24491]_ , \new_[24492]_ , \new_[24496]_ , \new_[24497]_ ,
    \new_[24501]_ , \new_[24502]_ , \new_[24503]_ , \new_[24507]_ ,
    \new_[24508]_ , \new_[24512]_ , \new_[24513]_ , \new_[24514]_ ,
    \new_[24518]_ , \new_[24519]_ , \new_[24523]_ , \new_[24524]_ ,
    \new_[24525]_ , \new_[24529]_ , \new_[24530]_ , \new_[24534]_ ,
    \new_[24535]_ , \new_[24536]_ , \new_[24540]_ , \new_[24541]_ ,
    \new_[24545]_ , \new_[24546]_ , \new_[24547]_ , \new_[24551]_ ,
    \new_[24552]_ , \new_[24556]_ , \new_[24557]_ , \new_[24558]_ ,
    \new_[24562]_ , \new_[24563]_ , \new_[24567]_ , \new_[24568]_ ,
    \new_[24569]_ , \new_[24573]_ , \new_[24574]_ , \new_[24578]_ ,
    \new_[24579]_ , \new_[24580]_ , \new_[24584]_ , \new_[24585]_ ,
    \new_[24589]_ , \new_[24590]_ , \new_[24591]_ , \new_[24595]_ ,
    \new_[24596]_ , \new_[24600]_ , \new_[24601]_ , \new_[24602]_ ,
    \new_[24606]_ , \new_[24607]_ , \new_[24611]_ , \new_[24612]_ ,
    \new_[24613]_ , \new_[24617]_ , \new_[24618]_ , \new_[24622]_ ,
    \new_[24623]_ , \new_[24624]_ , \new_[24628]_ , \new_[24629]_ ,
    \new_[24633]_ , \new_[24634]_ , \new_[24635]_ , \new_[24639]_ ,
    \new_[24640]_ , \new_[24644]_ , \new_[24645]_ , \new_[24646]_ ,
    \new_[24650]_ , \new_[24651]_ , \new_[24655]_ , \new_[24656]_ ,
    \new_[24657]_ , \new_[24661]_ , \new_[24662]_ , \new_[24666]_ ,
    \new_[24667]_ , \new_[24668]_ , \new_[24672]_ , \new_[24673]_ ,
    \new_[24677]_ , \new_[24678]_ , \new_[24679]_ , \new_[24683]_ ,
    \new_[24684]_ , \new_[24688]_ , \new_[24689]_ , \new_[24690]_ ,
    \new_[24694]_ , \new_[24695]_ , \new_[24699]_ , \new_[24700]_ ,
    \new_[24701]_ , \new_[24705]_ , \new_[24706]_ , \new_[24710]_ ,
    \new_[24711]_ , \new_[24712]_ , \new_[24716]_ , \new_[24717]_ ,
    \new_[24721]_ , \new_[24722]_ , \new_[24723]_ , \new_[24727]_ ,
    \new_[24728]_ , \new_[24732]_ , \new_[24733]_ , \new_[24734]_ ,
    \new_[24738]_ , \new_[24739]_ , \new_[24743]_ , \new_[24744]_ ,
    \new_[24745]_ , \new_[24749]_ , \new_[24750]_ , \new_[24754]_ ,
    \new_[24755]_ , \new_[24756]_ , \new_[24760]_ , \new_[24761]_ ,
    \new_[24765]_ , \new_[24766]_ , \new_[24767]_ , \new_[24771]_ ,
    \new_[24772]_ , \new_[24776]_ , \new_[24777]_ , \new_[24778]_ ,
    \new_[24782]_ , \new_[24783]_ , \new_[24787]_ , \new_[24788]_ ,
    \new_[24789]_ , \new_[24793]_ , \new_[24794]_ , \new_[24798]_ ,
    \new_[24799]_ , \new_[24800]_ , \new_[24804]_ , \new_[24805]_ ,
    \new_[24809]_ , \new_[24810]_ , \new_[24811]_ , \new_[24815]_ ,
    \new_[24816]_ , \new_[24820]_ , \new_[24821]_ , \new_[24822]_ ,
    \new_[24826]_ , \new_[24827]_ , \new_[24831]_ , \new_[24832]_ ,
    \new_[24833]_ , \new_[24837]_ , \new_[24838]_ , \new_[24842]_ ,
    \new_[24843]_ , \new_[24844]_ , \new_[24848]_ , \new_[24849]_ ,
    \new_[24853]_ , \new_[24854]_ , \new_[24855]_ , \new_[24859]_ ,
    \new_[24860]_ , \new_[24864]_ , \new_[24865]_ , \new_[24866]_ ,
    \new_[24870]_ , \new_[24871]_ , \new_[24875]_ , \new_[24876]_ ,
    \new_[24877]_ , \new_[24881]_ , \new_[24882]_ , \new_[24886]_ ,
    \new_[24887]_ , \new_[24888]_ , \new_[24892]_ , \new_[24893]_ ,
    \new_[24897]_ , \new_[24898]_ , \new_[24899]_ , \new_[24903]_ ,
    \new_[24904]_ , \new_[24908]_ , \new_[24909]_ , \new_[24910]_ ,
    \new_[24914]_ , \new_[24915]_ , \new_[24919]_ , \new_[24920]_ ,
    \new_[24921]_ , \new_[24925]_ , \new_[24926]_ , \new_[24930]_ ,
    \new_[24931]_ , \new_[24932]_ , \new_[24936]_ , \new_[24937]_ ,
    \new_[24941]_ , \new_[24942]_ , \new_[24943]_ , \new_[24947]_ ,
    \new_[24948]_ , \new_[24952]_ , \new_[24953]_ , \new_[24954]_ ,
    \new_[24958]_ , \new_[24959]_ , \new_[24963]_ , \new_[24964]_ ,
    \new_[24965]_ , \new_[24969]_ , \new_[24970]_ , \new_[24974]_ ,
    \new_[24975]_ , \new_[24976]_ , \new_[24980]_ , \new_[24981]_ ,
    \new_[24985]_ , \new_[24986]_ , \new_[24987]_ , \new_[24991]_ ,
    \new_[24992]_ , \new_[24996]_ , \new_[24997]_ , \new_[24998]_ ,
    \new_[25002]_ , \new_[25003]_ , \new_[25007]_ , \new_[25008]_ ,
    \new_[25009]_ , \new_[25013]_ , \new_[25014]_ , \new_[25018]_ ,
    \new_[25019]_ , \new_[25020]_ , \new_[25024]_ , \new_[25025]_ ,
    \new_[25029]_ , \new_[25030]_ , \new_[25031]_ , \new_[25035]_ ,
    \new_[25036]_ , \new_[25040]_ , \new_[25041]_ , \new_[25042]_ ,
    \new_[25046]_ , \new_[25047]_ , \new_[25051]_ , \new_[25052]_ ,
    \new_[25053]_ , \new_[25057]_ , \new_[25058]_ , \new_[25062]_ ,
    \new_[25063]_ , \new_[25064]_ , \new_[25068]_ , \new_[25069]_ ,
    \new_[25073]_ , \new_[25074]_ , \new_[25075]_ , \new_[25079]_ ,
    \new_[25080]_ , \new_[25084]_ , \new_[25085]_ , \new_[25086]_ ,
    \new_[25090]_ , \new_[25091]_ , \new_[25095]_ , \new_[25096]_ ,
    \new_[25097]_ , \new_[25101]_ , \new_[25102]_ , \new_[25106]_ ,
    \new_[25107]_ , \new_[25108]_ , \new_[25112]_ , \new_[25113]_ ,
    \new_[25117]_ , \new_[25118]_ , \new_[25119]_ , \new_[25123]_ ,
    \new_[25124]_ , \new_[25128]_ , \new_[25129]_ , \new_[25130]_ ,
    \new_[25134]_ , \new_[25135]_ , \new_[25139]_ , \new_[25140]_ ,
    \new_[25141]_ , \new_[25145]_ , \new_[25146]_ , \new_[25150]_ ,
    \new_[25151]_ , \new_[25152]_ , \new_[25156]_ , \new_[25157]_ ,
    \new_[25161]_ , \new_[25162]_ , \new_[25163]_ , \new_[25167]_ ,
    \new_[25168]_ , \new_[25172]_ , \new_[25173]_ , \new_[25174]_ ,
    \new_[25178]_ , \new_[25179]_ , \new_[25183]_ , \new_[25184]_ ,
    \new_[25185]_ , \new_[25189]_ , \new_[25190]_ , \new_[25194]_ ,
    \new_[25195]_ , \new_[25196]_ , \new_[25200]_ , \new_[25201]_ ,
    \new_[25205]_ , \new_[25206]_ , \new_[25207]_ , \new_[25211]_ ,
    \new_[25212]_ , \new_[25216]_ , \new_[25217]_ , \new_[25218]_ ,
    \new_[25222]_ , \new_[25223]_ , \new_[25227]_ , \new_[25228]_ ,
    \new_[25229]_ , \new_[25233]_ , \new_[25234]_ , \new_[25238]_ ,
    \new_[25239]_ , \new_[25240]_ , \new_[25244]_ , \new_[25245]_ ,
    \new_[25249]_ , \new_[25250]_ , \new_[25251]_ , \new_[25255]_ ,
    \new_[25256]_ , \new_[25260]_ , \new_[25261]_ , \new_[25262]_ ,
    \new_[25266]_ , \new_[25267]_ , \new_[25271]_ , \new_[25272]_ ,
    \new_[25273]_ , \new_[25277]_ , \new_[25278]_ , \new_[25282]_ ,
    \new_[25283]_ , \new_[25284]_ , \new_[25288]_ , \new_[25289]_ ,
    \new_[25293]_ , \new_[25294]_ , \new_[25295]_ , \new_[25299]_ ,
    \new_[25300]_ , \new_[25304]_ , \new_[25305]_ , \new_[25306]_ ,
    \new_[25310]_ , \new_[25311]_ , \new_[25315]_ , \new_[25316]_ ,
    \new_[25317]_ , \new_[25321]_ , \new_[25322]_ , \new_[25326]_ ,
    \new_[25327]_ , \new_[25328]_ , \new_[25332]_ , \new_[25333]_ ,
    \new_[25337]_ , \new_[25338]_ , \new_[25339]_ , \new_[25343]_ ,
    \new_[25344]_ , \new_[25348]_ , \new_[25349]_ , \new_[25350]_ ,
    \new_[25354]_ , \new_[25355]_ , \new_[25359]_ , \new_[25360]_ ,
    \new_[25361]_ , \new_[25365]_ , \new_[25366]_ , \new_[25370]_ ,
    \new_[25371]_ , \new_[25372]_ , \new_[25376]_ , \new_[25377]_ ,
    \new_[25381]_ , \new_[25382]_ , \new_[25383]_ , \new_[25387]_ ,
    \new_[25388]_ , \new_[25392]_ , \new_[25393]_ , \new_[25394]_ ,
    \new_[25398]_ , \new_[25399]_ , \new_[25403]_ , \new_[25404]_ ,
    \new_[25405]_ , \new_[25409]_ , \new_[25410]_ , \new_[25414]_ ,
    \new_[25415]_ , \new_[25416]_ , \new_[25420]_ , \new_[25421]_ ,
    \new_[25425]_ , \new_[25426]_ , \new_[25427]_ , \new_[25431]_ ,
    \new_[25432]_ , \new_[25436]_ , \new_[25437]_ , \new_[25438]_ ,
    \new_[25442]_ , \new_[25443]_ , \new_[25447]_ , \new_[25448]_ ,
    \new_[25449]_ , \new_[25453]_ , \new_[25454]_ , \new_[25458]_ ,
    \new_[25459]_ , \new_[25460]_ , \new_[25464]_ , \new_[25465]_ ,
    \new_[25469]_ , \new_[25470]_ , \new_[25471]_ , \new_[25475]_ ,
    \new_[25476]_ , \new_[25480]_ , \new_[25481]_ , \new_[25482]_ ,
    \new_[25486]_ , \new_[25487]_ , \new_[25491]_ , \new_[25492]_ ,
    \new_[25493]_ , \new_[25497]_ , \new_[25498]_ , \new_[25502]_ ,
    \new_[25503]_ , \new_[25504]_ , \new_[25508]_ , \new_[25509]_ ,
    \new_[25513]_ , \new_[25514]_ , \new_[25515]_ , \new_[25519]_ ,
    \new_[25520]_ , \new_[25524]_ , \new_[25525]_ , \new_[25526]_ ,
    \new_[25530]_ , \new_[25531]_ , \new_[25535]_ , \new_[25536]_ ,
    \new_[25537]_ , \new_[25541]_ , \new_[25542]_ , \new_[25546]_ ,
    \new_[25547]_ , \new_[25548]_ , \new_[25552]_ , \new_[25553]_ ,
    \new_[25557]_ , \new_[25558]_ , \new_[25559]_ , \new_[25563]_ ,
    \new_[25564]_ , \new_[25568]_ , \new_[25569]_ , \new_[25570]_ ,
    \new_[25574]_ , \new_[25575]_ , \new_[25579]_ , \new_[25580]_ ,
    \new_[25581]_ , \new_[25585]_ , \new_[25586]_ , \new_[25590]_ ,
    \new_[25591]_ , \new_[25592]_ , \new_[25596]_ , \new_[25597]_ ,
    \new_[25601]_ , \new_[25602]_ , \new_[25603]_ , \new_[25607]_ ,
    \new_[25608]_ , \new_[25612]_ , \new_[25613]_ , \new_[25614]_ ,
    \new_[25618]_ , \new_[25619]_ , \new_[25623]_ , \new_[25624]_ ,
    \new_[25625]_ , \new_[25629]_ , \new_[25630]_ , \new_[25634]_ ,
    \new_[25635]_ , \new_[25636]_ , \new_[25640]_ , \new_[25641]_ ,
    \new_[25645]_ , \new_[25646]_ , \new_[25647]_ , \new_[25651]_ ,
    \new_[25652]_ , \new_[25656]_ , \new_[25657]_ , \new_[25658]_ ,
    \new_[25662]_ , \new_[25663]_ , \new_[25667]_ , \new_[25668]_ ,
    \new_[25669]_ , \new_[25673]_ , \new_[25674]_ , \new_[25678]_ ,
    \new_[25679]_ , \new_[25680]_ , \new_[25684]_ , \new_[25685]_ ,
    \new_[25689]_ , \new_[25690]_ , \new_[25691]_ , \new_[25695]_ ,
    \new_[25696]_ , \new_[25700]_ , \new_[25701]_ , \new_[25702]_ ,
    \new_[25706]_ , \new_[25707]_ , \new_[25711]_ , \new_[25712]_ ,
    \new_[25713]_ , \new_[25717]_ , \new_[25718]_ , \new_[25722]_ ,
    \new_[25723]_ , \new_[25724]_ , \new_[25728]_ , \new_[25729]_ ,
    \new_[25733]_ , \new_[25734]_ , \new_[25735]_ , \new_[25739]_ ,
    \new_[25740]_ , \new_[25744]_ , \new_[25745]_ , \new_[25746]_ ,
    \new_[25750]_ , \new_[25751]_ , \new_[25755]_ , \new_[25756]_ ,
    \new_[25757]_ , \new_[25761]_ , \new_[25762]_ , \new_[25766]_ ,
    \new_[25767]_ , \new_[25768]_ , \new_[25772]_ , \new_[25773]_ ,
    \new_[25777]_ , \new_[25778]_ , \new_[25779]_ , \new_[25783]_ ,
    \new_[25784]_ , \new_[25788]_ , \new_[25789]_ , \new_[25790]_ ,
    \new_[25794]_ , \new_[25795]_ , \new_[25799]_ , \new_[25800]_ ,
    \new_[25801]_ , \new_[25805]_ , \new_[25806]_ , \new_[25810]_ ,
    \new_[25811]_ , \new_[25812]_ , \new_[25816]_ , \new_[25817]_ ,
    \new_[25821]_ , \new_[25822]_ , \new_[25823]_ , \new_[25827]_ ,
    \new_[25828]_ , \new_[25832]_ , \new_[25833]_ , \new_[25834]_ ,
    \new_[25838]_ , \new_[25839]_ , \new_[25843]_ , \new_[25844]_ ,
    \new_[25845]_ , \new_[25849]_ , \new_[25850]_ , \new_[25854]_ ,
    \new_[25855]_ , \new_[25856]_ , \new_[25860]_ , \new_[25861]_ ,
    \new_[25865]_ , \new_[25866]_ , \new_[25867]_ , \new_[25871]_ ,
    \new_[25872]_ , \new_[25876]_ , \new_[25877]_ , \new_[25878]_ ,
    \new_[25882]_ , \new_[25883]_ , \new_[25887]_ , \new_[25888]_ ,
    \new_[25889]_ , \new_[25893]_ , \new_[25894]_ , \new_[25898]_ ,
    \new_[25899]_ , \new_[25900]_ , \new_[25904]_ , \new_[25905]_ ,
    \new_[25909]_ , \new_[25910]_ , \new_[25911]_ , \new_[25915]_ ,
    \new_[25916]_ , \new_[25920]_ , \new_[25921]_ , \new_[25922]_ ,
    \new_[25926]_ , \new_[25927]_ , \new_[25931]_ , \new_[25932]_ ,
    \new_[25933]_ , \new_[25937]_ , \new_[25938]_ , \new_[25942]_ ,
    \new_[25943]_ , \new_[25944]_ , \new_[25948]_ , \new_[25949]_ ,
    \new_[25953]_ , \new_[25954]_ , \new_[25955]_ , \new_[25959]_ ,
    \new_[25960]_ , \new_[25964]_ , \new_[25965]_ , \new_[25966]_ ,
    \new_[25970]_ , \new_[25971]_ , \new_[25975]_ , \new_[25976]_ ,
    \new_[25977]_ , \new_[25981]_ , \new_[25982]_ , \new_[25986]_ ,
    \new_[25987]_ , \new_[25988]_ , \new_[25992]_ , \new_[25993]_ ,
    \new_[25997]_ , \new_[25998]_ , \new_[25999]_ , \new_[26003]_ ,
    \new_[26004]_ , \new_[26008]_ , \new_[26009]_ , \new_[26010]_ ,
    \new_[26014]_ , \new_[26015]_ , \new_[26019]_ , \new_[26020]_ ,
    \new_[26021]_ , \new_[26025]_ , \new_[26026]_ , \new_[26030]_ ,
    \new_[26031]_ , \new_[26032]_ , \new_[26036]_ , \new_[26037]_ ,
    \new_[26041]_ , \new_[26042]_ , \new_[26043]_ , \new_[26047]_ ,
    \new_[26048]_ , \new_[26052]_ , \new_[26053]_ , \new_[26054]_ ,
    \new_[26058]_ , \new_[26059]_ , \new_[26063]_ , \new_[26064]_ ,
    \new_[26065]_ , \new_[26069]_ , \new_[26070]_ , \new_[26074]_ ,
    \new_[26075]_ , \new_[26076]_ , \new_[26080]_ , \new_[26081]_ ,
    \new_[26085]_ , \new_[26086]_ , \new_[26087]_ , \new_[26091]_ ,
    \new_[26092]_ , \new_[26096]_ , \new_[26097]_ , \new_[26098]_ ,
    \new_[26102]_ , \new_[26103]_ , \new_[26107]_ , \new_[26108]_ ,
    \new_[26109]_ , \new_[26113]_ , \new_[26114]_ , \new_[26118]_ ,
    \new_[26119]_ , \new_[26120]_ , \new_[26124]_ , \new_[26125]_ ,
    \new_[26129]_ , \new_[26130]_ , \new_[26131]_ , \new_[26135]_ ,
    \new_[26136]_ , \new_[26140]_ , \new_[26141]_ , \new_[26142]_ ,
    \new_[26146]_ , \new_[26147]_ , \new_[26151]_ , \new_[26152]_ ,
    \new_[26153]_ , \new_[26157]_ , \new_[26158]_ , \new_[26162]_ ,
    \new_[26163]_ , \new_[26164]_ , \new_[26168]_ , \new_[26169]_ ,
    \new_[26173]_ , \new_[26174]_ , \new_[26175]_ , \new_[26179]_ ,
    \new_[26180]_ , \new_[26184]_ , \new_[26185]_ , \new_[26186]_ ,
    \new_[26190]_ , \new_[26191]_ , \new_[26195]_ , \new_[26196]_ ,
    \new_[26197]_ , \new_[26201]_ , \new_[26202]_ , \new_[26206]_ ,
    \new_[26207]_ , \new_[26208]_ , \new_[26212]_ , \new_[26213]_ ,
    \new_[26217]_ , \new_[26218]_ , \new_[26219]_ , \new_[26223]_ ,
    \new_[26224]_ , \new_[26228]_ , \new_[26229]_ , \new_[26230]_ ,
    \new_[26234]_ , \new_[26235]_ , \new_[26239]_ , \new_[26240]_ ,
    \new_[26241]_ , \new_[26245]_ , \new_[26246]_ , \new_[26250]_ ,
    \new_[26251]_ , \new_[26252]_ , \new_[26256]_ , \new_[26257]_ ,
    \new_[26261]_ , \new_[26262]_ , \new_[26263]_ , \new_[26267]_ ,
    \new_[26268]_ , \new_[26272]_ , \new_[26273]_ , \new_[26274]_ ,
    \new_[26278]_ , \new_[26279]_ , \new_[26283]_ , \new_[26284]_ ,
    \new_[26285]_ , \new_[26289]_ , \new_[26290]_ , \new_[26294]_ ,
    \new_[26295]_ , \new_[26296]_ , \new_[26300]_ , \new_[26301]_ ,
    \new_[26305]_ , \new_[26306]_ , \new_[26307]_ , \new_[26311]_ ,
    \new_[26312]_ , \new_[26316]_ , \new_[26317]_ , \new_[26318]_ ,
    \new_[26322]_ , \new_[26323]_ , \new_[26327]_ , \new_[26328]_ ,
    \new_[26329]_ , \new_[26333]_ , \new_[26334]_ , \new_[26338]_ ,
    \new_[26339]_ , \new_[26340]_ , \new_[26344]_ , \new_[26345]_ ,
    \new_[26349]_ , \new_[26350]_ , \new_[26351]_ , \new_[26355]_ ,
    \new_[26356]_ , \new_[26360]_ , \new_[26361]_ , \new_[26362]_ ,
    \new_[26366]_ , \new_[26367]_ , \new_[26371]_ , \new_[26372]_ ,
    \new_[26373]_ , \new_[26377]_ , \new_[26378]_ , \new_[26382]_ ,
    \new_[26383]_ , \new_[26384]_ , \new_[26388]_ , \new_[26389]_ ,
    \new_[26393]_ , \new_[26394]_ , \new_[26395]_ , \new_[26399]_ ,
    \new_[26400]_ , \new_[26404]_ , \new_[26405]_ , \new_[26406]_ ,
    \new_[26410]_ , \new_[26411]_ , \new_[26415]_ , \new_[26416]_ ,
    \new_[26417]_ , \new_[26421]_ , \new_[26422]_ , \new_[26426]_ ,
    \new_[26427]_ , \new_[26428]_ , \new_[26432]_ , \new_[26433]_ ,
    \new_[26437]_ , \new_[26438]_ , \new_[26439]_ , \new_[26443]_ ,
    \new_[26444]_ , \new_[26448]_ , \new_[26449]_ , \new_[26450]_ ,
    \new_[26454]_ , \new_[26455]_ , \new_[26459]_ , \new_[26460]_ ,
    \new_[26461]_ , \new_[26465]_ , \new_[26466]_ , \new_[26470]_ ,
    \new_[26471]_ , \new_[26472]_ , \new_[26476]_ , \new_[26477]_ ,
    \new_[26481]_ , \new_[26482]_ , \new_[26483]_ , \new_[26487]_ ,
    \new_[26488]_ , \new_[26492]_ , \new_[26493]_ , \new_[26494]_ ,
    \new_[26498]_ , \new_[26499]_ , \new_[26503]_ , \new_[26504]_ ,
    \new_[26505]_ , \new_[26509]_ , \new_[26510]_ , \new_[26514]_ ,
    \new_[26515]_ , \new_[26516]_ , \new_[26520]_ , \new_[26521]_ ,
    \new_[26525]_ , \new_[26526]_ , \new_[26527]_ , \new_[26531]_ ,
    \new_[26532]_ , \new_[26536]_ , \new_[26537]_ , \new_[26538]_ ,
    \new_[26542]_ , \new_[26543]_ , \new_[26547]_ , \new_[26548]_ ,
    \new_[26549]_ , \new_[26553]_ , \new_[26554]_ , \new_[26558]_ ,
    \new_[26559]_ , \new_[26560]_ , \new_[26564]_ , \new_[26565]_ ,
    \new_[26569]_ , \new_[26570]_ , \new_[26571]_ , \new_[26575]_ ,
    \new_[26576]_ , \new_[26580]_ , \new_[26581]_ , \new_[26582]_ ,
    \new_[26586]_ , \new_[26587]_ , \new_[26591]_ , \new_[26592]_ ,
    \new_[26593]_ , \new_[26597]_ , \new_[26598]_ , \new_[26602]_ ,
    \new_[26603]_ , \new_[26604]_ , \new_[26608]_ , \new_[26609]_ ,
    \new_[26613]_ , \new_[26614]_ , \new_[26615]_ , \new_[26619]_ ,
    \new_[26620]_ , \new_[26624]_ , \new_[26625]_ , \new_[26626]_ ,
    \new_[26630]_ , \new_[26631]_ , \new_[26635]_ , \new_[26636]_ ,
    \new_[26637]_ , \new_[26641]_ , \new_[26642]_ , \new_[26646]_ ,
    \new_[26647]_ , \new_[26648]_ , \new_[26652]_ , \new_[26653]_ ,
    \new_[26657]_ , \new_[26658]_ , \new_[26659]_ , \new_[26663]_ ,
    \new_[26664]_ , \new_[26668]_ , \new_[26669]_ , \new_[26670]_ ,
    \new_[26674]_ , \new_[26675]_ , \new_[26679]_ , \new_[26680]_ ,
    \new_[26681]_ , \new_[26685]_ , \new_[26686]_ , \new_[26690]_ ,
    \new_[26691]_ , \new_[26692]_ , \new_[26696]_ , \new_[26697]_ ,
    \new_[26701]_ , \new_[26702]_ , \new_[26703]_ , \new_[26707]_ ,
    \new_[26708]_ , \new_[26712]_ , \new_[26713]_ , \new_[26714]_ ,
    \new_[26718]_ , \new_[26719]_ , \new_[26723]_ , \new_[26724]_ ,
    \new_[26725]_ , \new_[26729]_ , \new_[26730]_ , \new_[26734]_ ,
    \new_[26735]_ , \new_[26736]_ , \new_[26740]_ , \new_[26741]_ ,
    \new_[26745]_ , \new_[26746]_ , \new_[26747]_ , \new_[26751]_ ,
    \new_[26752]_ , \new_[26756]_ , \new_[26757]_ , \new_[26758]_ ,
    \new_[26762]_ , \new_[26763]_ , \new_[26767]_ , \new_[26768]_ ,
    \new_[26769]_ , \new_[26773]_ , \new_[26774]_ , \new_[26778]_ ,
    \new_[26779]_ , \new_[26780]_ , \new_[26784]_ , \new_[26785]_ ,
    \new_[26789]_ , \new_[26790]_ , \new_[26791]_ , \new_[26795]_ ,
    \new_[26796]_ , \new_[26800]_ , \new_[26801]_ , \new_[26802]_ ,
    \new_[26806]_ , \new_[26807]_ , \new_[26811]_ , \new_[26812]_ ,
    \new_[26813]_ , \new_[26817]_ , \new_[26818]_ , \new_[26822]_ ,
    \new_[26823]_ , \new_[26824]_ , \new_[26828]_ , \new_[26829]_ ,
    \new_[26833]_ , \new_[26834]_ , \new_[26835]_ , \new_[26839]_ ,
    \new_[26840]_ , \new_[26844]_ , \new_[26845]_ , \new_[26846]_ ,
    \new_[26850]_ , \new_[26851]_ , \new_[26855]_ , \new_[26856]_ ,
    \new_[26857]_ , \new_[26861]_ , \new_[26862]_ , \new_[26866]_ ,
    \new_[26867]_ , \new_[26868]_ , \new_[26872]_ , \new_[26873]_ ,
    \new_[26877]_ , \new_[26878]_ , \new_[26879]_ , \new_[26883]_ ,
    \new_[26884]_ , \new_[26888]_ , \new_[26889]_ , \new_[26890]_ ,
    \new_[26894]_ , \new_[26895]_ , \new_[26899]_ , \new_[26900]_ ,
    \new_[26901]_ , \new_[26905]_ , \new_[26906]_ , \new_[26910]_ ,
    \new_[26911]_ , \new_[26912]_ , \new_[26916]_ , \new_[26917]_ ,
    \new_[26921]_ , \new_[26922]_ , \new_[26923]_ , \new_[26927]_ ,
    \new_[26928]_ , \new_[26932]_ , \new_[26933]_ , \new_[26934]_ ,
    \new_[26938]_ , \new_[26939]_ , \new_[26943]_ , \new_[26944]_ ,
    \new_[26945]_ , \new_[26949]_ , \new_[26950]_ , \new_[26954]_ ,
    \new_[26955]_ , \new_[26956]_ , \new_[26960]_ , \new_[26961]_ ,
    \new_[26965]_ , \new_[26966]_ , \new_[26967]_ , \new_[26971]_ ,
    \new_[26972]_ , \new_[26976]_ , \new_[26977]_ , \new_[26978]_ ,
    \new_[26982]_ , \new_[26983]_ , \new_[26987]_ , \new_[26988]_ ,
    \new_[26989]_ , \new_[26993]_ , \new_[26994]_ , \new_[26998]_ ,
    \new_[26999]_ , \new_[27000]_ , \new_[27004]_ , \new_[27005]_ ,
    \new_[27009]_ , \new_[27010]_ , \new_[27011]_ , \new_[27015]_ ,
    \new_[27016]_ , \new_[27020]_ , \new_[27021]_ , \new_[27022]_ ,
    \new_[27026]_ , \new_[27027]_ , \new_[27031]_ , \new_[27032]_ ,
    \new_[27033]_ , \new_[27037]_ , \new_[27038]_ , \new_[27042]_ ,
    \new_[27043]_ , \new_[27044]_ , \new_[27048]_ , \new_[27049]_ ,
    \new_[27053]_ , \new_[27054]_ , \new_[27055]_ , \new_[27059]_ ,
    \new_[27060]_ , \new_[27064]_ , \new_[27065]_ , \new_[27066]_ ,
    \new_[27070]_ , \new_[27071]_ , \new_[27075]_ , \new_[27076]_ ,
    \new_[27077]_ , \new_[27081]_ , \new_[27082]_ , \new_[27086]_ ,
    \new_[27087]_ , \new_[27088]_ , \new_[27092]_ , \new_[27093]_ ,
    \new_[27097]_ , \new_[27098]_ , \new_[27099]_ , \new_[27103]_ ,
    \new_[27104]_ , \new_[27108]_ , \new_[27109]_ , \new_[27110]_ ,
    \new_[27114]_ , \new_[27115]_ , \new_[27119]_ , \new_[27120]_ ,
    \new_[27121]_ , \new_[27125]_ , \new_[27126]_ , \new_[27130]_ ,
    \new_[27131]_ , \new_[27132]_ , \new_[27136]_ , \new_[27137]_ ,
    \new_[27141]_ , \new_[27142]_ , \new_[27143]_ , \new_[27147]_ ,
    \new_[27148]_ , \new_[27152]_ , \new_[27153]_ , \new_[27154]_ ,
    \new_[27158]_ , \new_[27159]_ , \new_[27163]_ , \new_[27164]_ ,
    \new_[27165]_ , \new_[27169]_ , \new_[27170]_ , \new_[27174]_ ,
    \new_[27175]_ , \new_[27176]_ , \new_[27180]_ , \new_[27181]_ ,
    \new_[27185]_ , \new_[27186]_ , \new_[27187]_ , \new_[27191]_ ,
    \new_[27192]_ , \new_[27196]_ , \new_[27197]_ , \new_[27198]_ ,
    \new_[27202]_ , \new_[27203]_ , \new_[27207]_ , \new_[27208]_ ,
    \new_[27209]_ , \new_[27213]_ , \new_[27214]_ , \new_[27218]_ ,
    \new_[27219]_ , \new_[27220]_ , \new_[27224]_ , \new_[27225]_ ,
    \new_[27229]_ , \new_[27230]_ , \new_[27231]_ , \new_[27235]_ ,
    \new_[27236]_ , \new_[27240]_ , \new_[27241]_ , \new_[27242]_ ,
    \new_[27246]_ , \new_[27247]_ , \new_[27251]_ , \new_[27252]_ ,
    \new_[27253]_ , \new_[27257]_ , \new_[27258]_ , \new_[27262]_ ,
    \new_[27263]_ , \new_[27264]_ , \new_[27268]_ , \new_[27269]_ ,
    \new_[27273]_ , \new_[27274]_ , \new_[27275]_ , \new_[27279]_ ,
    \new_[27280]_ , \new_[27284]_ , \new_[27285]_ , \new_[27286]_ ,
    \new_[27290]_ , \new_[27291]_ , \new_[27295]_ , \new_[27296]_ ,
    \new_[27297]_ , \new_[27301]_ , \new_[27302]_ , \new_[27306]_ ,
    \new_[27307]_ , \new_[27308]_ , \new_[27312]_ , \new_[27313]_ ,
    \new_[27317]_ , \new_[27318]_ , \new_[27319]_ , \new_[27323]_ ,
    \new_[27324]_ , \new_[27328]_ , \new_[27329]_ , \new_[27330]_ ,
    \new_[27334]_ , \new_[27335]_ , \new_[27339]_ , \new_[27340]_ ,
    \new_[27341]_ , \new_[27345]_ , \new_[27346]_ , \new_[27350]_ ,
    \new_[27351]_ , \new_[27352]_ , \new_[27356]_ , \new_[27357]_ ,
    \new_[27361]_ , \new_[27362]_ , \new_[27363]_ , \new_[27367]_ ,
    \new_[27368]_ , \new_[27372]_ , \new_[27373]_ , \new_[27374]_ ,
    \new_[27378]_ , \new_[27379]_ , \new_[27383]_ , \new_[27384]_ ,
    \new_[27385]_ , \new_[27389]_ , \new_[27390]_ , \new_[27394]_ ,
    \new_[27395]_ , \new_[27396]_ , \new_[27400]_ , \new_[27401]_ ,
    \new_[27405]_ , \new_[27406]_ , \new_[27407]_ , \new_[27411]_ ,
    \new_[27412]_ , \new_[27416]_ , \new_[27417]_ , \new_[27418]_ ,
    \new_[27422]_ , \new_[27423]_ , \new_[27427]_ , \new_[27428]_ ,
    \new_[27429]_ , \new_[27433]_ , \new_[27434]_ , \new_[27438]_ ,
    \new_[27439]_ , \new_[27440]_ , \new_[27444]_ , \new_[27445]_ ,
    \new_[27449]_ , \new_[27450]_ , \new_[27451]_ , \new_[27455]_ ,
    \new_[27456]_ , \new_[27460]_ , \new_[27461]_ , \new_[27462]_ ,
    \new_[27466]_ , \new_[27467]_ , \new_[27471]_ , \new_[27472]_ ,
    \new_[27473]_ , \new_[27477]_ , \new_[27478]_ , \new_[27482]_ ,
    \new_[27483]_ , \new_[27484]_ , \new_[27488]_ , \new_[27489]_ ,
    \new_[27493]_ , \new_[27494]_ , \new_[27495]_ , \new_[27499]_ ,
    \new_[27500]_ , \new_[27504]_ , \new_[27505]_ , \new_[27506]_ ,
    \new_[27510]_ , \new_[27511]_ , \new_[27515]_ , \new_[27516]_ ,
    \new_[27517]_ , \new_[27521]_ , \new_[27522]_ , \new_[27526]_ ,
    \new_[27527]_ , \new_[27528]_ , \new_[27532]_ , \new_[27533]_ ,
    \new_[27537]_ , \new_[27538]_ , \new_[27539]_ , \new_[27543]_ ,
    \new_[27544]_ , \new_[27548]_ , \new_[27549]_ , \new_[27550]_ ,
    \new_[27554]_ , \new_[27555]_ , \new_[27559]_ , \new_[27560]_ ,
    \new_[27561]_ , \new_[27565]_ , \new_[27566]_ , \new_[27570]_ ,
    \new_[27571]_ , \new_[27572]_ , \new_[27576]_ , \new_[27577]_ ,
    \new_[27581]_ , \new_[27582]_ , \new_[27583]_ , \new_[27587]_ ,
    \new_[27588]_ , \new_[27592]_ , \new_[27593]_ , \new_[27594]_ ,
    \new_[27598]_ , \new_[27599]_ , \new_[27603]_ , \new_[27604]_ ,
    \new_[27605]_ , \new_[27609]_ , \new_[27610]_ , \new_[27614]_ ,
    \new_[27615]_ , \new_[27616]_ , \new_[27620]_ , \new_[27621]_ ,
    \new_[27625]_ , \new_[27626]_ , \new_[27627]_ , \new_[27631]_ ,
    \new_[27632]_ , \new_[27636]_ , \new_[27637]_ , \new_[27638]_ ,
    \new_[27642]_ , \new_[27643]_ , \new_[27647]_ , \new_[27648]_ ,
    \new_[27649]_ , \new_[27653]_ , \new_[27654]_ , \new_[27658]_ ,
    \new_[27659]_ , \new_[27660]_ , \new_[27664]_ , \new_[27665]_ ,
    \new_[27669]_ , \new_[27670]_ , \new_[27671]_ , \new_[27675]_ ,
    \new_[27676]_ , \new_[27680]_ , \new_[27681]_ , \new_[27682]_ ,
    \new_[27686]_ , \new_[27687]_ , \new_[27691]_ , \new_[27692]_ ,
    \new_[27693]_ , \new_[27697]_ , \new_[27698]_ , \new_[27702]_ ,
    \new_[27703]_ , \new_[27704]_ , \new_[27708]_ , \new_[27709]_ ,
    \new_[27713]_ , \new_[27714]_ , \new_[27715]_ , \new_[27719]_ ,
    \new_[27720]_ , \new_[27724]_ , \new_[27725]_ , \new_[27726]_ ,
    \new_[27730]_ , \new_[27731]_ , \new_[27735]_ , \new_[27736]_ ,
    \new_[27737]_ , \new_[27741]_ , \new_[27742]_ , \new_[27746]_ ,
    \new_[27747]_ , \new_[27748]_ , \new_[27752]_ , \new_[27753]_ ,
    \new_[27757]_ , \new_[27758]_ , \new_[27759]_ , \new_[27763]_ ,
    \new_[27764]_ , \new_[27768]_ , \new_[27769]_ , \new_[27770]_ ,
    \new_[27774]_ , \new_[27775]_ , \new_[27779]_ , \new_[27780]_ ,
    \new_[27781]_ , \new_[27785]_ , \new_[27786]_ , \new_[27790]_ ,
    \new_[27791]_ , \new_[27792]_ , \new_[27796]_ , \new_[27797]_ ,
    \new_[27801]_ , \new_[27802]_ , \new_[27803]_ , \new_[27807]_ ,
    \new_[27808]_ , \new_[27812]_ , \new_[27813]_ , \new_[27814]_ ,
    \new_[27818]_ , \new_[27819]_ , \new_[27823]_ , \new_[27824]_ ,
    \new_[27825]_ , \new_[27829]_ , \new_[27830]_ , \new_[27834]_ ,
    \new_[27835]_ , \new_[27836]_ , \new_[27840]_ , \new_[27841]_ ,
    \new_[27845]_ , \new_[27846]_ , \new_[27847]_ , \new_[27851]_ ,
    \new_[27852]_ , \new_[27856]_ , \new_[27857]_ , \new_[27858]_ ,
    \new_[27862]_ , \new_[27863]_ , \new_[27867]_ , \new_[27868]_ ,
    \new_[27869]_ , \new_[27873]_ , \new_[27874]_ , \new_[27878]_ ,
    \new_[27879]_ , \new_[27880]_ , \new_[27884]_ , \new_[27885]_ ,
    \new_[27889]_ , \new_[27890]_ , \new_[27891]_ , \new_[27895]_ ,
    \new_[27896]_ , \new_[27900]_ , \new_[27901]_ , \new_[27902]_ ,
    \new_[27906]_ , \new_[27907]_ , \new_[27911]_ , \new_[27912]_ ,
    \new_[27913]_ , \new_[27917]_ , \new_[27918]_ , \new_[27922]_ ,
    \new_[27923]_ , \new_[27924]_ , \new_[27928]_ , \new_[27929]_ ,
    \new_[27933]_ , \new_[27934]_ , \new_[27935]_ , \new_[27939]_ ,
    \new_[27940]_ , \new_[27944]_ , \new_[27945]_ , \new_[27946]_ ,
    \new_[27950]_ , \new_[27951]_ , \new_[27955]_ , \new_[27956]_ ,
    \new_[27957]_ , \new_[27961]_ , \new_[27962]_ , \new_[27966]_ ,
    \new_[27967]_ , \new_[27968]_ , \new_[27972]_ , \new_[27973]_ ,
    \new_[27977]_ , \new_[27978]_ , \new_[27979]_ , \new_[27983]_ ,
    \new_[27984]_ , \new_[27988]_ , \new_[27989]_ , \new_[27990]_ ,
    \new_[27994]_ , \new_[27995]_ , \new_[27999]_ , \new_[28000]_ ,
    \new_[28001]_ , \new_[28005]_ , \new_[28006]_ , \new_[28010]_ ,
    \new_[28011]_ , \new_[28012]_ , \new_[28016]_ , \new_[28017]_ ,
    \new_[28021]_ , \new_[28022]_ , \new_[28023]_ , \new_[28027]_ ,
    \new_[28028]_ , \new_[28032]_ , \new_[28033]_ , \new_[28034]_ ,
    \new_[28038]_ , \new_[28039]_ , \new_[28043]_ , \new_[28044]_ ,
    \new_[28045]_ , \new_[28049]_ , \new_[28050]_ , \new_[28054]_ ,
    \new_[28055]_ , \new_[28056]_ , \new_[28060]_ , \new_[28061]_ ,
    \new_[28065]_ , \new_[28066]_ , \new_[28067]_ , \new_[28071]_ ,
    \new_[28072]_ , \new_[28076]_ , \new_[28077]_ , \new_[28078]_ ,
    \new_[28082]_ , \new_[28083]_ , \new_[28087]_ , \new_[28088]_ ,
    \new_[28089]_ , \new_[28093]_ , \new_[28094]_ , \new_[28098]_ ,
    \new_[28099]_ , \new_[28100]_ , \new_[28104]_ , \new_[28105]_ ,
    \new_[28109]_ , \new_[28110]_ , \new_[28111]_ , \new_[28115]_ ,
    \new_[28116]_ , \new_[28120]_ , \new_[28121]_ , \new_[28122]_ ,
    \new_[28126]_ , \new_[28127]_ , \new_[28131]_ , \new_[28132]_ ,
    \new_[28133]_ , \new_[28137]_ , \new_[28138]_ , \new_[28142]_ ,
    \new_[28143]_ , \new_[28144]_ , \new_[28148]_ , \new_[28149]_ ,
    \new_[28153]_ , \new_[28154]_ , \new_[28155]_ , \new_[28159]_ ,
    \new_[28160]_ , \new_[28164]_ , \new_[28165]_ , \new_[28166]_ ,
    \new_[28170]_ , \new_[28171]_ , \new_[28175]_ , \new_[28176]_ ,
    \new_[28177]_ , \new_[28181]_ , \new_[28182]_ , \new_[28186]_ ,
    \new_[28187]_ , \new_[28188]_ , \new_[28192]_ , \new_[28193]_ ,
    \new_[28197]_ , \new_[28198]_ , \new_[28199]_ , \new_[28203]_ ,
    \new_[28204]_ , \new_[28208]_ , \new_[28209]_ , \new_[28210]_ ,
    \new_[28214]_ , \new_[28215]_ , \new_[28219]_ , \new_[28220]_ ,
    \new_[28221]_ , \new_[28225]_ , \new_[28226]_ , \new_[28230]_ ,
    \new_[28231]_ , \new_[28232]_ , \new_[28236]_ , \new_[28237]_ ,
    \new_[28241]_ , \new_[28242]_ , \new_[28243]_ , \new_[28247]_ ,
    \new_[28248]_ , \new_[28252]_ , \new_[28253]_ , \new_[28254]_ ,
    \new_[28258]_ , \new_[28259]_ , \new_[28263]_ , \new_[28264]_ ,
    \new_[28265]_ , \new_[28269]_ , \new_[28270]_ , \new_[28274]_ ,
    \new_[28275]_ , \new_[28276]_ , \new_[28280]_ , \new_[28281]_ ,
    \new_[28285]_ , \new_[28286]_ , \new_[28287]_ , \new_[28291]_ ,
    \new_[28292]_ , \new_[28296]_ , \new_[28297]_ , \new_[28298]_ ,
    \new_[28302]_ , \new_[28303]_ , \new_[28307]_ , \new_[28308]_ ,
    \new_[28309]_ , \new_[28313]_ , \new_[28314]_ , \new_[28318]_ ,
    \new_[28319]_ , \new_[28320]_ , \new_[28324]_ , \new_[28325]_ ,
    \new_[28329]_ , \new_[28330]_ , \new_[28331]_ , \new_[28335]_ ,
    \new_[28336]_ , \new_[28340]_ , \new_[28341]_ , \new_[28342]_ ,
    \new_[28346]_ , \new_[28347]_ , \new_[28351]_ , \new_[28352]_ ,
    \new_[28353]_ , \new_[28357]_ , \new_[28358]_ , \new_[28362]_ ,
    \new_[28363]_ , \new_[28364]_ , \new_[28368]_ , \new_[28369]_ ,
    \new_[28373]_ , \new_[28374]_ , \new_[28375]_ , \new_[28379]_ ,
    \new_[28380]_ , \new_[28384]_ , \new_[28385]_ , \new_[28386]_ ,
    \new_[28390]_ , \new_[28391]_ , \new_[28395]_ , \new_[28396]_ ,
    \new_[28397]_ , \new_[28401]_ , \new_[28402]_ , \new_[28406]_ ,
    \new_[28407]_ , \new_[28408]_ , \new_[28412]_ , \new_[28413]_ ,
    \new_[28417]_ , \new_[28418]_ , \new_[28419]_ , \new_[28423]_ ,
    \new_[28424]_ , \new_[28428]_ , \new_[28429]_ , \new_[28430]_ ,
    \new_[28434]_ , \new_[28435]_ , \new_[28439]_ , \new_[28440]_ ,
    \new_[28441]_ , \new_[28445]_ , \new_[28446]_ , \new_[28450]_ ,
    \new_[28451]_ , \new_[28452]_ , \new_[28456]_ , \new_[28457]_ ,
    \new_[28461]_ , \new_[28462]_ , \new_[28463]_ , \new_[28467]_ ,
    \new_[28468]_ , \new_[28472]_ , \new_[28473]_ , \new_[28474]_ ,
    \new_[28478]_ , \new_[28479]_ , \new_[28483]_ , \new_[28484]_ ,
    \new_[28485]_ , \new_[28489]_ , \new_[28490]_ , \new_[28494]_ ,
    \new_[28495]_ , \new_[28496]_ , \new_[28500]_ , \new_[28501]_ ,
    \new_[28505]_ , \new_[28506]_ , \new_[28507]_ , \new_[28511]_ ,
    \new_[28512]_ , \new_[28516]_ , \new_[28517]_ , \new_[28518]_ ,
    \new_[28522]_ , \new_[28523]_ , \new_[28527]_ , \new_[28528]_ ,
    \new_[28529]_ , \new_[28533]_ , \new_[28534]_ , \new_[28538]_ ,
    \new_[28539]_ , \new_[28540]_ , \new_[28544]_ , \new_[28545]_ ,
    \new_[28549]_ , \new_[28550]_ , \new_[28551]_ , \new_[28555]_ ,
    \new_[28556]_ , \new_[28560]_ , \new_[28561]_ , \new_[28562]_ ,
    \new_[28566]_ , \new_[28567]_ , \new_[28571]_ , \new_[28572]_ ,
    \new_[28573]_ , \new_[28577]_ , \new_[28578]_ , \new_[28582]_ ,
    \new_[28583]_ , \new_[28584]_ , \new_[28588]_ , \new_[28589]_ ,
    \new_[28593]_ , \new_[28594]_ , \new_[28595]_ , \new_[28599]_ ,
    \new_[28600]_ , \new_[28604]_ , \new_[28605]_ , \new_[28606]_ ,
    \new_[28610]_ , \new_[28611]_ , \new_[28615]_ , \new_[28616]_ ,
    \new_[28617]_ , \new_[28621]_ , \new_[28622]_ , \new_[28626]_ ,
    \new_[28627]_ , \new_[28628]_ , \new_[28632]_ , \new_[28633]_ ,
    \new_[28637]_ , \new_[28638]_ , \new_[28639]_ , \new_[28643]_ ,
    \new_[28644]_ , \new_[28648]_ , \new_[28649]_ , \new_[28650]_ ,
    \new_[28654]_ , \new_[28655]_ , \new_[28659]_ , \new_[28660]_ ,
    \new_[28661]_ , \new_[28665]_ , \new_[28666]_ , \new_[28670]_ ,
    \new_[28671]_ , \new_[28672]_ , \new_[28676]_ , \new_[28677]_ ,
    \new_[28681]_ , \new_[28682]_ , \new_[28683]_ , \new_[28687]_ ,
    \new_[28688]_ , \new_[28692]_ , \new_[28693]_ , \new_[28694]_ ,
    \new_[28698]_ , \new_[28699]_ , \new_[28703]_ , \new_[28704]_ ,
    \new_[28705]_ , \new_[28709]_ , \new_[28710]_ , \new_[28714]_ ,
    \new_[28715]_ , \new_[28716]_ , \new_[28720]_ , \new_[28721]_ ,
    \new_[28725]_ , \new_[28726]_ , \new_[28727]_ , \new_[28731]_ ,
    \new_[28732]_ , \new_[28736]_ , \new_[28737]_ , \new_[28738]_ ,
    \new_[28742]_ , \new_[28743]_ , \new_[28747]_ , \new_[28748]_ ,
    \new_[28749]_ , \new_[28753]_ , \new_[28754]_ , \new_[28758]_ ,
    \new_[28759]_ , \new_[28760]_ , \new_[28764]_ , \new_[28765]_ ,
    \new_[28769]_ , \new_[28770]_ , \new_[28771]_ , \new_[28775]_ ,
    \new_[28776]_ , \new_[28780]_ , \new_[28781]_ , \new_[28782]_ ,
    \new_[28786]_ , \new_[28787]_ , \new_[28791]_ , \new_[28792]_ ,
    \new_[28793]_ , \new_[28797]_ , \new_[28798]_ , \new_[28802]_ ,
    \new_[28803]_ , \new_[28804]_ , \new_[28808]_ , \new_[28809]_ ,
    \new_[28813]_ , \new_[28814]_ , \new_[28815]_ , \new_[28819]_ ,
    \new_[28820]_ , \new_[28824]_ , \new_[28825]_ , \new_[28826]_ ,
    \new_[28830]_ , \new_[28831]_ , \new_[28835]_ , \new_[28836]_ ,
    \new_[28837]_ , \new_[28841]_ , \new_[28842]_ , \new_[28846]_ ,
    \new_[28847]_ , \new_[28848]_ , \new_[28852]_ , \new_[28853]_ ,
    \new_[28857]_ , \new_[28858]_ , \new_[28859]_ , \new_[28863]_ ,
    \new_[28864]_ , \new_[28868]_ , \new_[28869]_ , \new_[28870]_ ,
    \new_[28874]_ , \new_[28875]_ , \new_[28879]_ , \new_[28880]_ ,
    \new_[28881]_ , \new_[28885]_ , \new_[28886]_ , \new_[28890]_ ,
    \new_[28891]_ , \new_[28892]_ , \new_[28896]_ , \new_[28897]_ ,
    \new_[28901]_ , \new_[28902]_ , \new_[28903]_ , \new_[28907]_ ,
    \new_[28908]_ , \new_[28912]_ , \new_[28913]_ , \new_[28914]_ ,
    \new_[28918]_ , \new_[28919]_ , \new_[28923]_ , \new_[28924]_ ,
    \new_[28925]_ , \new_[28929]_ , \new_[28930]_ , \new_[28934]_ ,
    \new_[28935]_ , \new_[28936]_ , \new_[28940]_ , \new_[28941]_ ,
    \new_[28945]_ , \new_[28946]_ , \new_[28947]_ , \new_[28951]_ ,
    \new_[28952]_ , \new_[28956]_ , \new_[28957]_ , \new_[28958]_ ,
    \new_[28962]_ , \new_[28963]_ , \new_[28967]_ , \new_[28968]_ ,
    \new_[28969]_ , \new_[28973]_ , \new_[28974]_ , \new_[28978]_ ,
    \new_[28979]_ , \new_[28980]_ , \new_[28984]_ , \new_[28985]_ ,
    \new_[28989]_ , \new_[28990]_ , \new_[28991]_ , \new_[28995]_ ,
    \new_[28996]_ , \new_[29000]_ , \new_[29001]_ , \new_[29002]_ ,
    \new_[29006]_ , \new_[29007]_ , \new_[29011]_ , \new_[29012]_ ,
    \new_[29013]_ , \new_[29017]_ , \new_[29018]_ , \new_[29022]_ ,
    \new_[29023]_ , \new_[29024]_ , \new_[29028]_ , \new_[29029]_ ,
    \new_[29033]_ , \new_[29034]_ , \new_[29035]_ , \new_[29039]_ ,
    \new_[29040]_ , \new_[29044]_ , \new_[29045]_ , \new_[29046]_ ,
    \new_[29050]_ , \new_[29051]_ , \new_[29055]_ , \new_[29056]_ ,
    \new_[29057]_ , \new_[29061]_ , \new_[29062]_ , \new_[29066]_ ,
    \new_[29067]_ , \new_[29068]_ , \new_[29072]_ , \new_[29073]_ ,
    \new_[29077]_ , \new_[29078]_ , \new_[29079]_ , \new_[29083]_ ,
    \new_[29084]_ , \new_[29088]_ , \new_[29089]_ , \new_[29090]_ ,
    \new_[29094]_ , \new_[29095]_ , \new_[29099]_ , \new_[29100]_ ,
    \new_[29101]_ , \new_[29105]_ , \new_[29106]_ , \new_[29110]_ ,
    \new_[29111]_ , \new_[29112]_ , \new_[29116]_ , \new_[29117]_ ,
    \new_[29121]_ , \new_[29122]_ , \new_[29123]_ , \new_[29127]_ ,
    \new_[29128]_ , \new_[29132]_ , \new_[29133]_ , \new_[29134]_ ,
    \new_[29138]_ , \new_[29139]_ , \new_[29143]_ , \new_[29144]_ ,
    \new_[29145]_ , \new_[29149]_ , \new_[29150]_ , \new_[29154]_ ,
    \new_[29155]_ , \new_[29156]_ , \new_[29160]_ , \new_[29161]_ ,
    \new_[29165]_ , \new_[29166]_ , \new_[29167]_ , \new_[29171]_ ,
    \new_[29172]_ , \new_[29176]_ , \new_[29177]_ , \new_[29178]_ ,
    \new_[29182]_ , \new_[29183]_ , \new_[29187]_ , \new_[29188]_ ,
    \new_[29189]_ , \new_[29193]_ , \new_[29194]_ , \new_[29198]_ ,
    \new_[29199]_ , \new_[29200]_ , \new_[29204]_ , \new_[29205]_ ,
    \new_[29209]_ , \new_[29210]_ , \new_[29211]_ , \new_[29215]_ ,
    \new_[29216]_ , \new_[29220]_ , \new_[29221]_ , \new_[29222]_ ,
    \new_[29226]_ , \new_[29227]_ , \new_[29231]_ , \new_[29232]_ ,
    \new_[29233]_ , \new_[29237]_ , \new_[29238]_ , \new_[29242]_ ,
    \new_[29243]_ , \new_[29244]_ , \new_[29248]_ , \new_[29249]_ ,
    \new_[29253]_ , \new_[29254]_ , \new_[29255]_ , \new_[29259]_ ,
    \new_[29260]_ , \new_[29264]_ , \new_[29265]_ , \new_[29266]_ ,
    \new_[29270]_ , \new_[29271]_ , \new_[29275]_ , \new_[29276]_ ,
    \new_[29277]_ , \new_[29281]_ , \new_[29282]_ , \new_[29286]_ ,
    \new_[29287]_ , \new_[29288]_ , \new_[29292]_ , \new_[29293]_ ,
    \new_[29297]_ , \new_[29298]_ , \new_[29299]_ , \new_[29303]_ ,
    \new_[29304]_ , \new_[29308]_ , \new_[29309]_ , \new_[29310]_ ,
    \new_[29314]_ , \new_[29315]_ , \new_[29319]_ , \new_[29320]_ ,
    \new_[29321]_ , \new_[29325]_ , \new_[29326]_ , \new_[29330]_ ,
    \new_[29331]_ , \new_[29332]_ , \new_[29336]_ , \new_[29337]_ ,
    \new_[29341]_ , \new_[29342]_ , \new_[29343]_ , \new_[29347]_ ,
    \new_[29348]_ , \new_[29352]_ , \new_[29353]_ , \new_[29354]_ ,
    \new_[29358]_ , \new_[29359]_ , \new_[29363]_ , \new_[29364]_ ,
    \new_[29365]_ , \new_[29369]_ , \new_[29370]_ , \new_[29374]_ ,
    \new_[29375]_ , \new_[29376]_ , \new_[29380]_ , \new_[29381]_ ,
    \new_[29385]_ , \new_[29386]_ , \new_[29387]_ , \new_[29391]_ ,
    \new_[29392]_ , \new_[29396]_ , \new_[29397]_ , \new_[29398]_ ,
    \new_[29402]_ , \new_[29403]_ , \new_[29407]_ , \new_[29408]_ ,
    \new_[29409]_ , \new_[29413]_ , \new_[29414]_ , \new_[29418]_ ,
    \new_[29419]_ , \new_[29420]_ , \new_[29424]_ , \new_[29425]_ ,
    \new_[29429]_ , \new_[29430]_ , \new_[29431]_ , \new_[29435]_ ,
    \new_[29436]_ , \new_[29440]_ , \new_[29441]_ , \new_[29442]_ ,
    \new_[29446]_ , \new_[29447]_ , \new_[29451]_ , \new_[29452]_ ,
    \new_[29453]_ , \new_[29457]_ , \new_[29458]_ , \new_[29462]_ ,
    \new_[29463]_ , \new_[29464]_ , \new_[29468]_ , \new_[29469]_ ,
    \new_[29473]_ , \new_[29474]_ , \new_[29475]_ , \new_[29479]_ ,
    \new_[29480]_ , \new_[29484]_ , \new_[29485]_ , \new_[29486]_ ,
    \new_[29490]_ , \new_[29491]_ , \new_[29495]_ , \new_[29496]_ ,
    \new_[29497]_ , \new_[29501]_ , \new_[29502]_ , \new_[29506]_ ,
    \new_[29507]_ , \new_[29508]_ , \new_[29512]_ , \new_[29513]_ ,
    \new_[29517]_ , \new_[29518]_ , \new_[29519]_ , \new_[29523]_ ,
    \new_[29524]_ , \new_[29528]_ , \new_[29529]_ , \new_[29530]_ ,
    \new_[29534]_ , \new_[29535]_ , \new_[29539]_ , \new_[29540]_ ,
    \new_[29541]_ , \new_[29545]_ , \new_[29546]_ , \new_[29550]_ ,
    \new_[29551]_ , \new_[29552]_ , \new_[29556]_ , \new_[29557]_ ,
    \new_[29561]_ , \new_[29562]_ , \new_[29563]_ , \new_[29567]_ ,
    \new_[29568]_ , \new_[29572]_ , \new_[29573]_ , \new_[29574]_ ,
    \new_[29578]_ , \new_[29579]_ , \new_[29583]_ , \new_[29584]_ ,
    \new_[29585]_ , \new_[29589]_ , \new_[29590]_ , \new_[29594]_ ,
    \new_[29595]_ , \new_[29596]_ , \new_[29600]_ , \new_[29601]_ ,
    \new_[29605]_ , \new_[29606]_ , \new_[29607]_ , \new_[29611]_ ,
    \new_[29612]_ , \new_[29616]_ , \new_[29617]_ , \new_[29618]_ ,
    \new_[29622]_ , \new_[29623]_ , \new_[29627]_ , \new_[29628]_ ,
    \new_[29629]_ , \new_[29633]_ , \new_[29634]_ , \new_[29638]_ ,
    \new_[29639]_ , \new_[29640]_ , \new_[29644]_ , \new_[29645]_ ,
    \new_[29649]_ , \new_[29650]_ , \new_[29651]_ , \new_[29655]_ ,
    \new_[29656]_ , \new_[29660]_ , \new_[29661]_ , \new_[29662]_ ,
    \new_[29666]_ , \new_[29667]_ , \new_[29671]_ , \new_[29672]_ ,
    \new_[29673]_ , \new_[29677]_ , \new_[29678]_ , \new_[29682]_ ,
    \new_[29683]_ , \new_[29684]_ , \new_[29688]_ , \new_[29689]_ ,
    \new_[29693]_ , \new_[29694]_ , \new_[29695]_ , \new_[29699]_ ,
    \new_[29700]_ , \new_[29704]_ , \new_[29705]_ , \new_[29706]_ ,
    \new_[29710]_ , \new_[29711]_ , \new_[29715]_ , \new_[29716]_ ,
    \new_[29717]_ , \new_[29721]_ , \new_[29722]_ , \new_[29726]_ ,
    \new_[29727]_ , \new_[29728]_ , \new_[29732]_ , \new_[29733]_ ,
    \new_[29737]_ , \new_[29738]_ , \new_[29739]_ , \new_[29743]_ ,
    \new_[29744]_ , \new_[29748]_ , \new_[29749]_ , \new_[29750]_ ,
    \new_[29754]_ , \new_[29755]_ , \new_[29759]_ , \new_[29760]_ ,
    \new_[29761]_ , \new_[29765]_ , \new_[29766]_ , \new_[29770]_ ,
    \new_[29771]_ , \new_[29772]_ , \new_[29776]_ , \new_[29777]_ ,
    \new_[29781]_ , \new_[29782]_ , \new_[29783]_ , \new_[29787]_ ,
    \new_[29788]_ , \new_[29792]_ , \new_[29793]_ , \new_[29794]_ ,
    \new_[29798]_ , \new_[29799]_ , \new_[29803]_ , \new_[29804]_ ,
    \new_[29805]_ , \new_[29809]_ , \new_[29810]_ , \new_[29814]_ ,
    \new_[29815]_ , \new_[29816]_ , \new_[29820]_ , \new_[29821]_ ,
    \new_[29825]_ , \new_[29826]_ , \new_[29827]_ , \new_[29831]_ ,
    \new_[29832]_ , \new_[29836]_ , \new_[29837]_ , \new_[29838]_ ,
    \new_[29842]_ , \new_[29843]_ , \new_[29847]_ , \new_[29848]_ ,
    \new_[29849]_ , \new_[29853]_ , \new_[29854]_ , \new_[29858]_ ,
    \new_[29859]_ , \new_[29860]_ , \new_[29864]_ , \new_[29865]_ ,
    \new_[29869]_ , \new_[29870]_ , \new_[29871]_ , \new_[29875]_ ,
    \new_[29876]_ , \new_[29880]_ , \new_[29881]_ , \new_[29882]_ ,
    \new_[29886]_ , \new_[29887]_ , \new_[29891]_ , \new_[29892]_ ,
    \new_[29893]_ , \new_[29897]_ , \new_[29898]_ , \new_[29902]_ ,
    \new_[29903]_ , \new_[29904]_ , \new_[29908]_ , \new_[29909]_ ,
    \new_[29913]_ , \new_[29914]_ , \new_[29915]_ , \new_[29919]_ ,
    \new_[29920]_ , \new_[29924]_ , \new_[29925]_ , \new_[29926]_ ,
    \new_[29930]_ , \new_[29931]_ , \new_[29935]_ , \new_[29936]_ ,
    \new_[29937]_ , \new_[29941]_ , \new_[29942]_ , \new_[29946]_ ,
    \new_[29947]_ , \new_[29948]_ , \new_[29952]_ , \new_[29953]_ ,
    \new_[29957]_ , \new_[29958]_ , \new_[29959]_ , \new_[29963]_ ,
    \new_[29964]_ , \new_[29968]_ , \new_[29969]_ , \new_[29970]_ ,
    \new_[29974]_ , \new_[29975]_ , \new_[29979]_ , \new_[29980]_ ,
    \new_[29981]_ , \new_[29985]_ , \new_[29986]_ , \new_[29990]_ ,
    \new_[29991]_ , \new_[29992]_ , \new_[29996]_ , \new_[29997]_ ,
    \new_[30001]_ , \new_[30002]_ , \new_[30003]_ , \new_[30007]_ ,
    \new_[30008]_ , \new_[30012]_ , \new_[30013]_ , \new_[30014]_ ,
    \new_[30018]_ , \new_[30019]_ , \new_[30023]_ , \new_[30024]_ ,
    \new_[30025]_ , \new_[30029]_ , \new_[30030]_ , \new_[30034]_ ,
    \new_[30035]_ , \new_[30036]_ , \new_[30040]_ , \new_[30041]_ ,
    \new_[30045]_ , \new_[30046]_ , \new_[30047]_ , \new_[30051]_ ,
    \new_[30052]_ , \new_[30056]_ , \new_[30057]_ , \new_[30058]_ ,
    \new_[30062]_ , \new_[30063]_ , \new_[30067]_ , \new_[30068]_ ,
    \new_[30069]_ , \new_[30073]_ , \new_[30074]_ , \new_[30078]_ ,
    \new_[30079]_ , \new_[30080]_ , \new_[30084]_ , \new_[30085]_ ,
    \new_[30089]_ , \new_[30090]_ , \new_[30091]_ , \new_[30095]_ ,
    \new_[30096]_ , \new_[30100]_ , \new_[30101]_ , \new_[30102]_ ,
    \new_[30106]_ , \new_[30107]_ , \new_[30111]_ , \new_[30112]_ ,
    \new_[30113]_ , \new_[30117]_ , \new_[30118]_ , \new_[30122]_ ,
    \new_[30123]_ , \new_[30124]_ , \new_[30128]_ , \new_[30129]_ ,
    \new_[30133]_ , \new_[30134]_ , \new_[30135]_ , \new_[30139]_ ,
    \new_[30140]_ , \new_[30144]_ , \new_[30145]_ , \new_[30146]_ ,
    \new_[30150]_ , \new_[30151]_ , \new_[30155]_ , \new_[30156]_ ,
    \new_[30157]_ , \new_[30161]_ , \new_[30162]_ , \new_[30166]_ ,
    \new_[30167]_ , \new_[30168]_ , \new_[30172]_ , \new_[30173]_ ,
    \new_[30177]_ , \new_[30178]_ , \new_[30179]_ , \new_[30183]_ ,
    \new_[30184]_ , \new_[30188]_ , \new_[30189]_ , \new_[30190]_ ,
    \new_[30194]_ , \new_[30195]_ , \new_[30199]_ , \new_[30200]_ ,
    \new_[30201]_ , \new_[30205]_ , \new_[30206]_ , \new_[30210]_ ,
    \new_[30211]_ , \new_[30212]_ , \new_[30216]_ , \new_[30217]_ ,
    \new_[30221]_ , \new_[30222]_ , \new_[30223]_ , \new_[30227]_ ,
    \new_[30228]_ , \new_[30232]_ , \new_[30233]_ , \new_[30234]_ ,
    \new_[30238]_ , \new_[30239]_ , \new_[30243]_ , \new_[30244]_ ,
    \new_[30245]_ , \new_[30249]_ , \new_[30250]_ , \new_[30254]_ ,
    \new_[30255]_ , \new_[30256]_ , \new_[30260]_ , \new_[30261]_ ,
    \new_[30265]_ , \new_[30266]_ , \new_[30267]_ , \new_[30271]_ ,
    \new_[30272]_ , \new_[30276]_ , \new_[30277]_ , \new_[30278]_ ,
    \new_[30282]_ , \new_[30283]_ , \new_[30287]_ , \new_[30288]_ ,
    \new_[30289]_ , \new_[30293]_ , \new_[30294]_ , \new_[30298]_ ,
    \new_[30299]_ , \new_[30300]_ , \new_[30304]_ , \new_[30305]_ ,
    \new_[30309]_ , \new_[30310]_ , \new_[30311]_ , \new_[30315]_ ,
    \new_[30316]_ , \new_[30320]_ , \new_[30321]_ , \new_[30322]_ ,
    \new_[30326]_ , \new_[30327]_ , \new_[30331]_ , \new_[30332]_ ,
    \new_[30333]_ , \new_[30337]_ , \new_[30338]_ , \new_[30342]_ ,
    \new_[30343]_ , \new_[30344]_ , \new_[30348]_ , \new_[30349]_ ,
    \new_[30353]_ , \new_[30354]_ , \new_[30355]_ , \new_[30359]_ ,
    \new_[30360]_ , \new_[30364]_ , \new_[30365]_ , \new_[30366]_ ,
    \new_[30370]_ , \new_[30371]_ , \new_[30375]_ , \new_[30376]_ ,
    \new_[30377]_ , \new_[30381]_ , \new_[30382]_ , \new_[30386]_ ,
    \new_[30387]_ , \new_[30388]_ , \new_[30392]_ , \new_[30393]_ ,
    \new_[30397]_ , \new_[30398]_ , \new_[30399]_ , \new_[30403]_ ,
    \new_[30404]_ , \new_[30408]_ , \new_[30409]_ , \new_[30410]_ ,
    \new_[30414]_ , \new_[30415]_ , \new_[30419]_ , \new_[30420]_ ,
    \new_[30421]_ , \new_[30425]_ , \new_[30426]_ , \new_[30430]_ ,
    \new_[30431]_ , \new_[30432]_ , \new_[30436]_ , \new_[30437]_ ,
    \new_[30441]_ , \new_[30442]_ , \new_[30443]_ , \new_[30447]_ ,
    \new_[30448]_ , \new_[30452]_ , \new_[30453]_ , \new_[30454]_ ,
    \new_[30458]_ , \new_[30459]_ , \new_[30463]_ , \new_[30464]_ ,
    \new_[30465]_ , \new_[30469]_ , \new_[30470]_ , \new_[30474]_ ,
    \new_[30475]_ , \new_[30476]_ , \new_[30480]_ , \new_[30481]_ ,
    \new_[30485]_ , \new_[30486]_ , \new_[30487]_ , \new_[30491]_ ,
    \new_[30492]_ , \new_[30496]_ , \new_[30497]_ , \new_[30498]_ ,
    \new_[30502]_ , \new_[30503]_ , \new_[30507]_ , \new_[30508]_ ,
    \new_[30509]_ , \new_[30513]_ , \new_[30514]_ , \new_[30518]_ ,
    \new_[30519]_ , \new_[30520]_ , \new_[30524]_ , \new_[30525]_ ,
    \new_[30529]_ , \new_[30530]_ , \new_[30531]_ , \new_[30535]_ ,
    \new_[30536]_ , \new_[30540]_ , \new_[30541]_ , \new_[30542]_ ,
    \new_[30546]_ , \new_[30547]_ , \new_[30551]_ , \new_[30552]_ ,
    \new_[30553]_ , \new_[30557]_ , \new_[30558]_ , \new_[30562]_ ,
    \new_[30563]_ , \new_[30564]_ , \new_[30568]_ , \new_[30569]_ ,
    \new_[30573]_ , \new_[30574]_ , \new_[30575]_ , \new_[30579]_ ,
    \new_[30580]_ , \new_[30584]_ , \new_[30585]_ , \new_[30586]_ ,
    \new_[30590]_ , \new_[30591]_ , \new_[30595]_ , \new_[30596]_ ,
    \new_[30597]_ , \new_[30601]_ , \new_[30602]_ , \new_[30606]_ ,
    \new_[30607]_ , \new_[30608]_ , \new_[30612]_ , \new_[30613]_ ,
    \new_[30617]_ , \new_[30618]_ , \new_[30619]_ , \new_[30623]_ ,
    \new_[30624]_ , \new_[30628]_ , \new_[30629]_ , \new_[30630]_ ,
    \new_[30634]_ , \new_[30635]_ , \new_[30639]_ , \new_[30640]_ ,
    \new_[30641]_ , \new_[30645]_ , \new_[30646]_ , \new_[30650]_ ,
    \new_[30651]_ , \new_[30652]_ , \new_[30656]_ , \new_[30657]_ ,
    \new_[30661]_ , \new_[30662]_ , \new_[30663]_ , \new_[30667]_ ,
    \new_[30668]_ , \new_[30672]_ , \new_[30673]_ , \new_[30674]_ ,
    \new_[30678]_ , \new_[30679]_ , \new_[30683]_ , \new_[30684]_ ,
    \new_[30685]_ , \new_[30689]_ , \new_[30690]_ , \new_[30694]_ ,
    \new_[30695]_ , \new_[30696]_ , \new_[30700]_ , \new_[30701]_ ,
    \new_[30705]_ , \new_[30706]_ , \new_[30707]_ , \new_[30711]_ ,
    \new_[30712]_ , \new_[30716]_ , \new_[30717]_ , \new_[30718]_ ,
    \new_[30722]_ , \new_[30723]_ , \new_[30727]_ , \new_[30728]_ ,
    \new_[30729]_ , \new_[30733]_ , \new_[30734]_ , \new_[30738]_ ,
    \new_[30739]_ , \new_[30740]_ , \new_[30744]_ , \new_[30745]_ ,
    \new_[30749]_ , \new_[30750]_ , \new_[30751]_ , \new_[30755]_ ,
    \new_[30756]_ , \new_[30760]_ , \new_[30761]_ , \new_[30762]_ ,
    \new_[30766]_ , \new_[30767]_ , \new_[30771]_ , \new_[30772]_ ,
    \new_[30773]_ , \new_[30777]_ , \new_[30778]_ , \new_[30782]_ ,
    \new_[30783]_ , \new_[30784]_ , \new_[30788]_ , \new_[30789]_ ,
    \new_[30793]_ , \new_[30794]_ , \new_[30795]_ , \new_[30799]_ ,
    \new_[30800]_ , \new_[30804]_ , \new_[30805]_ , \new_[30806]_ ,
    \new_[30810]_ , \new_[30811]_ , \new_[30815]_ , \new_[30816]_ ,
    \new_[30817]_ , \new_[30821]_ , \new_[30822]_ , \new_[30826]_ ,
    \new_[30827]_ , \new_[30828]_ , \new_[30832]_ , \new_[30833]_ ,
    \new_[30837]_ , \new_[30838]_ , \new_[30839]_ , \new_[30843]_ ,
    \new_[30844]_ , \new_[30848]_ , \new_[30849]_ , \new_[30850]_ ,
    \new_[30854]_ , \new_[30855]_ , \new_[30859]_ , \new_[30860]_ ,
    \new_[30861]_ , \new_[30865]_ , \new_[30866]_ , \new_[30870]_ ,
    \new_[30871]_ , \new_[30872]_ , \new_[30876]_ , \new_[30877]_ ,
    \new_[30881]_ , \new_[30882]_ , \new_[30883]_ , \new_[30887]_ ,
    \new_[30888]_ , \new_[30892]_ , \new_[30893]_ , \new_[30894]_ ,
    \new_[30898]_ , \new_[30899]_ , \new_[30903]_ , \new_[30904]_ ,
    \new_[30905]_ , \new_[30909]_ , \new_[30910]_ , \new_[30914]_ ,
    \new_[30915]_ , \new_[30916]_ , \new_[30920]_ , \new_[30921]_ ,
    \new_[30925]_ , \new_[30926]_ , \new_[30927]_ , \new_[30931]_ ,
    \new_[30932]_ , \new_[30936]_ , \new_[30937]_ , \new_[30938]_ ,
    \new_[30942]_ , \new_[30943]_ , \new_[30947]_ , \new_[30948]_ ,
    \new_[30949]_ , \new_[30953]_ , \new_[30954]_ , \new_[30958]_ ,
    \new_[30959]_ , \new_[30960]_ , \new_[30964]_ , \new_[30965]_ ,
    \new_[30969]_ , \new_[30970]_ , \new_[30971]_ , \new_[30975]_ ,
    \new_[30976]_ , \new_[30980]_ , \new_[30981]_ , \new_[30982]_ ,
    \new_[30986]_ , \new_[30987]_ , \new_[30991]_ , \new_[30992]_ ,
    \new_[30993]_ , \new_[30997]_ , \new_[30998]_ , \new_[31002]_ ,
    \new_[31003]_ , \new_[31004]_ , \new_[31008]_ , \new_[31009]_ ,
    \new_[31013]_ , \new_[31014]_ , \new_[31015]_ , \new_[31019]_ ,
    \new_[31020]_ , \new_[31024]_ , \new_[31025]_ , \new_[31026]_ ,
    \new_[31030]_ , \new_[31031]_ , \new_[31035]_ , \new_[31036]_ ,
    \new_[31037]_ , \new_[31041]_ , \new_[31042]_ , \new_[31046]_ ,
    \new_[31047]_ , \new_[31048]_ , \new_[31052]_ , \new_[31053]_ ,
    \new_[31057]_ , \new_[31058]_ , \new_[31059]_ , \new_[31063]_ ,
    \new_[31064]_ , \new_[31068]_ , \new_[31069]_ , \new_[31070]_ ,
    \new_[31074]_ , \new_[31075]_ , \new_[31079]_ , \new_[31080]_ ,
    \new_[31081]_ , \new_[31085]_ , \new_[31086]_ , \new_[31090]_ ,
    \new_[31091]_ , \new_[31092]_ , \new_[31096]_ , \new_[31097]_ ,
    \new_[31101]_ , \new_[31102]_ , \new_[31103]_ , \new_[31107]_ ,
    \new_[31108]_ , \new_[31112]_ , \new_[31113]_ , \new_[31114]_ ,
    \new_[31118]_ , \new_[31119]_ , \new_[31123]_ , \new_[31124]_ ,
    \new_[31125]_ , \new_[31129]_ , \new_[31130]_ , \new_[31134]_ ,
    \new_[31135]_ , \new_[31136]_ , \new_[31140]_ , \new_[31141]_ ,
    \new_[31145]_ , \new_[31146]_ , \new_[31147]_ , \new_[31151]_ ,
    \new_[31152]_ , \new_[31156]_ , \new_[31157]_ , \new_[31158]_ ,
    \new_[31162]_ , \new_[31163]_ , \new_[31167]_ , \new_[31168]_ ,
    \new_[31169]_ , \new_[31173]_ , \new_[31174]_ , \new_[31178]_ ,
    \new_[31179]_ , \new_[31180]_ , \new_[31184]_ , \new_[31185]_ ,
    \new_[31189]_ , \new_[31190]_ , \new_[31191]_ , \new_[31195]_ ,
    \new_[31196]_ , \new_[31200]_ , \new_[31201]_ , \new_[31202]_ ,
    \new_[31206]_ , \new_[31207]_ , \new_[31211]_ , \new_[31212]_ ,
    \new_[31213]_ , \new_[31217]_ , \new_[31218]_ , \new_[31222]_ ,
    \new_[31223]_ , \new_[31224]_ , \new_[31228]_ , \new_[31229]_ ,
    \new_[31233]_ , \new_[31234]_ , \new_[31235]_ , \new_[31239]_ ,
    \new_[31240]_ , \new_[31244]_ , \new_[31245]_ , \new_[31246]_ ,
    \new_[31250]_ , \new_[31251]_ , \new_[31255]_ , \new_[31256]_ ,
    \new_[31257]_ , \new_[31261]_ , \new_[31262]_ , \new_[31266]_ ,
    \new_[31267]_ , \new_[31268]_ , \new_[31272]_ , \new_[31273]_ ,
    \new_[31277]_ , \new_[31278]_ , \new_[31279]_ , \new_[31283]_ ,
    \new_[31284]_ , \new_[31288]_ , \new_[31289]_ , \new_[31290]_ ,
    \new_[31294]_ , \new_[31295]_ , \new_[31299]_ , \new_[31300]_ ,
    \new_[31301]_ , \new_[31305]_ , \new_[31306]_ , \new_[31310]_ ,
    \new_[31311]_ , \new_[31312]_ , \new_[31316]_ , \new_[31317]_ ,
    \new_[31321]_ , \new_[31322]_ , \new_[31323]_ , \new_[31327]_ ,
    \new_[31328]_ , \new_[31332]_ , \new_[31333]_ , \new_[31334]_ ,
    \new_[31338]_ , \new_[31339]_ , \new_[31343]_ , \new_[31344]_ ,
    \new_[31345]_ , \new_[31349]_ , \new_[31350]_ , \new_[31354]_ ,
    \new_[31355]_ , \new_[31356]_ , \new_[31360]_ , \new_[31361]_ ,
    \new_[31365]_ , \new_[31366]_ , \new_[31367]_ , \new_[31371]_ ,
    \new_[31372]_ , \new_[31376]_ , \new_[31377]_ , \new_[31378]_ ,
    \new_[31382]_ , \new_[31383]_ , \new_[31387]_ , \new_[31388]_ ,
    \new_[31389]_ , \new_[31393]_ , \new_[31394]_ , \new_[31398]_ ,
    \new_[31399]_ , \new_[31400]_ , \new_[31404]_ , \new_[31405]_ ,
    \new_[31409]_ , \new_[31410]_ , \new_[31411]_ , \new_[31415]_ ,
    \new_[31416]_ , \new_[31420]_ , \new_[31421]_ , \new_[31422]_ ,
    \new_[31426]_ , \new_[31427]_ , \new_[31431]_ , \new_[31432]_ ,
    \new_[31433]_ , \new_[31437]_ , \new_[31438]_ , \new_[31442]_ ,
    \new_[31443]_ , \new_[31444]_ , \new_[31448]_ , \new_[31449]_ ,
    \new_[31453]_ , \new_[31454]_ , \new_[31455]_ , \new_[31459]_ ,
    \new_[31460]_ , \new_[31464]_ , \new_[31465]_ , \new_[31466]_ ,
    \new_[31470]_ , \new_[31471]_ , \new_[31475]_ , \new_[31476]_ ,
    \new_[31477]_ , \new_[31481]_ , \new_[31482]_ , \new_[31486]_ ,
    \new_[31487]_ , \new_[31488]_ , \new_[31492]_ , \new_[31493]_ ,
    \new_[31497]_ , \new_[31498]_ , \new_[31499]_ , \new_[31503]_ ,
    \new_[31504]_ , \new_[31508]_ , \new_[31509]_ , \new_[31510]_ ,
    \new_[31514]_ , \new_[31515]_ , \new_[31519]_ , \new_[31520]_ ,
    \new_[31521]_ , \new_[31525]_ , \new_[31526]_ , \new_[31530]_ ,
    \new_[31531]_ , \new_[31532]_ , \new_[31536]_ , \new_[31537]_ ,
    \new_[31541]_ , \new_[31542]_ , \new_[31543]_ , \new_[31547]_ ,
    \new_[31548]_ , \new_[31552]_ , \new_[31553]_ , \new_[31554]_ ,
    \new_[31558]_ , \new_[31559]_ , \new_[31563]_ , \new_[31564]_ ,
    \new_[31565]_ , \new_[31569]_ , \new_[31570]_ , \new_[31574]_ ,
    \new_[31575]_ , \new_[31576]_ , \new_[31580]_ , \new_[31581]_ ,
    \new_[31585]_ , \new_[31586]_ , \new_[31587]_ , \new_[31591]_ ,
    \new_[31592]_ , \new_[31596]_ , \new_[31597]_ , \new_[31598]_ ,
    \new_[31602]_ , \new_[31603]_ , \new_[31607]_ , \new_[31608]_ ,
    \new_[31609]_ , \new_[31613]_ , \new_[31614]_ , \new_[31618]_ ,
    \new_[31619]_ , \new_[31620]_ , \new_[31624]_ , \new_[31625]_ ,
    \new_[31629]_ , \new_[31630]_ , \new_[31631]_ , \new_[31635]_ ,
    \new_[31636]_ , \new_[31640]_ , \new_[31641]_ , \new_[31642]_ ,
    \new_[31646]_ , \new_[31647]_ , \new_[31651]_ , \new_[31652]_ ,
    \new_[31653]_ , \new_[31657]_ , \new_[31658]_ , \new_[31662]_ ,
    \new_[31663]_ , \new_[31664]_ , \new_[31668]_ , \new_[31669]_ ,
    \new_[31673]_ , \new_[31674]_ , \new_[31675]_ , \new_[31679]_ ,
    \new_[31680]_ , \new_[31684]_ , \new_[31685]_ , \new_[31686]_ ,
    \new_[31690]_ , \new_[31691]_ , \new_[31695]_ , \new_[31696]_ ,
    \new_[31697]_ , \new_[31701]_ , \new_[31702]_ , \new_[31706]_ ,
    \new_[31707]_ , \new_[31708]_ , \new_[31712]_ , \new_[31713]_ ,
    \new_[31717]_ , \new_[31718]_ , \new_[31719]_ , \new_[31723]_ ,
    \new_[31724]_ , \new_[31728]_ , \new_[31729]_ , \new_[31730]_ ,
    \new_[31734]_ , \new_[31735]_ , \new_[31739]_ , \new_[31740]_ ,
    \new_[31741]_ , \new_[31745]_ , \new_[31746]_ , \new_[31750]_ ,
    \new_[31751]_ , \new_[31752]_ , \new_[31756]_ , \new_[31757]_ ,
    \new_[31761]_ , \new_[31762]_ , \new_[31763]_ , \new_[31767]_ ,
    \new_[31768]_ , \new_[31772]_ , \new_[31773]_ , \new_[31774]_ ,
    \new_[31778]_ , \new_[31779]_ , \new_[31783]_ , \new_[31784]_ ,
    \new_[31785]_ , \new_[31789]_ , \new_[31790]_ , \new_[31794]_ ,
    \new_[31795]_ , \new_[31796]_ , \new_[31800]_ , \new_[31801]_ ,
    \new_[31805]_ , \new_[31806]_ , \new_[31807]_ , \new_[31811]_ ,
    \new_[31812]_ , \new_[31816]_ , \new_[31817]_ , \new_[31818]_ ,
    \new_[31822]_ , \new_[31823]_ , \new_[31827]_ , \new_[31828]_ ,
    \new_[31829]_ , \new_[31833]_ , \new_[31834]_ , \new_[31838]_ ,
    \new_[31839]_ , \new_[31840]_ , \new_[31844]_ , \new_[31845]_ ,
    \new_[31849]_ , \new_[31850]_ , \new_[31851]_ , \new_[31855]_ ,
    \new_[31856]_ , \new_[31860]_ , \new_[31861]_ , \new_[31862]_ ,
    \new_[31866]_ , \new_[31867]_ , \new_[31871]_ , \new_[31872]_ ,
    \new_[31873]_ , \new_[31877]_ , \new_[31878]_ , \new_[31882]_ ,
    \new_[31883]_ , \new_[31884]_ , \new_[31888]_ , \new_[31889]_ ,
    \new_[31893]_ , \new_[31894]_ , \new_[31895]_ , \new_[31899]_ ,
    \new_[31900]_ , \new_[31904]_ , \new_[31905]_ , \new_[31906]_ ,
    \new_[31910]_ , \new_[31911]_ , \new_[31915]_ , \new_[31916]_ ,
    \new_[31917]_ , \new_[31921]_ , \new_[31922]_ , \new_[31926]_ ,
    \new_[31927]_ , \new_[31928]_ , \new_[31932]_ , \new_[31933]_ ,
    \new_[31937]_ , \new_[31938]_ , \new_[31939]_ , \new_[31943]_ ,
    \new_[31944]_ , \new_[31948]_ , \new_[31949]_ , \new_[31950]_ ,
    \new_[31954]_ , \new_[31955]_ , \new_[31959]_ , \new_[31960]_ ,
    \new_[31961]_ , \new_[31965]_ , \new_[31966]_ , \new_[31970]_ ,
    \new_[31971]_ , \new_[31972]_ , \new_[31976]_ , \new_[31977]_ ,
    \new_[31981]_ , \new_[31982]_ , \new_[31983]_ , \new_[31987]_ ,
    \new_[31988]_ , \new_[31992]_ , \new_[31993]_ , \new_[31994]_ ,
    \new_[31998]_ , \new_[31999]_ , \new_[32003]_ , \new_[32004]_ ,
    \new_[32005]_ , \new_[32009]_ , \new_[32010]_ , \new_[32014]_ ,
    \new_[32015]_ , \new_[32016]_ , \new_[32020]_ , \new_[32021]_ ,
    \new_[32025]_ , \new_[32026]_ , \new_[32027]_ , \new_[32031]_ ,
    \new_[32032]_ , \new_[32036]_ , \new_[32037]_ , \new_[32038]_ ,
    \new_[32042]_ , \new_[32043]_ , \new_[32047]_ , \new_[32048]_ ,
    \new_[32049]_ , \new_[32053]_ , \new_[32054]_ , \new_[32058]_ ,
    \new_[32059]_ , \new_[32060]_ , \new_[32064]_ , \new_[32065]_ ,
    \new_[32069]_ , \new_[32070]_ , \new_[32071]_ , \new_[32075]_ ,
    \new_[32076]_ , \new_[32080]_ , \new_[32081]_ , \new_[32082]_ ,
    \new_[32086]_ , \new_[32087]_ , \new_[32091]_ , \new_[32092]_ ,
    \new_[32093]_ , \new_[32097]_ , \new_[32098]_ , \new_[32102]_ ,
    \new_[32103]_ , \new_[32104]_ , \new_[32108]_ , \new_[32109]_ ,
    \new_[32113]_ , \new_[32114]_ , \new_[32115]_ , \new_[32119]_ ,
    \new_[32120]_ , \new_[32124]_ , \new_[32125]_ , \new_[32126]_ ,
    \new_[32130]_ , \new_[32131]_ , \new_[32135]_ , \new_[32136]_ ,
    \new_[32137]_ , \new_[32141]_ , \new_[32142]_ , \new_[32146]_ ,
    \new_[32147]_ , \new_[32148]_ , \new_[32152]_ , \new_[32153]_ ,
    \new_[32157]_ , \new_[32158]_ , \new_[32159]_ , \new_[32163]_ ,
    \new_[32164]_ , \new_[32168]_ , \new_[32169]_ , \new_[32170]_ ,
    \new_[32174]_ , \new_[32175]_ , \new_[32179]_ , \new_[32180]_ ,
    \new_[32181]_ , \new_[32185]_ , \new_[32186]_ , \new_[32190]_ ,
    \new_[32191]_ , \new_[32192]_ , \new_[32196]_ , \new_[32197]_ ,
    \new_[32201]_ , \new_[32202]_ , \new_[32203]_ , \new_[32207]_ ,
    \new_[32208]_ , \new_[32212]_ , \new_[32213]_ , \new_[32214]_ ,
    \new_[32218]_ , \new_[32219]_ , \new_[32223]_ , \new_[32224]_ ,
    \new_[32225]_ , \new_[32229]_ , \new_[32230]_ , \new_[32234]_ ,
    \new_[32235]_ , \new_[32236]_ , \new_[32240]_ , \new_[32241]_ ,
    \new_[32245]_ , \new_[32246]_ , \new_[32247]_ , \new_[32251]_ ,
    \new_[32252]_ , \new_[32256]_ , \new_[32257]_ , \new_[32258]_ ,
    \new_[32262]_ , \new_[32263]_ , \new_[32267]_ , \new_[32268]_ ,
    \new_[32269]_ , \new_[32273]_ , \new_[32274]_ , \new_[32278]_ ,
    \new_[32279]_ , \new_[32280]_ , \new_[32284]_ , \new_[32285]_ ,
    \new_[32289]_ , \new_[32290]_ , \new_[32291]_ , \new_[32295]_ ,
    \new_[32296]_ , \new_[32300]_ , \new_[32301]_ , \new_[32302]_ ,
    \new_[32306]_ , \new_[32307]_ , \new_[32311]_ , \new_[32312]_ ,
    \new_[32313]_ , \new_[32317]_ , \new_[32318]_ , \new_[32322]_ ,
    \new_[32323]_ , \new_[32324]_ , \new_[32328]_ , \new_[32329]_ ,
    \new_[32333]_ , \new_[32334]_ , \new_[32335]_ , \new_[32339]_ ,
    \new_[32340]_ , \new_[32344]_ , \new_[32345]_ , \new_[32346]_ ,
    \new_[32350]_ , \new_[32351]_ , \new_[32355]_ , \new_[32356]_ ,
    \new_[32357]_ , \new_[32361]_ , \new_[32362]_ , \new_[32366]_ ,
    \new_[32367]_ , \new_[32368]_ , \new_[32372]_ , \new_[32373]_ ,
    \new_[32377]_ , \new_[32378]_ , \new_[32379]_ , \new_[32383]_ ,
    \new_[32384]_ , \new_[32388]_ , \new_[32389]_ , \new_[32390]_ ,
    \new_[32394]_ , \new_[32395]_ , \new_[32399]_ , \new_[32400]_ ,
    \new_[32401]_ , \new_[32405]_ , \new_[32406]_ , \new_[32410]_ ,
    \new_[32411]_ , \new_[32412]_ , \new_[32416]_ , \new_[32417]_ ,
    \new_[32421]_ , \new_[32422]_ , \new_[32423]_ , \new_[32427]_ ,
    \new_[32428]_ , \new_[32432]_ , \new_[32433]_ , \new_[32434]_ ,
    \new_[32438]_ , \new_[32439]_ , \new_[32443]_ , \new_[32444]_ ,
    \new_[32445]_ , \new_[32449]_ , \new_[32450]_ , \new_[32454]_ ,
    \new_[32455]_ , \new_[32456]_ , \new_[32460]_ , \new_[32461]_ ,
    \new_[32465]_ , \new_[32466]_ , \new_[32467]_ , \new_[32471]_ ,
    \new_[32472]_ , \new_[32476]_ , \new_[32477]_ , \new_[32478]_ ,
    \new_[32482]_ , \new_[32483]_ , \new_[32487]_ , \new_[32488]_ ,
    \new_[32489]_ , \new_[32493]_ , \new_[32494]_ , \new_[32498]_ ,
    \new_[32499]_ , \new_[32500]_ , \new_[32504]_ , \new_[32505]_ ,
    \new_[32509]_ , \new_[32510]_ , \new_[32511]_ , \new_[32515]_ ,
    \new_[32516]_ , \new_[32520]_ , \new_[32521]_ , \new_[32522]_ ,
    \new_[32526]_ , \new_[32527]_ , \new_[32531]_ , \new_[32532]_ ,
    \new_[32533]_ , \new_[32537]_ , \new_[32538]_ , \new_[32542]_ ,
    \new_[32543]_ , \new_[32544]_ , \new_[32548]_ , \new_[32549]_ ,
    \new_[32553]_ , \new_[32554]_ , \new_[32555]_ , \new_[32559]_ ,
    \new_[32560]_ , \new_[32564]_ , \new_[32565]_ , \new_[32566]_ ,
    \new_[32570]_ , \new_[32571]_ , \new_[32575]_ , \new_[32576]_ ,
    \new_[32577]_ , \new_[32581]_ , \new_[32582]_ , \new_[32586]_ ,
    \new_[32587]_ , \new_[32588]_ , \new_[32592]_ , \new_[32593]_ ,
    \new_[32597]_ , \new_[32598]_ , \new_[32599]_ , \new_[32603]_ ,
    \new_[32604]_ , \new_[32608]_ , \new_[32609]_ , \new_[32610]_ ,
    \new_[32614]_ , \new_[32615]_ , \new_[32619]_ , \new_[32620]_ ,
    \new_[32621]_ , \new_[32625]_ , \new_[32626]_ , \new_[32630]_ ,
    \new_[32631]_ , \new_[32632]_ , \new_[32636]_ , \new_[32637]_ ,
    \new_[32641]_ , \new_[32642]_ , \new_[32643]_ , \new_[32647]_ ,
    \new_[32648]_ , \new_[32652]_ , \new_[32653]_ , \new_[32654]_ ,
    \new_[32658]_ , \new_[32659]_ , \new_[32663]_ , \new_[32664]_ ,
    \new_[32665]_ , \new_[32669]_ , \new_[32670]_ , \new_[32674]_ ,
    \new_[32675]_ , \new_[32676]_ , \new_[32680]_ , \new_[32681]_ ,
    \new_[32685]_ , \new_[32686]_ , \new_[32687]_ , \new_[32691]_ ,
    \new_[32692]_ , \new_[32696]_ , \new_[32697]_ , \new_[32698]_ ,
    \new_[32702]_ , \new_[32703]_ , \new_[32707]_ , \new_[32708]_ ,
    \new_[32709]_ , \new_[32713]_ , \new_[32714]_ , \new_[32718]_ ,
    \new_[32719]_ , \new_[32720]_ , \new_[32724]_ , \new_[32725]_ ,
    \new_[32729]_ , \new_[32730]_ , \new_[32731]_ , \new_[32735]_ ,
    \new_[32736]_ , \new_[32740]_ , \new_[32741]_ , \new_[32742]_ ,
    \new_[32746]_ , \new_[32747]_ , \new_[32751]_ , \new_[32752]_ ,
    \new_[32753]_ , \new_[32757]_ , \new_[32758]_ , \new_[32762]_ ,
    \new_[32763]_ , \new_[32764]_ , \new_[32768]_ , \new_[32769]_ ,
    \new_[32773]_ , \new_[32774]_ , \new_[32775]_ , \new_[32779]_ ,
    \new_[32780]_ , \new_[32784]_ , \new_[32785]_ , \new_[32786]_ ,
    \new_[32790]_ , \new_[32791]_ , \new_[32795]_ , \new_[32796]_ ,
    \new_[32797]_ , \new_[32801]_ , \new_[32802]_ , \new_[32806]_ ,
    \new_[32807]_ , \new_[32808]_ , \new_[32812]_ , \new_[32813]_ ,
    \new_[32817]_ , \new_[32818]_ , \new_[32819]_ , \new_[32823]_ ,
    \new_[32824]_ , \new_[32828]_ , \new_[32829]_ , \new_[32830]_ ,
    \new_[32834]_ , \new_[32835]_ , \new_[32839]_ , \new_[32840]_ ,
    \new_[32841]_ , \new_[32845]_ , \new_[32846]_ , \new_[32850]_ ,
    \new_[32851]_ , \new_[32852]_ , \new_[32856]_ , \new_[32857]_ ,
    \new_[32861]_ , \new_[32862]_ , \new_[32863]_ , \new_[32867]_ ,
    \new_[32868]_ , \new_[32872]_ , \new_[32873]_ , \new_[32874]_ ,
    \new_[32878]_ , \new_[32879]_ , \new_[32883]_ , \new_[32884]_ ,
    \new_[32885]_ , \new_[32889]_ , \new_[32890]_ , \new_[32894]_ ,
    \new_[32895]_ , \new_[32896]_ , \new_[32900]_ , \new_[32901]_ ,
    \new_[32905]_ , \new_[32906]_ , \new_[32907]_ , \new_[32911]_ ,
    \new_[32912]_ , \new_[32916]_ , \new_[32917]_ , \new_[32918]_ ,
    \new_[32922]_ , \new_[32923]_ , \new_[32927]_ , \new_[32928]_ ,
    \new_[32929]_ , \new_[32933]_ , \new_[32934]_ , \new_[32938]_ ,
    \new_[32939]_ , \new_[32940]_ , \new_[32944]_ , \new_[32945]_ ,
    \new_[32949]_ , \new_[32950]_ , \new_[32951]_ , \new_[32955]_ ,
    \new_[32956]_ , \new_[32960]_ , \new_[32961]_ , \new_[32962]_ ,
    \new_[32966]_ , \new_[32967]_ , \new_[32971]_ , \new_[32972]_ ,
    \new_[32973]_ , \new_[32977]_ , \new_[32978]_ , \new_[32982]_ ,
    \new_[32983]_ , \new_[32984]_ , \new_[32988]_ , \new_[32989]_ ,
    \new_[32993]_ , \new_[32994]_ , \new_[32995]_ , \new_[32999]_ ,
    \new_[33000]_ , \new_[33004]_ , \new_[33005]_ , \new_[33006]_ ,
    \new_[33010]_ , \new_[33011]_ , \new_[33015]_ , \new_[33016]_ ,
    \new_[33017]_ , \new_[33021]_ , \new_[33022]_ , \new_[33026]_ ,
    \new_[33027]_ , \new_[33028]_ , \new_[33032]_ , \new_[33033]_ ,
    \new_[33037]_ , \new_[33038]_ , \new_[33039]_ , \new_[33043]_ ,
    \new_[33044]_ , \new_[33048]_ , \new_[33049]_ , \new_[33050]_ ,
    \new_[33054]_ , \new_[33055]_ , \new_[33059]_ , \new_[33060]_ ,
    \new_[33061]_ , \new_[33065]_ , \new_[33066]_ , \new_[33070]_ ,
    \new_[33071]_ , \new_[33072]_ , \new_[33076]_ , \new_[33077]_ ,
    \new_[33081]_ , \new_[33082]_ , \new_[33083]_ , \new_[33087]_ ,
    \new_[33088]_ , \new_[33092]_ , \new_[33093]_ , \new_[33094]_ ,
    \new_[33098]_ , \new_[33099]_ , \new_[33103]_ , \new_[33104]_ ,
    \new_[33105]_ , \new_[33109]_ , \new_[33110]_ , \new_[33114]_ ,
    \new_[33115]_ , \new_[33116]_ , \new_[33120]_ , \new_[33121]_ ,
    \new_[33125]_ , \new_[33126]_ , \new_[33127]_ , \new_[33131]_ ,
    \new_[33132]_ , \new_[33136]_ , \new_[33137]_ , \new_[33138]_ ,
    \new_[33142]_ , \new_[33143]_ , \new_[33147]_ , \new_[33148]_ ,
    \new_[33149]_ , \new_[33153]_ , \new_[33154]_ , \new_[33158]_ ,
    \new_[33159]_ , \new_[33160]_ , \new_[33164]_ , \new_[33165]_ ,
    \new_[33169]_ , \new_[33170]_ , \new_[33171]_ , \new_[33175]_ ,
    \new_[33176]_ , \new_[33180]_ , \new_[33181]_ , \new_[33182]_ ,
    \new_[33186]_ , \new_[33187]_ , \new_[33191]_ , \new_[33192]_ ,
    \new_[33193]_ , \new_[33197]_ , \new_[33198]_ , \new_[33202]_ ,
    \new_[33203]_ , \new_[33204]_ , \new_[33208]_ , \new_[33209]_ ,
    \new_[33213]_ , \new_[33214]_ , \new_[33215]_ , \new_[33219]_ ,
    \new_[33220]_ , \new_[33224]_ , \new_[33225]_ , \new_[33226]_ ,
    \new_[33230]_ , \new_[33231]_ , \new_[33235]_ , \new_[33236]_ ,
    \new_[33237]_ , \new_[33241]_ , \new_[33242]_ , \new_[33246]_ ,
    \new_[33247]_ , \new_[33248]_ , \new_[33252]_ , \new_[33253]_ ,
    \new_[33257]_ , \new_[33258]_ , \new_[33259]_ , \new_[33263]_ ,
    \new_[33264]_ , \new_[33268]_ , \new_[33269]_ , \new_[33270]_ ,
    \new_[33274]_ , \new_[33275]_ , \new_[33279]_ , \new_[33280]_ ,
    \new_[33281]_ , \new_[33285]_ , \new_[33286]_ , \new_[33290]_ ,
    \new_[33291]_ , \new_[33292]_ , \new_[33296]_ , \new_[33297]_ ,
    \new_[33301]_ , \new_[33302]_ , \new_[33303]_ , \new_[33307]_ ,
    \new_[33308]_ , \new_[33312]_ , \new_[33313]_ , \new_[33314]_ ,
    \new_[33318]_ , \new_[33319]_ , \new_[33323]_ , \new_[33324]_ ,
    \new_[33325]_ , \new_[33329]_ , \new_[33330]_ , \new_[33334]_ ,
    \new_[33335]_ , \new_[33336]_ , \new_[33340]_ , \new_[33341]_ ,
    \new_[33345]_ , \new_[33346]_ , \new_[33347]_ , \new_[33351]_ ,
    \new_[33352]_ , \new_[33356]_ , \new_[33357]_ , \new_[33358]_ ,
    \new_[33362]_ , \new_[33363]_ , \new_[33367]_ , \new_[33368]_ ,
    \new_[33369]_ , \new_[33373]_ , \new_[33374]_ , \new_[33378]_ ,
    \new_[33379]_ , \new_[33380]_ , \new_[33384]_ , \new_[33385]_ ,
    \new_[33389]_ , \new_[33390]_ , \new_[33391]_ , \new_[33395]_ ,
    \new_[33396]_ , \new_[33400]_ , \new_[33401]_ , \new_[33402]_ ,
    \new_[33406]_ , \new_[33407]_ , \new_[33411]_ , \new_[33412]_ ,
    \new_[33413]_ , \new_[33417]_ , \new_[33418]_ , \new_[33422]_ ,
    \new_[33423]_ , \new_[33424]_ , \new_[33428]_ , \new_[33429]_ ,
    \new_[33433]_ , \new_[33434]_ , \new_[33435]_ , \new_[33439]_ ,
    \new_[33440]_ , \new_[33444]_ , \new_[33445]_ , \new_[33446]_ ,
    \new_[33450]_ , \new_[33451]_ , \new_[33455]_ , \new_[33456]_ ,
    \new_[33457]_ , \new_[33461]_ , \new_[33462]_ , \new_[33466]_ ,
    \new_[33467]_ , \new_[33468]_ , \new_[33472]_ , \new_[33473]_ ,
    \new_[33477]_ , \new_[33478]_ , \new_[33479]_ , \new_[33483]_ ,
    \new_[33484]_ , \new_[33488]_ , \new_[33489]_ , \new_[33490]_ ,
    \new_[33494]_ , \new_[33495]_ , \new_[33499]_ , \new_[33500]_ ,
    \new_[33501]_ , \new_[33505]_ , \new_[33506]_ , \new_[33510]_ ,
    \new_[33511]_ , \new_[33512]_ , \new_[33516]_ , \new_[33517]_ ,
    \new_[33521]_ , \new_[33522]_ , \new_[33523]_ , \new_[33527]_ ,
    \new_[33528]_ , \new_[33532]_ , \new_[33533]_ , \new_[33534]_ ,
    \new_[33538]_ , \new_[33539]_ , \new_[33543]_ , \new_[33544]_ ,
    \new_[33545]_ , \new_[33549]_ , \new_[33550]_ , \new_[33554]_ ,
    \new_[33555]_ , \new_[33556]_ , \new_[33560]_ , \new_[33561]_ ,
    \new_[33565]_ , \new_[33566]_ , \new_[33567]_ , \new_[33571]_ ,
    \new_[33572]_ , \new_[33576]_ , \new_[33577]_ , \new_[33578]_ ,
    \new_[33582]_ , \new_[33583]_ , \new_[33587]_ , \new_[33588]_ ,
    \new_[33589]_ , \new_[33593]_ , \new_[33594]_ , \new_[33598]_ ,
    \new_[33599]_ , \new_[33600]_ , \new_[33604]_ , \new_[33605]_ ,
    \new_[33609]_ , \new_[33610]_ , \new_[33611]_ , \new_[33615]_ ,
    \new_[33616]_ , \new_[33620]_ , \new_[33621]_ , \new_[33622]_ ,
    \new_[33626]_ , \new_[33627]_ , \new_[33631]_ , \new_[33632]_ ,
    \new_[33633]_ , \new_[33637]_ , \new_[33638]_ , \new_[33642]_ ,
    \new_[33643]_ , \new_[33644]_ , \new_[33648]_ , \new_[33649]_ ,
    \new_[33653]_ , \new_[33654]_ , \new_[33655]_ , \new_[33659]_ ,
    \new_[33660]_ , \new_[33664]_ , \new_[33665]_ , \new_[33666]_ ,
    \new_[33670]_ , \new_[33671]_ , \new_[33675]_ , \new_[33676]_ ,
    \new_[33677]_ , \new_[33681]_ , \new_[33682]_ , \new_[33686]_ ,
    \new_[33687]_ , \new_[33688]_ , \new_[33692]_ , \new_[33693]_ ,
    \new_[33697]_ , \new_[33698]_ , \new_[33699]_ , \new_[33703]_ ,
    \new_[33704]_ , \new_[33708]_ , \new_[33709]_ , \new_[33710]_ ,
    \new_[33714]_ , \new_[33715]_ , \new_[33719]_ , \new_[33720]_ ,
    \new_[33721]_ , \new_[33725]_ , \new_[33726]_ , \new_[33730]_ ,
    \new_[33731]_ , \new_[33732]_ , \new_[33736]_ , \new_[33737]_ ,
    \new_[33741]_ , \new_[33742]_ , \new_[33743]_ , \new_[33747]_ ,
    \new_[33748]_ , \new_[33752]_ , \new_[33753]_ , \new_[33754]_ ,
    \new_[33758]_ , \new_[33759]_ , \new_[33763]_ , \new_[33764]_ ,
    \new_[33765]_ , \new_[33769]_ , \new_[33770]_ , \new_[33774]_ ,
    \new_[33775]_ , \new_[33776]_ , \new_[33780]_ , \new_[33781]_ ,
    \new_[33785]_ , \new_[33786]_ , \new_[33787]_ , \new_[33791]_ ,
    \new_[33792]_ , \new_[33796]_ , \new_[33797]_ , \new_[33798]_ ,
    \new_[33802]_ , \new_[33803]_ , \new_[33807]_ , \new_[33808]_ ,
    \new_[33809]_ , \new_[33813]_ , \new_[33814]_ , \new_[33818]_ ,
    \new_[33819]_ , \new_[33820]_ , \new_[33824]_ , \new_[33825]_ ,
    \new_[33829]_ , \new_[33830]_ , \new_[33831]_ , \new_[33835]_ ,
    \new_[33836]_ , \new_[33840]_ , \new_[33841]_ , \new_[33842]_ ,
    \new_[33846]_ , \new_[33847]_ , \new_[33851]_ , \new_[33852]_ ,
    \new_[33853]_ , \new_[33857]_ , \new_[33858]_ , \new_[33862]_ ,
    \new_[33863]_ , \new_[33864]_ , \new_[33868]_ , \new_[33869]_ ,
    \new_[33873]_ , \new_[33874]_ , \new_[33875]_ , \new_[33879]_ ,
    \new_[33880]_ , \new_[33884]_ , \new_[33885]_ , \new_[33886]_ ,
    \new_[33890]_ , \new_[33891]_ , \new_[33895]_ , \new_[33896]_ ,
    \new_[33897]_ , \new_[33901]_ , \new_[33902]_ , \new_[33906]_ ,
    \new_[33907]_ , \new_[33908]_ , \new_[33912]_ , \new_[33913]_ ,
    \new_[33917]_ , \new_[33918]_ , \new_[33919]_ , \new_[33923]_ ,
    \new_[33924]_ , \new_[33928]_ , \new_[33929]_ , \new_[33930]_ ,
    \new_[33934]_ , \new_[33935]_ , \new_[33939]_ , \new_[33940]_ ,
    \new_[33941]_ , \new_[33945]_ , \new_[33946]_ , \new_[33950]_ ,
    \new_[33951]_ , \new_[33952]_ , \new_[33956]_ , \new_[33957]_ ,
    \new_[33961]_ , \new_[33962]_ , \new_[33963]_ , \new_[33967]_ ,
    \new_[33968]_ , \new_[33972]_ , \new_[33973]_ , \new_[33974]_ ,
    \new_[33978]_ , \new_[33979]_ , \new_[33983]_ , \new_[33984]_ ,
    \new_[33985]_ , \new_[33989]_ , \new_[33990]_ , \new_[33994]_ ,
    \new_[33995]_ , \new_[33996]_ , \new_[34000]_ , \new_[34001]_ ,
    \new_[34005]_ , \new_[34006]_ , \new_[34007]_ , \new_[34011]_ ,
    \new_[34012]_ , \new_[34016]_ , \new_[34017]_ , \new_[34018]_ ,
    \new_[34022]_ , \new_[34023]_ , \new_[34027]_ , \new_[34028]_ ,
    \new_[34029]_ , \new_[34033]_ , \new_[34034]_ , \new_[34038]_ ,
    \new_[34039]_ , \new_[34040]_ , \new_[34044]_ , \new_[34045]_ ,
    \new_[34049]_ , \new_[34050]_ , \new_[34051]_ , \new_[34055]_ ,
    \new_[34056]_ , \new_[34060]_ , \new_[34061]_ , \new_[34062]_ ,
    \new_[34066]_ , \new_[34067]_ , \new_[34071]_ , \new_[34072]_ ,
    \new_[34073]_ , \new_[34077]_ , \new_[34078]_ , \new_[34082]_ ,
    \new_[34083]_ , \new_[34084]_ , \new_[34088]_ , \new_[34089]_ ,
    \new_[34093]_ , \new_[34094]_ , \new_[34095]_ , \new_[34099]_ ,
    \new_[34100]_ , \new_[34104]_ , \new_[34105]_ , \new_[34106]_ ,
    \new_[34110]_ , \new_[34111]_ , \new_[34115]_ , \new_[34116]_ ,
    \new_[34117]_ , \new_[34121]_ , \new_[34122]_ , \new_[34126]_ ,
    \new_[34127]_ , \new_[34128]_ , \new_[34132]_ , \new_[34133]_ ,
    \new_[34137]_ , \new_[34138]_ , \new_[34139]_ , \new_[34143]_ ,
    \new_[34144]_ , \new_[34148]_ , \new_[34149]_ , \new_[34150]_ ,
    \new_[34154]_ , \new_[34155]_ , \new_[34159]_ , \new_[34160]_ ,
    \new_[34161]_ , \new_[34165]_ , \new_[34166]_ , \new_[34170]_ ,
    \new_[34171]_ , \new_[34172]_ , \new_[34176]_ , \new_[34177]_ ,
    \new_[34181]_ , \new_[34182]_ , \new_[34183]_ , \new_[34187]_ ,
    \new_[34188]_ , \new_[34192]_ , \new_[34193]_ , \new_[34194]_ ,
    \new_[34198]_ , \new_[34199]_ , \new_[34203]_ , \new_[34204]_ ,
    \new_[34205]_ , \new_[34209]_ , \new_[34210]_ , \new_[34214]_ ,
    \new_[34215]_ , \new_[34216]_ , \new_[34220]_ , \new_[34221]_ ,
    \new_[34225]_ , \new_[34226]_ , \new_[34227]_ , \new_[34231]_ ,
    \new_[34232]_ , \new_[34236]_ , \new_[34237]_ , \new_[34238]_ ,
    \new_[34242]_ , \new_[34243]_ , \new_[34247]_ , \new_[34248]_ ,
    \new_[34249]_ , \new_[34253]_ , \new_[34254]_ , \new_[34258]_ ,
    \new_[34259]_ , \new_[34260]_ , \new_[34264]_ , \new_[34265]_ ,
    \new_[34269]_ , \new_[34270]_ , \new_[34271]_ , \new_[34275]_ ,
    \new_[34276]_ , \new_[34280]_ , \new_[34281]_ , \new_[34282]_ ,
    \new_[34286]_ , \new_[34287]_ , \new_[34291]_ , \new_[34292]_ ,
    \new_[34293]_ , \new_[34297]_ , \new_[34298]_ , \new_[34302]_ ,
    \new_[34303]_ , \new_[34304]_ , \new_[34308]_ , \new_[34309]_ ,
    \new_[34313]_ , \new_[34314]_ , \new_[34315]_ , \new_[34319]_ ,
    \new_[34320]_ , \new_[34324]_ , \new_[34325]_ , \new_[34326]_ ,
    \new_[34330]_ , \new_[34331]_ , \new_[34335]_ , \new_[34336]_ ,
    \new_[34337]_ , \new_[34341]_ , \new_[34342]_ , \new_[34346]_ ,
    \new_[34347]_ , \new_[34348]_ , \new_[34352]_ , \new_[34353]_ ,
    \new_[34357]_ , \new_[34358]_ , \new_[34359]_ , \new_[34363]_ ,
    \new_[34364]_ , \new_[34368]_ , \new_[34369]_ , \new_[34370]_ ,
    \new_[34374]_ , \new_[34375]_ , \new_[34379]_ , \new_[34380]_ ,
    \new_[34381]_ , \new_[34385]_ , \new_[34386]_ , \new_[34390]_ ,
    \new_[34391]_ , \new_[34392]_ , \new_[34396]_ , \new_[34397]_ ,
    \new_[34401]_ , \new_[34402]_ , \new_[34403]_ , \new_[34407]_ ,
    \new_[34408]_ , \new_[34412]_ , \new_[34413]_ , \new_[34414]_ ,
    \new_[34418]_ , \new_[34419]_ , \new_[34423]_ , \new_[34424]_ ,
    \new_[34425]_ , \new_[34429]_ , \new_[34430]_ , \new_[34434]_ ,
    \new_[34435]_ , \new_[34436]_ , \new_[34440]_ , \new_[34441]_ ,
    \new_[34445]_ , \new_[34446]_ , \new_[34447]_ , \new_[34451]_ ,
    \new_[34452]_ , \new_[34456]_ , \new_[34457]_ , \new_[34458]_ ,
    \new_[34462]_ , \new_[34463]_ , \new_[34467]_ , \new_[34468]_ ,
    \new_[34469]_ , \new_[34473]_ , \new_[34474]_ , \new_[34478]_ ,
    \new_[34479]_ , \new_[34480]_ , \new_[34484]_ , \new_[34485]_ ,
    \new_[34489]_ , \new_[34490]_ , \new_[34491]_ , \new_[34495]_ ,
    \new_[34496]_ , \new_[34500]_ , \new_[34501]_ , \new_[34502]_ ,
    \new_[34506]_ , \new_[34507]_ , \new_[34511]_ , \new_[34512]_ ,
    \new_[34513]_ , \new_[34517]_ , \new_[34518]_ , \new_[34522]_ ,
    \new_[34523]_ , \new_[34524]_ , \new_[34528]_ , \new_[34529]_ ,
    \new_[34533]_ , \new_[34534]_ , \new_[34535]_ , \new_[34539]_ ,
    \new_[34540]_ , \new_[34544]_ , \new_[34545]_ , \new_[34546]_ ,
    \new_[34550]_ , \new_[34551]_ , \new_[34555]_ , \new_[34556]_ ,
    \new_[34557]_ , \new_[34561]_ , \new_[34562]_ , \new_[34566]_ ,
    \new_[34567]_ , \new_[34568]_ , \new_[34572]_ , \new_[34573]_ ,
    \new_[34577]_ , \new_[34578]_ , \new_[34579]_ , \new_[34583]_ ,
    \new_[34584]_ , \new_[34588]_ , \new_[34589]_ , \new_[34590]_ ,
    \new_[34594]_ , \new_[34595]_ , \new_[34599]_ , \new_[34600]_ ,
    \new_[34601]_ , \new_[34605]_ , \new_[34606]_ , \new_[34610]_ ,
    \new_[34611]_ , \new_[34612]_ , \new_[34616]_ , \new_[34617]_ ,
    \new_[34621]_ , \new_[34622]_ , \new_[34623]_ , \new_[34627]_ ,
    \new_[34628]_ , \new_[34632]_ , \new_[34633]_ , \new_[34634]_ ,
    \new_[34638]_ , \new_[34639]_ , \new_[34643]_ , \new_[34644]_ ,
    \new_[34645]_ , \new_[34649]_ , \new_[34650]_ , \new_[34654]_ ,
    \new_[34655]_ , \new_[34656]_ , \new_[34660]_ , \new_[34661]_ ,
    \new_[34665]_ , \new_[34666]_ , \new_[34667]_ , \new_[34671]_ ,
    \new_[34672]_ , \new_[34676]_ , \new_[34677]_ , \new_[34678]_ ,
    \new_[34682]_ , \new_[34683]_ , \new_[34687]_ , \new_[34688]_ ,
    \new_[34689]_ , \new_[34693]_ , \new_[34694]_ , \new_[34698]_ ,
    \new_[34699]_ , \new_[34700]_ , \new_[34704]_ , \new_[34705]_ ,
    \new_[34709]_ , \new_[34710]_ , \new_[34711]_ , \new_[34715]_ ,
    \new_[34716]_ , \new_[34720]_ , \new_[34721]_ , \new_[34722]_ ,
    \new_[34726]_ , \new_[34727]_ , \new_[34731]_ , \new_[34732]_ ,
    \new_[34733]_ , \new_[34737]_ , \new_[34738]_ , \new_[34742]_ ,
    \new_[34743]_ , \new_[34744]_ , \new_[34748]_ , \new_[34749]_ ,
    \new_[34753]_ , \new_[34754]_ , \new_[34755]_ , \new_[34759]_ ,
    \new_[34760]_ , \new_[34764]_ , \new_[34765]_ , \new_[34766]_ ,
    \new_[34770]_ , \new_[34771]_ , \new_[34775]_ , \new_[34776]_ ,
    \new_[34777]_ , \new_[34781]_ , \new_[34782]_ , \new_[34786]_ ,
    \new_[34787]_ , \new_[34788]_ , \new_[34792]_ , \new_[34793]_ ,
    \new_[34797]_ , \new_[34798]_ , \new_[34799]_ , \new_[34803]_ ,
    \new_[34804]_ , \new_[34808]_ , \new_[34809]_ , \new_[34810]_ ,
    \new_[34814]_ , \new_[34815]_ , \new_[34819]_ , \new_[34820]_ ,
    \new_[34821]_ , \new_[34825]_ , \new_[34826]_ , \new_[34830]_ ,
    \new_[34831]_ , \new_[34832]_ , \new_[34836]_ , \new_[34837]_ ,
    \new_[34841]_ , \new_[34842]_ , \new_[34843]_ , \new_[34847]_ ,
    \new_[34848]_ , \new_[34852]_ , \new_[34853]_ , \new_[34854]_ ,
    \new_[34858]_ , \new_[34859]_ , \new_[34863]_ , \new_[34864]_ ,
    \new_[34865]_ , \new_[34869]_ , \new_[34870]_ , \new_[34874]_ ,
    \new_[34875]_ , \new_[34876]_ , \new_[34880]_ , \new_[34881]_ ,
    \new_[34885]_ , \new_[34886]_ , \new_[34887]_ , \new_[34891]_ ,
    \new_[34892]_ , \new_[34896]_ , \new_[34897]_ , \new_[34898]_ ,
    \new_[34902]_ , \new_[34903]_ , \new_[34907]_ , \new_[34908]_ ,
    \new_[34909]_ , \new_[34913]_ , \new_[34914]_ , \new_[34918]_ ,
    \new_[34919]_ , \new_[34920]_ , \new_[34924]_ , \new_[34925]_ ,
    \new_[34929]_ , \new_[34930]_ , \new_[34931]_ , \new_[34935]_ ,
    \new_[34936]_ , \new_[34940]_ , \new_[34941]_ , \new_[34942]_ ,
    \new_[34946]_ , \new_[34947]_ , \new_[34951]_ , \new_[34952]_ ,
    \new_[34953]_ , \new_[34957]_ , \new_[34958]_ , \new_[34962]_ ,
    \new_[34963]_ , \new_[34964]_ , \new_[34968]_ , \new_[34969]_ ,
    \new_[34973]_ , \new_[34974]_ , \new_[34975]_ , \new_[34979]_ ,
    \new_[34980]_ , \new_[34984]_ , \new_[34985]_ , \new_[34986]_ ,
    \new_[34990]_ , \new_[34991]_ , \new_[34995]_ , \new_[34996]_ ,
    \new_[34997]_ , \new_[35001]_ , \new_[35002]_ , \new_[35006]_ ,
    \new_[35007]_ , \new_[35008]_ , \new_[35012]_ , \new_[35013]_ ,
    \new_[35017]_ , \new_[35018]_ , \new_[35019]_ , \new_[35023]_ ,
    \new_[35024]_ , \new_[35028]_ , \new_[35029]_ , \new_[35030]_ ,
    \new_[35034]_ , \new_[35035]_ , \new_[35039]_ , \new_[35040]_ ,
    \new_[35041]_ , \new_[35045]_ , \new_[35046]_ , \new_[35050]_ ,
    \new_[35051]_ , \new_[35052]_ , \new_[35056]_ , \new_[35057]_ ,
    \new_[35061]_ , \new_[35062]_ , \new_[35063]_ , \new_[35067]_ ,
    \new_[35068]_ , \new_[35072]_ , \new_[35073]_ , \new_[35074]_ ,
    \new_[35078]_ , \new_[35079]_ , \new_[35083]_ , \new_[35084]_ ,
    \new_[35085]_ , \new_[35089]_ , \new_[35090]_ , \new_[35094]_ ,
    \new_[35095]_ , \new_[35096]_ , \new_[35100]_ , \new_[35101]_ ,
    \new_[35105]_ , \new_[35106]_ , \new_[35107]_ , \new_[35111]_ ,
    \new_[35112]_ , \new_[35116]_ , \new_[35117]_ , \new_[35118]_ ,
    \new_[35122]_ , \new_[35123]_ , \new_[35127]_ , \new_[35128]_ ,
    \new_[35129]_ , \new_[35133]_ , \new_[35134]_ , \new_[35138]_ ,
    \new_[35139]_ , \new_[35140]_ , \new_[35144]_ , \new_[35145]_ ,
    \new_[35149]_ , \new_[35150]_ , \new_[35151]_ , \new_[35155]_ ,
    \new_[35156]_ , \new_[35160]_ , \new_[35161]_ , \new_[35162]_ ,
    \new_[35166]_ , \new_[35167]_ , \new_[35171]_ , \new_[35172]_ ,
    \new_[35173]_ , \new_[35177]_ , \new_[35178]_ , \new_[35182]_ ,
    \new_[35183]_ , \new_[35184]_ , \new_[35188]_ , \new_[35189]_ ,
    \new_[35193]_ , \new_[35194]_ , \new_[35195]_ , \new_[35199]_ ,
    \new_[35200]_ , \new_[35204]_ , \new_[35205]_ , \new_[35206]_ ,
    \new_[35210]_ , \new_[35211]_ , \new_[35215]_ , \new_[35216]_ ,
    \new_[35217]_ , \new_[35221]_ , \new_[35222]_ , \new_[35226]_ ,
    \new_[35227]_ , \new_[35228]_ , \new_[35232]_ , \new_[35233]_ ,
    \new_[35237]_ , \new_[35238]_ , \new_[35239]_ , \new_[35243]_ ,
    \new_[35244]_ , \new_[35248]_ , \new_[35249]_ , \new_[35250]_ ,
    \new_[35254]_ , \new_[35255]_ , \new_[35259]_ , \new_[35260]_ ,
    \new_[35261]_ , \new_[35265]_ , \new_[35266]_ , \new_[35270]_ ,
    \new_[35271]_ , \new_[35272]_ , \new_[35276]_ , \new_[35277]_ ,
    \new_[35281]_ , \new_[35282]_ , \new_[35283]_ , \new_[35287]_ ,
    \new_[35288]_ , \new_[35292]_ , \new_[35293]_ , \new_[35294]_ ,
    \new_[35298]_ , \new_[35299]_ , \new_[35303]_ , \new_[35304]_ ,
    \new_[35305]_ , \new_[35309]_ , \new_[35310]_ , \new_[35314]_ ,
    \new_[35315]_ , \new_[35316]_ , \new_[35320]_ , \new_[35321]_ ,
    \new_[35325]_ , \new_[35326]_ , \new_[35327]_ , \new_[35331]_ ,
    \new_[35332]_ , \new_[35336]_ , \new_[35337]_ , \new_[35338]_ ,
    \new_[35342]_ , \new_[35343]_ , \new_[35347]_ , \new_[35348]_ ,
    \new_[35349]_ , \new_[35353]_ , \new_[35354]_ , \new_[35358]_ ,
    \new_[35359]_ , \new_[35360]_ , \new_[35364]_ , \new_[35365]_ ,
    \new_[35369]_ , \new_[35370]_ , \new_[35371]_ , \new_[35375]_ ,
    \new_[35376]_ , \new_[35380]_ , \new_[35381]_ , \new_[35382]_ ,
    \new_[35386]_ , \new_[35387]_ , \new_[35391]_ , \new_[35392]_ ,
    \new_[35393]_ , \new_[35397]_ , \new_[35398]_ , \new_[35402]_ ,
    \new_[35403]_ , \new_[35404]_ , \new_[35408]_ , \new_[35409]_ ,
    \new_[35413]_ , \new_[35414]_ , \new_[35415]_ , \new_[35419]_ ,
    \new_[35420]_ , \new_[35424]_ , \new_[35425]_ , \new_[35426]_ ,
    \new_[35430]_ , \new_[35431]_ , \new_[35435]_ , \new_[35436]_ ,
    \new_[35437]_ , \new_[35441]_ , \new_[35442]_ , \new_[35446]_ ,
    \new_[35447]_ , \new_[35448]_ , \new_[35452]_ , \new_[35453]_ ,
    \new_[35457]_ , \new_[35458]_ , \new_[35459]_ , \new_[35463]_ ,
    \new_[35464]_ , \new_[35468]_ , \new_[35469]_ , \new_[35470]_ ,
    \new_[35474]_ , \new_[35475]_ , \new_[35479]_ , \new_[35480]_ ,
    \new_[35481]_ , \new_[35485]_ , \new_[35486]_ , \new_[35490]_ ,
    \new_[35491]_ , \new_[35492]_ , \new_[35496]_ , \new_[35497]_ ,
    \new_[35501]_ , \new_[35502]_ , \new_[35503]_ , \new_[35507]_ ,
    \new_[35508]_ , \new_[35512]_ , \new_[35513]_ , \new_[35514]_ ,
    \new_[35518]_ , \new_[35519]_ , \new_[35523]_ , \new_[35524]_ ,
    \new_[35525]_ , \new_[35529]_ , \new_[35530]_ , \new_[35534]_ ,
    \new_[35535]_ , \new_[35536]_ , \new_[35540]_ , \new_[35541]_ ,
    \new_[35545]_ , \new_[35546]_ , \new_[35547]_ , \new_[35551]_ ,
    \new_[35552]_ , \new_[35556]_ , \new_[35557]_ , \new_[35558]_ ,
    \new_[35562]_ , \new_[35563]_ , \new_[35567]_ , \new_[35568]_ ,
    \new_[35569]_ , \new_[35573]_ , \new_[35574]_ , \new_[35578]_ ,
    \new_[35579]_ , \new_[35580]_ , \new_[35584]_ , \new_[35585]_ ,
    \new_[35589]_ , \new_[35590]_ , \new_[35591]_ , \new_[35595]_ ,
    \new_[35596]_ , \new_[35600]_ , \new_[35601]_ , \new_[35602]_ ,
    \new_[35606]_ , \new_[35607]_ , \new_[35611]_ , \new_[35612]_ ,
    \new_[35613]_ , \new_[35617]_ , \new_[35618]_ , \new_[35622]_ ,
    \new_[35623]_ , \new_[35624]_ , \new_[35628]_ , \new_[35629]_ ,
    \new_[35633]_ , \new_[35634]_ , \new_[35635]_ , \new_[35639]_ ,
    \new_[35640]_ , \new_[35644]_ , \new_[35645]_ , \new_[35646]_ ,
    \new_[35650]_ , \new_[35651]_ , \new_[35655]_ , \new_[35656]_ ,
    \new_[35657]_ , \new_[35661]_ , \new_[35662]_ , \new_[35666]_ ,
    \new_[35667]_ , \new_[35668]_ , \new_[35672]_ , \new_[35673]_ ,
    \new_[35677]_ , \new_[35678]_ , \new_[35679]_ , \new_[35683]_ ,
    \new_[35684]_ , \new_[35688]_ , \new_[35689]_ , \new_[35690]_ ,
    \new_[35694]_ , \new_[35695]_ , \new_[35699]_ , \new_[35700]_ ,
    \new_[35701]_ , \new_[35705]_ , \new_[35706]_ , \new_[35710]_ ,
    \new_[35711]_ , \new_[35712]_ , \new_[35716]_ , \new_[35717]_ ,
    \new_[35721]_ , \new_[35722]_ , \new_[35723]_ , \new_[35727]_ ,
    \new_[35728]_ , \new_[35732]_ , \new_[35733]_ , \new_[35734]_ ,
    \new_[35738]_ , \new_[35739]_ , \new_[35743]_ , \new_[35744]_ ,
    \new_[35745]_ , \new_[35749]_ , \new_[35750]_ , \new_[35754]_ ,
    \new_[35755]_ , \new_[35756]_ , \new_[35760]_ , \new_[35761]_ ,
    \new_[35765]_ , \new_[35766]_ , \new_[35767]_ , \new_[35771]_ ,
    \new_[35772]_ , \new_[35776]_ , \new_[35777]_ , \new_[35778]_ ,
    \new_[35782]_ , \new_[35783]_ , \new_[35787]_ , \new_[35788]_ ,
    \new_[35789]_ , \new_[35793]_ , \new_[35794]_ , \new_[35798]_ ,
    \new_[35799]_ , \new_[35800]_ , \new_[35804]_ , \new_[35805]_ ,
    \new_[35809]_ , \new_[35810]_ , \new_[35811]_ , \new_[35815]_ ,
    \new_[35816]_ , \new_[35820]_ , \new_[35821]_ , \new_[35822]_ ,
    \new_[35826]_ , \new_[35827]_ , \new_[35831]_ , \new_[35832]_ ,
    \new_[35833]_ , \new_[35837]_ , \new_[35838]_ , \new_[35842]_ ,
    \new_[35843]_ , \new_[35844]_ , \new_[35848]_ , \new_[35849]_ ,
    \new_[35853]_ , \new_[35854]_ , \new_[35855]_ , \new_[35859]_ ,
    \new_[35860]_ , \new_[35864]_ , \new_[35865]_ , \new_[35866]_ ,
    \new_[35870]_ , \new_[35871]_ , \new_[35875]_ , \new_[35876]_ ,
    \new_[35877]_ , \new_[35881]_ , \new_[35882]_ , \new_[35886]_ ,
    \new_[35887]_ , \new_[35888]_ , \new_[35892]_ , \new_[35893]_ ,
    \new_[35897]_ , \new_[35898]_ , \new_[35899]_ , \new_[35903]_ ,
    \new_[35904]_ , \new_[35908]_ , \new_[35909]_ , \new_[35910]_ ,
    \new_[35914]_ , \new_[35915]_ , \new_[35919]_ , \new_[35920]_ ,
    \new_[35921]_ , \new_[35925]_ , \new_[35926]_ , \new_[35930]_ ,
    \new_[35931]_ , \new_[35932]_ , \new_[35936]_ , \new_[35937]_ ,
    \new_[35941]_ , \new_[35942]_ , \new_[35943]_ , \new_[35947]_ ,
    \new_[35948]_ , \new_[35952]_ , \new_[35953]_ , \new_[35954]_ ,
    \new_[35958]_ , \new_[35959]_ , \new_[35963]_ , \new_[35964]_ ,
    \new_[35965]_ , \new_[35969]_ , \new_[35970]_ , \new_[35974]_ ,
    \new_[35975]_ , \new_[35976]_ , \new_[35980]_ , \new_[35981]_ ,
    \new_[35985]_ , \new_[35986]_ , \new_[35987]_ , \new_[35991]_ ,
    \new_[35992]_ , \new_[35996]_ , \new_[35997]_ , \new_[35998]_ ,
    \new_[36002]_ , \new_[36003]_ , \new_[36007]_ , \new_[36008]_ ,
    \new_[36009]_ , \new_[36013]_ , \new_[36014]_ , \new_[36018]_ ,
    \new_[36019]_ , \new_[36020]_ , \new_[36024]_ , \new_[36025]_ ,
    \new_[36029]_ , \new_[36030]_ , \new_[36031]_ , \new_[36035]_ ,
    \new_[36036]_ , \new_[36040]_ , \new_[36041]_ , \new_[36042]_ ,
    \new_[36046]_ , \new_[36047]_ , \new_[36051]_ , \new_[36052]_ ,
    \new_[36053]_ , \new_[36057]_ , \new_[36058]_ , \new_[36062]_ ,
    \new_[36063]_ , \new_[36064]_ , \new_[36068]_ , \new_[36069]_ ,
    \new_[36073]_ , \new_[36074]_ , \new_[36075]_ , \new_[36079]_ ,
    \new_[36080]_ , \new_[36084]_ , \new_[36085]_ , \new_[36086]_ ,
    \new_[36090]_ , \new_[36091]_ , \new_[36095]_ , \new_[36096]_ ,
    \new_[36097]_ , \new_[36101]_ , \new_[36102]_ , \new_[36106]_ ,
    \new_[36107]_ , \new_[36108]_ , \new_[36112]_ , \new_[36113]_ ,
    \new_[36117]_ , \new_[36118]_ , \new_[36119]_ , \new_[36123]_ ,
    \new_[36124]_ , \new_[36128]_ , \new_[36129]_ , \new_[36130]_ ,
    \new_[36134]_ , \new_[36135]_ , \new_[36139]_ , \new_[36140]_ ,
    \new_[36141]_ , \new_[36145]_ , \new_[36146]_ , \new_[36150]_ ,
    \new_[36151]_ , \new_[36152]_ , \new_[36156]_ , \new_[36157]_ ,
    \new_[36161]_ , \new_[36162]_ , \new_[36163]_ , \new_[36167]_ ,
    \new_[36168]_ , \new_[36172]_ , \new_[36173]_ , \new_[36174]_ ,
    \new_[36178]_ , \new_[36179]_ , \new_[36183]_ , \new_[36184]_ ,
    \new_[36185]_ , \new_[36189]_ , \new_[36190]_ , \new_[36194]_ ,
    \new_[36195]_ , \new_[36196]_ , \new_[36200]_ , \new_[36201]_ ,
    \new_[36205]_ , \new_[36206]_ , \new_[36207]_ , \new_[36211]_ ,
    \new_[36212]_ , \new_[36216]_ , \new_[36217]_ , \new_[36218]_ ,
    \new_[36222]_ , \new_[36223]_ , \new_[36227]_ , \new_[36228]_ ,
    \new_[36229]_ , \new_[36233]_ , \new_[36234]_ , \new_[36238]_ ,
    \new_[36239]_ , \new_[36240]_ , \new_[36244]_ , \new_[36245]_ ,
    \new_[36249]_ , \new_[36250]_ , \new_[36251]_ , \new_[36255]_ ,
    \new_[36256]_ , \new_[36260]_ , \new_[36261]_ , \new_[36262]_ ,
    \new_[36266]_ , \new_[36267]_ , \new_[36271]_ , \new_[36272]_ ,
    \new_[36273]_ , \new_[36277]_ , \new_[36278]_ , \new_[36282]_ ,
    \new_[36283]_ , \new_[36284]_ , \new_[36288]_ , \new_[36289]_ ,
    \new_[36293]_ , \new_[36294]_ , \new_[36295]_ , \new_[36299]_ ,
    \new_[36300]_ , \new_[36304]_ , \new_[36305]_ , \new_[36306]_ ,
    \new_[36310]_ , \new_[36311]_ , \new_[36315]_ , \new_[36316]_ ,
    \new_[36317]_ , \new_[36321]_ , \new_[36322]_ , \new_[36326]_ ,
    \new_[36327]_ , \new_[36328]_ , \new_[36332]_ , \new_[36333]_ ,
    \new_[36337]_ , \new_[36338]_ , \new_[36339]_ , \new_[36343]_ ,
    \new_[36344]_ , \new_[36348]_ , \new_[36349]_ , \new_[36350]_ ,
    \new_[36354]_ , \new_[36355]_ , \new_[36359]_ , \new_[36360]_ ,
    \new_[36361]_ , \new_[36365]_ , \new_[36366]_ , \new_[36370]_ ,
    \new_[36371]_ , \new_[36372]_ , \new_[36376]_ , \new_[36377]_ ,
    \new_[36381]_ , \new_[36382]_ , \new_[36383]_ , \new_[36387]_ ,
    \new_[36388]_ , \new_[36392]_ , \new_[36393]_ , \new_[36394]_ ,
    \new_[36398]_ , \new_[36399]_ , \new_[36403]_ , \new_[36404]_ ,
    \new_[36405]_ , \new_[36409]_ , \new_[36410]_ , \new_[36414]_ ,
    \new_[36415]_ , \new_[36416]_ , \new_[36420]_ , \new_[36421]_ ,
    \new_[36425]_ , \new_[36426]_ , \new_[36427]_ , \new_[36431]_ ,
    \new_[36432]_ , \new_[36436]_ , \new_[36437]_ , \new_[36438]_ ,
    \new_[36442]_ , \new_[36443]_ , \new_[36447]_ , \new_[36448]_ ,
    \new_[36449]_ , \new_[36453]_ , \new_[36454]_ , \new_[36458]_ ,
    \new_[36459]_ , \new_[36460]_ , \new_[36464]_ , \new_[36465]_ ,
    \new_[36469]_ , \new_[36470]_ , \new_[36471]_ , \new_[36475]_ ,
    \new_[36476]_ , \new_[36480]_ , \new_[36481]_ , \new_[36482]_ ,
    \new_[36486]_ , \new_[36487]_ , \new_[36491]_ , \new_[36492]_ ,
    \new_[36493]_ , \new_[36497]_ , \new_[36498]_ , \new_[36502]_ ,
    \new_[36503]_ , \new_[36504]_ , \new_[36508]_ , \new_[36509]_ ,
    \new_[36513]_ , \new_[36514]_ , \new_[36515]_ , \new_[36519]_ ,
    \new_[36520]_ , \new_[36524]_ , \new_[36525]_ , \new_[36526]_ ,
    \new_[36530]_ , \new_[36531]_ , \new_[36535]_ , \new_[36536]_ ,
    \new_[36537]_ , \new_[36541]_ , \new_[36542]_ , \new_[36546]_ ,
    \new_[36547]_ , \new_[36548]_ , \new_[36552]_ , \new_[36553]_ ,
    \new_[36557]_ , \new_[36558]_ , \new_[36559]_ , \new_[36563]_ ,
    \new_[36564]_ , \new_[36568]_ , \new_[36569]_ , \new_[36570]_ ,
    \new_[36574]_ , \new_[36575]_ , \new_[36579]_ , \new_[36580]_ ,
    \new_[36581]_ , \new_[36585]_ , \new_[36586]_ , \new_[36590]_ ,
    \new_[36591]_ , \new_[36592]_ , \new_[36596]_ , \new_[36597]_ ,
    \new_[36601]_ , \new_[36602]_ , \new_[36603]_ , \new_[36607]_ ,
    \new_[36608]_ , \new_[36612]_ , \new_[36613]_ , \new_[36614]_ ,
    \new_[36618]_ , \new_[36619]_ , \new_[36623]_ , \new_[36624]_ ,
    \new_[36625]_ , \new_[36629]_ , \new_[36630]_ , \new_[36634]_ ,
    \new_[36635]_ , \new_[36636]_ , \new_[36640]_ , \new_[36641]_ ,
    \new_[36645]_ , \new_[36646]_ , \new_[36647]_ , \new_[36651]_ ,
    \new_[36652]_ , \new_[36656]_ , \new_[36657]_ , \new_[36658]_ ,
    \new_[36662]_ , \new_[36663]_ , \new_[36667]_ , \new_[36668]_ ,
    \new_[36669]_ , \new_[36673]_ , \new_[36674]_ , \new_[36678]_ ,
    \new_[36679]_ , \new_[36680]_ , \new_[36684]_ , \new_[36685]_ ,
    \new_[36689]_ , \new_[36690]_ , \new_[36691]_ , \new_[36695]_ ,
    \new_[36696]_ , \new_[36700]_ , \new_[36701]_ , \new_[36702]_ ,
    \new_[36706]_ , \new_[36707]_ , \new_[36711]_ , \new_[36712]_ ,
    \new_[36713]_ , \new_[36717]_ , \new_[36718]_ , \new_[36722]_ ,
    \new_[36723]_ , \new_[36724]_ , \new_[36728]_ , \new_[36729]_ ,
    \new_[36733]_ , \new_[36734]_ , \new_[36735]_ , \new_[36739]_ ,
    \new_[36740]_ , \new_[36744]_ , \new_[36745]_ , \new_[36746]_ ,
    \new_[36750]_ , \new_[36751]_ , \new_[36755]_ , \new_[36756]_ ,
    \new_[36757]_ , \new_[36761]_ , \new_[36762]_ , \new_[36766]_ ,
    \new_[36767]_ , \new_[36768]_ , \new_[36772]_ , \new_[36773]_ ,
    \new_[36777]_ , \new_[36778]_ , \new_[36779]_ , \new_[36783]_ ,
    \new_[36784]_ , \new_[36788]_ , \new_[36789]_ , \new_[36790]_ ,
    \new_[36794]_ , \new_[36795]_ , \new_[36799]_ , \new_[36800]_ ,
    \new_[36801]_ , \new_[36805]_ , \new_[36806]_ , \new_[36810]_ ,
    \new_[36811]_ , \new_[36812]_ , \new_[36816]_ , \new_[36817]_ ,
    \new_[36821]_ , \new_[36822]_ , \new_[36823]_ , \new_[36827]_ ,
    \new_[36828]_ , \new_[36832]_ , \new_[36833]_ , \new_[36834]_ ,
    \new_[36838]_ , \new_[36839]_ , \new_[36843]_ , \new_[36844]_ ,
    \new_[36845]_ , \new_[36849]_ , \new_[36850]_ , \new_[36854]_ ,
    \new_[36855]_ , \new_[36856]_ , \new_[36860]_ , \new_[36861]_ ,
    \new_[36865]_ , \new_[36866]_ , \new_[36867]_ , \new_[36871]_ ,
    \new_[36872]_ , \new_[36876]_ , \new_[36877]_ , \new_[36878]_ ,
    \new_[36882]_ , \new_[36883]_ , \new_[36887]_ , \new_[36888]_ ,
    \new_[36889]_ , \new_[36893]_ , \new_[36894]_ , \new_[36898]_ ,
    \new_[36899]_ , \new_[36900]_ , \new_[36904]_ , \new_[36905]_ ,
    \new_[36909]_ , \new_[36910]_ , \new_[36911]_ , \new_[36915]_ ,
    \new_[36916]_ , \new_[36920]_ , \new_[36921]_ , \new_[36922]_ ,
    \new_[36926]_ , \new_[36927]_ , \new_[36931]_ , \new_[36932]_ ,
    \new_[36933]_ , \new_[36937]_ , \new_[36938]_ , \new_[36942]_ ,
    \new_[36943]_ , \new_[36944]_ , \new_[36948]_ , \new_[36949]_ ,
    \new_[36953]_ , \new_[36954]_ , \new_[36955]_ , \new_[36959]_ ,
    \new_[36960]_ , \new_[36964]_ , \new_[36965]_ , \new_[36966]_ ,
    \new_[36970]_ , \new_[36971]_ , \new_[36975]_ , \new_[36976]_ ,
    \new_[36977]_ , \new_[36981]_ , \new_[36982]_ , \new_[36986]_ ,
    \new_[36987]_ , \new_[36988]_ , \new_[36992]_ , \new_[36993]_ ,
    \new_[36997]_ , \new_[36998]_ , \new_[36999]_ , \new_[37003]_ ,
    \new_[37004]_ , \new_[37008]_ , \new_[37009]_ , \new_[37010]_ ,
    \new_[37014]_ , \new_[37015]_ , \new_[37019]_ , \new_[37020]_ ,
    \new_[37021]_ , \new_[37025]_ , \new_[37026]_ , \new_[37030]_ ,
    \new_[37031]_ , \new_[37032]_ , \new_[37036]_ , \new_[37037]_ ,
    \new_[37041]_ , \new_[37042]_ , \new_[37043]_ , \new_[37047]_ ,
    \new_[37048]_ , \new_[37052]_ , \new_[37053]_ , \new_[37054]_ ,
    \new_[37058]_ , \new_[37059]_ , \new_[37063]_ , \new_[37064]_ ,
    \new_[37065]_ , \new_[37069]_ , \new_[37070]_ , \new_[37074]_ ,
    \new_[37075]_ , \new_[37076]_ , \new_[37080]_ , \new_[37081]_ ,
    \new_[37085]_ , \new_[37086]_ , \new_[37087]_ , \new_[37091]_ ,
    \new_[37092]_ , \new_[37096]_ , \new_[37097]_ , \new_[37098]_ ,
    \new_[37102]_ , \new_[37103]_ , \new_[37107]_ , \new_[37108]_ ,
    \new_[37109]_ , \new_[37113]_ , \new_[37114]_ , \new_[37118]_ ,
    \new_[37119]_ , \new_[37120]_ , \new_[37124]_ , \new_[37125]_ ,
    \new_[37129]_ , \new_[37130]_ , \new_[37131]_ , \new_[37135]_ ,
    \new_[37136]_ , \new_[37140]_ , \new_[37141]_ , \new_[37142]_ ,
    \new_[37146]_ , \new_[37147]_ , \new_[37151]_ , \new_[37152]_ ,
    \new_[37153]_ , \new_[37157]_ , \new_[37158]_ , \new_[37162]_ ,
    \new_[37163]_ , \new_[37164]_ , \new_[37168]_ , \new_[37169]_ ,
    \new_[37173]_ , \new_[37174]_ , \new_[37175]_ , \new_[37179]_ ,
    \new_[37180]_ , \new_[37184]_ , \new_[37185]_ , \new_[37186]_ ,
    \new_[37190]_ , \new_[37191]_ , \new_[37195]_ , \new_[37196]_ ,
    \new_[37197]_ , \new_[37201]_ , \new_[37202]_ , \new_[37206]_ ,
    \new_[37207]_ , \new_[37208]_ , \new_[37212]_ , \new_[37213]_ ,
    \new_[37217]_ , \new_[37218]_ , \new_[37219]_ , \new_[37223]_ ,
    \new_[37224]_ , \new_[37228]_ , \new_[37229]_ , \new_[37230]_ ,
    \new_[37234]_ , \new_[37235]_ , \new_[37239]_ , \new_[37240]_ ,
    \new_[37241]_ , \new_[37245]_ , \new_[37246]_ , \new_[37250]_ ,
    \new_[37251]_ , \new_[37252]_ , \new_[37256]_ , \new_[37257]_ ,
    \new_[37261]_ , \new_[37262]_ , \new_[37263]_ , \new_[37267]_ ,
    \new_[37268]_ , \new_[37272]_ , \new_[37273]_ , \new_[37274]_ ,
    \new_[37278]_ , \new_[37279]_ , \new_[37283]_ , \new_[37284]_ ,
    \new_[37285]_ , \new_[37289]_ , \new_[37290]_ , \new_[37294]_ ,
    \new_[37295]_ , \new_[37296]_ , \new_[37300]_ , \new_[37301]_ ,
    \new_[37305]_ , \new_[37306]_ , \new_[37307]_ , \new_[37311]_ ,
    \new_[37312]_ , \new_[37316]_ , \new_[37317]_ , \new_[37318]_ ,
    \new_[37322]_ , \new_[37323]_ , \new_[37327]_ , \new_[37328]_ ,
    \new_[37329]_ , \new_[37333]_ , \new_[37334]_ , \new_[37338]_ ,
    \new_[37339]_ , \new_[37340]_ , \new_[37344]_ , \new_[37345]_ ,
    \new_[37349]_ , \new_[37350]_ , \new_[37351]_ , \new_[37355]_ ,
    \new_[37356]_ , \new_[37360]_ , \new_[37361]_ , \new_[37362]_ ,
    \new_[37366]_ , \new_[37367]_ , \new_[37371]_ , \new_[37372]_ ,
    \new_[37373]_ , \new_[37377]_ , \new_[37378]_ , \new_[37382]_ ,
    \new_[37383]_ , \new_[37384]_ , \new_[37388]_ , \new_[37389]_ ,
    \new_[37393]_ , \new_[37394]_ , \new_[37395]_ , \new_[37399]_ ,
    \new_[37400]_ , \new_[37404]_ , \new_[37405]_ , \new_[37406]_ ,
    \new_[37410]_ , \new_[37411]_ , \new_[37415]_ , \new_[37416]_ ,
    \new_[37417]_ , \new_[37421]_ , \new_[37422]_ , \new_[37426]_ ,
    \new_[37427]_ , \new_[37428]_ , \new_[37432]_ , \new_[37433]_ ,
    \new_[37437]_ , \new_[37438]_ , \new_[37439]_ , \new_[37443]_ ,
    \new_[37444]_ , \new_[37448]_ , \new_[37449]_ , \new_[37450]_ ,
    \new_[37454]_ , \new_[37455]_ , \new_[37459]_ , \new_[37460]_ ,
    \new_[37461]_ , \new_[37465]_ , \new_[37466]_ , \new_[37470]_ ,
    \new_[37471]_ , \new_[37472]_ , \new_[37476]_ , \new_[37477]_ ,
    \new_[37481]_ , \new_[37482]_ , \new_[37483]_ , \new_[37487]_ ,
    \new_[37488]_ , \new_[37492]_ , \new_[37493]_ , \new_[37494]_ ,
    \new_[37498]_ , \new_[37499]_ , \new_[37503]_ , \new_[37504]_ ,
    \new_[37505]_ , \new_[37509]_ , \new_[37510]_ , \new_[37514]_ ,
    \new_[37515]_ , \new_[37516]_ , \new_[37520]_ , \new_[37521]_ ,
    \new_[37525]_ , \new_[37526]_ , \new_[37527]_ , \new_[37531]_ ,
    \new_[37532]_ , \new_[37536]_ , \new_[37537]_ , \new_[37538]_ ,
    \new_[37542]_ , \new_[37543]_ , \new_[37547]_ , \new_[37548]_ ,
    \new_[37549]_ , \new_[37553]_ , \new_[37554]_ , \new_[37558]_ ,
    \new_[37559]_ , \new_[37560]_ , \new_[37564]_ , \new_[37565]_ ,
    \new_[37569]_ , \new_[37570]_ , \new_[37571]_ , \new_[37575]_ ,
    \new_[37576]_ , \new_[37580]_ , \new_[37581]_ , \new_[37582]_ ,
    \new_[37586]_ , \new_[37587]_ , \new_[37591]_ , \new_[37592]_ ,
    \new_[37593]_ , \new_[37597]_ , \new_[37598]_ , \new_[37602]_ ,
    \new_[37603]_ , \new_[37604]_ , \new_[37608]_ , \new_[37609]_ ,
    \new_[37613]_ , \new_[37614]_ , \new_[37615]_ , \new_[37619]_ ,
    \new_[37620]_ , \new_[37624]_ , \new_[37625]_ , \new_[37626]_ ,
    \new_[37630]_ , \new_[37631]_ , \new_[37635]_ , \new_[37636]_ ,
    \new_[37637]_ , \new_[37641]_ , \new_[37642]_ , \new_[37646]_ ,
    \new_[37647]_ , \new_[37648]_ , \new_[37652]_ , \new_[37653]_ ,
    \new_[37657]_ , \new_[37658]_ , \new_[37659]_ , \new_[37663]_ ,
    \new_[37664]_ , \new_[37667]_ , \new_[37670]_ , \new_[37671]_ ,
    \new_[37672]_ , \new_[37676]_ , \new_[37677]_ , \new_[37681]_ ,
    \new_[37682]_ , \new_[37683]_ , \new_[37687]_ , \new_[37688]_ ,
    \new_[37691]_ , \new_[37694]_ , \new_[37695]_ , \new_[37696]_ ,
    \new_[37700]_ , \new_[37701]_ , \new_[37705]_ , \new_[37706]_ ,
    \new_[37707]_ , \new_[37711]_ , \new_[37712]_ , \new_[37715]_ ,
    \new_[37718]_ , \new_[37719]_ , \new_[37720]_ , \new_[37724]_ ,
    \new_[37725]_ , \new_[37729]_ , \new_[37730]_ , \new_[37731]_ ,
    \new_[37735]_ , \new_[37736]_ , \new_[37739]_ , \new_[37742]_ ,
    \new_[37743]_ , \new_[37744]_ , \new_[37748]_ , \new_[37749]_ ,
    \new_[37753]_ , \new_[37754]_ , \new_[37755]_ , \new_[37759]_ ,
    \new_[37760]_ , \new_[37763]_ , \new_[37766]_ , \new_[37767]_ ,
    \new_[37768]_ , \new_[37772]_ , \new_[37773]_ , \new_[37777]_ ,
    \new_[37778]_ , \new_[37779]_ , \new_[37783]_ , \new_[37784]_ ,
    \new_[37787]_ , \new_[37790]_ , \new_[37791]_ , \new_[37792]_ ,
    \new_[37796]_ , \new_[37797]_ , \new_[37801]_ , \new_[37802]_ ,
    \new_[37803]_ , \new_[37807]_ , \new_[37808]_ , \new_[37811]_ ,
    \new_[37814]_ , \new_[37815]_ , \new_[37816]_ , \new_[37820]_ ,
    \new_[37821]_ , \new_[37825]_ , \new_[37826]_ , \new_[37827]_ ,
    \new_[37831]_ , \new_[37832]_ , \new_[37835]_ , \new_[37838]_ ,
    \new_[37839]_ , \new_[37840]_ , \new_[37844]_ , \new_[37845]_ ,
    \new_[37849]_ , \new_[37850]_ , \new_[37851]_ , \new_[37855]_ ,
    \new_[37856]_ , \new_[37859]_ , \new_[37862]_ , \new_[37863]_ ,
    \new_[37864]_ , \new_[37868]_ , \new_[37869]_ , \new_[37873]_ ,
    \new_[37874]_ , \new_[37875]_ , \new_[37879]_ , \new_[37880]_ ,
    \new_[37883]_ , \new_[37886]_ , \new_[37887]_ , \new_[37888]_ ,
    \new_[37892]_ , \new_[37893]_ , \new_[37897]_ , \new_[37898]_ ,
    \new_[37899]_ , \new_[37903]_ , \new_[37904]_ , \new_[37907]_ ,
    \new_[37910]_ , \new_[37911]_ , \new_[37912]_ , \new_[37916]_ ,
    \new_[37917]_ , \new_[37921]_ , \new_[37922]_ , \new_[37923]_ ,
    \new_[37927]_ , \new_[37928]_ , \new_[37931]_ , \new_[37934]_ ,
    \new_[37935]_ , \new_[37936]_ , \new_[37940]_ , \new_[37941]_ ,
    \new_[37945]_ , \new_[37946]_ , \new_[37947]_ , \new_[37951]_ ,
    \new_[37952]_ , \new_[37955]_ , \new_[37958]_ , \new_[37959]_ ,
    \new_[37960]_ , \new_[37964]_ , \new_[37965]_ , \new_[37969]_ ,
    \new_[37970]_ , \new_[37971]_ , \new_[37975]_ , \new_[37976]_ ,
    \new_[37979]_ , \new_[37982]_ , \new_[37983]_ , \new_[37984]_ ,
    \new_[37988]_ , \new_[37989]_ , \new_[37993]_ , \new_[37994]_ ,
    \new_[37995]_ , \new_[37999]_ , \new_[38000]_ , \new_[38003]_ ,
    \new_[38006]_ , \new_[38007]_ , \new_[38008]_ , \new_[38012]_ ,
    \new_[38013]_ , \new_[38017]_ , \new_[38018]_ , \new_[38019]_ ,
    \new_[38023]_ , \new_[38024]_ , \new_[38027]_ , \new_[38030]_ ,
    \new_[38031]_ , \new_[38032]_ , \new_[38036]_ , \new_[38037]_ ,
    \new_[38041]_ , \new_[38042]_ , \new_[38043]_ , \new_[38047]_ ,
    \new_[38048]_ , \new_[38051]_ , \new_[38054]_ , \new_[38055]_ ,
    \new_[38056]_ , \new_[38060]_ , \new_[38061]_ , \new_[38065]_ ,
    \new_[38066]_ , \new_[38067]_ , \new_[38071]_ , \new_[38072]_ ,
    \new_[38075]_ , \new_[38078]_ , \new_[38079]_ , \new_[38080]_ ,
    \new_[38084]_ , \new_[38085]_ , \new_[38089]_ , \new_[38090]_ ,
    \new_[38091]_ , \new_[38095]_ , \new_[38096]_ , \new_[38099]_ ,
    \new_[38102]_ , \new_[38103]_ , \new_[38104]_ , \new_[38108]_ ,
    \new_[38109]_ , \new_[38113]_ , \new_[38114]_ , \new_[38115]_ ,
    \new_[38119]_ , \new_[38120]_ , \new_[38123]_ , \new_[38126]_ ,
    \new_[38127]_ , \new_[38128]_ , \new_[38132]_ , \new_[38133]_ ,
    \new_[38137]_ , \new_[38138]_ , \new_[38139]_ , \new_[38143]_ ,
    \new_[38144]_ , \new_[38147]_ , \new_[38150]_ , \new_[38151]_ ,
    \new_[38152]_ , \new_[38156]_ , \new_[38157]_ , \new_[38161]_ ,
    \new_[38162]_ , \new_[38163]_ , \new_[38167]_ , \new_[38168]_ ,
    \new_[38171]_ , \new_[38174]_ , \new_[38175]_ , \new_[38176]_ ,
    \new_[38180]_ , \new_[38181]_ , \new_[38185]_ , \new_[38186]_ ,
    \new_[38187]_ , \new_[38191]_ , \new_[38192]_ , \new_[38195]_ ,
    \new_[38198]_ , \new_[38199]_ , \new_[38200]_ , \new_[38204]_ ,
    \new_[38205]_ , \new_[38209]_ , \new_[38210]_ , \new_[38211]_ ,
    \new_[38215]_ , \new_[38216]_ , \new_[38219]_ , \new_[38222]_ ,
    \new_[38223]_ , \new_[38224]_ , \new_[38228]_ , \new_[38229]_ ,
    \new_[38233]_ , \new_[38234]_ , \new_[38235]_ , \new_[38239]_ ,
    \new_[38240]_ , \new_[38243]_ , \new_[38246]_ , \new_[38247]_ ,
    \new_[38248]_ , \new_[38252]_ , \new_[38253]_ , \new_[38257]_ ,
    \new_[38258]_ , \new_[38259]_ , \new_[38263]_ , \new_[38264]_ ,
    \new_[38267]_ , \new_[38270]_ , \new_[38271]_ , \new_[38272]_ ,
    \new_[38276]_ , \new_[38277]_ , \new_[38281]_ , \new_[38282]_ ,
    \new_[38283]_ , \new_[38287]_ , \new_[38288]_ , \new_[38291]_ ,
    \new_[38294]_ , \new_[38295]_ , \new_[38296]_ , \new_[38300]_ ,
    \new_[38301]_ , \new_[38305]_ , \new_[38306]_ , \new_[38307]_ ,
    \new_[38311]_ , \new_[38312]_ , \new_[38315]_ , \new_[38318]_ ,
    \new_[38319]_ , \new_[38320]_ , \new_[38324]_ , \new_[38325]_ ,
    \new_[38329]_ , \new_[38330]_ , \new_[38331]_ , \new_[38335]_ ,
    \new_[38336]_ , \new_[38339]_ , \new_[38342]_ , \new_[38343]_ ,
    \new_[38344]_ , \new_[38348]_ , \new_[38349]_ , \new_[38353]_ ,
    \new_[38354]_ , \new_[38355]_ , \new_[38359]_ , \new_[38360]_ ,
    \new_[38363]_ , \new_[38366]_ , \new_[38367]_ , \new_[38368]_ ,
    \new_[38372]_ , \new_[38373]_ , \new_[38377]_ , \new_[38378]_ ,
    \new_[38379]_ , \new_[38383]_ , \new_[38384]_ , \new_[38387]_ ,
    \new_[38390]_ , \new_[38391]_ , \new_[38392]_ , \new_[38396]_ ,
    \new_[38397]_ , \new_[38401]_ , \new_[38402]_ , \new_[38403]_ ,
    \new_[38407]_ , \new_[38408]_ , \new_[38411]_ , \new_[38414]_ ,
    \new_[38415]_ , \new_[38416]_ , \new_[38420]_ , \new_[38421]_ ,
    \new_[38425]_ , \new_[38426]_ , \new_[38427]_ , \new_[38431]_ ,
    \new_[38432]_ , \new_[38435]_ , \new_[38438]_ , \new_[38439]_ ,
    \new_[38440]_ , \new_[38444]_ , \new_[38445]_ , \new_[38449]_ ,
    \new_[38450]_ , \new_[38451]_ , \new_[38455]_ , \new_[38456]_ ,
    \new_[38459]_ , \new_[38462]_ , \new_[38463]_ , \new_[38464]_ ,
    \new_[38468]_ , \new_[38469]_ , \new_[38473]_ , \new_[38474]_ ,
    \new_[38475]_ , \new_[38479]_ , \new_[38480]_ , \new_[38483]_ ,
    \new_[38486]_ , \new_[38487]_ , \new_[38488]_ , \new_[38492]_ ,
    \new_[38493]_ , \new_[38497]_ , \new_[38498]_ , \new_[38499]_ ,
    \new_[38503]_ , \new_[38504]_ , \new_[38507]_ , \new_[38510]_ ,
    \new_[38511]_ , \new_[38512]_ , \new_[38516]_ , \new_[38517]_ ,
    \new_[38521]_ , \new_[38522]_ , \new_[38523]_ , \new_[38527]_ ,
    \new_[38528]_ , \new_[38531]_ , \new_[38534]_ , \new_[38535]_ ,
    \new_[38536]_ , \new_[38540]_ , \new_[38541]_ , \new_[38545]_ ,
    \new_[38546]_ , \new_[38547]_ , \new_[38551]_ , \new_[38552]_ ,
    \new_[38555]_ , \new_[38558]_ , \new_[38559]_ , \new_[38560]_ ,
    \new_[38564]_ , \new_[38565]_ , \new_[38569]_ , \new_[38570]_ ,
    \new_[38571]_ , \new_[38575]_ , \new_[38576]_ , \new_[38579]_ ,
    \new_[38582]_ , \new_[38583]_ , \new_[38584]_ , \new_[38588]_ ,
    \new_[38589]_ , \new_[38593]_ , \new_[38594]_ , \new_[38595]_ ,
    \new_[38599]_ , \new_[38600]_ , \new_[38603]_ , \new_[38606]_ ,
    \new_[38607]_ , \new_[38608]_ , \new_[38612]_ , \new_[38613]_ ,
    \new_[38617]_ , \new_[38618]_ , \new_[38619]_ , \new_[38623]_ ,
    \new_[38624]_ , \new_[38627]_ , \new_[38630]_ , \new_[38631]_ ,
    \new_[38632]_ , \new_[38636]_ , \new_[38637]_ , \new_[38641]_ ,
    \new_[38642]_ , \new_[38643]_ , \new_[38647]_ , \new_[38648]_ ,
    \new_[38651]_ , \new_[38654]_ , \new_[38655]_ , \new_[38656]_ ,
    \new_[38660]_ , \new_[38661]_ , \new_[38665]_ , \new_[38666]_ ,
    \new_[38667]_ , \new_[38671]_ , \new_[38672]_ , \new_[38675]_ ,
    \new_[38678]_ , \new_[38679]_ , \new_[38680]_ , \new_[38684]_ ,
    \new_[38685]_ , \new_[38689]_ , \new_[38690]_ , \new_[38691]_ ,
    \new_[38695]_ , \new_[38696]_ , \new_[38699]_ , \new_[38702]_ ,
    \new_[38703]_ , \new_[38704]_ , \new_[38708]_ , \new_[38709]_ ,
    \new_[38713]_ , \new_[38714]_ , \new_[38715]_ , \new_[38719]_ ,
    \new_[38720]_ , \new_[38723]_ , \new_[38726]_ , \new_[38727]_ ,
    \new_[38728]_ , \new_[38732]_ , \new_[38733]_ , \new_[38737]_ ,
    \new_[38738]_ , \new_[38739]_ , \new_[38743]_ , \new_[38744]_ ,
    \new_[38747]_ , \new_[38750]_ , \new_[38751]_ , \new_[38752]_ ,
    \new_[38756]_ , \new_[38757]_ , \new_[38761]_ , \new_[38762]_ ,
    \new_[38763]_ , \new_[38767]_ , \new_[38768]_ , \new_[38771]_ ,
    \new_[38774]_ , \new_[38775]_ , \new_[38776]_ , \new_[38780]_ ,
    \new_[38781]_ , \new_[38785]_ , \new_[38786]_ , \new_[38787]_ ,
    \new_[38791]_ , \new_[38792]_ , \new_[38795]_ , \new_[38798]_ ,
    \new_[38799]_ , \new_[38800]_ , \new_[38804]_ , \new_[38805]_ ,
    \new_[38809]_ , \new_[38810]_ , \new_[38811]_ , \new_[38815]_ ,
    \new_[38816]_ , \new_[38819]_ , \new_[38822]_ , \new_[38823]_ ,
    \new_[38824]_ , \new_[38828]_ , \new_[38829]_ , \new_[38833]_ ,
    \new_[38834]_ , \new_[38835]_ , \new_[38839]_ , \new_[38840]_ ,
    \new_[38843]_ , \new_[38846]_ , \new_[38847]_ , \new_[38848]_ ,
    \new_[38852]_ , \new_[38853]_ , \new_[38857]_ , \new_[38858]_ ,
    \new_[38859]_ , \new_[38863]_ , \new_[38864]_ , \new_[38867]_ ,
    \new_[38870]_ , \new_[38871]_ , \new_[38872]_ , \new_[38876]_ ,
    \new_[38877]_ , \new_[38881]_ , \new_[38882]_ , \new_[38883]_ ,
    \new_[38887]_ , \new_[38888]_ , \new_[38891]_ , \new_[38894]_ ,
    \new_[38895]_ , \new_[38896]_ , \new_[38900]_ , \new_[38901]_ ,
    \new_[38905]_ , \new_[38906]_ , \new_[38907]_ , \new_[38911]_ ,
    \new_[38912]_ , \new_[38915]_ , \new_[38918]_ , \new_[38919]_ ,
    \new_[38920]_ , \new_[38924]_ , \new_[38925]_ , \new_[38929]_ ,
    \new_[38930]_ , \new_[38931]_ , \new_[38935]_ , \new_[38936]_ ,
    \new_[38939]_ , \new_[38942]_ , \new_[38943]_ , \new_[38944]_ ,
    \new_[38948]_ , \new_[38949]_ , \new_[38953]_ , \new_[38954]_ ,
    \new_[38955]_ , \new_[38959]_ , \new_[38960]_ , \new_[38963]_ ,
    \new_[38966]_ , \new_[38967]_ , \new_[38968]_ , \new_[38972]_ ,
    \new_[38973]_ , \new_[38977]_ , \new_[38978]_ , \new_[38979]_ ,
    \new_[38983]_ , \new_[38984]_ , \new_[38987]_ , \new_[38990]_ ,
    \new_[38991]_ , \new_[38992]_ , \new_[38996]_ , \new_[38997]_ ,
    \new_[39001]_ , \new_[39002]_ , \new_[39003]_ , \new_[39007]_ ,
    \new_[39008]_ , \new_[39011]_ , \new_[39014]_ , \new_[39015]_ ,
    \new_[39016]_ , \new_[39020]_ , \new_[39021]_ , \new_[39025]_ ,
    \new_[39026]_ , \new_[39027]_ , \new_[39031]_ , \new_[39032]_ ,
    \new_[39035]_ , \new_[39038]_ , \new_[39039]_ , \new_[39040]_ ,
    \new_[39044]_ , \new_[39045]_ , \new_[39049]_ , \new_[39050]_ ,
    \new_[39051]_ , \new_[39055]_ , \new_[39056]_ , \new_[39059]_ ,
    \new_[39062]_ , \new_[39063]_ , \new_[39064]_ , \new_[39068]_ ,
    \new_[39069]_ , \new_[39073]_ , \new_[39074]_ , \new_[39075]_ ,
    \new_[39079]_ , \new_[39080]_ , \new_[39083]_ , \new_[39086]_ ,
    \new_[39087]_ , \new_[39088]_ , \new_[39092]_ , \new_[39093]_ ,
    \new_[39097]_ , \new_[39098]_ , \new_[39099]_ , \new_[39103]_ ,
    \new_[39104]_ , \new_[39107]_ , \new_[39110]_ , \new_[39111]_ ,
    \new_[39112]_ , \new_[39116]_ , \new_[39117]_ , \new_[39121]_ ,
    \new_[39122]_ , \new_[39123]_ , \new_[39127]_ , \new_[39128]_ ,
    \new_[39131]_ , \new_[39134]_ , \new_[39135]_ , \new_[39136]_ ,
    \new_[39140]_ , \new_[39141]_ , \new_[39145]_ , \new_[39146]_ ,
    \new_[39147]_ , \new_[39151]_ , \new_[39152]_ , \new_[39155]_ ,
    \new_[39158]_ , \new_[39159]_ , \new_[39160]_ , \new_[39164]_ ,
    \new_[39165]_ , \new_[39169]_ , \new_[39170]_ , \new_[39171]_ ,
    \new_[39175]_ , \new_[39176]_ , \new_[39179]_ , \new_[39182]_ ,
    \new_[39183]_ , \new_[39184]_ , \new_[39188]_ , \new_[39189]_ ,
    \new_[39193]_ , \new_[39194]_ , \new_[39195]_ , \new_[39199]_ ,
    \new_[39200]_ , \new_[39203]_ , \new_[39206]_ , \new_[39207]_ ,
    \new_[39208]_ , \new_[39212]_ , \new_[39213]_ , \new_[39217]_ ,
    \new_[39218]_ , \new_[39219]_ , \new_[39223]_ , \new_[39224]_ ,
    \new_[39227]_ , \new_[39230]_ , \new_[39231]_ , \new_[39232]_ ,
    \new_[39236]_ , \new_[39237]_ , \new_[39241]_ , \new_[39242]_ ,
    \new_[39243]_ , \new_[39247]_ , \new_[39248]_ , \new_[39251]_ ,
    \new_[39254]_ , \new_[39255]_ , \new_[39256]_ , \new_[39260]_ ,
    \new_[39261]_ , \new_[39265]_ , \new_[39266]_ , \new_[39267]_ ,
    \new_[39271]_ , \new_[39272]_ , \new_[39275]_ , \new_[39278]_ ,
    \new_[39279]_ , \new_[39280]_ , \new_[39284]_ , \new_[39285]_ ,
    \new_[39289]_ , \new_[39290]_ , \new_[39291]_ , \new_[39295]_ ,
    \new_[39296]_ , \new_[39299]_ , \new_[39302]_ , \new_[39303]_ ,
    \new_[39304]_ , \new_[39308]_ , \new_[39309]_ , \new_[39313]_ ,
    \new_[39314]_ , \new_[39315]_ , \new_[39319]_ , \new_[39320]_ ,
    \new_[39323]_ , \new_[39326]_ , \new_[39327]_ , \new_[39328]_ ,
    \new_[39332]_ , \new_[39333]_ , \new_[39337]_ , \new_[39338]_ ,
    \new_[39339]_ , \new_[39343]_ , \new_[39344]_ , \new_[39347]_ ,
    \new_[39350]_ , \new_[39351]_ , \new_[39352]_ , \new_[39356]_ ,
    \new_[39357]_ , \new_[39361]_ , \new_[39362]_ , \new_[39363]_ ,
    \new_[39367]_ , \new_[39368]_ , \new_[39371]_ , \new_[39374]_ ,
    \new_[39375]_ , \new_[39376]_ , \new_[39380]_ , \new_[39381]_ ,
    \new_[39385]_ , \new_[39386]_ , \new_[39387]_ , \new_[39391]_ ,
    \new_[39392]_ , \new_[39395]_ , \new_[39398]_ , \new_[39399]_ ,
    \new_[39400]_ , \new_[39404]_ , \new_[39405]_ , \new_[39409]_ ,
    \new_[39410]_ , \new_[39411]_ , \new_[39415]_ , \new_[39416]_ ,
    \new_[39419]_ , \new_[39422]_ , \new_[39423]_ , \new_[39424]_ ,
    \new_[39428]_ , \new_[39429]_ , \new_[39433]_ , \new_[39434]_ ,
    \new_[39435]_ , \new_[39439]_ , \new_[39440]_ , \new_[39443]_ ,
    \new_[39446]_ , \new_[39447]_ , \new_[39448]_ , \new_[39452]_ ,
    \new_[39453]_ , \new_[39457]_ , \new_[39458]_ , \new_[39459]_ ,
    \new_[39463]_ , \new_[39464]_ , \new_[39467]_ , \new_[39470]_ ,
    \new_[39471]_ , \new_[39472]_ , \new_[39476]_ , \new_[39477]_ ,
    \new_[39481]_ , \new_[39482]_ , \new_[39483]_ , \new_[39487]_ ,
    \new_[39488]_ , \new_[39491]_ , \new_[39494]_ , \new_[39495]_ ,
    \new_[39496]_ , \new_[39500]_ , \new_[39501]_ , \new_[39505]_ ,
    \new_[39506]_ , \new_[39507]_ , \new_[39511]_ , \new_[39512]_ ,
    \new_[39515]_ , \new_[39518]_ , \new_[39519]_ , \new_[39520]_ ,
    \new_[39524]_ , \new_[39525]_ , \new_[39529]_ , \new_[39530]_ ,
    \new_[39531]_ , \new_[39535]_ , \new_[39536]_ , \new_[39539]_ ,
    \new_[39542]_ , \new_[39543]_ , \new_[39544]_ , \new_[39548]_ ,
    \new_[39549]_ , \new_[39553]_ , \new_[39554]_ , \new_[39555]_ ,
    \new_[39559]_ , \new_[39560]_ , \new_[39563]_ , \new_[39566]_ ,
    \new_[39567]_ , \new_[39568]_ , \new_[39572]_ , \new_[39573]_ ,
    \new_[39577]_ , \new_[39578]_ , \new_[39579]_ , \new_[39583]_ ,
    \new_[39584]_ , \new_[39587]_ , \new_[39590]_ , \new_[39591]_ ,
    \new_[39592]_ , \new_[39596]_ , \new_[39597]_ , \new_[39601]_ ,
    \new_[39602]_ , \new_[39603]_ , \new_[39607]_ , \new_[39608]_ ,
    \new_[39611]_ , \new_[39614]_ , \new_[39615]_ , \new_[39616]_ ,
    \new_[39620]_ , \new_[39621]_ , \new_[39625]_ , \new_[39626]_ ,
    \new_[39627]_ , \new_[39631]_ , \new_[39632]_ , \new_[39635]_ ,
    \new_[39638]_ , \new_[39639]_ , \new_[39640]_ , \new_[39644]_ ,
    \new_[39645]_ , \new_[39649]_ , \new_[39650]_ , \new_[39651]_ ,
    \new_[39655]_ , \new_[39656]_ , \new_[39659]_ , \new_[39662]_ ,
    \new_[39663]_ , \new_[39664]_ , \new_[39668]_ , \new_[39669]_ ,
    \new_[39673]_ , \new_[39674]_ , \new_[39675]_ , \new_[39679]_ ,
    \new_[39680]_ , \new_[39683]_ , \new_[39686]_ , \new_[39687]_ ,
    \new_[39688]_ , \new_[39692]_ , \new_[39693]_ , \new_[39697]_ ,
    \new_[39698]_ , \new_[39699]_ , \new_[39703]_ , \new_[39704]_ ,
    \new_[39707]_ , \new_[39710]_ , \new_[39711]_ , \new_[39712]_ ,
    \new_[39716]_ , \new_[39717]_ , \new_[39721]_ , \new_[39722]_ ,
    \new_[39723]_ , \new_[39727]_ , \new_[39728]_ , \new_[39731]_ ,
    \new_[39734]_ , \new_[39735]_ , \new_[39736]_ , \new_[39740]_ ,
    \new_[39741]_ , \new_[39745]_ , \new_[39746]_ , \new_[39747]_ ,
    \new_[39751]_ , \new_[39752]_ , \new_[39755]_ , \new_[39758]_ ,
    \new_[39759]_ , \new_[39760]_ , \new_[39764]_ , \new_[39765]_ ,
    \new_[39769]_ , \new_[39770]_ , \new_[39771]_ , \new_[39775]_ ,
    \new_[39776]_ , \new_[39779]_ , \new_[39782]_ , \new_[39783]_ ,
    \new_[39784]_ , \new_[39788]_ , \new_[39789]_ , \new_[39793]_ ,
    \new_[39794]_ , \new_[39795]_ , \new_[39799]_ , \new_[39800]_ ,
    \new_[39803]_ , \new_[39806]_ , \new_[39807]_ , \new_[39808]_ ,
    \new_[39812]_ , \new_[39813]_ , \new_[39817]_ , \new_[39818]_ ,
    \new_[39819]_ , \new_[39823]_ , \new_[39824]_ , \new_[39827]_ ,
    \new_[39830]_ , \new_[39831]_ , \new_[39832]_ , \new_[39836]_ ,
    \new_[39837]_ , \new_[39841]_ , \new_[39842]_ , \new_[39843]_ ,
    \new_[39847]_ , \new_[39848]_ , \new_[39851]_ , \new_[39854]_ ,
    \new_[39855]_ , \new_[39856]_ , \new_[39860]_ , \new_[39861]_ ,
    \new_[39865]_ , \new_[39866]_ , \new_[39867]_ , \new_[39871]_ ,
    \new_[39872]_ , \new_[39875]_ , \new_[39878]_ , \new_[39879]_ ,
    \new_[39880]_ , \new_[39884]_ , \new_[39885]_ , \new_[39889]_ ,
    \new_[39890]_ , \new_[39891]_ , \new_[39895]_ , \new_[39896]_ ,
    \new_[39899]_ , \new_[39902]_ , \new_[39903]_ , \new_[39904]_ ,
    \new_[39908]_ , \new_[39909]_ , \new_[39913]_ , \new_[39914]_ ,
    \new_[39915]_ , \new_[39919]_ , \new_[39920]_ , \new_[39923]_ ,
    \new_[39926]_ , \new_[39927]_ , \new_[39928]_ , \new_[39932]_ ,
    \new_[39933]_ , \new_[39937]_ , \new_[39938]_ , \new_[39939]_ ,
    \new_[39943]_ , \new_[39944]_ , \new_[39947]_ , \new_[39950]_ ,
    \new_[39951]_ , \new_[39952]_ , \new_[39956]_ , \new_[39957]_ ,
    \new_[39961]_ , \new_[39962]_ , \new_[39963]_ , \new_[39967]_ ,
    \new_[39968]_ , \new_[39971]_ , \new_[39974]_ , \new_[39975]_ ,
    \new_[39976]_ , \new_[39980]_ , \new_[39981]_ , \new_[39985]_ ,
    \new_[39986]_ , \new_[39987]_ , \new_[39991]_ , \new_[39992]_ ,
    \new_[39995]_ , \new_[39998]_ , \new_[39999]_ , \new_[40000]_ ,
    \new_[40004]_ , \new_[40005]_ , \new_[40009]_ , \new_[40010]_ ,
    \new_[40011]_ , \new_[40015]_ , \new_[40016]_ , \new_[40019]_ ,
    \new_[40022]_ , \new_[40023]_ , \new_[40024]_ , \new_[40028]_ ,
    \new_[40029]_ , \new_[40033]_ , \new_[40034]_ , \new_[40035]_ ,
    \new_[40039]_ , \new_[40040]_ , \new_[40043]_ , \new_[40046]_ ,
    \new_[40047]_ , \new_[40048]_ , \new_[40052]_ , \new_[40053]_ ,
    \new_[40057]_ , \new_[40058]_ , \new_[40059]_ , \new_[40063]_ ,
    \new_[40064]_ , \new_[40067]_ , \new_[40070]_ , \new_[40071]_ ,
    \new_[40072]_ , \new_[40076]_ , \new_[40077]_ , \new_[40081]_ ,
    \new_[40082]_ , \new_[40083]_ , \new_[40087]_ , \new_[40088]_ ,
    \new_[40091]_ , \new_[40094]_ , \new_[40095]_ , \new_[40096]_ ,
    \new_[40100]_ , \new_[40101]_ , \new_[40105]_ , \new_[40106]_ ,
    \new_[40107]_ , \new_[40111]_ , \new_[40112]_ , \new_[40115]_ ,
    \new_[40118]_ , \new_[40119]_ , \new_[40120]_ , \new_[40124]_ ,
    \new_[40125]_ , \new_[40129]_ , \new_[40130]_ , \new_[40131]_ ,
    \new_[40135]_ , \new_[40136]_ , \new_[40139]_ , \new_[40142]_ ,
    \new_[40143]_ , \new_[40144]_ , \new_[40148]_ , \new_[40149]_ ,
    \new_[40153]_ , \new_[40154]_ , \new_[40155]_ , \new_[40159]_ ,
    \new_[40160]_ , \new_[40163]_ , \new_[40166]_ , \new_[40167]_ ,
    \new_[40168]_ , \new_[40172]_ , \new_[40173]_ , \new_[40177]_ ,
    \new_[40178]_ , \new_[40179]_ , \new_[40183]_ , \new_[40184]_ ,
    \new_[40187]_ , \new_[40190]_ , \new_[40191]_ , \new_[40192]_ ,
    \new_[40196]_ , \new_[40197]_ , \new_[40201]_ , \new_[40202]_ ,
    \new_[40203]_ , \new_[40207]_ , \new_[40208]_ , \new_[40211]_ ,
    \new_[40214]_ , \new_[40215]_ , \new_[40216]_ , \new_[40220]_ ,
    \new_[40221]_ , \new_[40225]_ , \new_[40226]_ , \new_[40227]_ ,
    \new_[40231]_ , \new_[40232]_ , \new_[40235]_ , \new_[40238]_ ,
    \new_[40239]_ , \new_[40240]_ , \new_[40244]_ , \new_[40245]_ ,
    \new_[40249]_ , \new_[40250]_ , \new_[40251]_ , \new_[40255]_ ,
    \new_[40256]_ , \new_[40259]_ , \new_[40262]_ , \new_[40263]_ ,
    \new_[40264]_ , \new_[40268]_ , \new_[40269]_ , \new_[40273]_ ,
    \new_[40274]_ , \new_[40275]_ , \new_[40279]_ , \new_[40280]_ ,
    \new_[40283]_ , \new_[40286]_ , \new_[40287]_ , \new_[40288]_ ,
    \new_[40292]_ , \new_[40293]_ , \new_[40297]_ , \new_[40298]_ ,
    \new_[40299]_ , \new_[40303]_ , \new_[40304]_ , \new_[40307]_ ,
    \new_[40310]_ , \new_[40311]_ , \new_[40312]_ , \new_[40316]_ ,
    \new_[40317]_ , \new_[40321]_ , \new_[40322]_ , \new_[40323]_ ,
    \new_[40327]_ , \new_[40328]_ , \new_[40331]_ , \new_[40334]_ ,
    \new_[40335]_ , \new_[40336]_ , \new_[40340]_ , \new_[40341]_ ,
    \new_[40345]_ , \new_[40346]_ , \new_[40347]_ , \new_[40351]_ ,
    \new_[40352]_ , \new_[40355]_ , \new_[40358]_ , \new_[40359]_ ,
    \new_[40360]_ , \new_[40364]_ , \new_[40365]_ , \new_[40369]_ ,
    \new_[40370]_ , \new_[40371]_ , \new_[40375]_ , \new_[40376]_ ,
    \new_[40379]_ , \new_[40382]_ , \new_[40383]_ , \new_[40384]_ ,
    \new_[40388]_ , \new_[40389]_ , \new_[40393]_ , \new_[40394]_ ,
    \new_[40395]_ , \new_[40399]_ , \new_[40400]_ , \new_[40403]_ ,
    \new_[40406]_ , \new_[40407]_ , \new_[40408]_ , \new_[40412]_ ,
    \new_[40413]_ , \new_[40417]_ , \new_[40418]_ , \new_[40419]_ ,
    \new_[40423]_ , \new_[40424]_ , \new_[40427]_ , \new_[40430]_ ,
    \new_[40431]_ , \new_[40432]_ , \new_[40436]_ , \new_[40437]_ ,
    \new_[40441]_ , \new_[40442]_ , \new_[40443]_ , \new_[40447]_ ,
    \new_[40448]_ , \new_[40451]_ , \new_[40454]_ , \new_[40455]_ ,
    \new_[40456]_ , \new_[40460]_ , \new_[40461]_ , \new_[40465]_ ,
    \new_[40466]_ , \new_[40467]_ , \new_[40471]_ , \new_[40472]_ ,
    \new_[40475]_ , \new_[40478]_ , \new_[40479]_ , \new_[40480]_ ,
    \new_[40484]_ , \new_[40485]_ , \new_[40489]_ , \new_[40490]_ ,
    \new_[40491]_ , \new_[40495]_ , \new_[40496]_ , \new_[40499]_ ,
    \new_[40502]_ , \new_[40503]_ , \new_[40504]_ , \new_[40508]_ ,
    \new_[40509]_ , \new_[40513]_ , \new_[40514]_ , \new_[40515]_ ,
    \new_[40519]_ , \new_[40520]_ , \new_[40523]_ , \new_[40526]_ ,
    \new_[40527]_ , \new_[40528]_ , \new_[40532]_ , \new_[40533]_ ,
    \new_[40537]_ , \new_[40538]_ , \new_[40539]_ , \new_[40543]_ ,
    \new_[40544]_ , \new_[40547]_ , \new_[40550]_ , \new_[40551]_ ,
    \new_[40552]_ , \new_[40556]_ , \new_[40557]_ , \new_[40561]_ ,
    \new_[40562]_ , \new_[40563]_ , \new_[40567]_ , \new_[40568]_ ,
    \new_[40571]_ , \new_[40574]_ , \new_[40575]_ , \new_[40576]_ ,
    \new_[40580]_ , \new_[40581]_ , \new_[40585]_ , \new_[40586]_ ,
    \new_[40587]_ , \new_[40591]_ , \new_[40592]_ , \new_[40595]_ ,
    \new_[40598]_ , \new_[40599]_ , \new_[40600]_ , \new_[40604]_ ,
    \new_[40605]_ , \new_[40609]_ , \new_[40610]_ , \new_[40611]_ ,
    \new_[40615]_ , \new_[40616]_ , \new_[40619]_ , \new_[40622]_ ,
    \new_[40623]_ , \new_[40624]_ , \new_[40628]_ , \new_[40629]_ ,
    \new_[40633]_ , \new_[40634]_ , \new_[40635]_ , \new_[40639]_ ,
    \new_[40640]_ , \new_[40643]_ , \new_[40646]_ , \new_[40647]_ ,
    \new_[40648]_ , \new_[40652]_ , \new_[40653]_ , \new_[40657]_ ,
    \new_[40658]_ , \new_[40659]_ , \new_[40663]_ , \new_[40664]_ ,
    \new_[40667]_ , \new_[40670]_ , \new_[40671]_ , \new_[40672]_ ,
    \new_[40676]_ , \new_[40677]_ , \new_[40681]_ , \new_[40682]_ ,
    \new_[40683]_ , \new_[40687]_ , \new_[40688]_ , \new_[40691]_ ,
    \new_[40694]_ , \new_[40695]_ , \new_[40696]_ , \new_[40700]_ ,
    \new_[40701]_ , \new_[40705]_ , \new_[40706]_ , \new_[40707]_ ,
    \new_[40711]_ , \new_[40712]_ , \new_[40715]_ , \new_[40718]_ ,
    \new_[40719]_ , \new_[40720]_ , \new_[40724]_ , \new_[40725]_ ,
    \new_[40729]_ , \new_[40730]_ , \new_[40731]_ , \new_[40735]_ ,
    \new_[40736]_ , \new_[40739]_ , \new_[40742]_ , \new_[40743]_ ,
    \new_[40744]_ , \new_[40748]_ , \new_[40749]_ , \new_[40753]_ ,
    \new_[40754]_ , \new_[40755]_ , \new_[40759]_ , \new_[40760]_ ,
    \new_[40763]_ , \new_[40766]_ , \new_[40767]_ , \new_[40768]_ ,
    \new_[40772]_ , \new_[40773]_ , \new_[40777]_ , \new_[40778]_ ,
    \new_[40779]_ , \new_[40783]_ , \new_[40784]_ , \new_[40787]_ ,
    \new_[40790]_ , \new_[40791]_ , \new_[40792]_ , \new_[40796]_ ,
    \new_[40797]_ , \new_[40801]_ , \new_[40802]_ , \new_[40803]_ ,
    \new_[40807]_ , \new_[40808]_ , \new_[40811]_ , \new_[40814]_ ,
    \new_[40815]_ , \new_[40816]_ , \new_[40820]_ , \new_[40821]_ ,
    \new_[40825]_ , \new_[40826]_ , \new_[40827]_ , \new_[40831]_ ,
    \new_[40832]_ , \new_[40835]_ , \new_[40838]_ , \new_[40839]_ ,
    \new_[40840]_ , \new_[40844]_ , \new_[40845]_ , \new_[40849]_ ,
    \new_[40850]_ , \new_[40851]_ , \new_[40855]_ , \new_[40856]_ ,
    \new_[40859]_ , \new_[40862]_ , \new_[40863]_ , \new_[40864]_ ,
    \new_[40868]_ , \new_[40869]_ , \new_[40873]_ , \new_[40874]_ ,
    \new_[40875]_ , \new_[40879]_ , \new_[40880]_ , \new_[40883]_ ,
    \new_[40886]_ , \new_[40887]_ , \new_[40888]_ , \new_[40892]_ ,
    \new_[40893]_ , \new_[40897]_ , \new_[40898]_ , \new_[40899]_ ,
    \new_[40903]_ , \new_[40904]_ , \new_[40907]_ , \new_[40910]_ ,
    \new_[40911]_ , \new_[40912]_ , \new_[40916]_ , \new_[40917]_ ,
    \new_[40921]_ , \new_[40922]_ , \new_[40923]_ , \new_[40927]_ ,
    \new_[40928]_ , \new_[40931]_ , \new_[40934]_ , \new_[40935]_ ,
    \new_[40936]_ , \new_[40940]_ , \new_[40941]_ , \new_[40945]_ ,
    \new_[40946]_ , \new_[40947]_ , \new_[40951]_ , \new_[40952]_ ,
    \new_[40955]_ , \new_[40958]_ , \new_[40959]_ , \new_[40960]_ ,
    \new_[40964]_ , \new_[40965]_ , \new_[40969]_ , \new_[40970]_ ,
    \new_[40971]_ , \new_[40975]_ , \new_[40976]_ , \new_[40979]_ ,
    \new_[40982]_ , \new_[40983]_ , \new_[40984]_ , \new_[40988]_ ,
    \new_[40989]_ , \new_[40993]_ , \new_[40994]_ , \new_[40995]_ ,
    \new_[40999]_ , \new_[41000]_ , \new_[41003]_ , \new_[41006]_ ,
    \new_[41007]_ , \new_[41008]_ , \new_[41012]_ , \new_[41013]_ ,
    \new_[41017]_ , \new_[41018]_ , \new_[41019]_ , \new_[41023]_ ,
    \new_[41024]_ , \new_[41027]_ , \new_[41030]_ , \new_[41031]_ ,
    \new_[41032]_ , \new_[41036]_ , \new_[41037]_ , \new_[41041]_ ,
    \new_[41042]_ , \new_[41043]_ , \new_[41047]_ , \new_[41048]_ ,
    \new_[41051]_ , \new_[41054]_ , \new_[41055]_ , \new_[41056]_ ,
    \new_[41060]_ , \new_[41061]_ , \new_[41065]_ , \new_[41066]_ ,
    \new_[41067]_ , \new_[41071]_ , \new_[41072]_ , \new_[41075]_ ,
    \new_[41078]_ , \new_[41079]_ , \new_[41080]_ , \new_[41084]_ ,
    \new_[41085]_ , \new_[41089]_ , \new_[41090]_ , \new_[41091]_ ,
    \new_[41095]_ , \new_[41096]_ , \new_[41099]_ , \new_[41102]_ ,
    \new_[41103]_ , \new_[41104]_ , \new_[41108]_ , \new_[41109]_ ,
    \new_[41113]_ , \new_[41114]_ , \new_[41115]_ , \new_[41119]_ ,
    \new_[41120]_ , \new_[41123]_ , \new_[41126]_ , \new_[41127]_ ,
    \new_[41128]_ , \new_[41132]_ , \new_[41133]_ , \new_[41137]_ ,
    \new_[41138]_ , \new_[41139]_ , \new_[41143]_ , \new_[41144]_ ,
    \new_[41147]_ , \new_[41150]_ , \new_[41151]_ , \new_[41152]_ ,
    \new_[41156]_ , \new_[41157]_ , \new_[41161]_ , \new_[41162]_ ,
    \new_[41163]_ , \new_[41167]_ , \new_[41168]_ , \new_[41171]_ ,
    \new_[41174]_ , \new_[41175]_ , \new_[41176]_ , \new_[41180]_ ,
    \new_[41181]_ , \new_[41185]_ , \new_[41186]_ , \new_[41187]_ ,
    \new_[41191]_ , \new_[41192]_ , \new_[41195]_ , \new_[41198]_ ,
    \new_[41199]_ , \new_[41200]_ , \new_[41204]_ , \new_[41205]_ ,
    \new_[41209]_ , \new_[41210]_ , \new_[41211]_ , \new_[41215]_ ,
    \new_[41216]_ , \new_[41219]_ , \new_[41222]_ , \new_[41223]_ ,
    \new_[41224]_ , \new_[41228]_ , \new_[41229]_ , \new_[41233]_ ,
    \new_[41234]_ , \new_[41235]_ , \new_[41239]_ , \new_[41240]_ ,
    \new_[41243]_ , \new_[41246]_ , \new_[41247]_ , \new_[41248]_ ,
    \new_[41252]_ , \new_[41253]_ , \new_[41257]_ , \new_[41258]_ ,
    \new_[41259]_ , \new_[41263]_ , \new_[41264]_ , \new_[41267]_ ,
    \new_[41270]_ , \new_[41271]_ , \new_[41272]_ , \new_[41276]_ ,
    \new_[41277]_ , \new_[41281]_ , \new_[41282]_ , \new_[41283]_ ,
    \new_[41287]_ , \new_[41288]_ , \new_[41291]_ , \new_[41294]_ ,
    \new_[41295]_ , \new_[41296]_ , \new_[41300]_ , \new_[41301]_ ,
    \new_[41305]_ , \new_[41306]_ , \new_[41307]_ , \new_[41311]_ ,
    \new_[41312]_ , \new_[41315]_ , \new_[41318]_ , \new_[41319]_ ,
    \new_[41320]_ , \new_[41324]_ , \new_[41325]_ , \new_[41329]_ ,
    \new_[41330]_ , \new_[41331]_ , \new_[41335]_ , \new_[41336]_ ,
    \new_[41339]_ , \new_[41342]_ , \new_[41343]_ , \new_[41344]_ ,
    \new_[41348]_ , \new_[41349]_ , \new_[41353]_ , \new_[41354]_ ,
    \new_[41355]_ , \new_[41359]_ , \new_[41360]_ , \new_[41363]_ ,
    \new_[41366]_ , \new_[41367]_ , \new_[41368]_ , \new_[41372]_ ,
    \new_[41373]_ , \new_[41377]_ , \new_[41378]_ , \new_[41379]_ ,
    \new_[41383]_ , \new_[41384]_ , \new_[41387]_ , \new_[41390]_ ,
    \new_[41391]_ , \new_[41392]_ , \new_[41396]_ , \new_[41397]_ ,
    \new_[41401]_ , \new_[41402]_ , \new_[41403]_ , \new_[41407]_ ,
    \new_[41408]_ , \new_[41411]_ , \new_[41414]_ , \new_[41415]_ ,
    \new_[41416]_ , \new_[41420]_ , \new_[41421]_ , \new_[41425]_ ,
    \new_[41426]_ , \new_[41427]_ , \new_[41431]_ , \new_[41432]_ ,
    \new_[41435]_ , \new_[41438]_ , \new_[41439]_ , \new_[41440]_ ,
    \new_[41444]_ , \new_[41445]_ , \new_[41449]_ , \new_[41450]_ ,
    \new_[41451]_ , \new_[41455]_ , \new_[41456]_ , \new_[41459]_ ,
    \new_[41462]_ , \new_[41463]_ , \new_[41464]_ , \new_[41468]_ ,
    \new_[41469]_ , \new_[41473]_ , \new_[41474]_ , \new_[41475]_ ,
    \new_[41479]_ , \new_[41480]_ , \new_[41483]_ , \new_[41486]_ ,
    \new_[41487]_ , \new_[41488]_ , \new_[41492]_ , \new_[41493]_ ,
    \new_[41497]_ , \new_[41498]_ , \new_[41499]_ , \new_[41503]_ ,
    \new_[41504]_ , \new_[41507]_ , \new_[41510]_ , \new_[41511]_ ,
    \new_[41512]_ , \new_[41516]_ , \new_[41517]_ , \new_[41521]_ ,
    \new_[41522]_ , \new_[41523]_ , \new_[41527]_ , \new_[41528]_ ,
    \new_[41531]_ , \new_[41534]_ , \new_[41535]_ , \new_[41536]_ ,
    \new_[41540]_ , \new_[41541]_ , \new_[41545]_ , \new_[41546]_ ,
    \new_[41547]_ , \new_[41551]_ , \new_[41552]_ , \new_[41555]_ ,
    \new_[41558]_ , \new_[41559]_ , \new_[41560]_ , \new_[41564]_ ,
    \new_[41565]_ , \new_[41569]_ , \new_[41570]_ , \new_[41571]_ ,
    \new_[41575]_ , \new_[41576]_ , \new_[41579]_ , \new_[41582]_ ,
    \new_[41583]_ , \new_[41584]_ , \new_[41588]_ , \new_[41589]_ ,
    \new_[41593]_ , \new_[41594]_ , \new_[41595]_ , \new_[41599]_ ,
    \new_[41600]_ , \new_[41603]_ , \new_[41606]_ , \new_[41607]_ ,
    \new_[41608]_ , \new_[41612]_ , \new_[41613]_ , \new_[41617]_ ,
    \new_[41618]_ , \new_[41619]_ , \new_[41623]_ , \new_[41624]_ ,
    \new_[41627]_ , \new_[41630]_ , \new_[41631]_ , \new_[41632]_ ,
    \new_[41636]_ , \new_[41637]_ , \new_[41641]_ , \new_[41642]_ ,
    \new_[41643]_ , \new_[41647]_ , \new_[41648]_ , \new_[41651]_ ,
    \new_[41654]_ , \new_[41655]_ , \new_[41656]_ , \new_[41660]_ ,
    \new_[41661]_ , \new_[41665]_ , \new_[41666]_ , \new_[41667]_ ,
    \new_[41671]_ , \new_[41672]_ , \new_[41675]_ , \new_[41678]_ ,
    \new_[41679]_ , \new_[41680]_ , \new_[41684]_ , \new_[41685]_ ,
    \new_[41689]_ , \new_[41690]_ , \new_[41691]_ , \new_[41695]_ ,
    \new_[41696]_ , \new_[41699]_ , \new_[41702]_ , \new_[41703]_ ,
    \new_[41704]_ , \new_[41708]_ , \new_[41709]_ , \new_[41713]_ ,
    \new_[41714]_ , \new_[41715]_ , \new_[41719]_ , \new_[41720]_ ,
    \new_[41723]_ , \new_[41726]_ , \new_[41727]_ , \new_[41728]_ ,
    \new_[41732]_ , \new_[41733]_ , \new_[41737]_ , \new_[41738]_ ,
    \new_[41739]_ , \new_[41743]_ , \new_[41744]_ , \new_[41747]_ ,
    \new_[41750]_ , \new_[41751]_ , \new_[41752]_ , \new_[41756]_ ,
    \new_[41757]_ , \new_[41761]_ , \new_[41762]_ , \new_[41763]_ ,
    \new_[41767]_ , \new_[41768]_ , \new_[41771]_ , \new_[41774]_ ,
    \new_[41775]_ , \new_[41776]_ , \new_[41780]_ , \new_[41781]_ ,
    \new_[41785]_ , \new_[41786]_ , \new_[41787]_ , \new_[41791]_ ,
    \new_[41792]_ , \new_[41795]_ , \new_[41798]_ , \new_[41799]_ ,
    \new_[41800]_ , \new_[41804]_ , \new_[41805]_ , \new_[41809]_ ,
    \new_[41810]_ , \new_[41811]_ , \new_[41815]_ , \new_[41816]_ ,
    \new_[41819]_ , \new_[41822]_ , \new_[41823]_ , \new_[41824]_ ,
    \new_[41828]_ , \new_[41829]_ , \new_[41833]_ , \new_[41834]_ ,
    \new_[41835]_ , \new_[41839]_ , \new_[41840]_ , \new_[41843]_ ,
    \new_[41846]_ , \new_[41847]_ , \new_[41848]_ , \new_[41852]_ ,
    \new_[41853]_ , \new_[41857]_ , \new_[41858]_ , \new_[41859]_ ,
    \new_[41863]_ , \new_[41864]_ , \new_[41867]_ , \new_[41870]_ ,
    \new_[41871]_ , \new_[41872]_ , \new_[41876]_ , \new_[41877]_ ,
    \new_[41881]_ , \new_[41882]_ , \new_[41883]_ , \new_[41887]_ ,
    \new_[41888]_ , \new_[41891]_ , \new_[41894]_ , \new_[41895]_ ,
    \new_[41896]_ , \new_[41900]_ , \new_[41901]_ , \new_[41905]_ ,
    \new_[41906]_ , \new_[41907]_ , \new_[41911]_ , \new_[41912]_ ,
    \new_[41915]_ , \new_[41918]_ , \new_[41919]_ , \new_[41920]_ ,
    \new_[41924]_ , \new_[41925]_ , \new_[41929]_ , \new_[41930]_ ,
    \new_[41931]_ , \new_[41935]_ , \new_[41936]_ , \new_[41939]_ ,
    \new_[41942]_ , \new_[41943]_ , \new_[41944]_ , \new_[41948]_ ,
    \new_[41949]_ , \new_[41953]_ , \new_[41954]_ , \new_[41955]_ ,
    \new_[41959]_ , \new_[41960]_ , \new_[41963]_ , \new_[41966]_ ,
    \new_[41967]_ , \new_[41968]_ , \new_[41972]_ , \new_[41973]_ ,
    \new_[41977]_ , \new_[41978]_ , \new_[41979]_ , \new_[41983]_ ,
    \new_[41984]_ , \new_[41987]_ , \new_[41990]_ , \new_[41991]_ ,
    \new_[41992]_ , \new_[41996]_ , \new_[41997]_ , \new_[42001]_ ,
    \new_[42002]_ , \new_[42003]_ , \new_[42007]_ , \new_[42008]_ ,
    \new_[42011]_ , \new_[42014]_ , \new_[42015]_ , \new_[42016]_ ,
    \new_[42020]_ , \new_[42021]_ , \new_[42025]_ , \new_[42026]_ ,
    \new_[42027]_ , \new_[42031]_ , \new_[42032]_ , \new_[42035]_ ,
    \new_[42038]_ , \new_[42039]_ , \new_[42040]_ , \new_[42044]_ ,
    \new_[42045]_ , \new_[42049]_ , \new_[42050]_ , \new_[42051]_ ,
    \new_[42055]_ , \new_[42056]_ , \new_[42059]_ , \new_[42062]_ ,
    \new_[42063]_ , \new_[42064]_ , \new_[42068]_ , \new_[42069]_ ,
    \new_[42073]_ , \new_[42074]_ , \new_[42075]_ , \new_[42079]_ ,
    \new_[42080]_ , \new_[42083]_ , \new_[42086]_ , \new_[42087]_ ,
    \new_[42088]_ , \new_[42092]_ , \new_[42093]_ , \new_[42097]_ ,
    \new_[42098]_ , \new_[42099]_ , \new_[42103]_ , \new_[42104]_ ,
    \new_[42107]_ , \new_[42110]_ , \new_[42111]_ , \new_[42112]_ ,
    \new_[42116]_ , \new_[42117]_ , \new_[42121]_ , \new_[42122]_ ,
    \new_[42123]_ , \new_[42127]_ , \new_[42128]_ , \new_[42131]_ ,
    \new_[42134]_ , \new_[42135]_ , \new_[42136]_ , \new_[42140]_ ,
    \new_[42141]_ , \new_[42145]_ , \new_[42146]_ , \new_[42147]_ ,
    \new_[42151]_ , \new_[42152]_ , \new_[42155]_ , \new_[42158]_ ,
    \new_[42159]_ , \new_[42160]_ , \new_[42164]_ , \new_[42165]_ ,
    \new_[42169]_ , \new_[42170]_ , \new_[42171]_ , \new_[42175]_ ,
    \new_[42176]_ , \new_[42179]_ , \new_[42182]_ , \new_[42183]_ ,
    \new_[42184]_ , \new_[42188]_ , \new_[42189]_ , \new_[42193]_ ,
    \new_[42194]_ , \new_[42195]_ , \new_[42199]_ , \new_[42200]_ ,
    \new_[42203]_ , \new_[42206]_ , \new_[42207]_ , \new_[42208]_ ,
    \new_[42212]_ , \new_[42213]_ , \new_[42217]_ , \new_[42218]_ ,
    \new_[42219]_ , \new_[42223]_ , \new_[42224]_ , \new_[42227]_ ,
    \new_[42230]_ , \new_[42231]_ , \new_[42232]_ , \new_[42236]_ ,
    \new_[42237]_ , \new_[42241]_ , \new_[42242]_ , \new_[42243]_ ,
    \new_[42247]_ , \new_[42248]_ , \new_[42251]_ , \new_[42254]_ ,
    \new_[42255]_ , \new_[42256]_ , \new_[42260]_ , \new_[42261]_ ,
    \new_[42265]_ , \new_[42266]_ , \new_[42267]_ , \new_[42271]_ ,
    \new_[42272]_ , \new_[42275]_ , \new_[42278]_ , \new_[42279]_ ,
    \new_[42280]_ , \new_[42284]_ , \new_[42285]_ , \new_[42289]_ ,
    \new_[42290]_ , \new_[42291]_ , \new_[42295]_ , \new_[42296]_ ,
    \new_[42299]_ , \new_[42302]_ , \new_[42303]_ , \new_[42304]_ ,
    \new_[42308]_ , \new_[42309]_ , \new_[42313]_ , \new_[42314]_ ,
    \new_[42315]_ , \new_[42319]_ , \new_[42320]_ , \new_[42323]_ ,
    \new_[42326]_ , \new_[42327]_ , \new_[42328]_ , \new_[42332]_ ,
    \new_[42333]_ , \new_[42337]_ , \new_[42338]_ , \new_[42339]_ ,
    \new_[42343]_ , \new_[42344]_ , \new_[42347]_ , \new_[42350]_ ,
    \new_[42351]_ , \new_[42352]_ , \new_[42356]_ , \new_[42357]_ ,
    \new_[42361]_ , \new_[42362]_ , \new_[42363]_ , \new_[42367]_ ,
    \new_[42368]_ , \new_[42371]_ , \new_[42374]_ , \new_[42375]_ ,
    \new_[42376]_ , \new_[42380]_ , \new_[42381]_ , \new_[42385]_ ,
    \new_[42386]_ , \new_[42387]_ , \new_[42391]_ , \new_[42392]_ ,
    \new_[42395]_ , \new_[42398]_ , \new_[42399]_ , \new_[42400]_ ,
    \new_[42404]_ , \new_[42405]_ , \new_[42409]_ , \new_[42410]_ ,
    \new_[42411]_ , \new_[42415]_ , \new_[42416]_ , \new_[42419]_ ,
    \new_[42422]_ , \new_[42423]_ , \new_[42424]_ , \new_[42428]_ ,
    \new_[42429]_ , \new_[42433]_ , \new_[42434]_ , \new_[42435]_ ,
    \new_[42439]_ , \new_[42440]_ , \new_[42443]_ , \new_[42446]_ ,
    \new_[42447]_ , \new_[42448]_ , \new_[42452]_ , \new_[42453]_ ,
    \new_[42457]_ , \new_[42458]_ , \new_[42459]_ , \new_[42463]_ ,
    \new_[42464]_ , \new_[42467]_ , \new_[42470]_ , \new_[42471]_ ,
    \new_[42472]_ , \new_[42476]_ , \new_[42477]_ , \new_[42481]_ ,
    \new_[42482]_ , \new_[42483]_ , \new_[42487]_ , \new_[42488]_ ,
    \new_[42491]_ , \new_[42494]_ , \new_[42495]_ , \new_[42496]_ ,
    \new_[42500]_ , \new_[42501]_ , \new_[42505]_ , \new_[42506]_ ,
    \new_[42507]_ , \new_[42511]_ , \new_[42512]_ , \new_[42515]_ ,
    \new_[42518]_ , \new_[42519]_ , \new_[42520]_ , \new_[42524]_ ,
    \new_[42525]_ , \new_[42529]_ , \new_[42530]_ , \new_[42531]_ ,
    \new_[42535]_ , \new_[42536]_ , \new_[42539]_ , \new_[42542]_ ,
    \new_[42543]_ , \new_[42544]_ , \new_[42548]_ , \new_[42549]_ ,
    \new_[42553]_ , \new_[42554]_ , \new_[42555]_ , \new_[42559]_ ,
    \new_[42560]_ , \new_[42563]_ , \new_[42566]_ , \new_[42567]_ ,
    \new_[42568]_ , \new_[42572]_ , \new_[42573]_ , \new_[42577]_ ,
    \new_[42578]_ , \new_[42579]_ , \new_[42583]_ , \new_[42584]_ ,
    \new_[42587]_ , \new_[42590]_ , \new_[42591]_ , \new_[42592]_ ,
    \new_[42596]_ , \new_[42597]_ , \new_[42601]_ , \new_[42602]_ ,
    \new_[42603]_ , \new_[42607]_ , \new_[42608]_ , \new_[42611]_ ,
    \new_[42614]_ , \new_[42615]_ , \new_[42616]_ , \new_[42620]_ ,
    \new_[42621]_ , \new_[42625]_ , \new_[42626]_ , \new_[42627]_ ,
    \new_[42631]_ , \new_[42632]_ , \new_[42635]_ , \new_[42638]_ ,
    \new_[42639]_ , \new_[42640]_ , \new_[42644]_ , \new_[42645]_ ,
    \new_[42649]_ , \new_[42650]_ , \new_[42651]_ , \new_[42655]_ ,
    \new_[42656]_ , \new_[42659]_ , \new_[42662]_ , \new_[42663]_ ,
    \new_[42664]_ , \new_[42668]_ , \new_[42669]_ , \new_[42673]_ ,
    \new_[42674]_ , \new_[42675]_ , \new_[42679]_ , \new_[42680]_ ,
    \new_[42683]_ , \new_[42686]_ , \new_[42687]_ , \new_[42688]_ ,
    \new_[42692]_ , \new_[42693]_ , \new_[42697]_ , \new_[42698]_ ,
    \new_[42699]_ , \new_[42703]_ , \new_[42704]_ , \new_[42707]_ ,
    \new_[42710]_ , \new_[42711]_ , \new_[42712]_ , \new_[42716]_ ,
    \new_[42717]_ , \new_[42721]_ , \new_[42722]_ , \new_[42723]_ ,
    \new_[42727]_ , \new_[42728]_ , \new_[42731]_ , \new_[42734]_ ,
    \new_[42735]_ , \new_[42736]_ , \new_[42740]_ , \new_[42741]_ ,
    \new_[42745]_ , \new_[42746]_ , \new_[42747]_ , \new_[42751]_ ,
    \new_[42752]_ , \new_[42755]_ , \new_[42758]_ , \new_[42759]_ ,
    \new_[42760]_ , \new_[42764]_ , \new_[42765]_ , \new_[42769]_ ,
    \new_[42770]_ , \new_[42771]_ , \new_[42775]_ , \new_[42776]_ ,
    \new_[42779]_ , \new_[42782]_ , \new_[42783]_ , \new_[42784]_ ,
    \new_[42788]_ , \new_[42789]_ , \new_[42793]_ , \new_[42794]_ ,
    \new_[42795]_ , \new_[42799]_ , \new_[42800]_ , \new_[42803]_ ,
    \new_[42806]_ , \new_[42807]_ , \new_[42808]_ , \new_[42812]_ ,
    \new_[42813]_ , \new_[42817]_ , \new_[42818]_ , \new_[42819]_ ,
    \new_[42823]_ , \new_[42824]_ , \new_[42827]_ , \new_[42830]_ ,
    \new_[42831]_ , \new_[42832]_ , \new_[42836]_ , \new_[42837]_ ,
    \new_[42841]_ , \new_[42842]_ , \new_[42843]_ , \new_[42847]_ ,
    \new_[42848]_ , \new_[42851]_ , \new_[42854]_ , \new_[42855]_ ,
    \new_[42856]_ , \new_[42860]_ , \new_[42861]_ , \new_[42865]_ ,
    \new_[42866]_ , \new_[42867]_ , \new_[42871]_ , \new_[42872]_ ,
    \new_[42875]_ , \new_[42878]_ , \new_[42879]_ , \new_[42880]_ ,
    \new_[42884]_ , \new_[42885]_ , \new_[42889]_ , \new_[42890]_ ,
    \new_[42891]_ , \new_[42895]_ , \new_[42896]_ , \new_[42899]_ ,
    \new_[42902]_ , \new_[42903]_ , \new_[42904]_ , \new_[42908]_ ,
    \new_[42909]_ , \new_[42913]_ , \new_[42914]_ , \new_[42915]_ ,
    \new_[42919]_ , \new_[42920]_ , \new_[42923]_ , \new_[42926]_ ,
    \new_[42927]_ , \new_[42928]_ , \new_[42932]_ , \new_[42933]_ ,
    \new_[42937]_ , \new_[42938]_ , \new_[42939]_ , \new_[42943]_ ,
    \new_[42944]_ , \new_[42947]_ , \new_[42950]_ , \new_[42951]_ ,
    \new_[42952]_ , \new_[42956]_ , \new_[42957]_ , \new_[42961]_ ,
    \new_[42962]_ , \new_[42963]_ , \new_[42967]_ , \new_[42968]_ ,
    \new_[42971]_ , \new_[42974]_ , \new_[42975]_ , \new_[42976]_ ,
    \new_[42980]_ , \new_[42981]_ , \new_[42985]_ , \new_[42986]_ ,
    \new_[42987]_ , \new_[42991]_ , \new_[42992]_ , \new_[42995]_ ,
    \new_[42998]_ , \new_[42999]_ , \new_[43000]_ , \new_[43004]_ ,
    \new_[43005]_ , \new_[43009]_ , \new_[43010]_ , \new_[43011]_ ,
    \new_[43015]_ , \new_[43016]_ , \new_[43019]_ , \new_[43022]_ ,
    \new_[43023]_ , \new_[43024]_ , \new_[43028]_ , \new_[43029]_ ,
    \new_[43033]_ , \new_[43034]_ , \new_[43035]_ , \new_[43039]_ ,
    \new_[43040]_ , \new_[43043]_ , \new_[43046]_ , \new_[43047]_ ,
    \new_[43048]_ , \new_[43052]_ , \new_[43053]_ , \new_[43057]_ ,
    \new_[43058]_ , \new_[43059]_ , \new_[43063]_ , \new_[43064]_ ,
    \new_[43067]_ , \new_[43070]_ , \new_[43071]_ , \new_[43072]_ ,
    \new_[43076]_ , \new_[43077]_ , \new_[43081]_ , \new_[43082]_ ,
    \new_[43083]_ , \new_[43087]_ , \new_[43088]_ , \new_[43091]_ ,
    \new_[43094]_ , \new_[43095]_ , \new_[43096]_ , \new_[43100]_ ,
    \new_[43101]_ , \new_[43105]_ , \new_[43106]_ , \new_[43107]_ ,
    \new_[43111]_ , \new_[43112]_ , \new_[43115]_ , \new_[43118]_ ,
    \new_[43119]_ , \new_[43120]_ , \new_[43124]_ , \new_[43125]_ ,
    \new_[43129]_ , \new_[43130]_ , \new_[43131]_ , \new_[43135]_ ,
    \new_[43136]_ , \new_[43139]_ , \new_[43142]_ , \new_[43143]_ ,
    \new_[43144]_ , \new_[43148]_ , \new_[43149]_ , \new_[43153]_ ,
    \new_[43154]_ , \new_[43155]_ , \new_[43159]_ , \new_[43160]_ ,
    \new_[43163]_ , \new_[43166]_ , \new_[43167]_ , \new_[43168]_ ,
    \new_[43172]_ , \new_[43173]_ , \new_[43177]_ , \new_[43178]_ ,
    \new_[43179]_ , \new_[43183]_ , \new_[43184]_ , \new_[43187]_ ,
    \new_[43190]_ , \new_[43191]_ , \new_[43192]_ , \new_[43196]_ ,
    \new_[43197]_ , \new_[43201]_ , \new_[43202]_ , \new_[43203]_ ,
    \new_[43207]_ , \new_[43208]_ , \new_[43211]_ , \new_[43214]_ ,
    \new_[43215]_ , \new_[43216]_ , \new_[43220]_ , \new_[43221]_ ,
    \new_[43225]_ , \new_[43226]_ , \new_[43227]_ , \new_[43231]_ ,
    \new_[43232]_ , \new_[43235]_ , \new_[43238]_ , \new_[43239]_ ,
    \new_[43240]_ , \new_[43244]_ , \new_[43245]_ , \new_[43249]_ ,
    \new_[43250]_ , \new_[43251]_ , \new_[43255]_ , \new_[43256]_ ,
    \new_[43259]_ , \new_[43262]_ , \new_[43263]_ , \new_[43264]_ ,
    \new_[43268]_ , \new_[43269]_ , \new_[43273]_ , \new_[43274]_ ,
    \new_[43275]_ , \new_[43279]_ , \new_[43280]_ , \new_[43283]_ ,
    \new_[43286]_ , \new_[43287]_ , \new_[43288]_ , \new_[43292]_ ,
    \new_[43293]_ , \new_[43297]_ , \new_[43298]_ , \new_[43299]_ ,
    \new_[43303]_ , \new_[43304]_ , \new_[43307]_ , \new_[43310]_ ,
    \new_[43311]_ , \new_[43312]_ , \new_[43316]_ , \new_[43317]_ ,
    \new_[43321]_ , \new_[43322]_ , \new_[43323]_ , \new_[43327]_ ,
    \new_[43328]_ , \new_[43331]_ , \new_[43334]_ , \new_[43335]_ ,
    \new_[43336]_ , \new_[43340]_ , \new_[43341]_ , \new_[43345]_ ,
    \new_[43346]_ , \new_[43347]_ , \new_[43351]_ , \new_[43352]_ ,
    \new_[43355]_ , \new_[43358]_ , \new_[43359]_ , \new_[43360]_ ,
    \new_[43364]_ , \new_[43365]_ , \new_[43369]_ , \new_[43370]_ ,
    \new_[43371]_ , \new_[43375]_ , \new_[43376]_ , \new_[43379]_ ,
    \new_[43382]_ , \new_[43383]_ , \new_[43384]_ , \new_[43388]_ ,
    \new_[43389]_ , \new_[43393]_ , \new_[43394]_ , \new_[43395]_ ,
    \new_[43399]_ , \new_[43400]_ , \new_[43403]_ , \new_[43406]_ ,
    \new_[43407]_ , \new_[43408]_ , \new_[43412]_ , \new_[43413]_ ,
    \new_[43417]_ , \new_[43418]_ , \new_[43419]_ , \new_[43423]_ ,
    \new_[43424]_ , \new_[43427]_ , \new_[43430]_ , \new_[43431]_ ,
    \new_[43432]_ , \new_[43436]_ , \new_[43437]_ , \new_[43441]_ ,
    \new_[43442]_ , \new_[43443]_ , \new_[43447]_ , \new_[43448]_ ,
    \new_[43451]_ , \new_[43454]_ , \new_[43455]_ , \new_[43456]_ ,
    \new_[43460]_ , \new_[43461]_ , \new_[43465]_ , \new_[43466]_ ,
    \new_[43467]_ , \new_[43471]_ , \new_[43472]_ , \new_[43475]_ ,
    \new_[43478]_ , \new_[43479]_ , \new_[43480]_ , \new_[43484]_ ,
    \new_[43485]_ , \new_[43489]_ , \new_[43490]_ , \new_[43491]_ ,
    \new_[43495]_ , \new_[43496]_ , \new_[43499]_ , \new_[43502]_ ,
    \new_[43503]_ , \new_[43504]_ , \new_[43508]_ , \new_[43509]_ ,
    \new_[43513]_ , \new_[43514]_ , \new_[43515]_ , \new_[43519]_ ,
    \new_[43520]_ , \new_[43523]_ , \new_[43526]_ , \new_[43527]_ ,
    \new_[43528]_ , \new_[43532]_ , \new_[43533]_ , \new_[43537]_ ,
    \new_[43538]_ , \new_[43539]_ , \new_[43543]_ , \new_[43544]_ ,
    \new_[43547]_ , \new_[43550]_ , \new_[43551]_ , \new_[43552]_ ,
    \new_[43556]_ , \new_[43557]_ , \new_[43561]_ , \new_[43562]_ ,
    \new_[43563]_ , \new_[43567]_ , \new_[43568]_ , \new_[43571]_ ,
    \new_[43574]_ , \new_[43575]_ , \new_[43576]_ , \new_[43580]_ ,
    \new_[43581]_ , \new_[43585]_ , \new_[43586]_ , \new_[43587]_ ,
    \new_[43591]_ , \new_[43592]_ , \new_[43595]_ , \new_[43598]_ ,
    \new_[43599]_ , \new_[43600]_ , \new_[43604]_ , \new_[43605]_ ,
    \new_[43609]_ , \new_[43610]_ , \new_[43611]_ , \new_[43615]_ ,
    \new_[43616]_ , \new_[43619]_ , \new_[43622]_ , \new_[43623]_ ,
    \new_[43624]_ , \new_[43628]_ , \new_[43629]_ , \new_[43633]_ ,
    \new_[43634]_ , \new_[43635]_ , \new_[43639]_ , \new_[43640]_ ,
    \new_[43643]_ , \new_[43646]_ , \new_[43647]_ , \new_[43648]_ ,
    \new_[43652]_ , \new_[43653]_ , \new_[43657]_ , \new_[43658]_ ,
    \new_[43659]_ , \new_[43663]_ , \new_[43664]_ , \new_[43667]_ ,
    \new_[43670]_ , \new_[43671]_ , \new_[43672]_ , \new_[43676]_ ,
    \new_[43677]_ , \new_[43681]_ , \new_[43682]_ , \new_[43683]_ ,
    \new_[43687]_ , \new_[43688]_ , \new_[43691]_ , \new_[43694]_ ,
    \new_[43695]_ , \new_[43696]_ , \new_[43700]_ , \new_[43701]_ ,
    \new_[43705]_ , \new_[43706]_ , \new_[43707]_ , \new_[43711]_ ,
    \new_[43712]_ , \new_[43715]_ , \new_[43718]_ , \new_[43719]_ ,
    \new_[43720]_ , \new_[43724]_ , \new_[43725]_ , \new_[43729]_ ,
    \new_[43730]_ , \new_[43731]_ , \new_[43735]_ , \new_[43736]_ ,
    \new_[43739]_ , \new_[43742]_ , \new_[43743]_ , \new_[43744]_ ,
    \new_[43748]_ , \new_[43749]_ , \new_[43753]_ , \new_[43754]_ ,
    \new_[43755]_ , \new_[43759]_ , \new_[43760]_ , \new_[43763]_ ,
    \new_[43766]_ , \new_[43767]_ , \new_[43768]_ , \new_[43772]_ ,
    \new_[43773]_ , \new_[43777]_ , \new_[43778]_ , \new_[43779]_ ,
    \new_[43783]_ , \new_[43784]_ , \new_[43787]_ , \new_[43790]_ ,
    \new_[43791]_ , \new_[43792]_ , \new_[43796]_ , \new_[43797]_ ,
    \new_[43801]_ , \new_[43802]_ , \new_[43803]_ , \new_[43807]_ ,
    \new_[43808]_ , \new_[43811]_ , \new_[43814]_ , \new_[43815]_ ,
    \new_[43816]_ , \new_[43820]_ , \new_[43821]_ , \new_[43825]_ ,
    \new_[43826]_ , \new_[43827]_ , \new_[43831]_ , \new_[43832]_ ,
    \new_[43835]_ , \new_[43838]_ , \new_[43839]_ , \new_[43840]_ ,
    \new_[43844]_ , \new_[43845]_ , \new_[43849]_ , \new_[43850]_ ,
    \new_[43851]_ , \new_[43855]_ , \new_[43856]_ , \new_[43859]_ ,
    \new_[43862]_ , \new_[43863]_ , \new_[43864]_ , \new_[43868]_ ,
    \new_[43869]_ , \new_[43873]_ , \new_[43874]_ , \new_[43875]_ ,
    \new_[43879]_ , \new_[43880]_ , \new_[43883]_ , \new_[43886]_ ,
    \new_[43887]_ , \new_[43888]_ , \new_[43892]_ , \new_[43893]_ ,
    \new_[43897]_ , \new_[43898]_ , \new_[43899]_ , \new_[43903]_ ,
    \new_[43904]_ , \new_[43907]_ , \new_[43910]_ , \new_[43911]_ ,
    \new_[43912]_ , \new_[43916]_ , \new_[43917]_ , \new_[43921]_ ,
    \new_[43922]_ , \new_[43923]_ , \new_[43927]_ , \new_[43928]_ ,
    \new_[43931]_ , \new_[43934]_ , \new_[43935]_ , \new_[43936]_ ,
    \new_[43940]_ , \new_[43941]_ , \new_[43945]_ , \new_[43946]_ ,
    \new_[43947]_ , \new_[43951]_ , \new_[43952]_ , \new_[43955]_ ,
    \new_[43958]_ , \new_[43959]_ , \new_[43960]_ , \new_[43964]_ ,
    \new_[43965]_ , \new_[43969]_ , \new_[43970]_ , \new_[43971]_ ,
    \new_[43975]_ , \new_[43976]_ , \new_[43979]_ , \new_[43982]_ ,
    \new_[43983]_ , \new_[43984]_ , \new_[43988]_ , \new_[43989]_ ,
    \new_[43993]_ , \new_[43994]_ , \new_[43995]_ , \new_[43999]_ ,
    \new_[44000]_ , \new_[44003]_ , \new_[44006]_ , \new_[44007]_ ,
    \new_[44008]_ , \new_[44012]_ , \new_[44013]_ , \new_[44017]_ ,
    \new_[44018]_ , \new_[44019]_ , \new_[44023]_ , \new_[44024]_ ,
    \new_[44027]_ , \new_[44030]_ , \new_[44031]_ , \new_[44032]_ ,
    \new_[44036]_ , \new_[44037]_ , \new_[44041]_ , \new_[44042]_ ,
    \new_[44043]_ , \new_[44047]_ , \new_[44048]_ , \new_[44051]_ ,
    \new_[44054]_ , \new_[44055]_ , \new_[44056]_ , \new_[44060]_ ,
    \new_[44061]_ , \new_[44065]_ , \new_[44066]_ , \new_[44067]_ ,
    \new_[44071]_ , \new_[44072]_ , \new_[44075]_ , \new_[44078]_ ,
    \new_[44079]_ , \new_[44080]_ , \new_[44084]_ , \new_[44085]_ ,
    \new_[44089]_ , \new_[44090]_ , \new_[44091]_ , \new_[44095]_ ,
    \new_[44096]_ , \new_[44099]_ , \new_[44102]_ , \new_[44103]_ ,
    \new_[44104]_ , \new_[44108]_ , \new_[44109]_ , \new_[44113]_ ,
    \new_[44114]_ , \new_[44115]_ , \new_[44119]_ , \new_[44120]_ ,
    \new_[44123]_ , \new_[44126]_ , \new_[44127]_ , \new_[44128]_ ,
    \new_[44132]_ , \new_[44133]_ , \new_[44137]_ , \new_[44138]_ ,
    \new_[44139]_ , \new_[44143]_ , \new_[44144]_ , \new_[44147]_ ,
    \new_[44150]_ , \new_[44151]_ , \new_[44152]_ , \new_[44156]_ ,
    \new_[44157]_ , \new_[44161]_ , \new_[44162]_ , \new_[44163]_ ,
    \new_[44167]_ , \new_[44168]_ , \new_[44171]_ , \new_[44174]_ ,
    \new_[44175]_ , \new_[44176]_ , \new_[44180]_ , \new_[44181]_ ,
    \new_[44185]_ , \new_[44186]_ , \new_[44187]_ , \new_[44191]_ ,
    \new_[44192]_ , \new_[44195]_ , \new_[44198]_ , \new_[44199]_ ,
    \new_[44200]_ , \new_[44204]_ , \new_[44205]_ , \new_[44209]_ ,
    \new_[44210]_ , \new_[44211]_ , \new_[44215]_ , \new_[44216]_ ,
    \new_[44219]_ , \new_[44222]_ , \new_[44223]_ , \new_[44224]_ ,
    \new_[44228]_ , \new_[44229]_ , \new_[44233]_ , \new_[44234]_ ,
    \new_[44235]_ , \new_[44239]_ , \new_[44240]_ , \new_[44243]_ ,
    \new_[44246]_ , \new_[44247]_ , \new_[44248]_ , \new_[44252]_ ,
    \new_[44253]_ , \new_[44257]_ , \new_[44258]_ , \new_[44259]_ ,
    \new_[44263]_ , \new_[44264]_ , \new_[44267]_ , \new_[44270]_ ,
    \new_[44271]_ , \new_[44272]_ , \new_[44276]_ , \new_[44277]_ ,
    \new_[44281]_ , \new_[44282]_ , \new_[44283]_ , \new_[44287]_ ,
    \new_[44288]_ , \new_[44291]_ , \new_[44294]_ , \new_[44295]_ ,
    \new_[44296]_ , \new_[44300]_ , \new_[44301]_ , \new_[44305]_ ,
    \new_[44306]_ , \new_[44307]_ , \new_[44311]_ , \new_[44312]_ ,
    \new_[44315]_ , \new_[44318]_ , \new_[44319]_ , \new_[44320]_ ,
    \new_[44324]_ , \new_[44325]_ , \new_[44329]_ , \new_[44330]_ ,
    \new_[44331]_ , \new_[44335]_ , \new_[44336]_ , \new_[44339]_ ,
    \new_[44342]_ , \new_[44343]_ , \new_[44344]_ , \new_[44348]_ ,
    \new_[44349]_ , \new_[44353]_ , \new_[44354]_ , \new_[44355]_ ,
    \new_[44359]_ , \new_[44360]_ , \new_[44363]_ , \new_[44366]_ ,
    \new_[44367]_ , \new_[44368]_ , \new_[44372]_ , \new_[44373]_ ,
    \new_[44377]_ , \new_[44378]_ , \new_[44379]_ , \new_[44383]_ ,
    \new_[44384]_ , \new_[44387]_ , \new_[44390]_ , \new_[44391]_ ,
    \new_[44392]_ , \new_[44396]_ , \new_[44397]_ , \new_[44401]_ ,
    \new_[44402]_ , \new_[44403]_ , \new_[44407]_ , \new_[44408]_ ,
    \new_[44411]_ , \new_[44414]_ , \new_[44415]_ , \new_[44416]_ ,
    \new_[44420]_ , \new_[44421]_ , \new_[44425]_ , \new_[44426]_ ,
    \new_[44427]_ , \new_[44431]_ , \new_[44432]_ , \new_[44435]_ ,
    \new_[44438]_ , \new_[44439]_ , \new_[44440]_ , \new_[44444]_ ,
    \new_[44445]_ , \new_[44449]_ , \new_[44450]_ , \new_[44451]_ ,
    \new_[44455]_ , \new_[44456]_ , \new_[44459]_ , \new_[44462]_ ,
    \new_[44463]_ , \new_[44464]_ , \new_[44468]_ , \new_[44469]_ ,
    \new_[44473]_ , \new_[44474]_ , \new_[44475]_ , \new_[44479]_ ,
    \new_[44480]_ , \new_[44483]_ , \new_[44486]_ , \new_[44487]_ ,
    \new_[44488]_ , \new_[44492]_ , \new_[44493]_ , \new_[44497]_ ,
    \new_[44498]_ , \new_[44499]_ , \new_[44503]_ , \new_[44504]_ ,
    \new_[44507]_ , \new_[44510]_ , \new_[44511]_ , \new_[44512]_ ,
    \new_[44516]_ , \new_[44517]_ , \new_[44521]_ , \new_[44522]_ ,
    \new_[44523]_ , \new_[44527]_ , \new_[44528]_ , \new_[44531]_ ,
    \new_[44534]_ , \new_[44535]_ , \new_[44536]_ , \new_[44540]_ ,
    \new_[44541]_ , \new_[44545]_ , \new_[44546]_ , \new_[44547]_ ,
    \new_[44551]_ , \new_[44552]_ , \new_[44555]_ , \new_[44558]_ ,
    \new_[44559]_ , \new_[44560]_ , \new_[44564]_ , \new_[44565]_ ,
    \new_[44569]_ , \new_[44570]_ , \new_[44571]_ , \new_[44575]_ ,
    \new_[44576]_ , \new_[44579]_ , \new_[44582]_ , \new_[44583]_ ,
    \new_[44584]_ , \new_[44588]_ , \new_[44589]_ , \new_[44593]_ ,
    \new_[44594]_ , \new_[44595]_ , \new_[44599]_ , \new_[44600]_ ,
    \new_[44603]_ , \new_[44606]_ , \new_[44607]_ , \new_[44608]_ ,
    \new_[44612]_ , \new_[44613]_ , \new_[44617]_ , \new_[44618]_ ,
    \new_[44619]_ , \new_[44623]_ , \new_[44624]_ , \new_[44627]_ ,
    \new_[44630]_ , \new_[44631]_ , \new_[44632]_ , \new_[44636]_ ,
    \new_[44637]_ , \new_[44641]_ , \new_[44642]_ , \new_[44643]_ ,
    \new_[44647]_ , \new_[44648]_ , \new_[44651]_ , \new_[44654]_ ,
    \new_[44655]_ , \new_[44656]_ , \new_[44660]_ , \new_[44661]_ ,
    \new_[44665]_ , \new_[44666]_ , \new_[44667]_ , \new_[44671]_ ,
    \new_[44672]_ , \new_[44675]_ , \new_[44678]_ , \new_[44679]_ ,
    \new_[44680]_ , \new_[44684]_ , \new_[44685]_ , \new_[44689]_ ,
    \new_[44690]_ , \new_[44691]_ , \new_[44695]_ , \new_[44696]_ ,
    \new_[44699]_ , \new_[44702]_ , \new_[44703]_ , \new_[44704]_ ,
    \new_[44708]_ , \new_[44709]_ , \new_[44713]_ , \new_[44714]_ ,
    \new_[44715]_ , \new_[44719]_ , \new_[44720]_ , \new_[44723]_ ,
    \new_[44726]_ , \new_[44727]_ , \new_[44728]_ , \new_[44732]_ ,
    \new_[44733]_ , \new_[44737]_ , \new_[44738]_ , \new_[44739]_ ,
    \new_[44743]_ , \new_[44744]_ , \new_[44747]_ , \new_[44750]_ ,
    \new_[44751]_ , \new_[44752]_ , \new_[44756]_ , \new_[44757]_ ,
    \new_[44761]_ , \new_[44762]_ , \new_[44763]_ , \new_[44767]_ ,
    \new_[44768]_ , \new_[44771]_ , \new_[44774]_ , \new_[44775]_ ,
    \new_[44776]_ , \new_[44780]_ , \new_[44781]_ , \new_[44785]_ ,
    \new_[44786]_ , \new_[44787]_ , \new_[44791]_ , \new_[44792]_ ,
    \new_[44795]_ , \new_[44798]_ , \new_[44799]_ , \new_[44800]_ ,
    \new_[44804]_ , \new_[44805]_ , \new_[44809]_ , \new_[44810]_ ,
    \new_[44811]_ , \new_[44815]_ , \new_[44816]_ , \new_[44819]_ ,
    \new_[44822]_ , \new_[44823]_ , \new_[44824]_ , \new_[44828]_ ,
    \new_[44829]_ , \new_[44833]_ , \new_[44834]_ , \new_[44835]_ ,
    \new_[44839]_ , \new_[44840]_ , \new_[44843]_ , \new_[44846]_ ,
    \new_[44847]_ , \new_[44848]_ , \new_[44852]_ , \new_[44853]_ ,
    \new_[44857]_ , \new_[44858]_ , \new_[44859]_ , \new_[44863]_ ,
    \new_[44864]_ , \new_[44867]_ , \new_[44870]_ , \new_[44871]_ ,
    \new_[44872]_ , \new_[44876]_ , \new_[44877]_ , \new_[44881]_ ,
    \new_[44882]_ , \new_[44883]_ , \new_[44887]_ , \new_[44888]_ ,
    \new_[44891]_ , \new_[44894]_ , \new_[44895]_ , \new_[44896]_ ,
    \new_[44900]_ , \new_[44901]_ , \new_[44905]_ , \new_[44906]_ ,
    \new_[44907]_ , \new_[44911]_ , \new_[44912]_ , \new_[44915]_ ,
    \new_[44918]_ , \new_[44919]_ , \new_[44920]_ , \new_[44924]_ ,
    \new_[44925]_ , \new_[44929]_ , \new_[44930]_ , \new_[44931]_ ,
    \new_[44935]_ , \new_[44936]_ , \new_[44939]_ , \new_[44942]_ ,
    \new_[44943]_ , \new_[44944]_ , \new_[44948]_ , \new_[44949]_ ,
    \new_[44953]_ , \new_[44954]_ , \new_[44955]_ , \new_[44959]_ ,
    \new_[44960]_ , \new_[44963]_ , \new_[44966]_ , \new_[44967]_ ,
    \new_[44968]_ , \new_[44972]_ , \new_[44973]_ , \new_[44977]_ ,
    \new_[44978]_ , \new_[44979]_ , \new_[44983]_ , \new_[44984]_ ,
    \new_[44987]_ , \new_[44990]_ , \new_[44991]_ , \new_[44992]_ ,
    \new_[44996]_ , \new_[44997]_ , \new_[45001]_ , \new_[45002]_ ,
    \new_[45003]_ , \new_[45007]_ , \new_[45008]_ , \new_[45011]_ ,
    \new_[45014]_ , \new_[45015]_ , \new_[45016]_ , \new_[45020]_ ,
    \new_[45021]_ , \new_[45025]_ , \new_[45026]_ , \new_[45027]_ ,
    \new_[45031]_ , \new_[45032]_ , \new_[45035]_ , \new_[45038]_ ,
    \new_[45039]_ , \new_[45040]_ , \new_[45044]_ , \new_[45045]_ ,
    \new_[45049]_ , \new_[45050]_ , \new_[45051]_ , \new_[45055]_ ,
    \new_[45056]_ , \new_[45059]_ , \new_[45062]_ , \new_[45063]_ ,
    \new_[45064]_ , \new_[45068]_ , \new_[45069]_ , \new_[45073]_ ,
    \new_[45074]_ , \new_[45075]_ , \new_[45079]_ , \new_[45080]_ ,
    \new_[45083]_ , \new_[45086]_ , \new_[45087]_ , \new_[45088]_ ,
    \new_[45092]_ , \new_[45093]_ , \new_[45097]_ , \new_[45098]_ ,
    \new_[45099]_ , \new_[45103]_ , \new_[45104]_ , \new_[45107]_ ,
    \new_[45110]_ , \new_[45111]_ , \new_[45112]_ , \new_[45116]_ ,
    \new_[45117]_ , \new_[45121]_ , \new_[45122]_ , \new_[45123]_ ,
    \new_[45127]_ , \new_[45128]_ , \new_[45131]_ , \new_[45134]_ ,
    \new_[45135]_ , \new_[45136]_ , \new_[45140]_ , \new_[45141]_ ,
    \new_[45145]_ , \new_[45146]_ , \new_[45147]_ , \new_[45151]_ ,
    \new_[45152]_ , \new_[45155]_ , \new_[45158]_ , \new_[45159]_ ,
    \new_[45160]_ , \new_[45164]_ , \new_[45165]_ , \new_[45169]_ ,
    \new_[45170]_ , \new_[45171]_ , \new_[45175]_ , \new_[45176]_ ,
    \new_[45179]_ , \new_[45182]_ , \new_[45183]_ , \new_[45184]_ ,
    \new_[45188]_ , \new_[45189]_ , \new_[45193]_ , \new_[45194]_ ,
    \new_[45195]_ , \new_[45199]_ , \new_[45200]_ , \new_[45203]_ ,
    \new_[45206]_ , \new_[45207]_ , \new_[45208]_ , \new_[45212]_ ,
    \new_[45213]_ , \new_[45217]_ , \new_[45218]_ , \new_[45219]_ ,
    \new_[45223]_ , \new_[45224]_ , \new_[45227]_ , \new_[45230]_ ,
    \new_[45231]_ , \new_[45232]_ , \new_[45236]_ , \new_[45237]_ ,
    \new_[45241]_ , \new_[45242]_ , \new_[45243]_ , \new_[45247]_ ,
    \new_[45248]_ , \new_[45251]_ , \new_[45254]_ , \new_[45255]_ ,
    \new_[45256]_ , \new_[45260]_ , \new_[45261]_ , \new_[45265]_ ,
    \new_[45266]_ , \new_[45267]_ , \new_[45271]_ , \new_[45272]_ ,
    \new_[45275]_ , \new_[45278]_ , \new_[45279]_ , \new_[45280]_ ,
    \new_[45284]_ , \new_[45285]_ , \new_[45289]_ , \new_[45290]_ ,
    \new_[45291]_ , \new_[45295]_ , \new_[45296]_ , \new_[45299]_ ,
    \new_[45302]_ , \new_[45303]_ , \new_[45304]_ , \new_[45308]_ ,
    \new_[45309]_ , \new_[45313]_ , \new_[45314]_ , \new_[45315]_ ,
    \new_[45319]_ , \new_[45320]_ , \new_[45323]_ , \new_[45326]_ ,
    \new_[45327]_ , \new_[45328]_ , \new_[45332]_ , \new_[45333]_ ,
    \new_[45337]_ , \new_[45338]_ , \new_[45339]_ , \new_[45343]_ ,
    \new_[45344]_ , \new_[45347]_ , \new_[45350]_ , \new_[45351]_ ,
    \new_[45352]_ , \new_[45356]_ , \new_[45357]_ , \new_[45361]_ ,
    \new_[45362]_ , \new_[45363]_ , \new_[45367]_ , \new_[45368]_ ,
    \new_[45371]_ , \new_[45374]_ , \new_[45375]_ , \new_[45376]_ ,
    \new_[45380]_ , \new_[45381]_ , \new_[45385]_ , \new_[45386]_ ,
    \new_[45387]_ , \new_[45391]_ , \new_[45392]_ , \new_[45395]_ ,
    \new_[45398]_ , \new_[45399]_ , \new_[45400]_ , \new_[45404]_ ,
    \new_[45405]_ , \new_[45409]_ , \new_[45410]_ , \new_[45411]_ ,
    \new_[45415]_ , \new_[45416]_ , \new_[45419]_ , \new_[45422]_ ,
    \new_[45423]_ , \new_[45424]_ , \new_[45428]_ , \new_[45429]_ ,
    \new_[45433]_ , \new_[45434]_ , \new_[45435]_ , \new_[45439]_ ,
    \new_[45440]_ , \new_[45443]_ , \new_[45446]_ , \new_[45447]_ ,
    \new_[45448]_ , \new_[45452]_ , \new_[45453]_ , \new_[45457]_ ,
    \new_[45458]_ , \new_[45459]_ , \new_[45463]_ , \new_[45464]_ ,
    \new_[45467]_ , \new_[45470]_ , \new_[45471]_ , \new_[45472]_ ,
    \new_[45476]_ , \new_[45477]_ , \new_[45481]_ , \new_[45482]_ ,
    \new_[45483]_ , \new_[45487]_ , \new_[45488]_ , \new_[45491]_ ,
    \new_[45494]_ , \new_[45495]_ , \new_[45496]_ , \new_[45500]_ ,
    \new_[45501]_ , \new_[45505]_ , \new_[45506]_ , \new_[45507]_ ,
    \new_[45511]_ , \new_[45512]_ , \new_[45515]_ , \new_[45518]_ ,
    \new_[45519]_ , \new_[45520]_ , \new_[45524]_ , \new_[45525]_ ,
    \new_[45529]_ , \new_[45530]_ , \new_[45531]_ , \new_[45535]_ ,
    \new_[45536]_ , \new_[45539]_ , \new_[45542]_ , \new_[45543]_ ,
    \new_[45544]_ , \new_[45548]_ , \new_[45549]_ , \new_[45553]_ ,
    \new_[45554]_ , \new_[45555]_ , \new_[45559]_ , \new_[45560]_ ,
    \new_[45563]_ , \new_[45566]_ , \new_[45567]_ , \new_[45568]_ ,
    \new_[45572]_ , \new_[45573]_ , \new_[45577]_ , \new_[45578]_ ,
    \new_[45579]_ , \new_[45583]_ , \new_[45584]_ , \new_[45587]_ ,
    \new_[45590]_ , \new_[45591]_ , \new_[45592]_ , \new_[45596]_ ,
    \new_[45597]_ , \new_[45601]_ , \new_[45602]_ , \new_[45603]_ ,
    \new_[45607]_ , \new_[45608]_ , \new_[45611]_ , \new_[45614]_ ,
    \new_[45615]_ , \new_[45616]_ , \new_[45620]_ , \new_[45621]_ ,
    \new_[45625]_ , \new_[45626]_ , \new_[45627]_ , \new_[45631]_ ,
    \new_[45632]_ , \new_[45635]_ , \new_[45638]_ , \new_[45639]_ ,
    \new_[45640]_ , \new_[45644]_ , \new_[45645]_ , \new_[45649]_ ,
    \new_[45650]_ , \new_[45651]_ , \new_[45655]_ , \new_[45656]_ ,
    \new_[45659]_ , \new_[45662]_ , \new_[45663]_ , \new_[45664]_ ,
    \new_[45668]_ , \new_[45669]_ , \new_[45673]_ , \new_[45674]_ ,
    \new_[45675]_ , \new_[45679]_ , \new_[45680]_ , \new_[45683]_ ,
    \new_[45686]_ , \new_[45687]_ , \new_[45688]_ , \new_[45692]_ ,
    \new_[45693]_ , \new_[45697]_ , \new_[45698]_ , \new_[45699]_ ,
    \new_[45703]_ , \new_[45704]_ , \new_[45707]_ , \new_[45710]_ ,
    \new_[45711]_ , \new_[45712]_ , \new_[45716]_ , \new_[45717]_ ,
    \new_[45721]_ , \new_[45722]_ , \new_[45723]_ , \new_[45727]_ ,
    \new_[45728]_ , \new_[45731]_ , \new_[45734]_ , \new_[45735]_ ,
    \new_[45736]_ , \new_[45740]_ , \new_[45741]_ , \new_[45745]_ ,
    \new_[45746]_ , \new_[45747]_ , \new_[45751]_ , \new_[45752]_ ,
    \new_[45755]_ , \new_[45758]_ , \new_[45759]_ , \new_[45760]_ ,
    \new_[45764]_ , \new_[45765]_ , \new_[45769]_ , \new_[45770]_ ,
    \new_[45771]_ , \new_[45775]_ , \new_[45776]_ , \new_[45779]_ ,
    \new_[45782]_ , \new_[45783]_ , \new_[45784]_ , \new_[45788]_ ,
    \new_[45789]_ , \new_[45793]_ , \new_[45794]_ , \new_[45795]_ ,
    \new_[45799]_ , \new_[45800]_ , \new_[45803]_ , \new_[45806]_ ,
    \new_[45807]_ , \new_[45808]_ , \new_[45812]_ , \new_[45813]_ ,
    \new_[45817]_ , \new_[45818]_ , \new_[45819]_ , \new_[45823]_ ,
    \new_[45824]_ , \new_[45827]_ , \new_[45830]_ , \new_[45831]_ ,
    \new_[45832]_ , \new_[45836]_ , \new_[45837]_ , \new_[45841]_ ,
    \new_[45842]_ , \new_[45843]_ , \new_[45847]_ , \new_[45848]_ ,
    \new_[45851]_ , \new_[45854]_ , \new_[45855]_ , \new_[45856]_ ,
    \new_[45860]_ , \new_[45861]_ , \new_[45865]_ , \new_[45866]_ ,
    \new_[45867]_ , \new_[45871]_ , \new_[45872]_ , \new_[45875]_ ,
    \new_[45878]_ , \new_[45879]_ , \new_[45880]_ , \new_[45884]_ ,
    \new_[45885]_ , \new_[45889]_ , \new_[45890]_ , \new_[45891]_ ,
    \new_[45895]_ , \new_[45896]_ , \new_[45899]_ , \new_[45902]_ ,
    \new_[45903]_ , \new_[45904]_ , \new_[45908]_ , \new_[45909]_ ,
    \new_[45913]_ , \new_[45914]_ , \new_[45915]_ , \new_[45919]_ ,
    \new_[45920]_ , \new_[45923]_ , \new_[45926]_ , \new_[45927]_ ,
    \new_[45928]_ , \new_[45932]_ , \new_[45933]_ , \new_[45937]_ ,
    \new_[45938]_ , \new_[45939]_ , \new_[45943]_ , \new_[45944]_ ,
    \new_[45947]_ , \new_[45950]_ , \new_[45951]_ , \new_[45952]_ ,
    \new_[45956]_ , \new_[45957]_ , \new_[45961]_ , \new_[45962]_ ,
    \new_[45963]_ , \new_[45967]_ , \new_[45968]_ , \new_[45971]_ ,
    \new_[45974]_ , \new_[45975]_ , \new_[45976]_ , \new_[45980]_ ,
    \new_[45981]_ , \new_[45985]_ , \new_[45986]_ , \new_[45987]_ ,
    \new_[45991]_ , \new_[45992]_ , \new_[45995]_ , \new_[45998]_ ,
    \new_[45999]_ , \new_[46000]_ , \new_[46004]_ , \new_[46005]_ ,
    \new_[46009]_ , \new_[46010]_ , \new_[46011]_ , \new_[46015]_ ,
    \new_[46016]_ , \new_[46019]_ , \new_[46022]_ , \new_[46023]_ ,
    \new_[46024]_ , \new_[46028]_ , \new_[46029]_ , \new_[46033]_ ,
    \new_[46034]_ , \new_[46035]_ , \new_[46039]_ , \new_[46040]_ ,
    \new_[46043]_ , \new_[46046]_ , \new_[46047]_ , \new_[46048]_ ,
    \new_[46052]_ , \new_[46053]_ , \new_[46057]_ , \new_[46058]_ ,
    \new_[46059]_ , \new_[46063]_ , \new_[46064]_ , \new_[46067]_ ,
    \new_[46070]_ , \new_[46071]_ , \new_[46072]_ , \new_[46076]_ ,
    \new_[46077]_ , \new_[46081]_ , \new_[46082]_ , \new_[46083]_ ,
    \new_[46087]_ , \new_[46088]_ , \new_[46091]_ , \new_[46094]_ ,
    \new_[46095]_ , \new_[46096]_ , \new_[46100]_ , \new_[46101]_ ,
    \new_[46105]_ , \new_[46106]_ , \new_[46107]_ , \new_[46111]_ ,
    \new_[46112]_ , \new_[46115]_ , \new_[46118]_ , \new_[46119]_ ,
    \new_[46120]_ , \new_[46124]_ , \new_[46125]_ , \new_[46129]_ ,
    \new_[46130]_ , \new_[46131]_ , \new_[46135]_ , \new_[46136]_ ,
    \new_[46139]_ , \new_[46142]_ , \new_[46143]_ , \new_[46144]_ ,
    \new_[46148]_ , \new_[46149]_ , \new_[46153]_ , \new_[46154]_ ,
    \new_[46155]_ , \new_[46159]_ , \new_[46160]_ , \new_[46163]_ ,
    \new_[46166]_ , \new_[46167]_ , \new_[46168]_ , \new_[46172]_ ,
    \new_[46173]_ , \new_[46177]_ , \new_[46178]_ , \new_[46179]_ ,
    \new_[46183]_ , \new_[46184]_ , \new_[46187]_ , \new_[46190]_ ,
    \new_[46191]_ , \new_[46192]_ , \new_[46196]_ , \new_[46197]_ ,
    \new_[46201]_ , \new_[46202]_ , \new_[46203]_ , \new_[46207]_ ,
    \new_[46208]_ , \new_[46211]_ , \new_[46214]_ , \new_[46215]_ ,
    \new_[46216]_ , \new_[46220]_ , \new_[46221]_ , \new_[46225]_ ,
    \new_[46226]_ , \new_[46227]_ , \new_[46231]_ , \new_[46232]_ ,
    \new_[46235]_ , \new_[46238]_ , \new_[46239]_ , \new_[46240]_ ,
    \new_[46244]_ , \new_[46245]_ , \new_[46249]_ , \new_[46250]_ ,
    \new_[46251]_ , \new_[46255]_ , \new_[46256]_ , \new_[46259]_ ,
    \new_[46262]_ , \new_[46263]_ , \new_[46264]_ , \new_[46268]_ ,
    \new_[46269]_ , \new_[46273]_ , \new_[46274]_ , \new_[46275]_ ,
    \new_[46279]_ , \new_[46280]_ , \new_[46283]_ , \new_[46286]_ ,
    \new_[46287]_ , \new_[46288]_ , \new_[46292]_ , \new_[46293]_ ,
    \new_[46297]_ , \new_[46298]_ , \new_[46299]_ , \new_[46303]_ ,
    \new_[46304]_ , \new_[46307]_ , \new_[46310]_ , \new_[46311]_ ,
    \new_[46312]_ , \new_[46316]_ , \new_[46317]_ , \new_[46321]_ ,
    \new_[46322]_ , \new_[46323]_ , \new_[46327]_ , \new_[46328]_ ,
    \new_[46331]_ , \new_[46334]_ , \new_[46335]_ , \new_[46336]_ ,
    \new_[46340]_ , \new_[46341]_ , \new_[46345]_ , \new_[46346]_ ,
    \new_[46347]_ , \new_[46351]_ , \new_[46352]_ , \new_[46355]_ ,
    \new_[46358]_ , \new_[46359]_ , \new_[46360]_ , \new_[46364]_ ,
    \new_[46365]_ , \new_[46369]_ , \new_[46370]_ , \new_[46371]_ ,
    \new_[46375]_ , \new_[46376]_ , \new_[46379]_ , \new_[46382]_ ,
    \new_[46383]_ , \new_[46384]_ , \new_[46388]_ , \new_[46389]_ ,
    \new_[46393]_ , \new_[46394]_ , \new_[46395]_ , \new_[46399]_ ,
    \new_[46400]_ , \new_[46403]_ , \new_[46406]_ , \new_[46407]_ ,
    \new_[46408]_ , \new_[46412]_ , \new_[46413]_ , \new_[46417]_ ,
    \new_[46418]_ , \new_[46419]_ , \new_[46423]_ , \new_[46424]_ ,
    \new_[46427]_ , \new_[46430]_ , \new_[46431]_ , \new_[46432]_ ,
    \new_[46436]_ , \new_[46437]_ , \new_[46441]_ , \new_[46442]_ ,
    \new_[46443]_ , \new_[46447]_ , \new_[46448]_ , \new_[46451]_ ,
    \new_[46454]_ , \new_[46455]_ , \new_[46456]_ , \new_[46460]_ ,
    \new_[46461]_ , \new_[46465]_ , \new_[46466]_ , \new_[46467]_ ,
    \new_[46471]_ , \new_[46472]_ , \new_[46475]_ , \new_[46478]_ ,
    \new_[46479]_ , \new_[46480]_ , \new_[46484]_ , \new_[46485]_ ,
    \new_[46489]_ , \new_[46490]_ , \new_[46491]_ , \new_[46495]_ ,
    \new_[46496]_ , \new_[46499]_ , \new_[46502]_ , \new_[46503]_ ,
    \new_[46504]_ , \new_[46508]_ , \new_[46509]_ , \new_[46513]_ ,
    \new_[46514]_ , \new_[46515]_ , \new_[46519]_ , \new_[46520]_ ,
    \new_[46523]_ , \new_[46526]_ , \new_[46527]_ , \new_[46528]_ ,
    \new_[46532]_ , \new_[46533]_ , \new_[46537]_ , \new_[46538]_ ,
    \new_[46539]_ , \new_[46543]_ , \new_[46544]_ , \new_[46547]_ ,
    \new_[46550]_ , \new_[46551]_ , \new_[46552]_ , \new_[46556]_ ,
    \new_[46557]_ , \new_[46561]_ , \new_[46562]_ , \new_[46563]_ ,
    \new_[46567]_ , \new_[46568]_ , \new_[46571]_ , \new_[46574]_ ,
    \new_[46575]_ , \new_[46576]_ , \new_[46580]_ , \new_[46581]_ ,
    \new_[46585]_ , \new_[46586]_ , \new_[46587]_ , \new_[46591]_ ,
    \new_[46592]_ , \new_[46595]_ , \new_[46598]_ , \new_[46599]_ ,
    \new_[46600]_ , \new_[46604]_ , \new_[46605]_ , \new_[46609]_ ,
    \new_[46610]_ , \new_[46611]_ , \new_[46615]_ , \new_[46616]_ ,
    \new_[46619]_ , \new_[46622]_ , \new_[46623]_ , \new_[46624]_ ,
    \new_[46628]_ , \new_[46629]_ , \new_[46633]_ , \new_[46634]_ ,
    \new_[46635]_ , \new_[46639]_ , \new_[46640]_ , \new_[46643]_ ,
    \new_[46646]_ , \new_[46647]_ , \new_[46648]_ , \new_[46652]_ ,
    \new_[46653]_ , \new_[46657]_ , \new_[46658]_ , \new_[46659]_ ,
    \new_[46663]_ , \new_[46664]_ , \new_[46667]_ , \new_[46670]_ ,
    \new_[46671]_ , \new_[46672]_ , \new_[46676]_ , \new_[46677]_ ,
    \new_[46681]_ , \new_[46682]_ , \new_[46683]_ , \new_[46687]_ ,
    \new_[46688]_ , \new_[46691]_ , \new_[46694]_ , \new_[46695]_ ,
    \new_[46696]_ , \new_[46700]_ , \new_[46701]_ , \new_[46705]_ ,
    \new_[46706]_ , \new_[46707]_ , \new_[46711]_ , \new_[46712]_ ,
    \new_[46715]_ , \new_[46718]_ , \new_[46719]_ , \new_[46720]_ ,
    \new_[46724]_ , \new_[46725]_ , \new_[46729]_ , \new_[46730]_ ,
    \new_[46731]_ , \new_[46735]_ , \new_[46736]_ , \new_[46739]_ ,
    \new_[46742]_ , \new_[46743]_ , \new_[46744]_ , \new_[46748]_ ,
    \new_[46749]_ , \new_[46753]_ , \new_[46754]_ , \new_[46755]_ ,
    \new_[46759]_ , \new_[46760]_ , \new_[46763]_ , \new_[46766]_ ,
    \new_[46767]_ , \new_[46768]_ , \new_[46772]_ , \new_[46773]_ ,
    \new_[46777]_ , \new_[46778]_ , \new_[46779]_ , \new_[46783]_ ,
    \new_[46784]_ , \new_[46787]_ , \new_[46790]_ , \new_[46791]_ ,
    \new_[46792]_ , \new_[46796]_ , \new_[46797]_ , \new_[46801]_ ,
    \new_[46802]_ , \new_[46803]_ , \new_[46807]_ , \new_[46808]_ ,
    \new_[46811]_ , \new_[46814]_ , \new_[46815]_ , \new_[46816]_ ,
    \new_[46820]_ , \new_[46821]_ , \new_[46825]_ , \new_[46826]_ ,
    \new_[46827]_ , \new_[46831]_ , \new_[46832]_ , \new_[46835]_ ,
    \new_[46838]_ , \new_[46839]_ , \new_[46840]_ , \new_[46844]_ ,
    \new_[46845]_ , \new_[46849]_ , \new_[46850]_ , \new_[46851]_ ,
    \new_[46855]_ , \new_[46856]_ , \new_[46859]_ , \new_[46862]_ ,
    \new_[46863]_ , \new_[46864]_ , \new_[46868]_ , \new_[46869]_ ,
    \new_[46873]_ , \new_[46874]_ , \new_[46875]_ , \new_[46879]_ ,
    \new_[46880]_ , \new_[46883]_ , \new_[46886]_ , \new_[46887]_ ,
    \new_[46888]_ , \new_[46892]_ , \new_[46893]_ , \new_[46897]_ ,
    \new_[46898]_ , \new_[46899]_ , \new_[46903]_ , \new_[46904]_ ,
    \new_[46907]_ , \new_[46910]_ , \new_[46911]_ , \new_[46912]_ ,
    \new_[46916]_ , \new_[46917]_ , \new_[46921]_ , \new_[46922]_ ,
    \new_[46923]_ , \new_[46927]_ , \new_[46928]_ , \new_[46931]_ ,
    \new_[46934]_ , \new_[46935]_ , \new_[46936]_ , \new_[46940]_ ,
    \new_[46941]_ , \new_[46945]_ , \new_[46946]_ , \new_[46947]_ ,
    \new_[46951]_ , \new_[46952]_ , \new_[46955]_ , \new_[46958]_ ,
    \new_[46959]_ , \new_[46960]_ , \new_[46964]_ , \new_[46965]_ ,
    \new_[46969]_ , \new_[46970]_ , \new_[46971]_ , \new_[46975]_ ,
    \new_[46976]_ , \new_[46979]_ , \new_[46982]_ , \new_[46983]_ ,
    \new_[46984]_ , \new_[46988]_ , \new_[46989]_ , \new_[46993]_ ,
    \new_[46994]_ , \new_[46995]_ , \new_[46999]_ , \new_[47000]_ ,
    \new_[47003]_ , \new_[47006]_ , \new_[47007]_ , \new_[47008]_ ,
    \new_[47012]_ , \new_[47013]_ , \new_[47017]_ , \new_[47018]_ ,
    \new_[47019]_ , \new_[47023]_ , \new_[47024]_ , \new_[47027]_ ,
    \new_[47030]_ , \new_[47031]_ , \new_[47032]_ , \new_[47036]_ ,
    \new_[47037]_ , \new_[47041]_ , \new_[47042]_ , \new_[47043]_ ,
    \new_[47047]_ , \new_[47048]_ , \new_[47051]_ , \new_[47054]_ ,
    \new_[47055]_ , \new_[47056]_ , \new_[47060]_ , \new_[47061]_ ,
    \new_[47065]_ , \new_[47066]_ , \new_[47067]_ , \new_[47071]_ ,
    \new_[47072]_ , \new_[47075]_ , \new_[47078]_ , \new_[47079]_ ,
    \new_[47080]_ , \new_[47084]_ , \new_[47085]_ , \new_[47089]_ ,
    \new_[47090]_ , \new_[47091]_ , \new_[47095]_ , \new_[47096]_ ,
    \new_[47099]_ , \new_[47102]_ , \new_[47103]_ , \new_[47104]_ ,
    \new_[47108]_ , \new_[47109]_ , \new_[47113]_ , \new_[47114]_ ,
    \new_[47115]_ , \new_[47119]_ , \new_[47120]_ , \new_[47123]_ ,
    \new_[47126]_ , \new_[47127]_ , \new_[47128]_ , \new_[47132]_ ,
    \new_[47133]_ , \new_[47137]_ , \new_[47138]_ , \new_[47139]_ ,
    \new_[47143]_ , \new_[47144]_ , \new_[47147]_ , \new_[47150]_ ,
    \new_[47151]_ , \new_[47152]_ , \new_[47156]_ , \new_[47157]_ ,
    \new_[47161]_ , \new_[47162]_ , \new_[47163]_ , \new_[47167]_ ,
    \new_[47168]_ , \new_[47171]_ , \new_[47174]_ , \new_[47175]_ ,
    \new_[47176]_ , \new_[47180]_ , \new_[47181]_ , \new_[47185]_ ,
    \new_[47186]_ , \new_[47187]_ , \new_[47191]_ , \new_[47192]_ ,
    \new_[47195]_ , \new_[47198]_ , \new_[47199]_ , \new_[47200]_ ,
    \new_[47204]_ , \new_[47205]_ , \new_[47209]_ , \new_[47210]_ ,
    \new_[47211]_ , \new_[47215]_ , \new_[47216]_ , \new_[47219]_ ,
    \new_[47222]_ , \new_[47223]_ , \new_[47224]_ , \new_[47228]_ ,
    \new_[47229]_ , \new_[47233]_ , \new_[47234]_ , \new_[47235]_ ,
    \new_[47239]_ , \new_[47240]_ , \new_[47243]_ , \new_[47246]_ ,
    \new_[47247]_ , \new_[47248]_ , \new_[47252]_ , \new_[47253]_ ,
    \new_[47257]_ , \new_[47258]_ , \new_[47259]_ , \new_[47263]_ ,
    \new_[47264]_ , \new_[47267]_ , \new_[47270]_ , \new_[47271]_ ,
    \new_[47272]_ , \new_[47276]_ , \new_[47277]_ , \new_[47281]_ ,
    \new_[47282]_ , \new_[47283]_ , \new_[47287]_ , \new_[47288]_ ,
    \new_[47291]_ , \new_[47294]_ , \new_[47295]_ , \new_[47296]_ ,
    \new_[47300]_ , \new_[47301]_ , \new_[47305]_ , \new_[47306]_ ,
    \new_[47307]_ , \new_[47311]_ , \new_[47312]_ , \new_[47315]_ ,
    \new_[47318]_ , \new_[47319]_ , \new_[47320]_ , \new_[47324]_ ,
    \new_[47325]_ , \new_[47329]_ , \new_[47330]_ , \new_[47331]_ ,
    \new_[47335]_ , \new_[47336]_ , \new_[47339]_ , \new_[47342]_ ,
    \new_[47343]_ , \new_[47344]_ , \new_[47348]_ , \new_[47349]_ ,
    \new_[47353]_ , \new_[47354]_ , \new_[47355]_ , \new_[47359]_ ,
    \new_[47360]_ , \new_[47363]_ , \new_[47366]_ , \new_[47367]_ ,
    \new_[47368]_ , \new_[47372]_ , \new_[47373]_ , \new_[47377]_ ,
    \new_[47378]_ , \new_[47379]_ , \new_[47383]_ , \new_[47384]_ ,
    \new_[47387]_ , \new_[47390]_ , \new_[47391]_ , \new_[47392]_ ,
    \new_[47396]_ , \new_[47397]_ , \new_[47401]_ , \new_[47402]_ ,
    \new_[47403]_ , \new_[47407]_ , \new_[47408]_ , \new_[47411]_ ,
    \new_[47414]_ , \new_[47415]_ , \new_[47416]_ , \new_[47420]_ ,
    \new_[47421]_ , \new_[47425]_ , \new_[47426]_ , \new_[47427]_ ,
    \new_[47431]_ , \new_[47432]_ , \new_[47435]_ , \new_[47438]_ ,
    \new_[47439]_ , \new_[47440]_ , \new_[47444]_ , \new_[47445]_ ,
    \new_[47449]_ , \new_[47450]_ , \new_[47451]_ , \new_[47455]_ ,
    \new_[47456]_ , \new_[47459]_ , \new_[47462]_ , \new_[47463]_ ,
    \new_[47464]_ , \new_[47468]_ , \new_[47469]_ , \new_[47473]_ ,
    \new_[47474]_ , \new_[47475]_ , \new_[47479]_ , \new_[47480]_ ,
    \new_[47483]_ , \new_[47486]_ , \new_[47487]_ , \new_[47488]_ ,
    \new_[47492]_ , \new_[47493]_ , \new_[47497]_ , \new_[47498]_ ,
    \new_[47499]_ , \new_[47503]_ , \new_[47504]_ , \new_[47507]_ ,
    \new_[47510]_ , \new_[47511]_ , \new_[47512]_ , \new_[47516]_ ,
    \new_[47517]_ , \new_[47521]_ , \new_[47522]_ , \new_[47523]_ ,
    \new_[47527]_ , \new_[47528]_ , \new_[47531]_ , \new_[47534]_ ,
    \new_[47535]_ , \new_[47536]_ , \new_[47540]_ , \new_[47541]_ ,
    \new_[47545]_ , \new_[47546]_ , \new_[47547]_ , \new_[47551]_ ,
    \new_[47552]_ , \new_[47555]_ , \new_[47558]_ , \new_[47559]_ ,
    \new_[47560]_ , \new_[47564]_ , \new_[47565]_ , \new_[47569]_ ,
    \new_[47570]_ , \new_[47571]_ , \new_[47575]_ , \new_[47576]_ ,
    \new_[47579]_ , \new_[47582]_ , \new_[47583]_ , \new_[47584]_ ,
    \new_[47588]_ , \new_[47589]_ , \new_[47593]_ , \new_[47594]_ ,
    \new_[47595]_ , \new_[47599]_ , \new_[47600]_ , \new_[47603]_ ,
    \new_[47606]_ , \new_[47607]_ , \new_[47608]_ , \new_[47612]_ ,
    \new_[47613]_ , \new_[47617]_ , \new_[47618]_ , \new_[47619]_ ,
    \new_[47623]_ , \new_[47624]_ , \new_[47627]_ , \new_[47630]_ ,
    \new_[47631]_ , \new_[47632]_ , \new_[47636]_ , \new_[47637]_ ,
    \new_[47641]_ , \new_[47642]_ , \new_[47643]_ , \new_[47647]_ ,
    \new_[47648]_ , \new_[47651]_ , \new_[47654]_ , \new_[47655]_ ,
    \new_[47656]_ , \new_[47660]_ , \new_[47661]_ , \new_[47665]_ ,
    \new_[47666]_ , \new_[47667]_ , \new_[47671]_ , \new_[47672]_ ,
    \new_[47675]_ , \new_[47678]_ , \new_[47679]_ , \new_[47680]_ ,
    \new_[47684]_ , \new_[47685]_ , \new_[47689]_ , \new_[47690]_ ,
    \new_[47691]_ , \new_[47695]_ , \new_[47696]_ , \new_[47699]_ ,
    \new_[47702]_ , \new_[47703]_ , \new_[47704]_ , \new_[47708]_ ,
    \new_[47709]_ , \new_[47713]_ , \new_[47714]_ , \new_[47715]_ ,
    \new_[47719]_ , \new_[47720]_ , \new_[47723]_ , \new_[47726]_ ,
    \new_[47727]_ , \new_[47728]_ , \new_[47732]_ , \new_[47733]_ ,
    \new_[47737]_ , \new_[47738]_ , \new_[47739]_ , \new_[47743]_ ,
    \new_[47744]_ , \new_[47747]_ , \new_[47750]_ , \new_[47751]_ ,
    \new_[47752]_ , \new_[47756]_ , \new_[47757]_ , \new_[47761]_ ,
    \new_[47762]_ , \new_[47763]_ , \new_[47767]_ , \new_[47768]_ ,
    \new_[47771]_ , \new_[47774]_ , \new_[47775]_ , \new_[47776]_ ,
    \new_[47780]_ , \new_[47781]_ , \new_[47785]_ , \new_[47786]_ ,
    \new_[47787]_ , \new_[47791]_ , \new_[47792]_ , \new_[47795]_ ,
    \new_[47798]_ , \new_[47799]_ , \new_[47800]_ , \new_[47804]_ ,
    \new_[47805]_ , \new_[47809]_ , \new_[47810]_ , \new_[47811]_ ,
    \new_[47815]_ , \new_[47816]_ , \new_[47819]_ , \new_[47822]_ ,
    \new_[47823]_ , \new_[47824]_ , \new_[47828]_ , \new_[47829]_ ,
    \new_[47833]_ , \new_[47834]_ , \new_[47835]_ , \new_[47839]_ ,
    \new_[47840]_ , \new_[47843]_ , \new_[47846]_ , \new_[47847]_ ,
    \new_[47848]_ , \new_[47852]_ , \new_[47853]_ , \new_[47857]_ ,
    \new_[47858]_ , \new_[47859]_ , \new_[47863]_ , \new_[47864]_ ,
    \new_[47867]_ , \new_[47870]_ , \new_[47871]_ , \new_[47872]_ ,
    \new_[47876]_ , \new_[47877]_ , \new_[47881]_ , \new_[47882]_ ,
    \new_[47883]_ , \new_[47887]_ , \new_[47888]_ , \new_[47891]_ ,
    \new_[47894]_ , \new_[47895]_ , \new_[47896]_ , \new_[47900]_ ,
    \new_[47901]_ , \new_[47905]_ , \new_[47906]_ , \new_[47907]_ ,
    \new_[47911]_ , \new_[47912]_ , \new_[47915]_ , \new_[47918]_ ,
    \new_[47919]_ , \new_[47920]_ , \new_[47924]_ , \new_[47925]_ ,
    \new_[47929]_ , \new_[47930]_ , \new_[47931]_ , \new_[47935]_ ,
    \new_[47936]_ , \new_[47939]_ , \new_[47942]_ , \new_[47943]_ ,
    \new_[47944]_ , \new_[47948]_ , \new_[47949]_ , \new_[47953]_ ,
    \new_[47954]_ , \new_[47955]_ , \new_[47959]_ , \new_[47960]_ ,
    \new_[47963]_ , \new_[47966]_ , \new_[47967]_ , \new_[47968]_ ,
    \new_[47972]_ , \new_[47973]_ , \new_[47977]_ , \new_[47978]_ ,
    \new_[47979]_ , \new_[47983]_ , \new_[47984]_ , \new_[47987]_ ,
    \new_[47990]_ , \new_[47991]_ , \new_[47992]_ , \new_[47996]_ ,
    \new_[47997]_ , \new_[48001]_ , \new_[48002]_ , \new_[48003]_ ,
    \new_[48007]_ , \new_[48008]_ , \new_[48011]_ , \new_[48014]_ ,
    \new_[48015]_ , \new_[48016]_ , \new_[48020]_ , \new_[48021]_ ,
    \new_[48025]_ , \new_[48026]_ , \new_[48027]_ , \new_[48031]_ ,
    \new_[48032]_ , \new_[48035]_ , \new_[48038]_ , \new_[48039]_ ,
    \new_[48040]_ , \new_[48044]_ , \new_[48045]_ , \new_[48049]_ ,
    \new_[48050]_ , \new_[48051]_ , \new_[48055]_ , \new_[48056]_ ,
    \new_[48059]_ , \new_[48062]_ , \new_[48063]_ , \new_[48064]_ ,
    \new_[48068]_ , \new_[48069]_ , \new_[48073]_ , \new_[48074]_ ,
    \new_[48075]_ , \new_[48079]_ , \new_[48080]_ , \new_[48083]_ ,
    \new_[48086]_ , \new_[48087]_ , \new_[48088]_ , \new_[48092]_ ,
    \new_[48093]_ , \new_[48097]_ , \new_[48098]_ , \new_[48099]_ ,
    \new_[48103]_ , \new_[48104]_ , \new_[48107]_ , \new_[48110]_ ,
    \new_[48111]_ , \new_[48112]_ , \new_[48116]_ , \new_[48117]_ ,
    \new_[48121]_ , \new_[48122]_ , \new_[48123]_ , \new_[48127]_ ,
    \new_[48128]_ , \new_[48131]_ , \new_[48134]_ , \new_[48135]_ ,
    \new_[48136]_ , \new_[48140]_ , \new_[48141]_ , \new_[48145]_ ,
    \new_[48146]_ , \new_[48147]_ , \new_[48151]_ , \new_[48152]_ ,
    \new_[48155]_ , \new_[48158]_ , \new_[48159]_ , \new_[48160]_ ,
    \new_[48164]_ , \new_[48165]_ , \new_[48169]_ , \new_[48170]_ ,
    \new_[48171]_ , \new_[48175]_ , \new_[48176]_ , \new_[48179]_ ,
    \new_[48182]_ , \new_[48183]_ , \new_[48184]_ , \new_[48188]_ ,
    \new_[48189]_ , \new_[48193]_ , \new_[48194]_ , \new_[48195]_ ,
    \new_[48199]_ , \new_[48200]_ , \new_[48203]_ , \new_[48206]_ ,
    \new_[48207]_ , \new_[48208]_ , \new_[48212]_ , \new_[48213]_ ,
    \new_[48217]_ , \new_[48218]_ , \new_[48219]_ , \new_[48223]_ ,
    \new_[48224]_ , \new_[48227]_ , \new_[48230]_ , \new_[48231]_ ,
    \new_[48232]_ , \new_[48236]_ , \new_[48237]_ , \new_[48241]_ ,
    \new_[48242]_ , \new_[48243]_ , \new_[48247]_ , \new_[48248]_ ,
    \new_[48251]_ , \new_[48254]_ , \new_[48255]_ , \new_[48256]_ ,
    \new_[48260]_ , \new_[48261]_ , \new_[48265]_ , \new_[48266]_ ,
    \new_[48267]_ , \new_[48271]_ , \new_[48272]_ , \new_[48275]_ ,
    \new_[48278]_ , \new_[48279]_ , \new_[48280]_ , \new_[48284]_ ,
    \new_[48285]_ , \new_[48289]_ , \new_[48290]_ , \new_[48291]_ ,
    \new_[48295]_ , \new_[48296]_ , \new_[48299]_ , \new_[48302]_ ,
    \new_[48303]_ , \new_[48304]_ , \new_[48308]_ , \new_[48309]_ ,
    \new_[48313]_ , \new_[48314]_ , \new_[48315]_ , \new_[48319]_ ,
    \new_[48320]_ , \new_[48323]_ , \new_[48326]_ , \new_[48327]_ ,
    \new_[48328]_ , \new_[48332]_ , \new_[48333]_ , \new_[48337]_ ,
    \new_[48338]_ , \new_[48339]_ , \new_[48343]_ , \new_[48344]_ ,
    \new_[48347]_ , \new_[48350]_ , \new_[48351]_ , \new_[48352]_ ,
    \new_[48356]_ , \new_[48357]_ , \new_[48361]_ , \new_[48362]_ ,
    \new_[48363]_ , \new_[48367]_ , \new_[48368]_ , \new_[48371]_ ,
    \new_[48374]_ , \new_[48375]_ , \new_[48376]_ , \new_[48380]_ ,
    \new_[48381]_ , \new_[48385]_ , \new_[48386]_ , \new_[48387]_ ,
    \new_[48391]_ , \new_[48392]_ , \new_[48395]_ , \new_[48398]_ ,
    \new_[48399]_ , \new_[48400]_ , \new_[48404]_ , \new_[48405]_ ,
    \new_[48409]_ , \new_[48410]_ , \new_[48411]_ , \new_[48415]_ ,
    \new_[48416]_ , \new_[48419]_ , \new_[48422]_ , \new_[48423]_ ,
    \new_[48424]_ , \new_[48428]_ , \new_[48429]_ , \new_[48433]_ ,
    \new_[48434]_ , \new_[48435]_ , \new_[48439]_ , \new_[48440]_ ,
    \new_[48443]_ , \new_[48446]_ , \new_[48447]_ , \new_[48448]_ ,
    \new_[48452]_ , \new_[48453]_ , \new_[48457]_ , \new_[48458]_ ,
    \new_[48459]_ , \new_[48463]_ , \new_[48464]_ , \new_[48467]_ ,
    \new_[48470]_ , \new_[48471]_ , \new_[48472]_ , \new_[48476]_ ,
    \new_[48477]_ , \new_[48481]_ , \new_[48482]_ , \new_[48483]_ ,
    \new_[48487]_ , \new_[48488]_ , \new_[48491]_ , \new_[48494]_ ,
    \new_[48495]_ , \new_[48496]_ , \new_[48500]_ , \new_[48501]_ ,
    \new_[48505]_ , \new_[48506]_ , \new_[48507]_ , \new_[48511]_ ,
    \new_[48512]_ , \new_[48515]_ , \new_[48518]_ , \new_[48519]_ ,
    \new_[48520]_ , \new_[48524]_ , \new_[48525]_ , \new_[48529]_ ,
    \new_[48530]_ , \new_[48531]_ , \new_[48535]_ , \new_[48536]_ ,
    \new_[48539]_ , \new_[48542]_ , \new_[48543]_ , \new_[48544]_ ,
    \new_[48548]_ , \new_[48549]_ , \new_[48553]_ , \new_[48554]_ ,
    \new_[48555]_ , \new_[48559]_ , \new_[48560]_ , \new_[48563]_ ,
    \new_[48566]_ , \new_[48567]_ , \new_[48568]_ , \new_[48572]_ ,
    \new_[48573]_ , \new_[48577]_ , \new_[48578]_ , \new_[48579]_ ,
    \new_[48583]_ , \new_[48584]_ , \new_[48587]_ , \new_[48590]_ ,
    \new_[48591]_ , \new_[48592]_ , \new_[48596]_ , \new_[48597]_ ,
    \new_[48601]_ , \new_[48602]_ , \new_[48603]_ , \new_[48607]_ ,
    \new_[48608]_ , \new_[48611]_ , \new_[48614]_ , \new_[48615]_ ,
    \new_[48616]_ , \new_[48620]_ , \new_[48621]_ , \new_[48625]_ ,
    \new_[48626]_ , \new_[48627]_ , \new_[48631]_ , \new_[48632]_ ,
    \new_[48635]_ , \new_[48638]_ , \new_[48639]_ , \new_[48640]_ ,
    \new_[48644]_ , \new_[48645]_ , \new_[48649]_ , \new_[48650]_ ,
    \new_[48651]_ , \new_[48655]_ , \new_[48656]_ , \new_[48659]_ ,
    \new_[48662]_ , \new_[48663]_ , \new_[48664]_ , \new_[48668]_ ,
    \new_[48669]_ , \new_[48673]_ , \new_[48674]_ , \new_[48675]_ ,
    \new_[48679]_ , \new_[48680]_ , \new_[48683]_ , \new_[48686]_ ,
    \new_[48687]_ , \new_[48688]_ , \new_[48692]_ , \new_[48693]_ ,
    \new_[48697]_ , \new_[48698]_ , \new_[48699]_ , \new_[48703]_ ,
    \new_[48704]_ , \new_[48707]_ , \new_[48710]_ , \new_[48711]_ ,
    \new_[48712]_ , \new_[48716]_ , \new_[48717]_ , \new_[48721]_ ,
    \new_[48722]_ , \new_[48723]_ , \new_[48727]_ , \new_[48728]_ ,
    \new_[48731]_ , \new_[48734]_ , \new_[48735]_ , \new_[48736]_ ,
    \new_[48740]_ , \new_[48741]_ , \new_[48745]_ , \new_[48746]_ ,
    \new_[48747]_ , \new_[48751]_ , \new_[48752]_ , \new_[48755]_ ,
    \new_[48758]_ , \new_[48759]_ , \new_[48760]_ , \new_[48764]_ ,
    \new_[48765]_ , \new_[48769]_ , \new_[48770]_ , \new_[48771]_ ,
    \new_[48775]_ , \new_[48776]_ , \new_[48779]_ , \new_[48782]_ ,
    \new_[48783]_ , \new_[48784]_ , \new_[48788]_ , \new_[48789]_ ,
    \new_[48793]_ , \new_[48794]_ , \new_[48795]_ , \new_[48799]_ ,
    \new_[48800]_ , \new_[48803]_ , \new_[48806]_ , \new_[48807]_ ,
    \new_[48808]_ , \new_[48812]_ , \new_[48813]_ , \new_[48817]_ ,
    \new_[48818]_ , \new_[48819]_ , \new_[48823]_ , \new_[48824]_ ,
    \new_[48827]_ , \new_[48830]_ , \new_[48831]_ , \new_[48832]_ ,
    \new_[48836]_ , \new_[48837]_ , \new_[48841]_ , \new_[48842]_ ,
    \new_[48843]_ , \new_[48847]_ , \new_[48848]_ , \new_[48851]_ ,
    \new_[48854]_ , \new_[48855]_ , \new_[48856]_ , \new_[48860]_ ,
    \new_[48861]_ , \new_[48865]_ , \new_[48866]_ , \new_[48867]_ ,
    \new_[48871]_ , \new_[48872]_ , \new_[48875]_ , \new_[48878]_ ,
    \new_[48879]_ , \new_[48880]_ , \new_[48884]_ , \new_[48885]_ ,
    \new_[48889]_ , \new_[48890]_ , \new_[48891]_ , \new_[48895]_ ,
    \new_[48896]_ , \new_[48899]_ , \new_[48902]_ , \new_[48903]_ ,
    \new_[48904]_ , \new_[48908]_ , \new_[48909]_ , \new_[48913]_ ,
    \new_[48914]_ , \new_[48915]_ , \new_[48919]_ , \new_[48920]_ ,
    \new_[48923]_ , \new_[48926]_ , \new_[48927]_ , \new_[48928]_ ,
    \new_[48932]_ , \new_[48933]_ , \new_[48937]_ , \new_[48938]_ ,
    \new_[48939]_ , \new_[48943]_ , \new_[48944]_ , \new_[48947]_ ,
    \new_[48950]_ , \new_[48951]_ , \new_[48952]_ , \new_[48956]_ ,
    \new_[48957]_ , \new_[48961]_ , \new_[48962]_ , \new_[48963]_ ,
    \new_[48967]_ , \new_[48968]_ , \new_[48971]_ , \new_[48974]_ ,
    \new_[48975]_ , \new_[48976]_ , \new_[48980]_ , \new_[48981]_ ,
    \new_[48985]_ , \new_[48986]_ , \new_[48987]_ , \new_[48991]_ ,
    \new_[48992]_ , \new_[48995]_ , \new_[48998]_ , \new_[48999]_ ,
    \new_[49000]_ , \new_[49004]_ , \new_[49005]_ , \new_[49009]_ ,
    \new_[49010]_ , \new_[49011]_ , \new_[49015]_ , \new_[49016]_ ,
    \new_[49019]_ , \new_[49022]_ , \new_[49023]_ , \new_[49024]_ ,
    \new_[49028]_ , \new_[49029]_ , \new_[49033]_ , \new_[49034]_ ,
    \new_[49035]_ , \new_[49039]_ , \new_[49040]_ , \new_[49043]_ ,
    \new_[49046]_ , \new_[49047]_ , \new_[49048]_ , \new_[49052]_ ,
    \new_[49053]_ , \new_[49057]_ , \new_[49058]_ , \new_[49059]_ ,
    \new_[49063]_ , \new_[49064]_ , \new_[49067]_ , \new_[49070]_ ,
    \new_[49071]_ , \new_[49072]_ , \new_[49076]_ , \new_[49077]_ ,
    \new_[49081]_ , \new_[49082]_ , \new_[49083]_ , \new_[49087]_ ,
    \new_[49088]_ , \new_[49091]_ , \new_[49094]_ , \new_[49095]_ ,
    \new_[49096]_ , \new_[49100]_ , \new_[49101]_ , \new_[49105]_ ,
    \new_[49106]_ , \new_[49107]_ , \new_[49111]_ , \new_[49112]_ ,
    \new_[49115]_ , \new_[49118]_ , \new_[49119]_ , \new_[49120]_ ,
    \new_[49124]_ , \new_[49125]_ , \new_[49129]_ , \new_[49130]_ ,
    \new_[49131]_ , \new_[49135]_ , \new_[49136]_ , \new_[49139]_ ,
    \new_[49142]_ , \new_[49143]_ , \new_[49144]_ , \new_[49148]_ ,
    \new_[49149]_ , \new_[49153]_ , \new_[49154]_ , \new_[49155]_ ,
    \new_[49159]_ , \new_[49160]_ , \new_[49163]_ , \new_[49166]_ ,
    \new_[49167]_ , \new_[49168]_ , \new_[49172]_ , \new_[49173]_ ,
    \new_[49177]_ , \new_[49178]_ , \new_[49179]_ , \new_[49183]_ ,
    \new_[49184]_ , \new_[49187]_ , \new_[49190]_ , \new_[49191]_ ,
    \new_[49192]_ , \new_[49196]_ , \new_[49197]_ , \new_[49201]_ ,
    \new_[49202]_ , \new_[49203]_ , \new_[49207]_ , \new_[49208]_ ,
    \new_[49211]_ , \new_[49214]_ , \new_[49215]_ , \new_[49216]_ ,
    \new_[49220]_ , \new_[49221]_ , \new_[49225]_ , \new_[49226]_ ,
    \new_[49227]_ , \new_[49231]_ , \new_[49232]_ , \new_[49235]_ ,
    \new_[49238]_ , \new_[49239]_ , \new_[49240]_ , \new_[49244]_ ,
    \new_[49245]_ , \new_[49249]_ , \new_[49250]_ , \new_[49251]_ ,
    \new_[49255]_ , \new_[49256]_ , \new_[49259]_ , \new_[49262]_ ,
    \new_[49263]_ , \new_[49264]_ , \new_[49268]_ , \new_[49269]_ ,
    \new_[49273]_ , \new_[49274]_ , \new_[49275]_ , \new_[49279]_ ,
    \new_[49280]_ , \new_[49283]_ , \new_[49286]_ , \new_[49287]_ ,
    \new_[49288]_ , \new_[49292]_ , \new_[49293]_ , \new_[49297]_ ,
    \new_[49298]_ , \new_[49299]_ , \new_[49303]_ , \new_[49304]_ ,
    \new_[49307]_ , \new_[49310]_ , \new_[49311]_ , \new_[49312]_ ,
    \new_[49316]_ , \new_[49317]_ , \new_[49321]_ , \new_[49322]_ ,
    \new_[49323]_ , \new_[49327]_ , \new_[49328]_ , \new_[49331]_ ,
    \new_[49334]_ , \new_[49335]_ , \new_[49336]_ , \new_[49340]_ ,
    \new_[49341]_ , \new_[49345]_ , \new_[49346]_ , \new_[49347]_ ,
    \new_[49351]_ , \new_[49352]_ , \new_[49355]_ , \new_[49358]_ ,
    \new_[49359]_ , \new_[49360]_ , \new_[49364]_ , \new_[49365]_ ,
    \new_[49369]_ , \new_[49370]_ , \new_[49371]_ , \new_[49375]_ ,
    \new_[49376]_ , \new_[49379]_ , \new_[49382]_ , \new_[49383]_ ,
    \new_[49384]_ , \new_[49388]_ , \new_[49389]_ , \new_[49393]_ ,
    \new_[49394]_ , \new_[49395]_ , \new_[49399]_ , \new_[49400]_ ,
    \new_[49403]_ , \new_[49406]_ , \new_[49407]_ , \new_[49408]_ ,
    \new_[49412]_ , \new_[49413]_ , \new_[49417]_ , \new_[49418]_ ,
    \new_[49419]_ , \new_[49423]_ , \new_[49424]_ , \new_[49427]_ ,
    \new_[49430]_ , \new_[49431]_ , \new_[49432]_ , \new_[49436]_ ,
    \new_[49437]_ , \new_[49441]_ , \new_[49442]_ , \new_[49443]_ ,
    \new_[49447]_ , \new_[49448]_ , \new_[49451]_ , \new_[49454]_ ,
    \new_[49455]_ , \new_[49456]_ , \new_[49460]_ , \new_[49461]_ ,
    \new_[49465]_ , \new_[49466]_ , \new_[49467]_ , \new_[49471]_ ,
    \new_[49472]_ , \new_[49475]_ , \new_[49478]_ , \new_[49479]_ ,
    \new_[49480]_ , \new_[49484]_ , \new_[49485]_ , \new_[49489]_ ,
    \new_[49490]_ , \new_[49491]_ , \new_[49495]_ , \new_[49496]_ ,
    \new_[49499]_ , \new_[49502]_ , \new_[49503]_ , \new_[49504]_ ,
    \new_[49508]_ , \new_[49509]_ , \new_[49513]_ , \new_[49514]_ ,
    \new_[49515]_ , \new_[49519]_ , \new_[49520]_ , \new_[49523]_ ,
    \new_[49526]_ , \new_[49527]_ , \new_[49528]_ , \new_[49532]_ ,
    \new_[49533]_ , \new_[49537]_ , \new_[49538]_ , \new_[49539]_ ,
    \new_[49543]_ , \new_[49544]_ , \new_[49547]_ , \new_[49550]_ ,
    \new_[49551]_ , \new_[49552]_ , \new_[49556]_ , \new_[49557]_ ,
    \new_[49561]_ , \new_[49562]_ , \new_[49563]_ , \new_[49567]_ ,
    \new_[49568]_ , \new_[49571]_ , \new_[49574]_ , \new_[49575]_ ,
    \new_[49576]_ , \new_[49580]_ , \new_[49581]_ , \new_[49585]_ ,
    \new_[49586]_ , \new_[49587]_ , \new_[49591]_ , \new_[49592]_ ,
    \new_[49595]_ , \new_[49598]_ , \new_[49599]_ , \new_[49600]_ ,
    \new_[49604]_ , \new_[49605]_ , \new_[49609]_ , \new_[49610]_ ,
    \new_[49611]_ , \new_[49615]_ , \new_[49616]_ , \new_[49619]_ ,
    \new_[49622]_ , \new_[49623]_ , \new_[49624]_ , \new_[49628]_ ,
    \new_[49629]_ , \new_[49633]_ , \new_[49634]_ , \new_[49635]_ ,
    \new_[49639]_ , \new_[49640]_ , \new_[49643]_ , \new_[49646]_ ,
    \new_[49647]_ , \new_[49648]_ , \new_[49652]_ , \new_[49653]_ ,
    \new_[49657]_ , \new_[49658]_ , \new_[49659]_ , \new_[49663]_ ,
    \new_[49664]_ , \new_[49667]_ , \new_[49670]_ , \new_[49671]_ ,
    \new_[49672]_ , \new_[49676]_ , \new_[49677]_ , \new_[49681]_ ,
    \new_[49682]_ , \new_[49683]_ , \new_[49687]_ , \new_[49688]_ ,
    \new_[49691]_ , \new_[49694]_ , \new_[49695]_ , \new_[49696]_ ,
    \new_[49700]_ , \new_[49701]_ , \new_[49705]_ , \new_[49706]_ ,
    \new_[49707]_ , \new_[49711]_ , \new_[49712]_ , \new_[49715]_ ,
    \new_[49718]_ , \new_[49719]_ , \new_[49720]_ , \new_[49724]_ ,
    \new_[49725]_ , \new_[49729]_ , \new_[49730]_ , \new_[49731]_ ,
    \new_[49735]_ , \new_[49736]_ , \new_[49739]_ , \new_[49742]_ ,
    \new_[49743]_ , \new_[49744]_ , \new_[49748]_ , \new_[49749]_ ,
    \new_[49753]_ , \new_[49754]_ , \new_[49755]_ , \new_[49759]_ ,
    \new_[49760]_ , \new_[49763]_ , \new_[49766]_ , \new_[49767]_ ,
    \new_[49768]_ , \new_[49772]_ , \new_[49773]_ , \new_[49777]_ ,
    \new_[49778]_ , \new_[49779]_ , \new_[49783]_ , \new_[49784]_ ,
    \new_[49787]_ , \new_[49790]_ , \new_[49791]_ , \new_[49792]_ ,
    \new_[49796]_ , \new_[49797]_ , \new_[49801]_ , \new_[49802]_ ,
    \new_[49803]_ , \new_[49807]_ , \new_[49808]_ , \new_[49811]_ ,
    \new_[49814]_ , \new_[49815]_ , \new_[49816]_ , \new_[49820]_ ,
    \new_[49821]_ , \new_[49825]_ , \new_[49826]_ , \new_[49827]_ ,
    \new_[49831]_ , \new_[49832]_ , \new_[49835]_ , \new_[49838]_ ,
    \new_[49839]_ , \new_[49840]_ , \new_[49844]_ , \new_[49845]_ ,
    \new_[49849]_ , \new_[49850]_ , \new_[49851]_ , \new_[49855]_ ,
    \new_[49856]_ , \new_[49859]_ , \new_[49862]_ , \new_[49863]_ ,
    \new_[49864]_ , \new_[49868]_ , \new_[49869]_ , \new_[49873]_ ,
    \new_[49874]_ , \new_[49875]_ , \new_[49879]_ , \new_[49880]_ ,
    \new_[49883]_ , \new_[49886]_ , \new_[49887]_ , \new_[49888]_ ,
    \new_[49892]_ , \new_[49893]_ , \new_[49897]_ , \new_[49898]_ ,
    \new_[49899]_ , \new_[49903]_ , \new_[49904]_ , \new_[49907]_ ,
    \new_[49910]_ , \new_[49911]_ , \new_[49912]_ , \new_[49916]_ ,
    \new_[49917]_ , \new_[49921]_ , \new_[49922]_ , \new_[49923]_ ,
    \new_[49927]_ , \new_[49928]_ , \new_[49931]_ , \new_[49934]_ ,
    \new_[49935]_ , \new_[49936]_ , \new_[49940]_ , \new_[49941]_ ,
    \new_[49945]_ , \new_[49946]_ , \new_[49947]_ , \new_[49951]_ ,
    \new_[49952]_ , \new_[49955]_ , \new_[49958]_ , \new_[49959]_ ,
    \new_[49960]_ , \new_[49964]_ , \new_[49965]_ , \new_[49969]_ ,
    \new_[49970]_ , \new_[49971]_ , \new_[49975]_ , \new_[49976]_ ,
    \new_[49979]_ , \new_[49982]_ , \new_[49983]_ , \new_[49984]_ ,
    \new_[49988]_ , \new_[49989]_ , \new_[49993]_ , \new_[49994]_ ,
    \new_[49995]_ , \new_[49999]_ , \new_[50000]_ , \new_[50003]_ ,
    \new_[50006]_ , \new_[50007]_ , \new_[50008]_ , \new_[50012]_ ,
    \new_[50013]_ , \new_[50017]_ , \new_[50018]_ , \new_[50019]_ ,
    \new_[50023]_ , \new_[50024]_ , \new_[50027]_ , \new_[50030]_ ,
    \new_[50031]_ , \new_[50032]_ , \new_[50036]_ , \new_[50037]_ ,
    \new_[50041]_ , \new_[50042]_ , \new_[50043]_ , \new_[50047]_ ,
    \new_[50048]_ , \new_[50051]_ , \new_[50054]_ , \new_[50055]_ ,
    \new_[50056]_ , \new_[50060]_ , \new_[50061]_ , \new_[50065]_ ,
    \new_[50066]_ , \new_[50067]_ , \new_[50071]_ , \new_[50072]_ ,
    \new_[50075]_ , \new_[50078]_ , \new_[50079]_ , \new_[50080]_ ,
    \new_[50084]_ , \new_[50085]_ , \new_[50089]_ , \new_[50090]_ ,
    \new_[50091]_ , \new_[50095]_ , \new_[50096]_ , \new_[50099]_ ,
    \new_[50102]_ , \new_[50103]_ , \new_[50104]_ , \new_[50108]_ ,
    \new_[50109]_ , \new_[50113]_ , \new_[50114]_ , \new_[50115]_ ,
    \new_[50119]_ , \new_[50120]_ , \new_[50123]_ , \new_[50126]_ ,
    \new_[50127]_ , \new_[50128]_ , \new_[50132]_ , \new_[50133]_ ,
    \new_[50137]_ , \new_[50138]_ , \new_[50139]_ , \new_[50143]_ ,
    \new_[50144]_ , \new_[50147]_ , \new_[50150]_ , \new_[50151]_ ,
    \new_[50152]_ , \new_[50156]_ , \new_[50157]_ , \new_[50161]_ ,
    \new_[50162]_ , \new_[50163]_ , \new_[50167]_ , \new_[50168]_ ,
    \new_[50171]_ , \new_[50174]_ , \new_[50175]_ , \new_[50176]_ ,
    \new_[50180]_ , \new_[50181]_ , \new_[50185]_ , \new_[50186]_ ,
    \new_[50187]_ , \new_[50191]_ , \new_[50192]_ , \new_[50195]_ ,
    \new_[50198]_ , \new_[50199]_ , \new_[50200]_ , \new_[50204]_ ,
    \new_[50205]_ , \new_[50209]_ , \new_[50210]_ , \new_[50211]_ ,
    \new_[50215]_ , \new_[50216]_ , \new_[50219]_ , \new_[50222]_ ,
    \new_[50223]_ , \new_[50224]_ , \new_[50228]_ , \new_[50229]_ ,
    \new_[50233]_ , \new_[50234]_ , \new_[50235]_ , \new_[50239]_ ,
    \new_[50240]_ , \new_[50243]_ , \new_[50246]_ , \new_[50247]_ ,
    \new_[50248]_ , \new_[50252]_ , \new_[50253]_ , \new_[50257]_ ,
    \new_[50258]_ , \new_[50259]_ , \new_[50263]_ , \new_[50264]_ ,
    \new_[50267]_ , \new_[50270]_ , \new_[50271]_ , \new_[50272]_ ,
    \new_[50276]_ , \new_[50277]_ , \new_[50281]_ , \new_[50282]_ ,
    \new_[50283]_ , \new_[50287]_ , \new_[50288]_ , \new_[50291]_ ,
    \new_[50294]_ , \new_[50295]_ , \new_[50296]_ , \new_[50300]_ ,
    \new_[50301]_ , \new_[50305]_ , \new_[50306]_ , \new_[50307]_ ,
    \new_[50311]_ , \new_[50312]_ , \new_[50315]_ , \new_[50318]_ ,
    \new_[50319]_ , \new_[50320]_ , \new_[50324]_ , \new_[50325]_ ,
    \new_[50329]_ , \new_[50330]_ , \new_[50331]_ , \new_[50335]_ ,
    \new_[50336]_ , \new_[50339]_ , \new_[50342]_ , \new_[50343]_ ,
    \new_[50344]_ , \new_[50348]_ , \new_[50349]_ , \new_[50353]_ ,
    \new_[50354]_ , \new_[50355]_ , \new_[50359]_ , \new_[50360]_ ,
    \new_[50363]_ , \new_[50366]_ , \new_[50367]_ , \new_[50368]_ ,
    \new_[50372]_ , \new_[50373]_ , \new_[50377]_ , \new_[50378]_ ,
    \new_[50379]_ , \new_[50383]_ , \new_[50384]_ , \new_[50387]_ ,
    \new_[50390]_ , \new_[50391]_ , \new_[50392]_ , \new_[50396]_ ,
    \new_[50397]_ , \new_[50401]_ , \new_[50402]_ , \new_[50403]_ ,
    \new_[50407]_ , \new_[50408]_ , \new_[50411]_ , \new_[50414]_ ,
    \new_[50415]_ , \new_[50416]_ , \new_[50420]_ , \new_[50421]_ ,
    \new_[50425]_ , \new_[50426]_ , \new_[50427]_ , \new_[50431]_ ,
    \new_[50432]_ , \new_[50435]_ , \new_[50438]_ , \new_[50439]_ ,
    \new_[50440]_ , \new_[50444]_ , \new_[50445]_ , \new_[50449]_ ,
    \new_[50450]_ , \new_[50451]_ , \new_[50455]_ , \new_[50456]_ ,
    \new_[50459]_ , \new_[50462]_ , \new_[50463]_ , \new_[50464]_ ,
    \new_[50468]_ , \new_[50469]_ , \new_[50473]_ , \new_[50474]_ ,
    \new_[50475]_ , \new_[50479]_ , \new_[50480]_ , \new_[50483]_ ,
    \new_[50486]_ , \new_[50487]_ , \new_[50488]_ , \new_[50492]_ ,
    \new_[50493]_ , \new_[50497]_ , \new_[50498]_ , \new_[50499]_ ,
    \new_[50503]_ , \new_[50504]_ , \new_[50507]_ , \new_[50510]_ ,
    \new_[50511]_ , \new_[50512]_ , \new_[50516]_ , \new_[50517]_ ,
    \new_[50521]_ , \new_[50522]_ , \new_[50523]_ , \new_[50527]_ ,
    \new_[50528]_ , \new_[50531]_ , \new_[50534]_ , \new_[50535]_ ,
    \new_[50536]_ , \new_[50540]_ , \new_[50541]_ , \new_[50545]_ ,
    \new_[50546]_ , \new_[50547]_ , \new_[50551]_ , \new_[50552]_ ,
    \new_[50555]_ , \new_[50558]_ , \new_[50559]_ , \new_[50560]_ ,
    \new_[50564]_ , \new_[50565]_ , \new_[50569]_ , \new_[50570]_ ,
    \new_[50571]_ , \new_[50575]_ , \new_[50576]_ , \new_[50579]_ ,
    \new_[50582]_ , \new_[50583]_ , \new_[50584]_ , \new_[50588]_ ,
    \new_[50589]_ , \new_[50593]_ , \new_[50594]_ , \new_[50595]_ ,
    \new_[50599]_ , \new_[50600]_ , \new_[50603]_ , \new_[50606]_ ,
    \new_[50607]_ , \new_[50608]_ , \new_[50612]_ , \new_[50613]_ ,
    \new_[50617]_ , \new_[50618]_ , \new_[50619]_ , \new_[50623]_ ,
    \new_[50624]_ , \new_[50627]_ , \new_[50630]_ , \new_[50631]_ ,
    \new_[50632]_ , \new_[50636]_ , \new_[50637]_ , \new_[50641]_ ,
    \new_[50642]_ , \new_[50643]_ , \new_[50647]_ , \new_[50648]_ ,
    \new_[50651]_ , \new_[50654]_ , \new_[50655]_ , \new_[50656]_ ,
    \new_[50660]_ , \new_[50661]_ , \new_[50665]_ , \new_[50666]_ ,
    \new_[50667]_ , \new_[50671]_ , \new_[50672]_ , \new_[50675]_ ,
    \new_[50678]_ , \new_[50679]_ , \new_[50680]_ , \new_[50684]_ ,
    \new_[50685]_ , \new_[50689]_ , \new_[50690]_ , \new_[50691]_ ,
    \new_[50695]_ , \new_[50696]_ , \new_[50699]_ , \new_[50702]_ ,
    \new_[50703]_ , \new_[50704]_ , \new_[50708]_ , \new_[50709]_ ,
    \new_[50713]_ , \new_[50714]_ , \new_[50715]_ , \new_[50719]_ ,
    \new_[50720]_ , \new_[50723]_ , \new_[50726]_ , \new_[50727]_ ,
    \new_[50728]_ , \new_[50732]_ , \new_[50733]_ , \new_[50737]_ ,
    \new_[50738]_ , \new_[50739]_ , \new_[50743]_ , \new_[50744]_ ,
    \new_[50747]_ , \new_[50750]_ , \new_[50751]_ , \new_[50752]_ ,
    \new_[50756]_ , \new_[50757]_ , \new_[50761]_ , \new_[50762]_ ,
    \new_[50763]_ , \new_[50767]_ , \new_[50768]_ , \new_[50771]_ ,
    \new_[50774]_ , \new_[50775]_ , \new_[50776]_ , \new_[50780]_ ,
    \new_[50781]_ , \new_[50785]_ , \new_[50786]_ , \new_[50787]_ ,
    \new_[50791]_ , \new_[50792]_ , \new_[50795]_ , \new_[50798]_ ,
    \new_[50799]_ , \new_[50800]_ , \new_[50804]_ , \new_[50805]_ ,
    \new_[50809]_ , \new_[50810]_ , \new_[50811]_ , \new_[50815]_ ,
    \new_[50816]_ , \new_[50819]_ , \new_[50822]_ , \new_[50823]_ ,
    \new_[50824]_ , \new_[50828]_ , \new_[50829]_ , \new_[50833]_ ,
    \new_[50834]_ , \new_[50835]_ , \new_[50839]_ , \new_[50840]_ ,
    \new_[50843]_ , \new_[50846]_ , \new_[50847]_ , \new_[50848]_ ,
    \new_[50852]_ , \new_[50853]_ , \new_[50857]_ , \new_[50858]_ ,
    \new_[50859]_ , \new_[50863]_ , \new_[50864]_ , \new_[50867]_ ,
    \new_[50870]_ , \new_[50871]_ , \new_[50872]_ , \new_[50876]_ ,
    \new_[50877]_ , \new_[50881]_ , \new_[50882]_ , \new_[50883]_ ,
    \new_[50887]_ , \new_[50888]_ , \new_[50891]_ , \new_[50894]_ ,
    \new_[50895]_ , \new_[50896]_ , \new_[50900]_ , \new_[50901]_ ,
    \new_[50905]_ , \new_[50906]_ , \new_[50907]_ , \new_[50911]_ ,
    \new_[50912]_ , \new_[50915]_ , \new_[50918]_ , \new_[50919]_ ,
    \new_[50920]_ , \new_[50924]_ , \new_[50925]_ , \new_[50929]_ ,
    \new_[50930]_ , \new_[50931]_ , \new_[50935]_ , \new_[50936]_ ,
    \new_[50939]_ , \new_[50942]_ , \new_[50943]_ , \new_[50944]_ ,
    \new_[50948]_ , \new_[50949]_ , \new_[50953]_ , \new_[50954]_ ,
    \new_[50955]_ , \new_[50959]_ , \new_[50960]_ , \new_[50963]_ ,
    \new_[50966]_ , \new_[50967]_ , \new_[50968]_ , \new_[50972]_ ,
    \new_[50973]_ , \new_[50977]_ , \new_[50978]_ , \new_[50979]_ ,
    \new_[50983]_ , \new_[50984]_ , \new_[50987]_ , \new_[50990]_ ,
    \new_[50991]_ , \new_[50992]_ , \new_[50996]_ , \new_[50997]_ ,
    \new_[51001]_ , \new_[51002]_ , \new_[51003]_ , \new_[51007]_ ,
    \new_[51008]_ , \new_[51011]_ , \new_[51014]_ , \new_[51015]_ ,
    \new_[51016]_ , \new_[51020]_ , \new_[51021]_ , \new_[51025]_ ,
    \new_[51026]_ , \new_[51027]_ , \new_[51031]_ , \new_[51032]_ ,
    \new_[51035]_ , \new_[51038]_ , \new_[51039]_ , \new_[51040]_ ,
    \new_[51044]_ , \new_[51045]_ , \new_[51049]_ , \new_[51050]_ ,
    \new_[51051]_ , \new_[51055]_ , \new_[51056]_ , \new_[51059]_ ,
    \new_[51062]_ , \new_[51063]_ , \new_[51064]_ , \new_[51068]_ ,
    \new_[51069]_ , \new_[51073]_ , \new_[51074]_ , \new_[51075]_ ,
    \new_[51079]_ , \new_[51080]_ , \new_[51083]_ , \new_[51086]_ ,
    \new_[51087]_ , \new_[51088]_ , \new_[51092]_ , \new_[51093]_ ,
    \new_[51097]_ , \new_[51098]_ , \new_[51099]_ , \new_[51103]_ ,
    \new_[51104]_ , \new_[51107]_ , \new_[51110]_ , \new_[51111]_ ,
    \new_[51112]_ , \new_[51116]_ , \new_[51117]_ , \new_[51121]_ ,
    \new_[51122]_ , \new_[51123]_ , \new_[51127]_ , \new_[51128]_ ,
    \new_[51131]_ , \new_[51134]_ , \new_[51135]_ , \new_[51136]_ ,
    \new_[51140]_ , \new_[51141]_ , \new_[51145]_ , \new_[51146]_ ,
    \new_[51147]_ , \new_[51151]_ , \new_[51152]_ , \new_[51155]_ ,
    \new_[51158]_ , \new_[51159]_ , \new_[51160]_ , \new_[51164]_ ,
    \new_[51165]_ , \new_[51169]_ , \new_[51170]_ , \new_[51171]_ ,
    \new_[51175]_ , \new_[51176]_ , \new_[51179]_ , \new_[51182]_ ,
    \new_[51183]_ , \new_[51184]_ , \new_[51188]_ , \new_[51189]_ ,
    \new_[51193]_ , \new_[51194]_ , \new_[51195]_ , \new_[51199]_ ,
    \new_[51200]_ , \new_[51203]_ , \new_[51206]_ , \new_[51207]_ ,
    \new_[51208]_ , \new_[51212]_ , \new_[51213]_ , \new_[51217]_ ,
    \new_[51218]_ , \new_[51219]_ , \new_[51223]_ , \new_[51224]_ ,
    \new_[51227]_ , \new_[51230]_ , \new_[51231]_ , \new_[51232]_ ,
    \new_[51236]_ , \new_[51237]_ , \new_[51241]_ , \new_[51242]_ ,
    \new_[51243]_ , \new_[51247]_ , \new_[51248]_ , \new_[51251]_ ,
    \new_[51254]_ , \new_[51255]_ , \new_[51256]_ , \new_[51260]_ ,
    \new_[51261]_ , \new_[51265]_ , \new_[51266]_ , \new_[51267]_ ,
    \new_[51271]_ , \new_[51272]_ , \new_[51275]_ , \new_[51278]_ ,
    \new_[51279]_ , \new_[51280]_ , \new_[51284]_ , \new_[51285]_ ,
    \new_[51289]_ , \new_[51290]_ , \new_[51291]_ , \new_[51295]_ ,
    \new_[51296]_ , \new_[51299]_ , \new_[51302]_ , \new_[51303]_ ,
    \new_[51304]_ , \new_[51308]_ , \new_[51309]_ , \new_[51313]_ ,
    \new_[51314]_ , \new_[51315]_ , \new_[51319]_ , \new_[51320]_ ,
    \new_[51323]_ , \new_[51326]_ , \new_[51327]_ , \new_[51328]_ ,
    \new_[51332]_ , \new_[51333]_ , \new_[51337]_ , \new_[51338]_ ,
    \new_[51339]_ , \new_[51343]_ , \new_[51344]_ , \new_[51347]_ ,
    \new_[51350]_ , \new_[51351]_ , \new_[51352]_ , \new_[51356]_ ,
    \new_[51357]_ , \new_[51361]_ , \new_[51362]_ , \new_[51363]_ ,
    \new_[51367]_ , \new_[51368]_ , \new_[51371]_ , \new_[51374]_ ,
    \new_[51375]_ , \new_[51376]_ , \new_[51380]_ , \new_[51381]_ ,
    \new_[51385]_ , \new_[51386]_ , \new_[51387]_ , \new_[51391]_ ,
    \new_[51392]_ , \new_[51395]_ , \new_[51398]_ , \new_[51399]_ ,
    \new_[51400]_ , \new_[51404]_ , \new_[51405]_ , \new_[51409]_ ,
    \new_[51410]_ , \new_[51411]_ , \new_[51415]_ , \new_[51416]_ ,
    \new_[51419]_ , \new_[51422]_ , \new_[51423]_ , \new_[51424]_ ,
    \new_[51428]_ , \new_[51429]_ , \new_[51433]_ , \new_[51434]_ ,
    \new_[51435]_ , \new_[51439]_ , \new_[51440]_ , \new_[51443]_ ,
    \new_[51446]_ , \new_[51447]_ , \new_[51448]_ , \new_[51452]_ ,
    \new_[51453]_ , \new_[51457]_ , \new_[51458]_ , \new_[51459]_ ,
    \new_[51463]_ , \new_[51464]_ , \new_[51467]_ , \new_[51470]_ ,
    \new_[51471]_ , \new_[51472]_ , \new_[51476]_ , \new_[51477]_ ,
    \new_[51481]_ , \new_[51482]_ , \new_[51483]_ , \new_[51487]_ ,
    \new_[51488]_ , \new_[51491]_ , \new_[51494]_ , \new_[51495]_ ,
    \new_[51496]_ , \new_[51500]_ , \new_[51501]_ , \new_[51505]_ ,
    \new_[51506]_ , \new_[51507]_ , \new_[51511]_ , \new_[51512]_ ,
    \new_[51515]_ , \new_[51518]_ , \new_[51519]_ , \new_[51520]_ ,
    \new_[51524]_ , \new_[51525]_ , \new_[51529]_ , \new_[51530]_ ,
    \new_[51531]_ , \new_[51535]_ , \new_[51536]_ , \new_[51539]_ ,
    \new_[51542]_ , \new_[51543]_ , \new_[51544]_ , \new_[51548]_ ,
    \new_[51549]_ , \new_[51553]_ , \new_[51554]_ , \new_[51555]_ ,
    \new_[51559]_ , \new_[51560]_ , \new_[51563]_ , \new_[51566]_ ,
    \new_[51567]_ , \new_[51568]_ , \new_[51572]_ , \new_[51573]_ ,
    \new_[51577]_ , \new_[51578]_ , \new_[51579]_ , \new_[51583]_ ,
    \new_[51584]_ , \new_[51587]_ , \new_[51590]_ , \new_[51591]_ ,
    \new_[51592]_ , \new_[51596]_ , \new_[51597]_ , \new_[51601]_ ,
    \new_[51602]_ , \new_[51603]_ , \new_[51607]_ , \new_[51608]_ ,
    \new_[51611]_ , \new_[51614]_ , \new_[51615]_ , \new_[51616]_ ,
    \new_[51620]_ , \new_[51621]_ , \new_[51625]_ , \new_[51626]_ ,
    \new_[51627]_ , \new_[51631]_ , \new_[51632]_ , \new_[51635]_ ,
    \new_[51638]_ , \new_[51639]_ , \new_[51640]_ , \new_[51644]_ ,
    \new_[51645]_ , \new_[51649]_ , \new_[51650]_ , \new_[51651]_ ,
    \new_[51655]_ , \new_[51656]_ , \new_[51659]_ , \new_[51662]_ ,
    \new_[51663]_ , \new_[51664]_ , \new_[51668]_ , \new_[51669]_ ,
    \new_[51673]_ , \new_[51674]_ , \new_[51675]_ , \new_[51679]_ ,
    \new_[51680]_ , \new_[51683]_ , \new_[51686]_ , \new_[51687]_ ,
    \new_[51688]_ , \new_[51692]_ , \new_[51693]_ , \new_[51697]_ ,
    \new_[51698]_ , \new_[51699]_ , \new_[51703]_ , \new_[51704]_ ,
    \new_[51707]_ , \new_[51710]_ , \new_[51711]_ , \new_[51712]_ ,
    \new_[51716]_ , \new_[51717]_ , \new_[51721]_ , \new_[51722]_ ,
    \new_[51723]_ , \new_[51727]_ , \new_[51728]_ , \new_[51731]_ ,
    \new_[51734]_ , \new_[51735]_ , \new_[51736]_ , \new_[51740]_ ,
    \new_[51741]_ , \new_[51745]_ , \new_[51746]_ , \new_[51747]_ ,
    \new_[51751]_ , \new_[51752]_ , \new_[51755]_ , \new_[51758]_ ,
    \new_[51759]_ , \new_[51760]_ , \new_[51764]_ , \new_[51765]_ ,
    \new_[51769]_ , \new_[51770]_ , \new_[51771]_ , \new_[51775]_ ,
    \new_[51776]_ , \new_[51779]_ , \new_[51782]_ , \new_[51783]_ ,
    \new_[51784]_ , \new_[51788]_ , \new_[51789]_ , \new_[51793]_ ,
    \new_[51794]_ , \new_[51795]_ , \new_[51799]_ , \new_[51800]_ ,
    \new_[51803]_ , \new_[51806]_ , \new_[51807]_ , \new_[51808]_ ,
    \new_[51812]_ , \new_[51813]_ , \new_[51817]_ , \new_[51818]_ ,
    \new_[51819]_ , \new_[51823]_ , \new_[51824]_ , \new_[51827]_ ,
    \new_[51830]_ , \new_[51831]_ , \new_[51832]_ , \new_[51836]_ ,
    \new_[51837]_ , \new_[51841]_ , \new_[51842]_ , \new_[51843]_ ,
    \new_[51847]_ , \new_[51848]_ , \new_[51851]_ , \new_[51854]_ ,
    \new_[51855]_ , \new_[51856]_ , \new_[51860]_ , \new_[51861]_ ,
    \new_[51865]_ , \new_[51866]_ , \new_[51867]_ , \new_[51871]_ ,
    \new_[51872]_ , \new_[51875]_ , \new_[51878]_ , \new_[51879]_ ,
    \new_[51880]_ , \new_[51884]_ , \new_[51885]_ , \new_[51889]_ ,
    \new_[51890]_ , \new_[51891]_ , \new_[51895]_ , \new_[51896]_ ,
    \new_[51899]_ , \new_[51902]_ , \new_[51903]_ , \new_[51904]_ ,
    \new_[51908]_ , \new_[51909]_ , \new_[51913]_ , \new_[51914]_ ,
    \new_[51915]_ , \new_[51919]_ , \new_[51920]_ , \new_[51923]_ ,
    \new_[51926]_ , \new_[51927]_ , \new_[51928]_ , \new_[51932]_ ,
    \new_[51933]_ , \new_[51937]_ , \new_[51938]_ , \new_[51939]_ ,
    \new_[51943]_ , \new_[51944]_ , \new_[51947]_ , \new_[51950]_ ,
    \new_[51951]_ , \new_[51952]_ , \new_[51956]_ , \new_[51957]_ ,
    \new_[51961]_ , \new_[51962]_ , \new_[51963]_ , \new_[51967]_ ,
    \new_[51968]_ , \new_[51971]_ , \new_[51974]_ , \new_[51975]_ ,
    \new_[51976]_ , \new_[51980]_ , \new_[51981]_ , \new_[51985]_ ,
    \new_[51986]_ , \new_[51987]_ , \new_[51991]_ , \new_[51992]_ ,
    \new_[51995]_ , \new_[51998]_ , \new_[51999]_ , \new_[52000]_ ,
    \new_[52004]_ , \new_[52005]_ , \new_[52009]_ , \new_[52010]_ ,
    \new_[52011]_ , \new_[52015]_ , \new_[52016]_ , \new_[52019]_ ,
    \new_[52022]_ , \new_[52023]_ , \new_[52024]_ , \new_[52028]_ ,
    \new_[52029]_ , \new_[52033]_ , \new_[52034]_ , \new_[52035]_ ,
    \new_[52039]_ , \new_[52040]_ , \new_[52043]_ , \new_[52046]_ ,
    \new_[52047]_ , \new_[52048]_ , \new_[52052]_ , \new_[52053]_ ,
    \new_[52057]_ , \new_[52058]_ , \new_[52059]_ , \new_[52063]_ ,
    \new_[52064]_ , \new_[52067]_ , \new_[52070]_ , \new_[52071]_ ,
    \new_[52072]_ , \new_[52076]_ , \new_[52077]_ , \new_[52081]_ ,
    \new_[52082]_ , \new_[52083]_ , \new_[52087]_ , \new_[52088]_ ,
    \new_[52091]_ , \new_[52094]_ , \new_[52095]_ , \new_[52096]_ ,
    \new_[52100]_ , \new_[52101]_ , \new_[52105]_ , \new_[52106]_ ,
    \new_[52107]_ , \new_[52111]_ , \new_[52112]_ , \new_[52115]_ ,
    \new_[52118]_ , \new_[52119]_ , \new_[52120]_ , \new_[52124]_ ,
    \new_[52125]_ , \new_[52129]_ , \new_[52130]_ , \new_[52131]_ ,
    \new_[52135]_ , \new_[52136]_ , \new_[52139]_ , \new_[52142]_ ,
    \new_[52143]_ , \new_[52144]_ , \new_[52148]_ , \new_[52149]_ ,
    \new_[52153]_ , \new_[52154]_ , \new_[52155]_ , \new_[52159]_ ,
    \new_[52160]_ , \new_[52163]_ , \new_[52166]_ , \new_[52167]_ ,
    \new_[52168]_ , \new_[52172]_ , \new_[52173]_ , \new_[52177]_ ,
    \new_[52178]_ , \new_[52179]_ , \new_[52183]_ , \new_[52184]_ ,
    \new_[52187]_ , \new_[52190]_ , \new_[52191]_ , \new_[52192]_ ,
    \new_[52196]_ , \new_[52197]_ , \new_[52201]_ , \new_[52202]_ ,
    \new_[52203]_ , \new_[52207]_ , \new_[52208]_ , \new_[52211]_ ,
    \new_[52214]_ , \new_[52215]_ , \new_[52216]_ , \new_[52220]_ ,
    \new_[52221]_ , \new_[52225]_ , \new_[52226]_ , \new_[52227]_ ,
    \new_[52231]_ , \new_[52232]_ , \new_[52235]_ , \new_[52238]_ ,
    \new_[52239]_ , \new_[52240]_ , \new_[52244]_ , \new_[52245]_ ,
    \new_[52249]_ , \new_[52250]_ , \new_[52251]_ , \new_[52255]_ ,
    \new_[52256]_ , \new_[52259]_ , \new_[52262]_ , \new_[52263]_ ,
    \new_[52264]_ , \new_[52268]_ , \new_[52269]_ , \new_[52273]_ ,
    \new_[52274]_ , \new_[52275]_ , \new_[52279]_ , \new_[52280]_ ,
    \new_[52283]_ , \new_[52286]_ , \new_[52287]_ , \new_[52288]_ ,
    \new_[52292]_ , \new_[52293]_ , \new_[52297]_ , \new_[52298]_ ,
    \new_[52299]_ , \new_[52303]_ , \new_[52304]_ , \new_[52307]_ ,
    \new_[52310]_ , \new_[52311]_ , \new_[52312]_ , \new_[52316]_ ,
    \new_[52317]_ , \new_[52321]_ , \new_[52322]_ , \new_[52323]_ ,
    \new_[52327]_ , \new_[52328]_ , \new_[52331]_ , \new_[52334]_ ,
    \new_[52335]_ , \new_[52336]_ , \new_[52340]_ , \new_[52341]_ ,
    \new_[52345]_ , \new_[52346]_ , \new_[52347]_ , \new_[52351]_ ,
    \new_[52352]_ , \new_[52355]_ , \new_[52358]_ , \new_[52359]_ ,
    \new_[52360]_ , \new_[52364]_ , \new_[52365]_ , \new_[52369]_ ,
    \new_[52370]_ , \new_[52371]_ , \new_[52375]_ , \new_[52376]_ ,
    \new_[52379]_ , \new_[52382]_ , \new_[52383]_ , \new_[52384]_ ,
    \new_[52388]_ , \new_[52389]_ , \new_[52393]_ , \new_[52394]_ ,
    \new_[52395]_ , \new_[52399]_ , \new_[52400]_ , \new_[52403]_ ,
    \new_[52406]_ , \new_[52407]_ , \new_[52408]_ , \new_[52412]_ ,
    \new_[52413]_ , \new_[52417]_ , \new_[52418]_ , \new_[52419]_ ,
    \new_[52423]_ , \new_[52424]_ , \new_[52427]_ , \new_[52430]_ ,
    \new_[52431]_ , \new_[52432]_ , \new_[52436]_ , \new_[52437]_ ,
    \new_[52441]_ , \new_[52442]_ , \new_[52443]_ , \new_[52447]_ ,
    \new_[52448]_ , \new_[52451]_ , \new_[52454]_ , \new_[52455]_ ,
    \new_[52456]_ , \new_[52460]_ , \new_[52461]_ , \new_[52465]_ ,
    \new_[52466]_ , \new_[52467]_ , \new_[52471]_ , \new_[52472]_ ,
    \new_[52475]_ , \new_[52478]_ , \new_[52479]_ , \new_[52480]_ ,
    \new_[52484]_ , \new_[52485]_ , \new_[52489]_ , \new_[52490]_ ,
    \new_[52491]_ , \new_[52495]_ , \new_[52496]_ , \new_[52499]_ ,
    \new_[52502]_ , \new_[52503]_ , \new_[52504]_ , \new_[52508]_ ,
    \new_[52509]_ , \new_[52513]_ , \new_[52514]_ , \new_[52515]_ ,
    \new_[52519]_ , \new_[52520]_ , \new_[52523]_ , \new_[52526]_ ,
    \new_[52527]_ , \new_[52528]_ , \new_[52532]_ , \new_[52533]_ ,
    \new_[52537]_ , \new_[52538]_ , \new_[52539]_ , \new_[52543]_ ,
    \new_[52544]_ , \new_[52547]_ , \new_[52550]_ , \new_[52551]_ ,
    \new_[52552]_ , \new_[52556]_ , \new_[52557]_ , \new_[52561]_ ,
    \new_[52562]_ , \new_[52563]_ , \new_[52567]_ , \new_[52568]_ ,
    \new_[52571]_ , \new_[52574]_ , \new_[52575]_ , \new_[52576]_ ,
    \new_[52580]_ , \new_[52581]_ , \new_[52585]_ , \new_[52586]_ ,
    \new_[52587]_ , \new_[52591]_ , \new_[52592]_ , \new_[52595]_ ,
    \new_[52598]_ , \new_[52599]_ , \new_[52600]_ , \new_[52604]_ ,
    \new_[52605]_ , \new_[52609]_ , \new_[52610]_ , \new_[52611]_ ,
    \new_[52615]_ , \new_[52616]_ , \new_[52619]_ , \new_[52622]_ ,
    \new_[52623]_ , \new_[52624]_ , \new_[52628]_ , \new_[52629]_ ,
    \new_[52633]_ , \new_[52634]_ , \new_[52635]_ , \new_[52639]_ ,
    \new_[52640]_ , \new_[52643]_ , \new_[52646]_ , \new_[52647]_ ,
    \new_[52648]_ , \new_[52652]_ , \new_[52653]_ , \new_[52657]_ ,
    \new_[52658]_ , \new_[52659]_ , \new_[52663]_ , \new_[52664]_ ,
    \new_[52667]_ , \new_[52670]_ , \new_[52671]_ , \new_[52672]_ ,
    \new_[52676]_ , \new_[52677]_ , \new_[52681]_ , \new_[52682]_ ,
    \new_[52683]_ , \new_[52687]_ , \new_[52688]_ , \new_[52691]_ ,
    \new_[52694]_ , \new_[52695]_ , \new_[52696]_ , \new_[52700]_ ,
    \new_[52701]_ , \new_[52705]_ , \new_[52706]_ , \new_[52707]_ ,
    \new_[52711]_ , \new_[52712]_ , \new_[52715]_ , \new_[52718]_ ,
    \new_[52719]_ , \new_[52720]_ , \new_[52724]_ , \new_[52725]_ ,
    \new_[52729]_ , \new_[52730]_ , \new_[52731]_ , \new_[52735]_ ,
    \new_[52736]_ , \new_[52739]_ , \new_[52742]_ , \new_[52743]_ ,
    \new_[52744]_ , \new_[52748]_ , \new_[52749]_ , \new_[52753]_ ,
    \new_[52754]_ , \new_[52755]_ , \new_[52759]_ , \new_[52760]_ ,
    \new_[52763]_ , \new_[52766]_ , \new_[52767]_ , \new_[52768]_ ,
    \new_[52772]_ , \new_[52773]_ , \new_[52777]_ , \new_[52778]_ ,
    \new_[52779]_ , \new_[52783]_ , \new_[52784]_ , \new_[52787]_ ,
    \new_[52790]_ , \new_[52791]_ , \new_[52792]_ , \new_[52796]_ ,
    \new_[52797]_ , \new_[52801]_ , \new_[52802]_ , \new_[52803]_ ,
    \new_[52807]_ , \new_[52808]_ , \new_[52811]_ , \new_[52814]_ ,
    \new_[52815]_ , \new_[52816]_ , \new_[52820]_ , \new_[52821]_ ,
    \new_[52825]_ , \new_[52826]_ , \new_[52827]_ , \new_[52831]_ ,
    \new_[52832]_ , \new_[52835]_ , \new_[52838]_ , \new_[52839]_ ,
    \new_[52840]_ , \new_[52844]_ , \new_[52845]_ , \new_[52849]_ ,
    \new_[52850]_ , \new_[52851]_ , \new_[52855]_ , \new_[52856]_ ,
    \new_[52859]_ , \new_[52862]_ , \new_[52863]_ , \new_[52864]_ ,
    \new_[52868]_ , \new_[52869]_ , \new_[52873]_ , \new_[52874]_ ,
    \new_[52875]_ , \new_[52879]_ , \new_[52880]_ , \new_[52883]_ ,
    \new_[52886]_ , \new_[52887]_ , \new_[52888]_ , \new_[52892]_ ,
    \new_[52893]_ , \new_[52897]_ , \new_[52898]_ , \new_[52899]_ ,
    \new_[52903]_ , \new_[52904]_ , \new_[52907]_ , \new_[52910]_ ,
    \new_[52911]_ , \new_[52912]_ , \new_[52916]_ , \new_[52917]_ ,
    \new_[52921]_ , \new_[52922]_ , \new_[52923]_ , \new_[52927]_ ,
    \new_[52928]_ , \new_[52931]_ , \new_[52934]_ , \new_[52935]_ ,
    \new_[52936]_ , \new_[52940]_ , \new_[52941]_ , \new_[52945]_ ,
    \new_[52946]_ , \new_[52947]_ , \new_[52951]_ , \new_[52952]_ ,
    \new_[52955]_ , \new_[52958]_ , \new_[52959]_ , \new_[52960]_ ,
    \new_[52964]_ , \new_[52965]_ , \new_[52969]_ , \new_[52970]_ ,
    \new_[52971]_ , \new_[52975]_ , \new_[52976]_ , \new_[52979]_ ,
    \new_[52982]_ , \new_[52983]_ , \new_[52984]_ , \new_[52988]_ ,
    \new_[52989]_ , \new_[52993]_ , \new_[52994]_ , \new_[52995]_ ,
    \new_[52999]_ , \new_[53000]_ , \new_[53003]_ , \new_[53006]_ ,
    \new_[53007]_ , \new_[53008]_ , \new_[53012]_ , \new_[53013]_ ,
    \new_[53017]_ , \new_[53018]_ , \new_[53019]_ , \new_[53023]_ ,
    \new_[53024]_ , \new_[53027]_ , \new_[53030]_ , \new_[53031]_ ,
    \new_[53032]_ , \new_[53036]_ , \new_[53037]_ , \new_[53041]_ ,
    \new_[53042]_ , \new_[53043]_ , \new_[53047]_ , \new_[53048]_ ,
    \new_[53051]_ , \new_[53054]_ , \new_[53055]_ , \new_[53056]_ ,
    \new_[53060]_ , \new_[53061]_ , \new_[53065]_ , \new_[53066]_ ,
    \new_[53067]_ , \new_[53071]_ , \new_[53072]_ , \new_[53075]_ ,
    \new_[53078]_ , \new_[53079]_ , \new_[53080]_ , \new_[53084]_ ,
    \new_[53085]_ , \new_[53089]_ , \new_[53090]_ , \new_[53091]_ ,
    \new_[53095]_ , \new_[53096]_ , \new_[53099]_ , \new_[53102]_ ,
    \new_[53103]_ , \new_[53104]_ , \new_[53108]_ , \new_[53109]_ ,
    \new_[53113]_ , \new_[53114]_ , \new_[53115]_ , \new_[53119]_ ,
    \new_[53120]_ , \new_[53123]_ , \new_[53126]_ , \new_[53127]_ ,
    \new_[53128]_ , \new_[53132]_ , \new_[53133]_ , \new_[53137]_ ,
    \new_[53138]_ , \new_[53139]_ , \new_[53143]_ , \new_[53144]_ ,
    \new_[53147]_ , \new_[53150]_ , \new_[53151]_ , \new_[53152]_ ,
    \new_[53156]_ , \new_[53157]_ , \new_[53161]_ , \new_[53162]_ ,
    \new_[53163]_ , \new_[53167]_ , \new_[53168]_ , \new_[53171]_ ,
    \new_[53174]_ , \new_[53175]_ , \new_[53176]_ , \new_[53180]_ ,
    \new_[53181]_ , \new_[53185]_ , \new_[53186]_ , \new_[53187]_ ,
    \new_[53191]_ , \new_[53192]_ , \new_[53195]_ , \new_[53198]_ ,
    \new_[53199]_ , \new_[53200]_ , \new_[53204]_ , \new_[53205]_ ,
    \new_[53209]_ , \new_[53210]_ , \new_[53211]_ , \new_[53215]_ ,
    \new_[53216]_ , \new_[53219]_ , \new_[53222]_ , \new_[53223]_ ,
    \new_[53224]_ , \new_[53228]_ , \new_[53229]_ , \new_[53233]_ ,
    \new_[53234]_ , \new_[53235]_ , \new_[53239]_ , \new_[53240]_ ,
    \new_[53243]_ , \new_[53246]_ , \new_[53247]_ , \new_[53248]_ ,
    \new_[53252]_ , \new_[53253]_ , \new_[53257]_ , \new_[53258]_ ,
    \new_[53259]_ , \new_[53263]_ , \new_[53264]_ , \new_[53267]_ ,
    \new_[53270]_ , \new_[53271]_ , \new_[53272]_ , \new_[53276]_ ,
    \new_[53277]_ , \new_[53281]_ , \new_[53282]_ , \new_[53283]_ ,
    \new_[53287]_ , \new_[53288]_ , \new_[53291]_ , \new_[53294]_ ,
    \new_[53295]_ , \new_[53296]_ , \new_[53300]_ , \new_[53301]_ ,
    \new_[53305]_ , \new_[53306]_ , \new_[53307]_ , \new_[53311]_ ,
    \new_[53312]_ , \new_[53315]_ , \new_[53318]_ , \new_[53319]_ ,
    \new_[53320]_ , \new_[53324]_ , \new_[53325]_ , \new_[53329]_ ,
    \new_[53330]_ , \new_[53331]_ , \new_[53335]_ , \new_[53336]_ ,
    \new_[53339]_ , \new_[53342]_ , \new_[53343]_ , \new_[53344]_ ,
    \new_[53348]_ , \new_[53349]_ , \new_[53353]_ , \new_[53354]_ ,
    \new_[53355]_ , \new_[53359]_ , \new_[53360]_ , \new_[53363]_ ,
    \new_[53366]_ , \new_[53367]_ , \new_[53368]_ , \new_[53372]_ ,
    \new_[53373]_ , \new_[53377]_ , \new_[53378]_ , \new_[53379]_ ,
    \new_[53383]_ , \new_[53384]_ , \new_[53387]_ , \new_[53390]_ ,
    \new_[53391]_ , \new_[53392]_ , \new_[53396]_ , \new_[53397]_ ,
    \new_[53401]_ , \new_[53402]_ , \new_[53403]_ , \new_[53407]_ ,
    \new_[53408]_ , \new_[53411]_ , \new_[53414]_ , \new_[53415]_ ,
    \new_[53416]_ , \new_[53420]_ , \new_[53421]_ , \new_[53425]_ ,
    \new_[53426]_ , \new_[53427]_ , \new_[53431]_ , \new_[53432]_ ,
    \new_[53435]_ , \new_[53438]_ , \new_[53439]_ , \new_[53440]_ ,
    \new_[53444]_ , \new_[53445]_ , \new_[53449]_ , \new_[53450]_ ,
    \new_[53451]_ , \new_[53455]_ , \new_[53456]_ , \new_[53459]_ ,
    \new_[53462]_ , \new_[53463]_ , \new_[53464]_ , \new_[53468]_ ,
    \new_[53469]_ , \new_[53473]_ , \new_[53474]_ , \new_[53475]_ ,
    \new_[53479]_ , \new_[53480]_ , \new_[53483]_ , \new_[53486]_ ,
    \new_[53487]_ , \new_[53488]_ , \new_[53492]_ , \new_[53493]_ ,
    \new_[53497]_ , \new_[53498]_ , \new_[53499]_ , \new_[53503]_ ,
    \new_[53504]_ , \new_[53507]_ , \new_[53510]_ , \new_[53511]_ ,
    \new_[53512]_ , \new_[53516]_ , \new_[53517]_ , \new_[53521]_ ,
    \new_[53522]_ , \new_[53523]_ , \new_[53527]_ , \new_[53528]_ ,
    \new_[53531]_ , \new_[53534]_ , \new_[53535]_ , \new_[53536]_ ,
    \new_[53540]_ , \new_[53541]_ , \new_[53545]_ , \new_[53546]_ ,
    \new_[53547]_ , \new_[53551]_ , \new_[53552]_ , \new_[53555]_ ,
    \new_[53558]_ , \new_[53559]_ , \new_[53560]_ , \new_[53564]_ ,
    \new_[53565]_ , \new_[53569]_ , \new_[53570]_ , \new_[53571]_ ,
    \new_[53575]_ , \new_[53576]_ , \new_[53579]_ , \new_[53582]_ ,
    \new_[53583]_ , \new_[53584]_ , \new_[53588]_ , \new_[53589]_ ,
    \new_[53593]_ , \new_[53594]_ , \new_[53595]_ , \new_[53599]_ ,
    \new_[53600]_ , \new_[53603]_ , \new_[53606]_ , \new_[53607]_ ,
    \new_[53608]_ , \new_[53612]_ , \new_[53613]_ , \new_[53617]_ ,
    \new_[53618]_ , \new_[53619]_ , \new_[53623]_ , \new_[53624]_ ,
    \new_[53627]_ , \new_[53630]_ , \new_[53631]_ , \new_[53632]_ ,
    \new_[53636]_ , \new_[53637]_ , \new_[53641]_ , \new_[53642]_ ,
    \new_[53643]_ , \new_[53647]_ , \new_[53648]_ , \new_[53651]_ ,
    \new_[53654]_ , \new_[53655]_ , \new_[53656]_ , \new_[53660]_ ,
    \new_[53661]_ , \new_[53665]_ , \new_[53666]_ , \new_[53667]_ ,
    \new_[53671]_ , \new_[53672]_ , \new_[53675]_ , \new_[53678]_ ,
    \new_[53679]_ , \new_[53680]_ , \new_[53684]_ , \new_[53685]_ ,
    \new_[53689]_ , \new_[53690]_ , \new_[53691]_ , \new_[53695]_ ,
    \new_[53696]_ , \new_[53699]_ , \new_[53702]_ , \new_[53703]_ ,
    \new_[53704]_ , \new_[53708]_ , \new_[53709]_ , \new_[53713]_ ,
    \new_[53714]_ , \new_[53715]_ , \new_[53719]_ , \new_[53720]_ ,
    \new_[53723]_ , \new_[53726]_ , \new_[53727]_ , \new_[53728]_ ,
    \new_[53732]_ , \new_[53733]_ , \new_[53737]_ , \new_[53738]_ ,
    \new_[53739]_ , \new_[53743]_ , \new_[53744]_ , \new_[53747]_ ,
    \new_[53750]_ , \new_[53751]_ , \new_[53752]_ , \new_[53756]_ ,
    \new_[53757]_ , \new_[53761]_ , \new_[53762]_ , \new_[53763]_ ,
    \new_[53767]_ , \new_[53768]_ , \new_[53771]_ , \new_[53774]_ ,
    \new_[53775]_ , \new_[53776]_ , \new_[53780]_ , \new_[53781]_ ,
    \new_[53785]_ , \new_[53786]_ , \new_[53787]_ , \new_[53791]_ ,
    \new_[53792]_ , \new_[53795]_ , \new_[53798]_ , \new_[53799]_ ,
    \new_[53800]_ , \new_[53804]_ , \new_[53805]_ , \new_[53809]_ ,
    \new_[53810]_ , \new_[53811]_ , \new_[53815]_ , \new_[53816]_ ,
    \new_[53819]_ , \new_[53822]_ , \new_[53823]_ , \new_[53824]_ ,
    \new_[53828]_ , \new_[53829]_ , \new_[53833]_ , \new_[53834]_ ,
    \new_[53835]_ , \new_[53839]_ , \new_[53840]_ , \new_[53843]_ ,
    \new_[53846]_ , \new_[53847]_ , \new_[53848]_ , \new_[53852]_ ,
    \new_[53853]_ , \new_[53857]_ , \new_[53858]_ , \new_[53859]_ ,
    \new_[53863]_ , \new_[53864]_ , \new_[53867]_ , \new_[53870]_ ,
    \new_[53871]_ , \new_[53872]_ , \new_[53876]_ , \new_[53877]_ ,
    \new_[53881]_ , \new_[53882]_ , \new_[53883]_ , \new_[53887]_ ,
    \new_[53888]_ , \new_[53891]_ , \new_[53894]_ , \new_[53895]_ ,
    \new_[53896]_ , \new_[53900]_ , \new_[53901]_ , \new_[53905]_ ,
    \new_[53906]_ , \new_[53907]_ , \new_[53911]_ , \new_[53912]_ ,
    \new_[53915]_ , \new_[53918]_ , \new_[53919]_ , \new_[53920]_ ,
    \new_[53924]_ , \new_[53925]_ , \new_[53929]_ , \new_[53930]_ ,
    \new_[53931]_ , \new_[53935]_ , \new_[53936]_ , \new_[53939]_ ,
    \new_[53942]_ , \new_[53943]_ , \new_[53944]_ , \new_[53948]_ ,
    \new_[53949]_ , \new_[53953]_ , \new_[53954]_ , \new_[53955]_ ,
    \new_[53959]_ , \new_[53960]_ , \new_[53963]_ , \new_[53966]_ ,
    \new_[53967]_ , \new_[53968]_ , \new_[53972]_ , \new_[53973]_ ,
    \new_[53977]_ , \new_[53978]_ , \new_[53979]_ , \new_[53983]_ ,
    \new_[53984]_ , \new_[53987]_ , \new_[53990]_ , \new_[53991]_ ,
    \new_[53992]_ , \new_[53996]_ , \new_[53997]_ , \new_[54001]_ ,
    \new_[54002]_ , \new_[54003]_ , \new_[54007]_ , \new_[54008]_ ,
    \new_[54011]_ , \new_[54014]_ , \new_[54015]_ , \new_[54016]_ ,
    \new_[54020]_ , \new_[54021]_ , \new_[54025]_ , \new_[54026]_ ,
    \new_[54027]_ , \new_[54031]_ , \new_[54032]_ , \new_[54035]_ ,
    \new_[54038]_ , \new_[54039]_ , \new_[54040]_ , \new_[54044]_ ,
    \new_[54045]_ , \new_[54049]_ , \new_[54050]_ , \new_[54051]_ ,
    \new_[54055]_ , \new_[54056]_ , \new_[54059]_ , \new_[54062]_ ,
    \new_[54063]_ , \new_[54064]_ , \new_[54068]_ , \new_[54069]_ ,
    \new_[54073]_ , \new_[54074]_ , \new_[54075]_ , \new_[54079]_ ,
    \new_[54080]_ , \new_[54083]_ , \new_[54086]_ , \new_[54087]_ ,
    \new_[54088]_ , \new_[54092]_ , \new_[54093]_ , \new_[54097]_ ,
    \new_[54098]_ , \new_[54099]_ , \new_[54103]_ , \new_[54104]_ ,
    \new_[54107]_ , \new_[54110]_ , \new_[54111]_ , \new_[54112]_ ,
    \new_[54116]_ , \new_[54117]_ , \new_[54121]_ , \new_[54122]_ ,
    \new_[54123]_ , \new_[54127]_ , \new_[54128]_ , \new_[54131]_ ,
    \new_[54134]_ , \new_[54135]_ , \new_[54136]_ , \new_[54140]_ ,
    \new_[54141]_ , \new_[54145]_ , \new_[54146]_ , \new_[54147]_ ,
    \new_[54151]_ , \new_[54152]_ , \new_[54155]_ , \new_[54158]_ ,
    \new_[54159]_ , \new_[54160]_ , \new_[54164]_ , \new_[54165]_ ,
    \new_[54169]_ , \new_[54170]_ , \new_[54171]_ , \new_[54175]_ ,
    \new_[54176]_ , \new_[54179]_ , \new_[54182]_ , \new_[54183]_ ,
    \new_[54184]_ , \new_[54188]_ , \new_[54189]_ , \new_[54193]_ ,
    \new_[54194]_ , \new_[54195]_ , \new_[54199]_ , \new_[54200]_ ,
    \new_[54203]_ , \new_[54206]_ , \new_[54207]_ , \new_[54208]_ ,
    \new_[54212]_ , \new_[54213]_ , \new_[54217]_ , \new_[54218]_ ,
    \new_[54219]_ , \new_[54223]_ , \new_[54224]_ , \new_[54227]_ ,
    \new_[54230]_ , \new_[54231]_ , \new_[54232]_ , \new_[54236]_ ,
    \new_[54237]_ , \new_[54241]_ , \new_[54242]_ , \new_[54243]_ ,
    \new_[54247]_ , \new_[54248]_ , \new_[54251]_ , \new_[54254]_ ,
    \new_[54255]_ , \new_[54256]_ , \new_[54260]_ , \new_[54261]_ ,
    \new_[54265]_ , \new_[54266]_ , \new_[54267]_ , \new_[54271]_ ,
    \new_[54272]_ , \new_[54275]_ , \new_[54278]_ , \new_[54279]_ ,
    \new_[54280]_ , \new_[54284]_ , \new_[54285]_ , \new_[54289]_ ,
    \new_[54290]_ , \new_[54291]_ , \new_[54295]_ , \new_[54296]_ ,
    \new_[54299]_ , \new_[54302]_ , \new_[54303]_ , \new_[54304]_ ,
    \new_[54308]_ , \new_[54309]_ , \new_[54313]_ , \new_[54314]_ ,
    \new_[54315]_ , \new_[54319]_ , \new_[54320]_ , \new_[54323]_ ,
    \new_[54326]_ , \new_[54327]_ , \new_[54328]_ , \new_[54332]_ ,
    \new_[54333]_ , \new_[54337]_ , \new_[54338]_ , \new_[54339]_ ,
    \new_[54343]_ , \new_[54344]_ , \new_[54347]_ , \new_[54350]_ ,
    \new_[54351]_ , \new_[54352]_ , \new_[54356]_ , \new_[54357]_ ,
    \new_[54361]_ , \new_[54362]_ , \new_[54363]_ , \new_[54367]_ ,
    \new_[54368]_ , \new_[54371]_ , \new_[54374]_ , \new_[54375]_ ,
    \new_[54376]_ , \new_[54380]_ , \new_[54381]_ , \new_[54385]_ ,
    \new_[54386]_ , \new_[54387]_ , \new_[54391]_ , \new_[54392]_ ,
    \new_[54395]_ , \new_[54398]_ , \new_[54399]_ , \new_[54400]_ ,
    \new_[54404]_ , \new_[54405]_ , \new_[54409]_ , \new_[54410]_ ,
    \new_[54411]_ , \new_[54415]_ , \new_[54416]_ , \new_[54419]_ ,
    \new_[54422]_ , \new_[54423]_ , \new_[54424]_ , \new_[54428]_ ,
    \new_[54429]_ , \new_[54433]_ , \new_[54434]_ , \new_[54435]_ ,
    \new_[54439]_ , \new_[54440]_ , \new_[54443]_ , \new_[54446]_ ,
    \new_[54447]_ , \new_[54448]_ , \new_[54452]_ , \new_[54453]_ ,
    \new_[54457]_ , \new_[54458]_ , \new_[54459]_ , \new_[54463]_ ,
    \new_[54464]_ , \new_[54467]_ , \new_[54470]_ , \new_[54471]_ ,
    \new_[54472]_ , \new_[54476]_ , \new_[54477]_ , \new_[54481]_ ,
    \new_[54482]_ , \new_[54483]_ , \new_[54487]_ , \new_[54488]_ ,
    \new_[54491]_ , \new_[54494]_ , \new_[54495]_ , \new_[54496]_ ,
    \new_[54500]_ , \new_[54501]_ , \new_[54505]_ , \new_[54506]_ ,
    \new_[54507]_ , \new_[54511]_ , \new_[54512]_ , \new_[54515]_ ,
    \new_[54518]_ , \new_[54519]_ , \new_[54520]_ , \new_[54524]_ ,
    \new_[54525]_ , \new_[54529]_ , \new_[54530]_ , \new_[54531]_ ,
    \new_[54535]_ , \new_[54536]_ , \new_[54539]_ , \new_[54542]_ ,
    \new_[54543]_ , \new_[54544]_ , \new_[54548]_ , \new_[54549]_ ,
    \new_[54553]_ , \new_[54554]_ , \new_[54555]_ , \new_[54559]_ ,
    \new_[54560]_ , \new_[54563]_ , \new_[54566]_ , \new_[54567]_ ,
    \new_[54568]_ , \new_[54572]_ , \new_[54573]_ , \new_[54577]_ ,
    \new_[54578]_ , \new_[54579]_ , \new_[54583]_ , \new_[54584]_ ,
    \new_[54587]_ , \new_[54590]_ , \new_[54591]_ , \new_[54592]_ ,
    \new_[54596]_ , \new_[54597]_ , \new_[54601]_ , \new_[54602]_ ,
    \new_[54603]_ , \new_[54607]_ , \new_[54608]_ , \new_[54611]_ ,
    \new_[54614]_ , \new_[54615]_ , \new_[54616]_ , \new_[54620]_ ,
    \new_[54621]_ , \new_[54625]_ , \new_[54626]_ , \new_[54627]_ ,
    \new_[54631]_ , \new_[54632]_ , \new_[54635]_ , \new_[54638]_ ,
    \new_[54639]_ , \new_[54640]_ , \new_[54644]_ , \new_[54645]_ ,
    \new_[54649]_ , \new_[54650]_ , \new_[54651]_ , \new_[54655]_ ,
    \new_[54656]_ , \new_[54659]_ , \new_[54662]_ , \new_[54663]_ ,
    \new_[54664]_ , \new_[54668]_ , \new_[54669]_ , \new_[54673]_ ,
    \new_[54674]_ , \new_[54675]_ , \new_[54679]_ , \new_[54680]_ ,
    \new_[54683]_ , \new_[54686]_ , \new_[54687]_ , \new_[54688]_ ,
    \new_[54692]_ , \new_[54693]_ , \new_[54697]_ , \new_[54698]_ ,
    \new_[54699]_ , \new_[54703]_ , \new_[54704]_ , \new_[54707]_ ,
    \new_[54710]_ , \new_[54711]_ , \new_[54712]_ , \new_[54716]_ ,
    \new_[54717]_ , \new_[54721]_ , \new_[54722]_ , \new_[54723]_ ,
    \new_[54727]_ , \new_[54728]_ , \new_[54731]_ , \new_[54734]_ ,
    \new_[54735]_ , \new_[54736]_ , \new_[54740]_ , \new_[54741]_ ,
    \new_[54745]_ , \new_[54746]_ , \new_[54747]_ , \new_[54751]_ ,
    \new_[54752]_ , \new_[54755]_ , \new_[54758]_ , \new_[54759]_ ,
    \new_[54760]_ , \new_[54764]_ , \new_[54765]_ , \new_[54769]_ ,
    \new_[54770]_ , \new_[54771]_ , \new_[54775]_ , \new_[54776]_ ,
    \new_[54779]_ , \new_[54782]_ , \new_[54783]_ , \new_[54784]_ ,
    \new_[54788]_ , \new_[54789]_ , \new_[54793]_ , \new_[54794]_ ,
    \new_[54795]_ , \new_[54799]_ , \new_[54800]_ , \new_[54803]_ ,
    \new_[54806]_ , \new_[54807]_ , \new_[54808]_ , \new_[54812]_ ,
    \new_[54813]_ , \new_[54817]_ , \new_[54818]_ , \new_[54819]_ ,
    \new_[54823]_ , \new_[54824]_ , \new_[54827]_ , \new_[54830]_ ,
    \new_[54831]_ , \new_[54832]_ , \new_[54836]_ , \new_[54837]_ ,
    \new_[54841]_ , \new_[54842]_ , \new_[54843]_ , \new_[54847]_ ,
    \new_[54848]_ , \new_[54851]_ , \new_[54854]_ , \new_[54855]_ ,
    \new_[54856]_ , \new_[54860]_ , \new_[54861]_ , \new_[54865]_ ,
    \new_[54866]_ , \new_[54867]_ , \new_[54871]_ , \new_[54872]_ ,
    \new_[54875]_ , \new_[54878]_ , \new_[54879]_ , \new_[54880]_ ,
    \new_[54884]_ , \new_[54885]_ , \new_[54889]_ , \new_[54890]_ ,
    \new_[54891]_ , \new_[54895]_ , \new_[54896]_ , \new_[54899]_ ,
    \new_[54902]_ , \new_[54903]_ , \new_[54904]_ , \new_[54908]_ ,
    \new_[54909]_ , \new_[54913]_ , \new_[54914]_ , \new_[54915]_ ,
    \new_[54919]_ , \new_[54920]_ , \new_[54923]_ , \new_[54926]_ ,
    \new_[54927]_ , \new_[54928]_ , \new_[54932]_ , \new_[54933]_ ,
    \new_[54937]_ , \new_[54938]_ , \new_[54939]_ , \new_[54943]_ ,
    \new_[54944]_ , \new_[54947]_ , \new_[54950]_ , \new_[54951]_ ,
    \new_[54952]_ , \new_[54956]_ , \new_[54957]_ , \new_[54961]_ ,
    \new_[54962]_ , \new_[54963]_ , \new_[54967]_ , \new_[54968]_ ,
    \new_[54971]_ , \new_[54974]_ , \new_[54975]_ , \new_[54976]_ ,
    \new_[54980]_ , \new_[54981]_ , \new_[54985]_ , \new_[54986]_ ,
    \new_[54987]_ , \new_[54991]_ , \new_[54992]_ , \new_[54995]_ ,
    \new_[54998]_ , \new_[54999]_ , \new_[55000]_ , \new_[55004]_ ,
    \new_[55005]_ , \new_[55009]_ , \new_[55010]_ , \new_[55011]_ ,
    \new_[55015]_ , \new_[55016]_ , \new_[55019]_ , \new_[55022]_ ,
    \new_[55023]_ , \new_[55024]_ , \new_[55028]_ , \new_[55029]_ ,
    \new_[55033]_ , \new_[55034]_ , \new_[55035]_ , \new_[55039]_ ,
    \new_[55040]_ , \new_[55043]_ , \new_[55046]_ , \new_[55047]_ ,
    \new_[55048]_ , \new_[55052]_ , \new_[55053]_ , \new_[55057]_ ,
    \new_[55058]_ , \new_[55059]_ , \new_[55063]_ , \new_[55064]_ ,
    \new_[55067]_ , \new_[55070]_ , \new_[55071]_ , \new_[55072]_ ,
    \new_[55076]_ , \new_[55077]_ , \new_[55081]_ , \new_[55082]_ ,
    \new_[55083]_ , \new_[55087]_ , \new_[55088]_ , \new_[55091]_ ,
    \new_[55094]_ , \new_[55095]_ , \new_[55096]_ , \new_[55100]_ ,
    \new_[55101]_ , \new_[55105]_ , \new_[55106]_ , \new_[55107]_ ,
    \new_[55111]_ , \new_[55112]_ , \new_[55115]_ , \new_[55118]_ ,
    \new_[55119]_ , \new_[55120]_ , \new_[55124]_ , \new_[55125]_ ,
    \new_[55129]_ , \new_[55130]_ , \new_[55131]_ , \new_[55135]_ ,
    \new_[55136]_ , \new_[55139]_ , \new_[55142]_ , \new_[55143]_ ,
    \new_[55144]_ , \new_[55148]_ , \new_[55149]_ , \new_[55153]_ ,
    \new_[55154]_ , \new_[55155]_ , \new_[55159]_ , \new_[55160]_ ,
    \new_[55163]_ , \new_[55166]_ , \new_[55167]_ , \new_[55168]_ ,
    \new_[55172]_ , \new_[55173]_ , \new_[55177]_ , \new_[55178]_ ,
    \new_[55179]_ , \new_[55183]_ , \new_[55184]_ , \new_[55187]_ ,
    \new_[55190]_ , \new_[55191]_ , \new_[55192]_ , \new_[55196]_ ,
    \new_[55197]_ , \new_[55201]_ , \new_[55202]_ , \new_[55203]_ ,
    \new_[55207]_ , \new_[55208]_ , \new_[55211]_ , \new_[55214]_ ,
    \new_[55215]_ , \new_[55216]_ , \new_[55220]_ , \new_[55221]_ ,
    \new_[55225]_ , \new_[55226]_ , \new_[55227]_ , \new_[55231]_ ,
    \new_[55232]_ , \new_[55235]_ , \new_[55238]_ , \new_[55239]_ ,
    \new_[55240]_ , \new_[55244]_ , \new_[55245]_ , \new_[55249]_ ,
    \new_[55250]_ , \new_[55251]_ , \new_[55255]_ , \new_[55256]_ ,
    \new_[55259]_ , \new_[55262]_ , \new_[55263]_ , \new_[55264]_ ,
    \new_[55268]_ , \new_[55269]_ , \new_[55273]_ , \new_[55274]_ ,
    \new_[55275]_ , \new_[55279]_ , \new_[55280]_ , \new_[55283]_ ,
    \new_[55286]_ , \new_[55287]_ , \new_[55288]_ , \new_[55292]_ ,
    \new_[55293]_ , \new_[55297]_ , \new_[55298]_ , \new_[55299]_ ,
    \new_[55303]_ , \new_[55304]_ , \new_[55307]_ , \new_[55310]_ ,
    \new_[55311]_ , \new_[55312]_ , \new_[55316]_ , \new_[55317]_ ,
    \new_[55321]_ , \new_[55322]_ , \new_[55323]_ , \new_[55327]_ ,
    \new_[55328]_ , \new_[55331]_ , \new_[55334]_ , \new_[55335]_ ,
    \new_[55336]_ , \new_[55340]_ , \new_[55341]_ , \new_[55345]_ ,
    \new_[55346]_ , \new_[55347]_ , \new_[55351]_ , \new_[55352]_ ,
    \new_[55355]_ , \new_[55358]_ , \new_[55359]_ , \new_[55360]_ ,
    \new_[55364]_ , \new_[55365]_ , \new_[55369]_ , \new_[55370]_ ,
    \new_[55371]_ , \new_[55375]_ , \new_[55376]_ , \new_[55379]_ ,
    \new_[55382]_ , \new_[55383]_ , \new_[55384]_ , \new_[55388]_ ,
    \new_[55389]_ , \new_[55393]_ , \new_[55394]_ , \new_[55395]_ ,
    \new_[55399]_ , \new_[55400]_ , \new_[55403]_ , \new_[55406]_ ,
    \new_[55407]_ , \new_[55408]_ , \new_[55412]_ , \new_[55413]_ ,
    \new_[55417]_ , \new_[55418]_ , \new_[55419]_ , \new_[55423]_ ,
    \new_[55424]_ , \new_[55427]_ , \new_[55430]_ , \new_[55431]_ ,
    \new_[55432]_ , \new_[55436]_ , \new_[55437]_ , \new_[55441]_ ,
    \new_[55442]_ , \new_[55443]_ , \new_[55447]_ , \new_[55448]_ ,
    \new_[55451]_ , \new_[55454]_ , \new_[55455]_ , \new_[55456]_ ,
    \new_[55460]_ , \new_[55461]_ , \new_[55465]_ , \new_[55466]_ ,
    \new_[55467]_ , \new_[55471]_ , \new_[55472]_ , \new_[55475]_ ,
    \new_[55478]_ , \new_[55479]_ , \new_[55480]_ , \new_[55484]_ ,
    \new_[55485]_ , \new_[55489]_ , \new_[55490]_ , \new_[55491]_ ,
    \new_[55495]_ , \new_[55496]_ , \new_[55499]_ , \new_[55502]_ ,
    \new_[55503]_ , \new_[55504]_ , \new_[55508]_ , \new_[55509]_ ,
    \new_[55513]_ , \new_[55514]_ , \new_[55515]_ , \new_[55519]_ ,
    \new_[55520]_ , \new_[55523]_ , \new_[55526]_ , \new_[55527]_ ,
    \new_[55528]_ , \new_[55532]_ , \new_[55533]_ , \new_[55537]_ ,
    \new_[55538]_ , \new_[55539]_ , \new_[55543]_ , \new_[55544]_ ,
    \new_[55547]_ , \new_[55550]_ , \new_[55551]_ , \new_[55552]_ ,
    \new_[55556]_ , \new_[55557]_ , \new_[55561]_ , \new_[55562]_ ,
    \new_[55563]_ , \new_[55567]_ , \new_[55568]_ , \new_[55571]_ ,
    \new_[55574]_ , \new_[55575]_ , \new_[55576]_ , \new_[55580]_ ,
    \new_[55581]_ , \new_[55585]_ , \new_[55586]_ , \new_[55587]_ ,
    \new_[55591]_ , \new_[55592]_ , \new_[55595]_ , \new_[55598]_ ,
    \new_[55599]_ , \new_[55600]_ , \new_[55604]_ , \new_[55605]_ ,
    \new_[55609]_ , \new_[55610]_ , \new_[55611]_ , \new_[55615]_ ,
    \new_[55616]_ , \new_[55619]_ , \new_[55622]_ , \new_[55623]_ ,
    \new_[55624]_ , \new_[55628]_ , \new_[55629]_ , \new_[55633]_ ,
    \new_[55634]_ , \new_[55635]_ , \new_[55639]_ , \new_[55640]_ ,
    \new_[55643]_ , \new_[55646]_ , \new_[55647]_ , \new_[55648]_ ,
    \new_[55652]_ , \new_[55653]_ , \new_[55657]_ , \new_[55658]_ ,
    \new_[55659]_ , \new_[55663]_ , \new_[55664]_ , \new_[55667]_ ,
    \new_[55670]_ , \new_[55671]_ , \new_[55672]_ , \new_[55676]_ ,
    \new_[55677]_ , \new_[55681]_ , \new_[55682]_ , \new_[55683]_ ,
    \new_[55687]_ , \new_[55688]_ , \new_[55691]_ , \new_[55694]_ ,
    \new_[55695]_ , \new_[55696]_ , \new_[55700]_ , \new_[55701]_ ,
    \new_[55705]_ , \new_[55706]_ , \new_[55707]_ , \new_[55711]_ ,
    \new_[55712]_ , \new_[55715]_ , \new_[55718]_ , \new_[55719]_ ,
    \new_[55720]_ , \new_[55724]_ , \new_[55725]_ , \new_[55729]_ ,
    \new_[55730]_ , \new_[55731]_ , \new_[55735]_ , \new_[55736]_ ,
    \new_[55739]_ , \new_[55742]_ , \new_[55743]_ , \new_[55744]_ ,
    \new_[55748]_ , \new_[55749]_ , \new_[55753]_ , \new_[55754]_ ,
    \new_[55755]_ , \new_[55759]_ , \new_[55760]_ , \new_[55763]_ ,
    \new_[55766]_ , \new_[55767]_ , \new_[55768]_ , \new_[55772]_ ,
    \new_[55773]_ , \new_[55777]_ , \new_[55778]_ , \new_[55779]_ ,
    \new_[55783]_ , \new_[55784]_ , \new_[55787]_ , \new_[55790]_ ,
    \new_[55791]_ , \new_[55792]_ , \new_[55796]_ , \new_[55797]_ ,
    \new_[55801]_ , \new_[55802]_ , \new_[55803]_ , \new_[55807]_ ,
    \new_[55808]_ , \new_[55811]_ , \new_[55814]_ , \new_[55815]_ ,
    \new_[55816]_ , \new_[55820]_ , \new_[55821]_ , \new_[55825]_ ,
    \new_[55826]_ , \new_[55827]_ , \new_[55831]_ , \new_[55832]_ ,
    \new_[55835]_ , \new_[55838]_ , \new_[55839]_ , \new_[55840]_ ,
    \new_[55844]_ , \new_[55845]_ , \new_[55849]_ , \new_[55850]_ ,
    \new_[55851]_ , \new_[55855]_ , \new_[55856]_ , \new_[55859]_ ,
    \new_[55862]_ , \new_[55863]_ , \new_[55864]_ , \new_[55868]_ ,
    \new_[55869]_ , \new_[55873]_ , \new_[55874]_ , \new_[55875]_ ,
    \new_[55879]_ , \new_[55880]_ , \new_[55883]_ , \new_[55886]_ ,
    \new_[55887]_ , \new_[55888]_ , \new_[55892]_ , \new_[55893]_ ,
    \new_[55897]_ , \new_[55898]_ , \new_[55899]_ , \new_[55903]_ ,
    \new_[55904]_ , \new_[55907]_ , \new_[55910]_ , \new_[55911]_ ,
    \new_[55912]_ , \new_[55916]_ , \new_[55917]_ , \new_[55921]_ ,
    \new_[55922]_ , \new_[55923]_ , \new_[55927]_ , \new_[55928]_ ,
    \new_[55931]_ , \new_[55934]_ , \new_[55935]_ , \new_[55936]_ ,
    \new_[55940]_ , \new_[55941]_ , \new_[55945]_ , \new_[55946]_ ,
    \new_[55947]_ , \new_[55951]_ , \new_[55952]_ , \new_[55955]_ ,
    \new_[55958]_ , \new_[55959]_ , \new_[55960]_ , \new_[55964]_ ,
    \new_[55965]_ , \new_[55969]_ , \new_[55970]_ , \new_[55971]_ ,
    \new_[55975]_ , \new_[55976]_ , \new_[55979]_ , \new_[55982]_ ,
    \new_[55983]_ , \new_[55984]_ , \new_[55988]_ , \new_[55989]_ ,
    \new_[55993]_ , \new_[55994]_ , \new_[55995]_ , \new_[55999]_ ,
    \new_[56000]_ , \new_[56003]_ , \new_[56006]_ , \new_[56007]_ ,
    \new_[56008]_ , \new_[56012]_ , \new_[56013]_ , \new_[56017]_ ,
    \new_[56018]_ , \new_[56019]_ , \new_[56023]_ , \new_[56024]_ ,
    \new_[56027]_ , \new_[56030]_ , \new_[56031]_ , \new_[56032]_ ,
    \new_[56036]_ , \new_[56037]_ , \new_[56041]_ , \new_[56042]_ ,
    \new_[56043]_ , \new_[56047]_ , \new_[56048]_ , \new_[56051]_ ,
    \new_[56054]_ , \new_[56055]_ , \new_[56056]_ , \new_[56060]_ ,
    \new_[56061]_ , \new_[56065]_ , \new_[56066]_ , \new_[56067]_ ,
    \new_[56071]_ , \new_[56072]_ , \new_[56075]_ , \new_[56078]_ ,
    \new_[56079]_ , \new_[56080]_ , \new_[56084]_ , \new_[56085]_ ,
    \new_[56089]_ , \new_[56090]_ , \new_[56091]_ , \new_[56095]_ ,
    \new_[56096]_ , \new_[56099]_ , \new_[56102]_ , \new_[56103]_ ,
    \new_[56104]_ , \new_[56108]_ , \new_[56109]_ , \new_[56113]_ ,
    \new_[56114]_ , \new_[56115]_ , \new_[56119]_ , \new_[56120]_ ,
    \new_[56123]_ , \new_[56126]_ , \new_[56127]_ , \new_[56128]_ ,
    \new_[56132]_ , \new_[56133]_ , \new_[56137]_ , \new_[56138]_ ,
    \new_[56139]_ , \new_[56143]_ , \new_[56144]_ , \new_[56147]_ ,
    \new_[56150]_ , \new_[56151]_ , \new_[56152]_ , \new_[56156]_ ,
    \new_[56157]_ , \new_[56161]_ , \new_[56162]_ , \new_[56163]_ ,
    \new_[56167]_ , \new_[56168]_ , \new_[56171]_ , \new_[56174]_ ,
    \new_[56175]_ , \new_[56176]_ , \new_[56180]_ , \new_[56181]_ ,
    \new_[56185]_ , \new_[56186]_ , \new_[56187]_ , \new_[56191]_ ,
    \new_[56192]_ , \new_[56195]_ , \new_[56198]_ , \new_[56199]_ ,
    \new_[56200]_ , \new_[56204]_ , \new_[56205]_ , \new_[56209]_ ,
    \new_[56210]_ , \new_[56211]_ , \new_[56215]_ , \new_[56216]_ ,
    \new_[56219]_ , \new_[56222]_ , \new_[56223]_ , \new_[56224]_ ,
    \new_[56228]_ , \new_[56229]_ , \new_[56233]_ , \new_[56234]_ ,
    \new_[56235]_ , \new_[56239]_ , \new_[56240]_ , \new_[56243]_ ,
    \new_[56246]_ , \new_[56247]_ , \new_[56248]_ , \new_[56252]_ ,
    \new_[56253]_ , \new_[56257]_ , \new_[56258]_ , \new_[56259]_ ,
    \new_[56263]_ , \new_[56264]_ , \new_[56267]_ , \new_[56270]_ ,
    \new_[56271]_ , \new_[56272]_ , \new_[56276]_ , \new_[56277]_ ,
    \new_[56281]_ , \new_[56282]_ , \new_[56283]_ , \new_[56287]_ ,
    \new_[56288]_ , \new_[56291]_ , \new_[56294]_ , \new_[56295]_ ,
    \new_[56296]_ , \new_[56300]_ , \new_[56301]_ , \new_[56305]_ ,
    \new_[56306]_ , \new_[56307]_ , \new_[56311]_ , \new_[56312]_ ,
    \new_[56315]_ , \new_[56318]_ , \new_[56319]_ , \new_[56320]_ ,
    \new_[56324]_ , \new_[56325]_ , \new_[56329]_ , \new_[56330]_ ,
    \new_[56331]_ , \new_[56335]_ , \new_[56336]_ , \new_[56339]_ ,
    \new_[56342]_ , \new_[56343]_ , \new_[56344]_ , \new_[56348]_ ,
    \new_[56349]_ , \new_[56353]_ , \new_[56354]_ , \new_[56355]_ ,
    \new_[56359]_ , \new_[56360]_ , \new_[56363]_ , \new_[56366]_ ,
    \new_[56367]_ , \new_[56368]_ , \new_[56372]_ , \new_[56373]_ ,
    \new_[56377]_ , \new_[56378]_ , \new_[56379]_ , \new_[56383]_ ,
    \new_[56384]_ , \new_[56387]_ , \new_[56390]_ , \new_[56391]_ ,
    \new_[56392]_ , \new_[56396]_ , \new_[56397]_ , \new_[56401]_ ,
    \new_[56402]_ , \new_[56403]_ , \new_[56407]_ , \new_[56408]_ ,
    \new_[56411]_ , \new_[56414]_ , \new_[56415]_ , \new_[56416]_ ,
    \new_[56420]_ , \new_[56421]_ , \new_[56425]_ , \new_[56426]_ ,
    \new_[56427]_ , \new_[56431]_ , \new_[56432]_ , \new_[56435]_ ,
    \new_[56438]_ , \new_[56439]_ , \new_[56440]_ , \new_[56444]_ ,
    \new_[56445]_ , \new_[56449]_ , \new_[56450]_ , \new_[56451]_ ,
    \new_[56455]_ , \new_[56456]_ , \new_[56459]_ , \new_[56462]_ ,
    \new_[56463]_ , \new_[56464]_ , \new_[56468]_ , \new_[56469]_ ,
    \new_[56473]_ , \new_[56474]_ , \new_[56475]_ , \new_[56479]_ ,
    \new_[56480]_ , \new_[56483]_ , \new_[56486]_ , \new_[56487]_ ,
    \new_[56488]_ , \new_[56492]_ , \new_[56493]_ , \new_[56497]_ ,
    \new_[56498]_ , \new_[56499]_ , \new_[56503]_ , \new_[56504]_ ,
    \new_[56507]_ , \new_[56510]_ , \new_[56511]_ , \new_[56512]_ ,
    \new_[56516]_ , \new_[56517]_ , \new_[56521]_ , \new_[56522]_ ,
    \new_[56523]_ , \new_[56527]_ , \new_[56528]_ , \new_[56531]_ ,
    \new_[56534]_ , \new_[56535]_ , \new_[56536]_ , \new_[56540]_ ,
    \new_[56541]_ , \new_[56545]_ , \new_[56546]_ , \new_[56547]_ ,
    \new_[56551]_ , \new_[56552]_ , \new_[56555]_ , \new_[56558]_ ,
    \new_[56559]_ , \new_[56560]_ , \new_[56564]_ , \new_[56565]_ ,
    \new_[56569]_ , \new_[56570]_ , \new_[56571]_ , \new_[56575]_ ,
    \new_[56576]_ , \new_[56579]_ , \new_[56582]_ , \new_[56583]_ ,
    \new_[56584]_ , \new_[56588]_ , \new_[56589]_ , \new_[56593]_ ,
    \new_[56594]_ , \new_[56595]_ , \new_[56599]_ , \new_[56600]_ ,
    \new_[56603]_ , \new_[56606]_ , \new_[56607]_ , \new_[56608]_ ,
    \new_[56612]_ , \new_[56613]_ , \new_[56617]_ , \new_[56618]_ ,
    \new_[56619]_ , \new_[56623]_ , \new_[56624]_ , \new_[56627]_ ,
    \new_[56630]_ , \new_[56631]_ , \new_[56632]_ , \new_[56636]_ ,
    \new_[56637]_ , \new_[56641]_ , \new_[56642]_ , \new_[56643]_ ,
    \new_[56647]_ , \new_[56648]_ , \new_[56651]_ , \new_[56654]_ ,
    \new_[56655]_ , \new_[56656]_ , \new_[56660]_ , \new_[56661]_ ,
    \new_[56665]_ , \new_[56666]_ , \new_[56667]_ , \new_[56671]_ ,
    \new_[56672]_ , \new_[56675]_ , \new_[56678]_ , \new_[56679]_ ,
    \new_[56680]_ , \new_[56684]_ , \new_[56685]_ , \new_[56689]_ ,
    \new_[56690]_ , \new_[56691]_ , \new_[56695]_ , \new_[56696]_ ,
    \new_[56699]_ , \new_[56702]_ , \new_[56703]_ , \new_[56704]_ ,
    \new_[56708]_ , \new_[56709]_ , \new_[56713]_ , \new_[56714]_ ,
    \new_[56715]_ , \new_[56719]_ , \new_[56720]_ , \new_[56723]_ ,
    \new_[56726]_ , \new_[56727]_ , \new_[56728]_ , \new_[56732]_ ,
    \new_[56733]_ , \new_[56737]_ , \new_[56738]_ , \new_[56739]_ ,
    \new_[56743]_ , \new_[56744]_ , \new_[56747]_ , \new_[56750]_ ,
    \new_[56751]_ , \new_[56752]_ , \new_[56756]_ , \new_[56757]_ ,
    \new_[56760]_ , \new_[56763]_ , \new_[56764]_ , \new_[56765]_ ,
    \new_[56769]_ , \new_[56770]_ , \new_[56773]_ , \new_[56776]_ ,
    \new_[56777]_ , \new_[56778]_ , \new_[56782]_ , \new_[56783]_ ,
    \new_[56786]_ , \new_[56789]_ , \new_[56790]_ , \new_[56791]_ ,
    \new_[56795]_ , \new_[56796]_ , \new_[56799]_ , \new_[56802]_ ,
    \new_[56803]_ , \new_[56804]_ , \new_[56808]_ , \new_[56809]_ ,
    \new_[56812]_ , \new_[56815]_ , \new_[56816]_ , \new_[56817]_ ,
    \new_[56821]_ , \new_[56822]_ , \new_[56825]_ , \new_[56828]_ ,
    \new_[56829]_ , \new_[56830]_ , \new_[56834]_ , \new_[56835]_ ,
    \new_[56838]_ , \new_[56841]_ , \new_[56842]_ , \new_[56843]_ ,
    \new_[56847]_ , \new_[56848]_ , \new_[56851]_ , \new_[56854]_ ,
    \new_[56855]_ , \new_[56856]_ , \new_[56860]_ , \new_[56861]_ ,
    \new_[56864]_ , \new_[56867]_ , \new_[56868]_ , \new_[56869]_ ,
    \new_[56873]_ , \new_[56874]_ , \new_[56877]_ , \new_[56880]_ ,
    \new_[56881]_ , \new_[56882]_ , \new_[56886]_ , \new_[56887]_ ,
    \new_[56890]_ , \new_[56893]_ , \new_[56894]_ , \new_[56895]_ ,
    \new_[56899]_ , \new_[56900]_ , \new_[56903]_ , \new_[56906]_ ,
    \new_[56907]_ , \new_[56908]_ , \new_[56912]_ , \new_[56913]_ ,
    \new_[56916]_ , \new_[56919]_ , \new_[56920]_ , \new_[56921]_ ,
    \new_[56925]_ , \new_[56926]_ , \new_[56929]_ , \new_[56932]_ ,
    \new_[56933]_ , \new_[56934]_ , \new_[56938]_ , \new_[56939]_ ,
    \new_[56942]_ , \new_[56945]_ , \new_[56946]_ , \new_[56947]_ ,
    \new_[56951]_ , \new_[56952]_ , \new_[56955]_ , \new_[56958]_ ,
    \new_[56959]_ , \new_[56960]_ , \new_[56964]_ , \new_[56965]_ ,
    \new_[56968]_ , \new_[56971]_ , \new_[56972]_ , \new_[56973]_ ,
    \new_[56977]_ , \new_[56978]_ , \new_[56981]_ , \new_[56984]_ ,
    \new_[56985]_ , \new_[56986]_ , \new_[56990]_ , \new_[56991]_ ,
    \new_[56994]_ , \new_[56997]_ , \new_[56998]_ , \new_[56999]_ ,
    \new_[57003]_ , \new_[57004]_ , \new_[57007]_ , \new_[57010]_ ,
    \new_[57011]_ , \new_[57012]_ , \new_[57016]_ , \new_[57017]_ ,
    \new_[57020]_ , \new_[57023]_ , \new_[57024]_ , \new_[57025]_ ,
    \new_[57029]_ , \new_[57030]_ , \new_[57033]_ , \new_[57036]_ ,
    \new_[57037]_ , \new_[57038]_ , \new_[57042]_ , \new_[57043]_ ,
    \new_[57046]_ , \new_[57049]_ , \new_[57050]_ , \new_[57051]_ ,
    \new_[57055]_ , \new_[57056]_ , \new_[57059]_ , \new_[57062]_ ,
    \new_[57063]_ , \new_[57064]_ , \new_[57068]_ , \new_[57069]_ ,
    \new_[57072]_ , \new_[57075]_ , \new_[57076]_ , \new_[57077]_ ,
    \new_[57081]_ , \new_[57082]_ , \new_[57085]_ , \new_[57088]_ ,
    \new_[57089]_ , \new_[57090]_ , \new_[57094]_ , \new_[57095]_ ,
    \new_[57098]_ , \new_[57101]_ , \new_[57102]_ , \new_[57103]_ ,
    \new_[57107]_ , \new_[57108]_ , \new_[57111]_ , \new_[57114]_ ,
    \new_[57115]_ , \new_[57116]_ , \new_[57120]_ , \new_[57121]_ ,
    \new_[57124]_ , \new_[57127]_ , \new_[57128]_ , \new_[57129]_ ,
    \new_[57133]_ , \new_[57134]_ , \new_[57137]_ , \new_[57140]_ ,
    \new_[57141]_ , \new_[57142]_ , \new_[57146]_ , \new_[57147]_ ,
    \new_[57150]_ , \new_[57153]_ , \new_[57154]_ , \new_[57155]_ ,
    \new_[57159]_ , \new_[57160]_ , \new_[57163]_ , \new_[57166]_ ,
    \new_[57167]_ , \new_[57168]_ , \new_[57172]_ , \new_[57173]_ ,
    \new_[57176]_ , \new_[57179]_ , \new_[57180]_ , \new_[57181]_ ,
    \new_[57185]_ , \new_[57186]_ , \new_[57189]_ , \new_[57192]_ ,
    \new_[57193]_ , \new_[57194]_ , \new_[57198]_ , \new_[57199]_ ,
    \new_[57202]_ , \new_[57205]_ , \new_[57206]_ , \new_[57207]_ ,
    \new_[57211]_ , \new_[57212]_ , \new_[57215]_ , \new_[57218]_ ,
    \new_[57219]_ , \new_[57220]_ , \new_[57224]_ , \new_[57225]_ ,
    \new_[57228]_ , \new_[57231]_ , \new_[57232]_ , \new_[57233]_ ,
    \new_[57237]_ , \new_[57238]_ , \new_[57241]_ , \new_[57244]_ ,
    \new_[57245]_ , \new_[57246]_ , \new_[57250]_ , \new_[57251]_ ,
    \new_[57254]_ , \new_[57257]_ , \new_[57258]_ , \new_[57259]_ ,
    \new_[57263]_ , \new_[57264]_ , \new_[57267]_ , \new_[57270]_ ,
    \new_[57271]_ , \new_[57272]_ , \new_[57276]_ , \new_[57277]_ ,
    \new_[57280]_ , \new_[57283]_ , \new_[57284]_ , \new_[57285]_ ,
    \new_[57289]_ , \new_[57290]_ , \new_[57293]_ , \new_[57296]_ ,
    \new_[57297]_ , \new_[57298]_ , \new_[57302]_ , \new_[57303]_ ,
    \new_[57306]_ , \new_[57309]_ , \new_[57310]_ , \new_[57311]_ ,
    \new_[57315]_ , \new_[57316]_ , \new_[57319]_ , \new_[57322]_ ,
    \new_[57323]_ , \new_[57324]_ , \new_[57328]_ , \new_[57329]_ ,
    \new_[57332]_ , \new_[57335]_ , \new_[57336]_ , \new_[57337]_ ,
    \new_[57341]_ , \new_[57342]_ , \new_[57345]_ , \new_[57348]_ ,
    \new_[57349]_ , \new_[57350]_ , \new_[57354]_ , \new_[57355]_ ,
    \new_[57358]_ , \new_[57361]_ , \new_[57362]_ , \new_[57363]_ ,
    \new_[57367]_ , \new_[57368]_ , \new_[57371]_ , \new_[57374]_ ,
    \new_[57375]_ , \new_[57376]_ , \new_[57380]_ , \new_[57381]_ ,
    \new_[57384]_ , \new_[57387]_ , \new_[57388]_ , \new_[57389]_ ,
    \new_[57393]_ , \new_[57394]_ , \new_[57397]_ , \new_[57400]_ ,
    \new_[57401]_ , \new_[57402]_ , \new_[57406]_ , \new_[57407]_ ,
    \new_[57410]_ , \new_[57413]_ , \new_[57414]_ , \new_[57415]_ ,
    \new_[57419]_ , \new_[57420]_ , \new_[57423]_ , \new_[57426]_ ,
    \new_[57427]_ , \new_[57428]_ , \new_[57432]_ , \new_[57433]_ ,
    \new_[57436]_ , \new_[57439]_ , \new_[57440]_ , \new_[57441]_ ,
    \new_[57445]_ , \new_[57446]_ , \new_[57449]_ , \new_[57452]_ ,
    \new_[57453]_ , \new_[57454]_ , \new_[57458]_ , \new_[57459]_ ,
    \new_[57462]_ , \new_[57465]_ , \new_[57466]_ , \new_[57467]_ ,
    \new_[57471]_ , \new_[57472]_ , \new_[57475]_ , \new_[57478]_ ,
    \new_[57479]_ , \new_[57480]_ , \new_[57484]_ , \new_[57485]_ ,
    \new_[57488]_ , \new_[57491]_ , \new_[57492]_ , \new_[57493]_ ,
    \new_[57497]_ , \new_[57498]_ , \new_[57501]_ , \new_[57504]_ ,
    \new_[57505]_ , \new_[57506]_ , \new_[57510]_ , \new_[57511]_ ,
    \new_[57514]_ , \new_[57517]_ , \new_[57518]_ , \new_[57519]_ ,
    \new_[57523]_ , \new_[57524]_ , \new_[57527]_ , \new_[57530]_ ,
    \new_[57531]_ , \new_[57532]_ , \new_[57536]_ , \new_[57537]_ ,
    \new_[57540]_ , \new_[57543]_ , \new_[57544]_ , \new_[57545]_ ,
    \new_[57549]_ , \new_[57550]_ , \new_[57553]_ , \new_[57556]_ ,
    \new_[57557]_ , \new_[57558]_ , \new_[57562]_ , \new_[57563]_ ,
    \new_[57566]_ , \new_[57569]_ , \new_[57570]_ , \new_[57571]_ ,
    \new_[57575]_ , \new_[57576]_ , \new_[57579]_ , \new_[57582]_ ,
    \new_[57583]_ , \new_[57584]_ , \new_[57588]_ , \new_[57589]_ ,
    \new_[57592]_ , \new_[57595]_ , \new_[57596]_ , \new_[57597]_ ,
    \new_[57601]_ , \new_[57602]_ , \new_[57605]_ , \new_[57608]_ ,
    \new_[57609]_ , \new_[57610]_ , \new_[57614]_ , \new_[57615]_ ,
    \new_[57618]_ , \new_[57621]_ , \new_[57622]_ , \new_[57623]_ ,
    \new_[57627]_ , \new_[57628]_ , \new_[57631]_ , \new_[57634]_ ,
    \new_[57635]_ , \new_[57636]_ , \new_[57640]_ , \new_[57641]_ ,
    \new_[57644]_ , \new_[57647]_ , \new_[57648]_ , \new_[57649]_ ,
    \new_[57653]_ , \new_[57654]_ , \new_[57657]_ , \new_[57660]_ ,
    \new_[57661]_ , \new_[57662]_ , \new_[57666]_ , \new_[57667]_ ,
    \new_[57670]_ , \new_[57673]_ , \new_[57674]_ , \new_[57675]_ ,
    \new_[57679]_ , \new_[57680]_ , \new_[57683]_ , \new_[57686]_ ,
    \new_[57687]_ , \new_[57688]_ , \new_[57692]_ , \new_[57693]_ ,
    \new_[57696]_ , \new_[57699]_ , \new_[57700]_ , \new_[57701]_ ,
    \new_[57705]_ , \new_[57706]_ , \new_[57709]_ , \new_[57712]_ ,
    \new_[57713]_ , \new_[57714]_ , \new_[57718]_ , \new_[57719]_ ,
    \new_[57722]_ , \new_[57725]_ , \new_[57726]_ , \new_[57727]_ ,
    \new_[57731]_ , \new_[57732]_ , \new_[57735]_ , \new_[57738]_ ,
    \new_[57739]_ , \new_[57740]_ , \new_[57744]_ , \new_[57745]_ ,
    \new_[57748]_ , \new_[57751]_ , \new_[57752]_ , \new_[57753]_ ,
    \new_[57757]_ , \new_[57758]_ , \new_[57761]_ , \new_[57764]_ ,
    \new_[57765]_ , \new_[57766]_ , \new_[57770]_ , \new_[57771]_ ,
    \new_[57774]_ , \new_[57777]_ , \new_[57778]_ , \new_[57779]_ ,
    \new_[57783]_ , \new_[57784]_ , \new_[57787]_ , \new_[57790]_ ,
    \new_[57791]_ , \new_[57792]_ , \new_[57796]_ , \new_[57797]_ ,
    \new_[57800]_ , \new_[57803]_ , \new_[57804]_ , \new_[57805]_ ,
    \new_[57809]_ , \new_[57810]_ , \new_[57813]_ , \new_[57816]_ ,
    \new_[57817]_ , \new_[57818]_ , \new_[57822]_ , \new_[57823]_ ,
    \new_[57826]_ , \new_[57829]_ , \new_[57830]_ , \new_[57831]_ ,
    \new_[57835]_ , \new_[57836]_ , \new_[57839]_ , \new_[57842]_ ,
    \new_[57843]_ , \new_[57844]_ , \new_[57848]_ , \new_[57849]_ ,
    \new_[57852]_ , \new_[57855]_ , \new_[57856]_ , \new_[57857]_ ,
    \new_[57861]_ , \new_[57862]_ , \new_[57865]_ , \new_[57868]_ ,
    \new_[57869]_ , \new_[57870]_ , \new_[57874]_ , \new_[57875]_ ,
    \new_[57878]_ , \new_[57881]_ , \new_[57882]_ , \new_[57883]_ ,
    \new_[57887]_ , \new_[57888]_ , \new_[57891]_ , \new_[57894]_ ,
    \new_[57895]_ , \new_[57896]_ , \new_[57900]_ , \new_[57901]_ ,
    \new_[57904]_ , \new_[57907]_ , \new_[57908]_ , \new_[57909]_ ,
    \new_[57913]_ , \new_[57914]_ , \new_[57917]_ , \new_[57920]_ ,
    \new_[57921]_ , \new_[57922]_ , \new_[57926]_ , \new_[57927]_ ,
    \new_[57930]_ , \new_[57933]_ , \new_[57934]_ , \new_[57935]_ ,
    \new_[57939]_ , \new_[57940]_ , \new_[57943]_ , \new_[57946]_ ,
    \new_[57947]_ , \new_[57948]_ , \new_[57952]_ , \new_[57953]_ ,
    \new_[57956]_ , \new_[57959]_ , \new_[57960]_ , \new_[57961]_ ,
    \new_[57965]_ , \new_[57966]_ , \new_[57969]_ , \new_[57972]_ ,
    \new_[57973]_ , \new_[57974]_ , \new_[57978]_ , \new_[57979]_ ,
    \new_[57982]_ , \new_[57985]_ , \new_[57986]_ , \new_[57987]_ ,
    \new_[57991]_ , \new_[57992]_ , \new_[57995]_ , \new_[57998]_ ,
    \new_[57999]_ , \new_[58000]_ , \new_[58004]_ , \new_[58005]_ ,
    \new_[58008]_ , \new_[58011]_ , \new_[58012]_ , \new_[58013]_ ,
    \new_[58017]_ , \new_[58018]_ , \new_[58021]_ , \new_[58024]_ ,
    \new_[58025]_ , \new_[58026]_ , \new_[58030]_ , \new_[58031]_ ,
    \new_[58034]_ , \new_[58037]_ , \new_[58038]_ , \new_[58039]_ ,
    \new_[58043]_ , \new_[58044]_ , \new_[58047]_ , \new_[58050]_ ,
    \new_[58051]_ , \new_[58052]_ , \new_[58056]_ , \new_[58057]_ ,
    \new_[58060]_ , \new_[58063]_ , \new_[58064]_ , \new_[58065]_ ,
    \new_[58069]_ , \new_[58070]_ , \new_[58073]_ , \new_[58076]_ ,
    \new_[58077]_ , \new_[58078]_ , \new_[58082]_ , \new_[58083]_ ,
    \new_[58086]_ , \new_[58089]_ , \new_[58090]_ , \new_[58091]_ ,
    \new_[58095]_ , \new_[58096]_ , \new_[58099]_ , \new_[58102]_ ,
    \new_[58103]_ , \new_[58104]_ , \new_[58108]_ , \new_[58109]_ ,
    \new_[58112]_ , \new_[58115]_ , \new_[58116]_ , \new_[58117]_ ,
    \new_[58121]_ , \new_[58122]_ , \new_[58125]_ , \new_[58128]_ ,
    \new_[58129]_ , \new_[58130]_ , \new_[58134]_ , \new_[58135]_ ,
    \new_[58138]_ , \new_[58141]_ , \new_[58142]_ , \new_[58143]_ ,
    \new_[58147]_ , \new_[58148]_ , \new_[58151]_ , \new_[58154]_ ,
    \new_[58155]_ , \new_[58156]_ , \new_[58160]_ , \new_[58161]_ ,
    \new_[58164]_ , \new_[58167]_ , \new_[58168]_ , \new_[58169]_ ,
    \new_[58173]_ , \new_[58174]_ , \new_[58177]_ , \new_[58180]_ ,
    \new_[58181]_ , \new_[58182]_ , \new_[58186]_ , \new_[58187]_ ,
    \new_[58190]_ , \new_[58193]_ , \new_[58194]_ , \new_[58195]_ ,
    \new_[58199]_ , \new_[58200]_ , \new_[58203]_ , \new_[58206]_ ,
    \new_[58207]_ , \new_[58208]_ , \new_[58212]_ , \new_[58213]_ ,
    \new_[58216]_ , \new_[58219]_ , \new_[58220]_ , \new_[58221]_ ,
    \new_[58225]_ , \new_[58226]_ , \new_[58229]_ , \new_[58232]_ ,
    \new_[58233]_ , \new_[58234]_ , \new_[58238]_ , \new_[58239]_ ,
    \new_[58242]_ , \new_[58245]_ , \new_[58246]_ , \new_[58247]_ ,
    \new_[58251]_ , \new_[58252]_ , \new_[58255]_ , \new_[58258]_ ,
    \new_[58259]_ , \new_[58260]_ , \new_[58264]_ , \new_[58265]_ ,
    \new_[58268]_ , \new_[58271]_ , \new_[58272]_ , \new_[58273]_ ,
    \new_[58277]_ , \new_[58278]_ , \new_[58281]_ , \new_[58284]_ ,
    \new_[58285]_ , \new_[58286]_ , \new_[58290]_ , \new_[58291]_ ,
    \new_[58294]_ , \new_[58297]_ , \new_[58298]_ , \new_[58299]_ ,
    \new_[58303]_ , \new_[58304]_ , \new_[58307]_ , \new_[58310]_ ,
    \new_[58311]_ , \new_[58312]_ , \new_[58316]_ , \new_[58317]_ ,
    \new_[58320]_ , \new_[58323]_ , \new_[58324]_ , \new_[58325]_ ,
    \new_[58329]_ , \new_[58330]_ , \new_[58333]_ , \new_[58336]_ ,
    \new_[58337]_ , \new_[58338]_ , \new_[58342]_ , \new_[58343]_ ,
    \new_[58346]_ , \new_[58349]_ , \new_[58350]_ , \new_[58351]_ ,
    \new_[58355]_ , \new_[58356]_ , \new_[58359]_ , \new_[58362]_ ,
    \new_[58363]_ , \new_[58364]_ , \new_[58368]_ , \new_[58369]_ ,
    \new_[58372]_ , \new_[58375]_ , \new_[58376]_ , \new_[58377]_ ,
    \new_[58381]_ , \new_[58382]_ , \new_[58385]_ , \new_[58388]_ ,
    \new_[58389]_ , \new_[58390]_ , \new_[58394]_ , \new_[58395]_ ,
    \new_[58398]_ , \new_[58401]_ , \new_[58402]_ , \new_[58403]_ ,
    \new_[58407]_ , \new_[58408]_ , \new_[58411]_ , \new_[58414]_ ,
    \new_[58415]_ , \new_[58416]_ , \new_[58420]_ , \new_[58421]_ ,
    \new_[58424]_ , \new_[58427]_ , \new_[58428]_ , \new_[58429]_ ,
    \new_[58433]_ , \new_[58434]_ , \new_[58437]_ , \new_[58440]_ ,
    \new_[58441]_ , \new_[58442]_ , \new_[58446]_ , \new_[58447]_ ,
    \new_[58450]_ , \new_[58453]_ , \new_[58454]_ , \new_[58455]_ ,
    \new_[58459]_ , \new_[58460]_ , \new_[58463]_ , \new_[58466]_ ,
    \new_[58467]_ , \new_[58468]_ , \new_[58472]_ , \new_[58473]_ ,
    \new_[58476]_ , \new_[58479]_ , \new_[58480]_ , \new_[58481]_ ,
    \new_[58485]_ , \new_[58486]_ , \new_[58489]_ , \new_[58492]_ ,
    \new_[58493]_ , \new_[58494]_ , \new_[58498]_ , \new_[58499]_ ,
    \new_[58502]_ , \new_[58505]_ , \new_[58506]_ , \new_[58507]_ ,
    \new_[58511]_ , \new_[58512]_ , \new_[58515]_ , \new_[58518]_ ,
    \new_[58519]_ , \new_[58520]_ , \new_[58524]_ , \new_[58525]_ ,
    \new_[58528]_ , \new_[58531]_ , \new_[58532]_ , \new_[58533]_ ,
    \new_[58537]_ , \new_[58538]_ , \new_[58541]_ , \new_[58544]_ ,
    \new_[58545]_ , \new_[58546]_ , \new_[58550]_ , \new_[58551]_ ,
    \new_[58554]_ , \new_[58557]_ , \new_[58558]_ , \new_[58559]_ ,
    \new_[58563]_ , \new_[58564]_ , \new_[58567]_ , \new_[58570]_ ,
    \new_[58571]_ , \new_[58572]_ , \new_[58576]_ , \new_[58577]_ ,
    \new_[58580]_ , \new_[58583]_ , \new_[58584]_ , \new_[58585]_ ,
    \new_[58589]_ , \new_[58590]_ , \new_[58593]_ , \new_[58596]_ ,
    \new_[58597]_ , \new_[58598]_ , \new_[58602]_ , \new_[58603]_ ,
    \new_[58606]_ , \new_[58609]_ , \new_[58610]_ , \new_[58611]_ ,
    \new_[58615]_ , \new_[58616]_ , \new_[58619]_ , \new_[58622]_ ,
    \new_[58623]_ , \new_[58624]_ , \new_[58628]_ , \new_[58629]_ ,
    \new_[58632]_ , \new_[58635]_ , \new_[58636]_ , \new_[58637]_ ,
    \new_[58641]_ , \new_[58642]_ , \new_[58645]_ , \new_[58648]_ ,
    \new_[58649]_ , \new_[58650]_ , \new_[58654]_ , \new_[58655]_ ,
    \new_[58658]_ , \new_[58661]_ , \new_[58662]_ , \new_[58663]_ ,
    \new_[58667]_ , \new_[58668]_ , \new_[58671]_ , \new_[58674]_ ,
    \new_[58675]_ , \new_[58676]_ , \new_[58680]_ , \new_[58681]_ ,
    \new_[58684]_ , \new_[58687]_ , \new_[58688]_ , \new_[58689]_ ,
    \new_[58693]_ , \new_[58694]_ , \new_[58697]_ , \new_[58700]_ ,
    \new_[58701]_ , \new_[58702]_ , \new_[58706]_ , \new_[58707]_ ,
    \new_[58710]_ , \new_[58713]_ , \new_[58714]_ , \new_[58715]_ ,
    \new_[58719]_ , \new_[58720]_ , \new_[58723]_ , \new_[58726]_ ,
    \new_[58727]_ , \new_[58728]_ , \new_[58732]_ , \new_[58733]_ ,
    \new_[58736]_ , \new_[58739]_ , \new_[58740]_ , \new_[58741]_ ,
    \new_[58745]_ , \new_[58746]_ , \new_[58749]_ , \new_[58752]_ ,
    \new_[58753]_ , \new_[58754]_ , \new_[58758]_ , \new_[58759]_ ,
    \new_[58762]_ , \new_[58765]_ , \new_[58766]_ , \new_[58767]_ ,
    \new_[58771]_ , \new_[58772]_ , \new_[58775]_ , \new_[58778]_ ,
    \new_[58779]_ , \new_[58780]_ , \new_[58784]_ , \new_[58785]_ ,
    \new_[58788]_ , \new_[58791]_ , \new_[58792]_ , \new_[58793]_ ,
    \new_[58797]_ , \new_[58798]_ , \new_[58801]_ , \new_[58804]_ ,
    \new_[58805]_ , \new_[58806]_ , \new_[58810]_ , \new_[58811]_ ,
    \new_[58814]_ , \new_[58817]_ , \new_[58818]_ , \new_[58819]_ ,
    \new_[58823]_ , \new_[58824]_ , \new_[58827]_ , \new_[58830]_ ,
    \new_[58831]_ , \new_[58832]_ , \new_[58836]_ , \new_[58837]_ ,
    \new_[58840]_ , \new_[58843]_ , \new_[58844]_ , \new_[58845]_ ,
    \new_[58849]_ , \new_[58850]_ , \new_[58853]_ , \new_[58856]_ ,
    \new_[58857]_ , \new_[58858]_ , \new_[58862]_ , \new_[58863]_ ,
    \new_[58866]_ , \new_[58869]_ , \new_[58870]_ , \new_[58871]_ ,
    \new_[58875]_ , \new_[58876]_ , \new_[58879]_ , \new_[58882]_ ,
    \new_[58883]_ , \new_[58884]_ , \new_[58888]_ , \new_[58889]_ ,
    \new_[58892]_ , \new_[58895]_ , \new_[58896]_ , \new_[58897]_ ,
    \new_[58901]_ , \new_[58902]_ , \new_[58905]_ , \new_[58908]_ ,
    \new_[58909]_ , \new_[58910]_ , \new_[58914]_ , \new_[58915]_ ,
    \new_[58918]_ , \new_[58921]_ , \new_[58922]_ , \new_[58923]_ ,
    \new_[58927]_ , \new_[58928]_ , \new_[58931]_ , \new_[58934]_ ,
    \new_[58935]_ , \new_[58936]_ , \new_[58940]_ , \new_[58941]_ ,
    \new_[58944]_ , \new_[58947]_ , \new_[58948]_ , \new_[58949]_ ,
    \new_[58953]_ , \new_[58954]_ , \new_[58957]_ , \new_[58960]_ ,
    \new_[58961]_ , \new_[58962]_ , \new_[58966]_ , \new_[58967]_ ,
    \new_[58970]_ , \new_[58973]_ , \new_[58974]_ , \new_[58975]_ ,
    \new_[58979]_ , \new_[58980]_ , \new_[58983]_ , \new_[58986]_ ,
    \new_[58987]_ , \new_[58988]_ , \new_[58992]_ , \new_[58993]_ ,
    \new_[58996]_ , \new_[58999]_ , \new_[59000]_ , \new_[59001]_ ,
    \new_[59005]_ , \new_[59006]_ , \new_[59009]_ , \new_[59012]_ ,
    \new_[59013]_ , \new_[59014]_ , \new_[59018]_ , \new_[59019]_ ,
    \new_[59022]_ , \new_[59025]_ , \new_[59026]_ , \new_[59027]_ ,
    \new_[59031]_ , \new_[59032]_ , \new_[59035]_ , \new_[59038]_ ,
    \new_[59039]_ , \new_[59040]_ , \new_[59044]_ , \new_[59045]_ ,
    \new_[59048]_ , \new_[59051]_ , \new_[59052]_ , \new_[59053]_ ,
    \new_[59057]_ , \new_[59058]_ , \new_[59061]_ , \new_[59064]_ ,
    \new_[59065]_ , \new_[59066]_ , \new_[59070]_ , \new_[59071]_ ,
    \new_[59074]_ , \new_[59077]_ , \new_[59078]_ , \new_[59079]_ ,
    \new_[59083]_ , \new_[59084]_ , \new_[59087]_ , \new_[59090]_ ,
    \new_[59091]_ , \new_[59092]_ , \new_[59096]_ , \new_[59097]_ ,
    \new_[59100]_ , \new_[59103]_ , \new_[59104]_ , \new_[59105]_ ,
    \new_[59109]_ , \new_[59110]_ , \new_[59113]_ , \new_[59116]_ ,
    \new_[59117]_ , \new_[59118]_ , \new_[59122]_ , \new_[59123]_ ,
    \new_[59126]_ , \new_[59129]_ , \new_[59130]_ , \new_[59131]_ ,
    \new_[59135]_ , \new_[59136]_ , \new_[59139]_ , \new_[59142]_ ,
    \new_[59143]_ , \new_[59144]_ , \new_[59148]_ , \new_[59149]_ ,
    \new_[59152]_ , \new_[59155]_ , \new_[59156]_ , \new_[59157]_ ,
    \new_[59161]_ , \new_[59162]_ , \new_[59165]_ , \new_[59168]_ ,
    \new_[59169]_ , \new_[59170]_ , \new_[59174]_ , \new_[59175]_ ,
    \new_[59178]_ , \new_[59181]_ , \new_[59182]_ , \new_[59183]_ ,
    \new_[59187]_ , \new_[59188]_ , \new_[59191]_ , \new_[59194]_ ,
    \new_[59195]_ , \new_[59196]_ , \new_[59200]_ , \new_[59201]_ ,
    \new_[59204]_ , \new_[59207]_ , \new_[59208]_ , \new_[59209]_ ,
    \new_[59213]_ , \new_[59214]_ , \new_[59217]_ , \new_[59220]_ ,
    \new_[59221]_ , \new_[59222]_ , \new_[59226]_ , \new_[59227]_ ,
    \new_[59230]_ , \new_[59233]_ , \new_[59234]_ , \new_[59235]_ ,
    \new_[59239]_ , \new_[59240]_ , \new_[59243]_ , \new_[59246]_ ,
    \new_[59247]_ , \new_[59248]_ , \new_[59252]_ , \new_[59253]_ ,
    \new_[59256]_ , \new_[59259]_ , \new_[59260]_ , \new_[59261]_ ,
    \new_[59265]_ , \new_[59266]_ , \new_[59269]_ , \new_[59272]_ ,
    \new_[59273]_ , \new_[59274]_ , \new_[59278]_ , \new_[59279]_ ,
    \new_[59282]_ , \new_[59285]_ , \new_[59286]_ , \new_[59287]_ ,
    \new_[59291]_ , \new_[59292]_ , \new_[59295]_ , \new_[59298]_ ,
    \new_[59299]_ , \new_[59300]_ , \new_[59304]_ , \new_[59305]_ ,
    \new_[59308]_ , \new_[59311]_ , \new_[59312]_ , \new_[59313]_ ,
    \new_[59317]_ , \new_[59318]_ , \new_[59321]_ , \new_[59324]_ ,
    \new_[59325]_ , \new_[59326]_ , \new_[59330]_ , \new_[59331]_ ,
    \new_[59334]_ , \new_[59337]_ , \new_[59338]_ , \new_[59339]_ ,
    \new_[59343]_ , \new_[59344]_ , \new_[59347]_ , \new_[59350]_ ,
    \new_[59351]_ , \new_[59352]_ , \new_[59356]_ , \new_[59357]_ ,
    \new_[59360]_ , \new_[59363]_ , \new_[59364]_ , \new_[59365]_ ,
    \new_[59369]_ , \new_[59370]_ , \new_[59373]_ , \new_[59376]_ ,
    \new_[59377]_ , \new_[59378]_ , \new_[59382]_ , \new_[59383]_ ,
    \new_[59386]_ , \new_[59389]_ , \new_[59390]_ , \new_[59391]_ ,
    \new_[59395]_ , \new_[59396]_ , \new_[59399]_ , \new_[59402]_ ,
    \new_[59403]_ , \new_[59404]_ , \new_[59408]_ , \new_[59409]_ ,
    \new_[59412]_ , \new_[59415]_ , \new_[59416]_ , \new_[59417]_ ,
    \new_[59421]_ , \new_[59422]_ , \new_[59425]_ , \new_[59428]_ ,
    \new_[59429]_ , \new_[59430]_ , \new_[59434]_ , \new_[59435]_ ,
    \new_[59438]_ , \new_[59441]_ , \new_[59442]_ , \new_[59443]_ ,
    \new_[59447]_ , \new_[59448]_ , \new_[59451]_ , \new_[59454]_ ,
    \new_[59455]_ , \new_[59456]_ , \new_[59460]_ , \new_[59461]_ ,
    \new_[59464]_ , \new_[59467]_ , \new_[59468]_ , \new_[59469]_ ,
    \new_[59473]_ , \new_[59474]_ , \new_[59477]_ , \new_[59480]_ ,
    \new_[59481]_ , \new_[59482]_ , \new_[59486]_ , \new_[59487]_ ,
    \new_[59490]_ , \new_[59493]_ , \new_[59494]_ , \new_[59495]_ ,
    \new_[59499]_ , \new_[59500]_ , \new_[59503]_ , \new_[59506]_ ,
    \new_[59507]_ , \new_[59508]_ , \new_[59512]_ , \new_[59513]_ ,
    \new_[59516]_ , \new_[59519]_ , \new_[59520]_ , \new_[59521]_ ,
    \new_[59525]_ , \new_[59526]_ , \new_[59529]_ , \new_[59532]_ ,
    \new_[59533]_ , \new_[59534]_ , \new_[59538]_ , \new_[59539]_ ,
    \new_[59542]_ , \new_[59545]_ , \new_[59546]_ , \new_[59547]_ ,
    \new_[59551]_ , \new_[59552]_ , \new_[59555]_ , \new_[59558]_ ,
    \new_[59559]_ , \new_[59560]_ , \new_[59564]_ , \new_[59565]_ ,
    \new_[59568]_ , \new_[59571]_ , \new_[59572]_ , \new_[59573]_ ,
    \new_[59577]_ , \new_[59578]_ , \new_[59581]_ , \new_[59584]_ ,
    \new_[59585]_ , \new_[59586]_ , \new_[59590]_ , \new_[59591]_ ,
    \new_[59594]_ , \new_[59597]_ , \new_[59598]_ , \new_[59599]_ ,
    \new_[59603]_ , \new_[59604]_ , \new_[59607]_ , \new_[59610]_ ,
    \new_[59611]_ , \new_[59612]_ , \new_[59616]_ , \new_[59617]_ ,
    \new_[59620]_ , \new_[59623]_ , \new_[59624]_ , \new_[59625]_ ,
    \new_[59629]_ , \new_[59630]_ , \new_[59633]_ , \new_[59636]_ ,
    \new_[59637]_ , \new_[59638]_ , \new_[59642]_ , \new_[59643]_ ,
    \new_[59646]_ , \new_[59649]_ , \new_[59650]_ , \new_[59651]_ ,
    \new_[59655]_ , \new_[59656]_ , \new_[59659]_ , \new_[59662]_ ,
    \new_[59663]_ , \new_[59664]_ , \new_[59668]_ , \new_[59669]_ ,
    \new_[59672]_ , \new_[59675]_ , \new_[59676]_ , \new_[59677]_ ,
    \new_[59681]_ , \new_[59682]_ , \new_[59685]_ , \new_[59688]_ ,
    \new_[59689]_ , \new_[59690]_ , \new_[59694]_ , \new_[59695]_ ,
    \new_[59698]_ , \new_[59701]_ , \new_[59702]_ , \new_[59703]_ ,
    \new_[59707]_ , \new_[59708]_ , \new_[59711]_ , \new_[59714]_ ,
    \new_[59715]_ , \new_[59716]_ , \new_[59720]_ , \new_[59721]_ ,
    \new_[59724]_ , \new_[59727]_ , \new_[59728]_ , \new_[59729]_ ,
    \new_[59733]_ , \new_[59734]_ , \new_[59737]_ , \new_[59740]_ ,
    \new_[59741]_ , \new_[59742]_ , \new_[59746]_ , \new_[59747]_ ,
    \new_[59750]_ , \new_[59753]_ , \new_[59754]_ , \new_[59755]_ ,
    \new_[59759]_ , \new_[59760]_ , \new_[59763]_ , \new_[59766]_ ,
    \new_[59767]_ , \new_[59768]_ , \new_[59772]_ , \new_[59773]_ ,
    \new_[59776]_ , \new_[59779]_ , \new_[59780]_ , \new_[59781]_ ,
    \new_[59785]_ , \new_[59786]_ , \new_[59789]_ , \new_[59792]_ ,
    \new_[59793]_ , \new_[59794]_ , \new_[59798]_ , \new_[59799]_ ,
    \new_[59802]_ , \new_[59805]_ , \new_[59806]_ , \new_[59807]_ ,
    \new_[59811]_ , \new_[59812]_ , \new_[59815]_ , \new_[59818]_ ,
    \new_[59819]_ , \new_[59820]_ , \new_[59824]_ , \new_[59825]_ ,
    \new_[59828]_ , \new_[59831]_ , \new_[59832]_ , \new_[59833]_ ,
    \new_[59837]_ , \new_[59838]_ , \new_[59841]_ , \new_[59844]_ ,
    \new_[59845]_ , \new_[59846]_ , \new_[59850]_ , \new_[59851]_ ,
    \new_[59854]_ , \new_[59857]_ , \new_[59858]_ , \new_[59859]_ ,
    \new_[59863]_ , \new_[59864]_ , \new_[59867]_ , \new_[59870]_ ,
    \new_[59871]_ , \new_[59872]_ , \new_[59876]_ , \new_[59877]_ ,
    \new_[59880]_ , \new_[59883]_ , \new_[59884]_ , \new_[59885]_ ,
    \new_[59889]_ , \new_[59890]_ , \new_[59893]_ , \new_[59896]_ ,
    \new_[59897]_ , \new_[59898]_ , \new_[59902]_ , \new_[59903]_ ,
    \new_[59906]_ , \new_[59909]_ , \new_[59910]_ , \new_[59911]_ ,
    \new_[59915]_ , \new_[59916]_ , \new_[59919]_ , \new_[59922]_ ,
    \new_[59923]_ , \new_[59924]_ , \new_[59928]_ , \new_[59929]_ ,
    \new_[59932]_ , \new_[59935]_ , \new_[59936]_ , \new_[59937]_ ,
    \new_[59941]_ , \new_[59942]_ , \new_[59945]_ , \new_[59948]_ ,
    \new_[59949]_ , \new_[59950]_ , \new_[59954]_ , \new_[59955]_ ,
    \new_[59958]_ , \new_[59961]_ , \new_[59962]_ , \new_[59963]_ ,
    \new_[59967]_ , \new_[59968]_ , \new_[59971]_ , \new_[59974]_ ,
    \new_[59975]_ , \new_[59976]_ , \new_[59980]_ , \new_[59981]_ ,
    \new_[59984]_ , \new_[59987]_ , \new_[59988]_ , \new_[59989]_ ,
    \new_[59993]_ , \new_[59994]_ , \new_[59997]_ , \new_[60000]_ ,
    \new_[60001]_ , \new_[60002]_ , \new_[60006]_ , \new_[60007]_ ,
    \new_[60010]_ , \new_[60013]_ , \new_[60014]_ , \new_[60015]_ ,
    \new_[60019]_ , \new_[60020]_ , \new_[60023]_ , \new_[60026]_ ,
    \new_[60027]_ , \new_[60028]_ , \new_[60032]_ , \new_[60033]_ ,
    \new_[60036]_ , \new_[60039]_ , \new_[60040]_ , \new_[60041]_ ,
    \new_[60045]_ , \new_[60046]_ , \new_[60049]_ , \new_[60052]_ ,
    \new_[60053]_ , \new_[60054]_ , \new_[60058]_ , \new_[60059]_ ,
    \new_[60062]_ , \new_[60065]_ , \new_[60066]_ , \new_[60067]_ ,
    \new_[60071]_ , \new_[60072]_ , \new_[60075]_ , \new_[60078]_ ,
    \new_[60079]_ , \new_[60080]_ , \new_[60084]_ , \new_[60085]_ ,
    \new_[60088]_ , \new_[60091]_ , \new_[60092]_ , \new_[60093]_ ,
    \new_[60097]_ , \new_[60098]_ , \new_[60101]_ , \new_[60104]_ ,
    \new_[60105]_ , \new_[60106]_ , \new_[60110]_ , \new_[60111]_ ,
    \new_[60114]_ , \new_[60117]_ , \new_[60118]_ , \new_[60119]_ ,
    \new_[60123]_ , \new_[60124]_ , \new_[60127]_ , \new_[60130]_ ,
    \new_[60131]_ , \new_[60132]_ , \new_[60136]_ , \new_[60137]_ ,
    \new_[60140]_ , \new_[60143]_ , \new_[60144]_ , \new_[60145]_ ,
    \new_[60149]_ , \new_[60150]_ , \new_[60153]_ , \new_[60156]_ ,
    \new_[60157]_ , \new_[60158]_ , \new_[60162]_ , \new_[60163]_ ,
    \new_[60166]_ , \new_[60169]_ , \new_[60170]_ , \new_[60171]_ ,
    \new_[60175]_ , \new_[60176]_ , \new_[60179]_ , \new_[60182]_ ,
    \new_[60183]_ , \new_[60184]_ , \new_[60188]_ , \new_[60189]_ ,
    \new_[60192]_ , \new_[60195]_ , \new_[60196]_ , \new_[60197]_ ,
    \new_[60201]_ , \new_[60202]_ , \new_[60205]_ , \new_[60208]_ ,
    \new_[60209]_ , \new_[60210]_ , \new_[60214]_ , \new_[60215]_ ,
    \new_[60218]_ , \new_[60221]_ , \new_[60222]_ , \new_[60223]_ ,
    \new_[60227]_ , \new_[60228]_ , \new_[60231]_ , \new_[60234]_ ,
    \new_[60235]_ , \new_[60236]_ , \new_[60240]_ , \new_[60241]_ ,
    \new_[60244]_ , \new_[60247]_ , \new_[60248]_ , \new_[60249]_ ,
    \new_[60253]_ , \new_[60254]_ , \new_[60257]_ , \new_[60260]_ ,
    \new_[60261]_ , \new_[60262]_ , \new_[60266]_ , \new_[60267]_ ,
    \new_[60270]_ , \new_[60273]_ , \new_[60274]_ , \new_[60275]_ ,
    \new_[60279]_ , \new_[60280]_ , \new_[60283]_ , \new_[60286]_ ,
    \new_[60287]_ , \new_[60288]_ , \new_[60292]_ , \new_[60293]_ ,
    \new_[60296]_ , \new_[60299]_ , \new_[60300]_ , \new_[60301]_ ,
    \new_[60305]_ , \new_[60306]_ , \new_[60309]_ , \new_[60312]_ ,
    \new_[60313]_ , \new_[60314]_ , \new_[60318]_ , \new_[60319]_ ,
    \new_[60322]_ , \new_[60325]_ , \new_[60326]_ , \new_[60327]_ ,
    \new_[60331]_ , \new_[60332]_ , \new_[60335]_ , \new_[60338]_ ,
    \new_[60339]_ , \new_[60340]_ , \new_[60344]_ , \new_[60345]_ ,
    \new_[60348]_ , \new_[60351]_ , \new_[60352]_ , \new_[60353]_ ,
    \new_[60357]_ , \new_[60358]_ , \new_[60361]_ , \new_[60364]_ ,
    \new_[60365]_ , \new_[60366]_ , \new_[60370]_ , \new_[60371]_ ,
    \new_[60374]_ , \new_[60377]_ , \new_[60378]_ , \new_[60379]_ ,
    \new_[60383]_ , \new_[60384]_ , \new_[60387]_ , \new_[60390]_ ,
    \new_[60391]_ , \new_[60392]_ , \new_[60396]_ , \new_[60397]_ ,
    \new_[60400]_ , \new_[60403]_ , \new_[60404]_ , \new_[60405]_ ,
    \new_[60409]_ , \new_[60410]_ , \new_[60413]_ , \new_[60416]_ ,
    \new_[60417]_ , \new_[60418]_ , \new_[60422]_ , \new_[60423]_ ,
    \new_[60426]_ , \new_[60429]_ , \new_[60430]_ , \new_[60431]_ ,
    \new_[60435]_ , \new_[60436]_ , \new_[60439]_ , \new_[60442]_ ,
    \new_[60443]_ , \new_[60444]_ , \new_[60448]_ , \new_[60449]_ ,
    \new_[60452]_ , \new_[60455]_ , \new_[60456]_ , \new_[60457]_ ,
    \new_[60461]_ , \new_[60462]_ , \new_[60465]_ , \new_[60468]_ ,
    \new_[60469]_ , \new_[60470]_ , \new_[60474]_ , \new_[60475]_ ,
    \new_[60478]_ , \new_[60481]_ , \new_[60482]_ , \new_[60483]_ ,
    \new_[60487]_ , \new_[60488]_ , \new_[60491]_ , \new_[60494]_ ,
    \new_[60495]_ , \new_[60496]_ , \new_[60500]_ , \new_[60501]_ ,
    \new_[60504]_ , \new_[60507]_ , \new_[60508]_ , \new_[60509]_ ,
    \new_[60513]_ , \new_[60514]_ , \new_[60517]_ , \new_[60520]_ ,
    \new_[60521]_ , \new_[60522]_ , \new_[60526]_ , \new_[60527]_ ,
    \new_[60530]_ , \new_[60533]_ , \new_[60534]_ , \new_[60535]_ ,
    \new_[60539]_ , \new_[60540]_ , \new_[60543]_ , \new_[60546]_ ,
    \new_[60547]_ , \new_[60548]_ , \new_[60552]_ , \new_[60553]_ ,
    \new_[60556]_ , \new_[60559]_ , \new_[60560]_ , \new_[60561]_ ,
    \new_[60565]_ , \new_[60566]_ , \new_[60569]_ , \new_[60572]_ ,
    \new_[60573]_ , \new_[60574]_ , \new_[60578]_ , \new_[60579]_ ,
    \new_[60582]_ , \new_[60585]_ , \new_[60586]_ , \new_[60587]_ ,
    \new_[60591]_ , \new_[60592]_ , \new_[60595]_ , \new_[60598]_ ,
    \new_[60599]_ , \new_[60600]_ , \new_[60604]_ , \new_[60605]_ ,
    \new_[60608]_ , \new_[60611]_ , \new_[60612]_ , \new_[60613]_ ,
    \new_[60617]_ , \new_[60618]_ , \new_[60621]_ , \new_[60624]_ ,
    \new_[60625]_ , \new_[60626]_ , \new_[60630]_ , \new_[60631]_ ,
    \new_[60634]_ , \new_[60637]_ , \new_[60638]_ , \new_[60639]_ ,
    \new_[60643]_ , \new_[60644]_ , \new_[60647]_ , \new_[60650]_ ,
    \new_[60651]_ , \new_[60652]_ , \new_[60656]_ , \new_[60657]_ ,
    \new_[60660]_ , \new_[60663]_ , \new_[60664]_ , \new_[60665]_ ,
    \new_[60669]_ , \new_[60670]_ , \new_[60673]_ , \new_[60676]_ ,
    \new_[60677]_ , \new_[60678]_ , \new_[60682]_ , \new_[60683]_ ,
    \new_[60686]_ , \new_[60689]_ , \new_[60690]_ , \new_[60691]_ ,
    \new_[60695]_ , \new_[60696]_ , \new_[60699]_ , \new_[60702]_ ,
    \new_[60703]_ , \new_[60704]_ , \new_[60708]_ , \new_[60709]_ ,
    \new_[60712]_ , \new_[60715]_ , \new_[60716]_ , \new_[60717]_ ,
    \new_[60721]_ , \new_[60722]_ , \new_[60725]_ , \new_[60728]_ ,
    \new_[60729]_ , \new_[60730]_ , \new_[60734]_ , \new_[60735]_ ,
    \new_[60738]_ , \new_[60741]_ , \new_[60742]_ , \new_[60743]_ ,
    \new_[60747]_ , \new_[60748]_ , \new_[60751]_ , \new_[60754]_ ,
    \new_[60755]_ , \new_[60756]_ , \new_[60760]_ , \new_[60761]_ ,
    \new_[60764]_ , \new_[60767]_ , \new_[60768]_ , \new_[60769]_ ,
    \new_[60773]_ , \new_[60774]_ , \new_[60777]_ , \new_[60780]_ ,
    \new_[60781]_ , \new_[60782]_ , \new_[60786]_ , \new_[60787]_ ,
    \new_[60790]_ , \new_[60793]_ , \new_[60794]_ , \new_[60795]_ ,
    \new_[60799]_ , \new_[60800]_ , \new_[60803]_ , \new_[60806]_ ,
    \new_[60807]_ , \new_[60808]_ , \new_[60812]_ , \new_[60813]_ ,
    \new_[60816]_ , \new_[60819]_ , \new_[60820]_ , \new_[60821]_ ,
    \new_[60825]_ , \new_[60826]_ , \new_[60829]_ , \new_[60832]_ ,
    \new_[60833]_ , \new_[60834]_ , \new_[60838]_ , \new_[60839]_ ,
    \new_[60842]_ , \new_[60845]_ , \new_[60846]_ , \new_[60847]_ ,
    \new_[60851]_ , \new_[60852]_ , \new_[60855]_ , \new_[60858]_ ,
    \new_[60859]_ , \new_[60860]_ , \new_[60864]_ , \new_[60865]_ ,
    \new_[60868]_ , \new_[60871]_ , \new_[60872]_ , \new_[60873]_ ,
    \new_[60877]_ , \new_[60878]_ , \new_[60881]_ , \new_[60884]_ ,
    \new_[60885]_ , \new_[60886]_ , \new_[60890]_ , \new_[60891]_ ,
    \new_[60894]_ , \new_[60897]_ , \new_[60898]_ , \new_[60899]_ ,
    \new_[60903]_ , \new_[60904]_ , \new_[60907]_ , \new_[60910]_ ,
    \new_[60911]_ , \new_[60912]_ , \new_[60916]_ , \new_[60917]_ ,
    \new_[60920]_ , \new_[60923]_ , \new_[60924]_ , \new_[60925]_ ,
    \new_[60929]_ , \new_[60930]_ , \new_[60933]_ , \new_[60936]_ ,
    \new_[60937]_ , \new_[60938]_ , \new_[60942]_ , \new_[60943]_ ,
    \new_[60946]_ , \new_[60949]_ , \new_[60950]_ , \new_[60951]_ ,
    \new_[60955]_ , \new_[60956]_ , \new_[60959]_ , \new_[60962]_ ,
    \new_[60963]_ , \new_[60964]_ , \new_[60968]_ , \new_[60969]_ ,
    \new_[60972]_ , \new_[60975]_ , \new_[60976]_ , \new_[60977]_ ,
    \new_[60981]_ , \new_[60982]_ , \new_[60985]_ , \new_[60988]_ ,
    \new_[60989]_ , \new_[60990]_ , \new_[60994]_ , \new_[60995]_ ,
    \new_[60998]_ , \new_[61001]_ , \new_[61002]_ , \new_[61003]_ ,
    \new_[61007]_ , \new_[61008]_ , \new_[61011]_ , \new_[61014]_ ,
    \new_[61015]_ , \new_[61016]_ , \new_[61020]_ , \new_[61021]_ ,
    \new_[61024]_ , \new_[61027]_ , \new_[61028]_ , \new_[61029]_ ,
    \new_[61033]_ , \new_[61034]_ , \new_[61037]_ , \new_[61040]_ ,
    \new_[61041]_ , \new_[61042]_ , \new_[61046]_ , \new_[61047]_ ,
    \new_[61050]_ , \new_[61053]_ , \new_[61054]_ , \new_[61055]_ ,
    \new_[61059]_ , \new_[61060]_ , \new_[61063]_ , \new_[61066]_ ,
    \new_[61067]_ , \new_[61068]_ , \new_[61072]_ , \new_[61073]_ ,
    \new_[61076]_ , \new_[61079]_ , \new_[61080]_ , \new_[61081]_ ,
    \new_[61085]_ , \new_[61086]_ , \new_[61089]_ , \new_[61092]_ ,
    \new_[61093]_ , \new_[61094]_ , \new_[61098]_ , \new_[61099]_ ,
    \new_[61102]_ , \new_[61105]_ , \new_[61106]_ , \new_[61107]_ ,
    \new_[61111]_ , \new_[61112]_ , \new_[61115]_ , \new_[61118]_ ,
    \new_[61119]_ , \new_[61120]_ , \new_[61124]_ , \new_[61125]_ ,
    \new_[61128]_ , \new_[61131]_ , \new_[61132]_ , \new_[61133]_ ,
    \new_[61137]_ , \new_[61138]_ , \new_[61141]_ , \new_[61144]_ ,
    \new_[61145]_ , \new_[61146]_ , \new_[61150]_ , \new_[61151]_ ,
    \new_[61154]_ , \new_[61157]_ , \new_[61158]_ , \new_[61159]_ ,
    \new_[61163]_ , \new_[61164]_ , \new_[61167]_ , \new_[61170]_ ,
    \new_[61171]_ , \new_[61172]_ , \new_[61176]_ , \new_[61177]_ ,
    \new_[61180]_ , \new_[61183]_ , \new_[61184]_ , \new_[61185]_ ,
    \new_[61189]_ , \new_[61190]_ , \new_[61193]_ , \new_[61196]_ ,
    \new_[61197]_ , \new_[61198]_ , \new_[61202]_ , \new_[61203]_ ,
    \new_[61206]_ , \new_[61209]_ , \new_[61210]_ , \new_[61211]_ ,
    \new_[61215]_ , \new_[61216]_ , \new_[61219]_ , \new_[61222]_ ,
    \new_[61223]_ , \new_[61224]_ , \new_[61228]_ , \new_[61229]_ ,
    \new_[61232]_ , \new_[61235]_ , \new_[61236]_ , \new_[61237]_ ,
    \new_[61241]_ , \new_[61242]_ , \new_[61245]_ , \new_[61248]_ ,
    \new_[61249]_ , \new_[61250]_ , \new_[61254]_ , \new_[61255]_ ,
    \new_[61258]_ , \new_[61261]_ , \new_[61262]_ , \new_[61263]_ ,
    \new_[61267]_ , \new_[61268]_ , \new_[61271]_ , \new_[61274]_ ,
    \new_[61275]_ , \new_[61276]_ , \new_[61280]_ , \new_[61281]_ ,
    \new_[61284]_ , \new_[61287]_ , \new_[61288]_ , \new_[61289]_ ,
    \new_[61293]_ , \new_[61294]_ , \new_[61297]_ , \new_[61300]_ ,
    \new_[61301]_ , \new_[61302]_ , \new_[61306]_ , \new_[61307]_ ,
    \new_[61310]_ , \new_[61313]_ , \new_[61314]_ , \new_[61315]_ ,
    \new_[61319]_ , \new_[61320]_ , \new_[61323]_ , \new_[61326]_ ,
    \new_[61327]_ , \new_[61328]_ , \new_[61332]_ , \new_[61333]_ ,
    \new_[61336]_ , \new_[61339]_ , \new_[61340]_ , \new_[61341]_ ,
    \new_[61345]_ , \new_[61346]_ , \new_[61349]_ , \new_[61352]_ ,
    \new_[61353]_ , \new_[61354]_ , \new_[61358]_ , \new_[61359]_ ,
    \new_[61362]_ , \new_[61365]_ , \new_[61366]_ , \new_[61367]_ ,
    \new_[61371]_ , \new_[61372]_ , \new_[61375]_ , \new_[61378]_ ,
    \new_[61379]_ , \new_[61380]_ , \new_[61384]_ , \new_[61385]_ ,
    \new_[61388]_ , \new_[61391]_ , \new_[61392]_ , \new_[61393]_ ,
    \new_[61397]_ , \new_[61398]_ , \new_[61401]_ , \new_[61404]_ ,
    \new_[61405]_ , \new_[61406]_ , \new_[61410]_ , \new_[61411]_ ,
    \new_[61414]_ , \new_[61417]_ , \new_[61418]_ , \new_[61419]_ ,
    \new_[61423]_ , \new_[61424]_ , \new_[61427]_ , \new_[61430]_ ,
    \new_[61431]_ , \new_[61432]_ , \new_[61436]_ , \new_[61437]_ ,
    \new_[61440]_ , \new_[61443]_ , \new_[61444]_ , \new_[61445]_ ,
    \new_[61449]_ , \new_[61450]_ , \new_[61453]_ , \new_[61456]_ ,
    \new_[61457]_ , \new_[61458]_ , \new_[61462]_ , \new_[61463]_ ,
    \new_[61466]_ , \new_[61469]_ , \new_[61470]_ , \new_[61471]_ ,
    \new_[61475]_ , \new_[61476]_ , \new_[61479]_ , \new_[61482]_ ,
    \new_[61483]_ , \new_[61484]_ , \new_[61488]_ , \new_[61489]_ ,
    \new_[61492]_ , \new_[61495]_ , \new_[61496]_ , \new_[61497]_ ,
    \new_[61501]_ , \new_[61502]_ , \new_[61505]_ , \new_[61508]_ ,
    \new_[61509]_ , \new_[61510]_ , \new_[61514]_ , \new_[61515]_ ,
    \new_[61518]_ , \new_[61521]_ , \new_[61522]_ , \new_[61523]_ ,
    \new_[61527]_ , \new_[61528]_ , \new_[61531]_ , \new_[61534]_ ,
    \new_[61535]_ , \new_[61536]_ , \new_[61540]_ , \new_[61541]_ ,
    \new_[61544]_ , \new_[61547]_ , \new_[61548]_ , \new_[61549]_ ,
    \new_[61553]_ , \new_[61554]_ , \new_[61557]_ , \new_[61560]_ ,
    \new_[61561]_ , \new_[61562]_ , \new_[61566]_ , \new_[61567]_ ,
    \new_[61570]_ , \new_[61573]_ , \new_[61574]_ , \new_[61575]_ ,
    \new_[61579]_ , \new_[61580]_ , \new_[61583]_ , \new_[61586]_ ,
    \new_[61587]_ , \new_[61588]_ , \new_[61592]_ , \new_[61593]_ ,
    \new_[61596]_ , \new_[61599]_ , \new_[61600]_ , \new_[61601]_ ,
    \new_[61605]_ , \new_[61606]_ , \new_[61609]_ , \new_[61612]_ ,
    \new_[61613]_ , \new_[61614]_ , \new_[61618]_ , \new_[61619]_ ,
    \new_[61622]_ , \new_[61625]_ , \new_[61626]_ , \new_[61627]_ ,
    \new_[61631]_ , \new_[61632]_ , \new_[61635]_ , \new_[61638]_ ,
    \new_[61639]_ , \new_[61640]_ , \new_[61644]_ , \new_[61645]_ ,
    \new_[61648]_ , \new_[61651]_ , \new_[61652]_ , \new_[61653]_ ,
    \new_[61657]_ , \new_[61658]_ , \new_[61661]_ , \new_[61664]_ ,
    \new_[61665]_ , \new_[61666]_ , \new_[61670]_ , \new_[61671]_ ,
    \new_[61674]_ , \new_[61677]_ , \new_[61678]_ , \new_[61679]_ ,
    \new_[61683]_ , \new_[61684]_ , \new_[61687]_ , \new_[61690]_ ,
    \new_[61691]_ , \new_[61692]_ , \new_[61696]_ , \new_[61697]_ ,
    \new_[61700]_ , \new_[61703]_ , \new_[61704]_ , \new_[61705]_ ,
    \new_[61709]_ , \new_[61710]_ , \new_[61713]_ , \new_[61716]_ ,
    \new_[61717]_ , \new_[61718]_ , \new_[61722]_ , \new_[61723]_ ,
    \new_[61726]_ , \new_[61729]_ , \new_[61730]_ , \new_[61731]_ ,
    \new_[61735]_ , \new_[61736]_ , \new_[61739]_ , \new_[61742]_ ,
    \new_[61743]_ , \new_[61744]_ , \new_[61748]_ , \new_[61749]_ ,
    \new_[61752]_ , \new_[61755]_ , \new_[61756]_ , \new_[61757]_ ,
    \new_[61761]_ , \new_[61762]_ , \new_[61765]_ , \new_[61768]_ ,
    \new_[61769]_ , \new_[61770]_ , \new_[61774]_ , \new_[61775]_ ,
    \new_[61778]_ , \new_[61781]_ , \new_[61782]_ , \new_[61783]_ ,
    \new_[61787]_ , \new_[61788]_ , \new_[61791]_ , \new_[61794]_ ,
    \new_[61795]_ , \new_[61796]_ , \new_[61800]_ , \new_[61801]_ ,
    \new_[61804]_ , \new_[61807]_ , \new_[61808]_ , \new_[61809]_ ,
    \new_[61813]_ , \new_[61814]_ , \new_[61817]_ , \new_[61820]_ ,
    \new_[61821]_ , \new_[61822]_ , \new_[61826]_ , \new_[61827]_ ,
    \new_[61830]_ , \new_[61833]_ , \new_[61834]_ , \new_[61835]_ ,
    \new_[61839]_ , \new_[61840]_ , \new_[61843]_ , \new_[61846]_ ,
    \new_[61847]_ , \new_[61848]_ , \new_[61852]_ , \new_[61853]_ ,
    \new_[61856]_ , \new_[61859]_ , \new_[61860]_ , \new_[61861]_ ,
    \new_[61865]_ , \new_[61866]_ , \new_[61869]_ , \new_[61872]_ ,
    \new_[61873]_ , \new_[61874]_ , \new_[61878]_ , \new_[61879]_ ,
    \new_[61882]_ , \new_[61885]_ , \new_[61886]_ , \new_[61887]_ ,
    \new_[61891]_ , \new_[61892]_ , \new_[61895]_ , \new_[61898]_ ,
    \new_[61899]_ , \new_[61900]_ , \new_[61904]_ , \new_[61905]_ ,
    \new_[61908]_ , \new_[61911]_ , \new_[61912]_ , \new_[61913]_ ,
    \new_[61917]_ , \new_[61918]_ , \new_[61921]_ , \new_[61924]_ ,
    \new_[61925]_ , \new_[61926]_ , \new_[61930]_ , \new_[61931]_ ,
    \new_[61934]_ , \new_[61937]_ , \new_[61938]_ , \new_[61939]_ ,
    \new_[61943]_ , \new_[61944]_ , \new_[61947]_ , \new_[61950]_ ,
    \new_[61951]_ , \new_[61952]_ , \new_[61956]_ , \new_[61957]_ ,
    \new_[61960]_ , \new_[61963]_ , \new_[61964]_ , \new_[61965]_ ,
    \new_[61969]_ , \new_[61970]_ , \new_[61973]_ , \new_[61976]_ ,
    \new_[61977]_ , \new_[61978]_ , \new_[61982]_ , \new_[61983]_ ,
    \new_[61986]_ , \new_[61989]_ , \new_[61990]_ , \new_[61991]_ ,
    \new_[61995]_ , \new_[61996]_ , \new_[61999]_ , \new_[62002]_ ,
    \new_[62003]_ , \new_[62004]_ , \new_[62008]_ , \new_[62009]_ ,
    \new_[62012]_ , \new_[62015]_ , \new_[62016]_ , \new_[62017]_ ,
    \new_[62021]_ , \new_[62022]_ , \new_[62025]_ , \new_[62028]_ ,
    \new_[62029]_ , \new_[62030]_ , \new_[62034]_ , \new_[62035]_ ,
    \new_[62038]_ , \new_[62041]_ , \new_[62042]_ , \new_[62043]_ ,
    \new_[62047]_ , \new_[62048]_ , \new_[62051]_ , \new_[62054]_ ,
    \new_[62055]_ , \new_[62056]_ , \new_[62060]_ , \new_[62061]_ ,
    \new_[62064]_ , \new_[62067]_ , \new_[62068]_ , \new_[62069]_ ,
    \new_[62073]_ , \new_[62074]_ , \new_[62077]_ , \new_[62080]_ ,
    \new_[62081]_ , \new_[62082]_ , \new_[62086]_ , \new_[62087]_ ,
    \new_[62090]_ , \new_[62093]_ , \new_[62094]_ , \new_[62095]_ ,
    \new_[62099]_ , \new_[62100]_ , \new_[62103]_ , \new_[62106]_ ,
    \new_[62107]_ , \new_[62108]_ , \new_[62112]_ , \new_[62113]_ ,
    \new_[62116]_ , \new_[62119]_ , \new_[62120]_ , \new_[62121]_ ,
    \new_[62125]_ , \new_[62126]_ , \new_[62129]_ , \new_[62132]_ ,
    \new_[62133]_ , \new_[62134]_ , \new_[62138]_ , \new_[62139]_ ,
    \new_[62142]_ , \new_[62145]_ , \new_[62146]_ , \new_[62147]_ ,
    \new_[62151]_ , \new_[62152]_ , \new_[62155]_ , \new_[62158]_ ,
    \new_[62159]_ , \new_[62160]_ , \new_[62164]_ , \new_[62165]_ ,
    \new_[62168]_ , \new_[62171]_ , \new_[62172]_ , \new_[62173]_ ,
    \new_[62177]_ , \new_[62178]_ , \new_[62181]_ , \new_[62184]_ ,
    \new_[62185]_ , \new_[62186]_ , \new_[62190]_ , \new_[62191]_ ,
    \new_[62194]_ , \new_[62197]_ , \new_[62198]_ , \new_[62199]_ ,
    \new_[62203]_ , \new_[62204]_ , \new_[62207]_ , \new_[62210]_ ,
    \new_[62211]_ , \new_[62212]_ , \new_[62216]_ , \new_[62217]_ ,
    \new_[62220]_ , \new_[62223]_ , \new_[62224]_ , \new_[62225]_ ,
    \new_[62229]_ , \new_[62230]_ , \new_[62233]_ , \new_[62236]_ ,
    \new_[62237]_ , \new_[62238]_ , \new_[62242]_ , \new_[62243]_ ,
    \new_[62246]_ , \new_[62249]_ , \new_[62250]_ , \new_[62251]_ ,
    \new_[62255]_ , \new_[62256]_ , \new_[62259]_ , \new_[62262]_ ,
    \new_[62263]_ , \new_[62264]_ , \new_[62268]_ , \new_[62269]_ ,
    \new_[62272]_ , \new_[62275]_ , \new_[62276]_ , \new_[62277]_ ,
    \new_[62281]_ , \new_[62282]_ , \new_[62285]_ , \new_[62288]_ ,
    \new_[62289]_ , \new_[62290]_ , \new_[62294]_ , \new_[62295]_ ,
    \new_[62298]_ , \new_[62301]_ , \new_[62302]_ , \new_[62303]_ ,
    \new_[62307]_ , \new_[62308]_ , \new_[62311]_ , \new_[62314]_ ,
    \new_[62315]_ , \new_[62316]_ , \new_[62320]_ , \new_[62321]_ ,
    \new_[62324]_ , \new_[62327]_ , \new_[62328]_ , \new_[62329]_ ,
    \new_[62333]_ , \new_[62334]_ , \new_[62337]_ , \new_[62340]_ ,
    \new_[62341]_ , \new_[62342]_ , \new_[62346]_ , \new_[62347]_ ,
    \new_[62350]_ , \new_[62353]_ , \new_[62354]_ , \new_[62355]_ ,
    \new_[62359]_ , \new_[62360]_ , \new_[62363]_ , \new_[62366]_ ,
    \new_[62367]_ , \new_[62368]_ , \new_[62372]_ , \new_[62373]_ ,
    \new_[62376]_ , \new_[62379]_ , \new_[62380]_ , \new_[62381]_ ,
    \new_[62385]_ , \new_[62386]_ , \new_[62389]_ , \new_[62392]_ ,
    \new_[62393]_ , \new_[62394]_ , \new_[62398]_ , \new_[62399]_ ,
    \new_[62402]_ , \new_[62405]_ , \new_[62406]_ , \new_[62407]_ ,
    \new_[62411]_ , \new_[62412]_ , \new_[62415]_ , \new_[62418]_ ,
    \new_[62419]_ , \new_[62420]_ , \new_[62424]_ , \new_[62425]_ ,
    \new_[62428]_ , \new_[62431]_ , \new_[62432]_ , \new_[62433]_ ,
    \new_[62437]_ , \new_[62438]_ , \new_[62441]_ , \new_[62444]_ ,
    \new_[62445]_ , \new_[62446]_ , \new_[62450]_ , \new_[62451]_ ,
    \new_[62454]_ , \new_[62457]_ , \new_[62458]_ , \new_[62459]_ ,
    \new_[62463]_ , \new_[62464]_ , \new_[62467]_ , \new_[62470]_ ,
    \new_[62471]_ , \new_[62472]_ , \new_[62476]_ , \new_[62477]_ ,
    \new_[62480]_ , \new_[62483]_ , \new_[62484]_ , \new_[62485]_ ,
    \new_[62489]_ , \new_[62490]_ , \new_[62493]_ , \new_[62496]_ ,
    \new_[62497]_ , \new_[62498]_ , \new_[62502]_ , \new_[62503]_ ,
    \new_[62506]_ , \new_[62509]_ , \new_[62510]_ , \new_[62511]_ ,
    \new_[62515]_ , \new_[62516]_ , \new_[62519]_ , \new_[62522]_ ,
    \new_[62523]_ , \new_[62524]_ , \new_[62528]_ , \new_[62529]_ ,
    \new_[62532]_ , \new_[62535]_ , \new_[62536]_ , \new_[62537]_ ,
    \new_[62541]_ , \new_[62542]_ , \new_[62545]_ , \new_[62548]_ ,
    \new_[62549]_ , \new_[62550]_ , \new_[62554]_ , \new_[62555]_ ,
    \new_[62558]_ , \new_[62561]_ , \new_[62562]_ , \new_[62563]_ ,
    \new_[62567]_ , \new_[62568]_ , \new_[62571]_ , \new_[62574]_ ,
    \new_[62575]_ , \new_[62576]_ , \new_[62580]_ , \new_[62581]_ ,
    \new_[62584]_ , \new_[62587]_ , \new_[62588]_ , \new_[62589]_ ,
    \new_[62593]_ , \new_[62594]_ , \new_[62597]_ , \new_[62600]_ ,
    \new_[62601]_ , \new_[62602]_ , \new_[62606]_ , \new_[62607]_ ,
    \new_[62610]_ , \new_[62613]_ , \new_[62614]_ , \new_[62615]_ ,
    \new_[62619]_ , \new_[62620]_ , \new_[62623]_ , \new_[62626]_ ,
    \new_[62627]_ , \new_[62628]_ , \new_[62632]_ , \new_[62633]_ ,
    \new_[62636]_ , \new_[62639]_ , \new_[62640]_ , \new_[62641]_ ,
    \new_[62645]_ , \new_[62646]_ , \new_[62649]_ , \new_[62652]_ ,
    \new_[62653]_ , \new_[62654]_ , \new_[62658]_ , \new_[62659]_ ,
    \new_[62662]_ , \new_[62665]_ , \new_[62666]_ , \new_[62667]_ ,
    \new_[62671]_ , \new_[62672]_ , \new_[62675]_ , \new_[62678]_ ,
    \new_[62679]_ , \new_[62680]_ , \new_[62684]_ , \new_[62685]_ ,
    \new_[62688]_ , \new_[62691]_ , \new_[62692]_ , \new_[62693]_ ,
    \new_[62697]_ , \new_[62698]_ , \new_[62701]_ , \new_[62704]_ ,
    \new_[62705]_ , \new_[62706]_ , \new_[62710]_ , \new_[62711]_ ,
    \new_[62714]_ , \new_[62717]_ , \new_[62718]_ , \new_[62719]_ ,
    \new_[62723]_ , \new_[62724]_ , \new_[62727]_ , \new_[62730]_ ,
    \new_[62731]_ , \new_[62732]_ , \new_[62736]_ , \new_[62737]_ ,
    \new_[62740]_ , \new_[62743]_ , \new_[62744]_ , \new_[62745]_ ,
    \new_[62749]_ , \new_[62750]_ , \new_[62753]_ , \new_[62756]_ ,
    \new_[62757]_ , \new_[62758]_ , \new_[62762]_ , \new_[62763]_ ,
    \new_[62766]_ , \new_[62769]_ , \new_[62770]_ , \new_[62771]_ ,
    \new_[62775]_ , \new_[62776]_ , \new_[62779]_ , \new_[62782]_ ,
    \new_[62783]_ , \new_[62784]_ , \new_[62788]_ , \new_[62789]_ ,
    \new_[62792]_ , \new_[62795]_ , \new_[62796]_ , \new_[62797]_ ,
    \new_[62801]_ , \new_[62802]_ , \new_[62805]_ , \new_[62808]_ ,
    \new_[62809]_ , \new_[62810]_ , \new_[62814]_ , \new_[62815]_ ,
    \new_[62818]_ , \new_[62821]_ , \new_[62822]_ , \new_[62823]_ ,
    \new_[62827]_ , \new_[62828]_ , \new_[62831]_ , \new_[62834]_ ,
    \new_[62835]_ , \new_[62836]_ , \new_[62840]_ , \new_[62841]_ ,
    \new_[62844]_ , \new_[62847]_ , \new_[62848]_ , \new_[62849]_ ,
    \new_[62853]_ , \new_[62854]_ , \new_[62857]_ , \new_[62860]_ ,
    \new_[62861]_ , \new_[62862]_ , \new_[62866]_ , \new_[62867]_ ,
    \new_[62870]_ , \new_[62873]_ , \new_[62874]_ , \new_[62875]_ ,
    \new_[62879]_ , \new_[62880]_ , \new_[62883]_ , \new_[62886]_ ,
    \new_[62887]_ , \new_[62888]_ , \new_[62892]_ , \new_[62893]_ ,
    \new_[62896]_ , \new_[62899]_ , \new_[62900]_ , \new_[62901]_ ,
    \new_[62905]_ , \new_[62906]_ , \new_[62909]_ , \new_[62912]_ ,
    \new_[62913]_ , \new_[62914]_ , \new_[62918]_ , \new_[62919]_ ,
    \new_[62922]_ , \new_[62925]_ , \new_[62926]_ , \new_[62927]_ ,
    \new_[62931]_ , \new_[62932]_ , \new_[62935]_ , \new_[62938]_ ,
    \new_[62939]_ , \new_[62940]_ , \new_[62944]_ , \new_[62945]_ ,
    \new_[62948]_ , \new_[62951]_ , \new_[62952]_ , \new_[62953]_ ,
    \new_[62957]_ , \new_[62958]_ , \new_[62961]_ , \new_[62964]_ ,
    \new_[62965]_ , \new_[62966]_ , \new_[62970]_ , \new_[62971]_ ,
    \new_[62974]_ , \new_[62977]_ , \new_[62978]_ , \new_[62979]_ ,
    \new_[62983]_ , \new_[62984]_ , \new_[62987]_ , \new_[62990]_ ,
    \new_[62991]_ , \new_[62992]_ , \new_[62996]_ , \new_[62997]_ ,
    \new_[63000]_ , \new_[63003]_ , \new_[63004]_ , \new_[63005]_ ,
    \new_[63009]_ , \new_[63010]_ , \new_[63013]_ , \new_[63016]_ ,
    \new_[63017]_ , \new_[63018]_ , \new_[63022]_ , \new_[63023]_ ,
    \new_[63026]_ , \new_[63029]_ , \new_[63030]_ , \new_[63031]_ ,
    \new_[63035]_ , \new_[63036]_ , \new_[63039]_ , \new_[63042]_ ,
    \new_[63043]_ , \new_[63044]_ , \new_[63048]_ , \new_[63049]_ ,
    \new_[63052]_ , \new_[63055]_ , \new_[63056]_ , \new_[63057]_ ,
    \new_[63061]_ , \new_[63062]_ , \new_[63065]_ , \new_[63068]_ ,
    \new_[63069]_ , \new_[63070]_ , \new_[63074]_ , \new_[63075]_ ,
    \new_[63078]_ , \new_[63081]_ , \new_[63082]_ , \new_[63083]_ ,
    \new_[63087]_ , \new_[63088]_ , \new_[63091]_ , \new_[63094]_ ,
    \new_[63095]_ , \new_[63096]_ , \new_[63100]_ , \new_[63101]_ ,
    \new_[63104]_ , \new_[63107]_ , \new_[63108]_ , \new_[63109]_ ,
    \new_[63113]_ , \new_[63114]_ , \new_[63117]_ , \new_[63120]_ ,
    \new_[63121]_ , \new_[63122]_ , \new_[63126]_ , \new_[63127]_ ,
    \new_[63130]_ , \new_[63133]_ , \new_[63134]_ , \new_[63135]_ ,
    \new_[63139]_ , \new_[63140]_ , \new_[63143]_ , \new_[63146]_ ,
    \new_[63147]_ , \new_[63148]_ , \new_[63152]_ , \new_[63153]_ ,
    \new_[63156]_ , \new_[63159]_ , \new_[63160]_ , \new_[63161]_ ,
    \new_[63165]_ , \new_[63166]_ , \new_[63169]_ , \new_[63172]_ ,
    \new_[63173]_ , \new_[63174]_ , \new_[63178]_ , \new_[63179]_ ,
    \new_[63182]_ , \new_[63185]_ , \new_[63186]_ , \new_[63187]_ ,
    \new_[63191]_ , \new_[63192]_ , \new_[63195]_ , \new_[63198]_ ,
    \new_[63199]_ , \new_[63200]_ , \new_[63204]_ , \new_[63205]_ ,
    \new_[63208]_ , \new_[63211]_ , \new_[63212]_ , \new_[63213]_ ,
    \new_[63217]_ , \new_[63218]_ , \new_[63221]_ , \new_[63224]_ ,
    \new_[63225]_ , \new_[63226]_ , \new_[63230]_ , \new_[63231]_ ,
    \new_[63234]_ , \new_[63237]_ , \new_[63238]_ , \new_[63239]_ ,
    \new_[63243]_ , \new_[63244]_ , \new_[63247]_ , \new_[63250]_ ,
    \new_[63251]_ , \new_[63252]_ , \new_[63256]_ , \new_[63257]_ ,
    \new_[63260]_ , \new_[63263]_ , \new_[63264]_ , \new_[63265]_ ,
    \new_[63269]_ , \new_[63270]_ , \new_[63273]_ , \new_[63276]_ ,
    \new_[63277]_ , \new_[63278]_ , \new_[63282]_ , \new_[63283]_ ,
    \new_[63286]_ , \new_[63289]_ , \new_[63290]_ , \new_[63291]_ ,
    \new_[63295]_ , \new_[63296]_ , \new_[63299]_ , \new_[63302]_ ,
    \new_[63303]_ , \new_[63304]_ , \new_[63308]_ , \new_[63309]_ ,
    \new_[63312]_ , \new_[63315]_ , \new_[63316]_ , \new_[63317]_ ,
    \new_[63321]_ , \new_[63322]_ , \new_[63325]_ , \new_[63328]_ ,
    \new_[63329]_ , \new_[63330]_ , \new_[63334]_ , \new_[63335]_ ,
    \new_[63338]_ , \new_[63341]_ , \new_[63342]_ , \new_[63343]_ ,
    \new_[63347]_ , \new_[63348]_ , \new_[63351]_ , \new_[63354]_ ,
    \new_[63355]_ , \new_[63356]_ , \new_[63360]_ , \new_[63361]_ ,
    \new_[63364]_ , \new_[63367]_ , \new_[63368]_ , \new_[63369]_ ,
    \new_[63373]_ , \new_[63374]_ , \new_[63377]_ , \new_[63380]_ ,
    \new_[63381]_ , \new_[63382]_ , \new_[63386]_ , \new_[63387]_ ,
    \new_[63390]_ , \new_[63393]_ , \new_[63394]_ , \new_[63395]_ ,
    \new_[63399]_ , \new_[63400]_ , \new_[63403]_ , \new_[63406]_ ,
    \new_[63407]_ , \new_[63408]_ , \new_[63412]_ , \new_[63413]_ ,
    \new_[63416]_ , \new_[63419]_ , \new_[63420]_ , \new_[63421]_ ,
    \new_[63425]_ , \new_[63426]_ , \new_[63429]_ , \new_[63432]_ ,
    \new_[63433]_ , \new_[63434]_ , \new_[63438]_ , \new_[63439]_ ,
    \new_[63442]_ , \new_[63445]_ , \new_[63446]_ , \new_[63447]_ ,
    \new_[63451]_ , \new_[63452]_ , \new_[63455]_ , \new_[63458]_ ,
    \new_[63459]_ , \new_[63460]_ , \new_[63464]_ , \new_[63465]_ ,
    \new_[63468]_ , \new_[63471]_ , \new_[63472]_ , \new_[63473]_ ,
    \new_[63477]_ , \new_[63478]_ , \new_[63481]_ , \new_[63484]_ ,
    \new_[63485]_ , \new_[63486]_ , \new_[63490]_ , \new_[63491]_ ,
    \new_[63494]_ , \new_[63497]_ , \new_[63498]_ , \new_[63499]_ ,
    \new_[63503]_ , \new_[63504]_ , \new_[63507]_ , \new_[63510]_ ,
    \new_[63511]_ , \new_[63512]_ , \new_[63516]_ , \new_[63517]_ ,
    \new_[63520]_ , \new_[63523]_ , \new_[63524]_ , \new_[63525]_ ,
    \new_[63529]_ , \new_[63530]_ , \new_[63533]_ , \new_[63536]_ ,
    \new_[63537]_ , \new_[63538]_ , \new_[63542]_ , \new_[63543]_ ,
    \new_[63546]_ , \new_[63549]_ , \new_[63550]_ , \new_[63551]_ ,
    \new_[63555]_ , \new_[63556]_ , \new_[63559]_ , \new_[63562]_ ,
    \new_[63563]_ , \new_[63564]_ , \new_[63568]_ , \new_[63569]_ ,
    \new_[63572]_ , \new_[63575]_ , \new_[63576]_ , \new_[63577]_ ,
    \new_[63581]_ , \new_[63582]_ , \new_[63585]_ , \new_[63588]_ ,
    \new_[63589]_ , \new_[63590]_ , \new_[63594]_ , \new_[63595]_ ,
    \new_[63598]_ , \new_[63601]_ , \new_[63602]_ , \new_[63603]_ ,
    \new_[63607]_ , \new_[63608]_ , \new_[63611]_ , \new_[63614]_ ,
    \new_[63615]_ , \new_[63616]_ , \new_[63620]_ , \new_[63621]_ ,
    \new_[63624]_ , \new_[63627]_ , \new_[63628]_ , \new_[63629]_ ,
    \new_[63633]_ , \new_[63634]_ , \new_[63637]_ , \new_[63640]_ ,
    \new_[63641]_ , \new_[63642]_ , \new_[63646]_ , \new_[63647]_ ,
    \new_[63650]_ , \new_[63653]_ , \new_[63654]_ , \new_[63655]_ ,
    \new_[63659]_ , \new_[63660]_ , \new_[63663]_ , \new_[63666]_ ,
    \new_[63667]_ , \new_[63668]_ , \new_[63672]_ , \new_[63673]_ ,
    \new_[63676]_ , \new_[63679]_ , \new_[63680]_ , \new_[63681]_ ,
    \new_[63685]_ , \new_[63686]_ , \new_[63689]_ , \new_[63692]_ ,
    \new_[63693]_ , \new_[63694]_ , \new_[63698]_ , \new_[63699]_ ,
    \new_[63702]_ , \new_[63705]_ , \new_[63706]_ , \new_[63707]_ ,
    \new_[63711]_ , \new_[63712]_ , \new_[63715]_ , \new_[63718]_ ,
    \new_[63719]_ , \new_[63720]_ , \new_[63724]_ , \new_[63725]_ ,
    \new_[63728]_ , \new_[63731]_ , \new_[63732]_ , \new_[63733]_ ,
    \new_[63737]_ , \new_[63738]_ , \new_[63741]_ , \new_[63744]_ ,
    \new_[63745]_ , \new_[63746]_ , \new_[63750]_ , \new_[63751]_ ,
    \new_[63754]_ , \new_[63757]_ , \new_[63758]_ , \new_[63759]_ ,
    \new_[63763]_ , \new_[63764]_ , \new_[63767]_ , \new_[63770]_ ,
    \new_[63771]_ , \new_[63772]_ , \new_[63776]_ , \new_[63777]_ ,
    \new_[63780]_ , \new_[63783]_ , \new_[63784]_ , \new_[63785]_ ,
    \new_[63789]_ , \new_[63790]_ , \new_[63793]_ , \new_[63796]_ ,
    \new_[63797]_ , \new_[63798]_ , \new_[63802]_ , \new_[63803]_ ,
    \new_[63806]_ , \new_[63809]_ , \new_[63810]_ , \new_[63811]_ ,
    \new_[63815]_ , \new_[63816]_ , \new_[63819]_ , \new_[63822]_ ,
    \new_[63823]_ , \new_[63824]_ , \new_[63828]_ , \new_[63829]_ ,
    \new_[63832]_ , \new_[63835]_ , \new_[63836]_ , \new_[63837]_ ,
    \new_[63841]_ , \new_[63842]_ , \new_[63845]_ , \new_[63848]_ ,
    \new_[63849]_ , \new_[63850]_ , \new_[63854]_ , \new_[63855]_ ,
    \new_[63858]_ , \new_[63861]_ , \new_[63862]_ , \new_[63863]_ ,
    \new_[63867]_ , \new_[63868]_ , \new_[63871]_ , \new_[63874]_ ,
    \new_[63875]_ , \new_[63876]_ , \new_[63880]_ , \new_[63881]_ ,
    \new_[63884]_ , \new_[63887]_ , \new_[63888]_ , \new_[63889]_ ,
    \new_[63893]_ , \new_[63894]_ , \new_[63897]_ , \new_[63900]_ ,
    \new_[63901]_ , \new_[63902]_ , \new_[63906]_ , \new_[63907]_ ,
    \new_[63910]_ , \new_[63913]_ , \new_[63914]_ , \new_[63915]_ ,
    \new_[63919]_ , \new_[63920]_ , \new_[63923]_ , \new_[63926]_ ,
    \new_[63927]_ , \new_[63928]_ , \new_[63932]_ , \new_[63933]_ ,
    \new_[63936]_ , \new_[63939]_ , \new_[63940]_ , \new_[63941]_ ,
    \new_[63945]_ , \new_[63946]_ , \new_[63949]_ , \new_[63952]_ ,
    \new_[63953]_ , \new_[63954]_ , \new_[63958]_ , \new_[63959]_ ,
    \new_[63962]_ , \new_[63965]_ , \new_[63966]_ , \new_[63967]_ ,
    \new_[63971]_ , \new_[63972]_ , \new_[63975]_ , \new_[63978]_ ,
    \new_[63979]_ , \new_[63980]_ , \new_[63984]_ , \new_[63985]_ ,
    \new_[63988]_ , \new_[63991]_ , \new_[63992]_ , \new_[63993]_ ,
    \new_[63997]_ , \new_[63998]_ , \new_[64001]_ , \new_[64004]_ ,
    \new_[64005]_ , \new_[64006]_ , \new_[64010]_ , \new_[64011]_ ,
    \new_[64014]_ , \new_[64017]_ , \new_[64018]_ , \new_[64019]_ ,
    \new_[64023]_ , \new_[64024]_ , \new_[64027]_ , \new_[64030]_ ,
    \new_[64031]_ , \new_[64032]_ , \new_[64036]_ , \new_[64037]_ ,
    \new_[64040]_ , \new_[64043]_ , \new_[64044]_ , \new_[64045]_ ,
    \new_[64049]_ , \new_[64050]_ , \new_[64053]_ , \new_[64056]_ ,
    \new_[64057]_ , \new_[64058]_ , \new_[64062]_ , \new_[64063]_ ,
    \new_[64066]_ , \new_[64069]_ , \new_[64070]_ , \new_[64071]_ ,
    \new_[64075]_ , \new_[64076]_ , \new_[64079]_ , \new_[64082]_ ,
    \new_[64083]_ , \new_[64084]_ , \new_[64088]_ , \new_[64089]_ ,
    \new_[64092]_ , \new_[64095]_ , \new_[64096]_ , \new_[64097]_ ,
    \new_[64101]_ , \new_[64102]_ , \new_[64105]_ , \new_[64108]_ ,
    \new_[64109]_ , \new_[64110]_ , \new_[64114]_ , \new_[64115]_ ,
    \new_[64118]_ , \new_[64121]_ , \new_[64122]_ , \new_[64123]_ ,
    \new_[64127]_ , \new_[64128]_ , \new_[64131]_ , \new_[64134]_ ,
    \new_[64135]_ , \new_[64136]_ , \new_[64140]_ , \new_[64141]_ ,
    \new_[64144]_ , \new_[64147]_ , \new_[64148]_ , \new_[64149]_ ,
    \new_[64153]_ , \new_[64154]_ , \new_[64157]_ , \new_[64160]_ ,
    \new_[64161]_ , \new_[64162]_ , \new_[64166]_ , \new_[64167]_ ,
    \new_[64170]_ , \new_[64173]_ , \new_[64174]_ , \new_[64175]_ ,
    \new_[64179]_ , \new_[64180]_ , \new_[64183]_ , \new_[64186]_ ,
    \new_[64187]_ , \new_[64188]_ , \new_[64192]_ , \new_[64193]_ ,
    \new_[64196]_ , \new_[64199]_ , \new_[64200]_ , \new_[64201]_ ,
    \new_[64205]_ , \new_[64206]_ , \new_[64209]_ , \new_[64212]_ ,
    \new_[64213]_ , \new_[64214]_ , \new_[64218]_ , \new_[64219]_ ,
    \new_[64222]_ , \new_[64225]_ , \new_[64226]_ , \new_[64227]_ ,
    \new_[64231]_ , \new_[64232]_ , \new_[64235]_ , \new_[64238]_ ,
    \new_[64239]_ , \new_[64240]_ , \new_[64244]_ , \new_[64245]_ ,
    \new_[64248]_ , \new_[64251]_ , \new_[64252]_ , \new_[64253]_ ,
    \new_[64257]_ , \new_[64258]_ , \new_[64261]_ , \new_[64264]_ ,
    \new_[64265]_ , \new_[64266]_ , \new_[64270]_ , \new_[64271]_ ,
    \new_[64274]_ , \new_[64277]_ , \new_[64278]_ , \new_[64279]_ ,
    \new_[64283]_ , \new_[64284]_ , \new_[64287]_ , \new_[64290]_ ,
    \new_[64291]_ , \new_[64292]_ , \new_[64296]_ , \new_[64297]_ ,
    \new_[64300]_ , \new_[64303]_ , \new_[64304]_ , \new_[64305]_ ,
    \new_[64309]_ , \new_[64310]_ , \new_[64313]_ , \new_[64316]_ ,
    \new_[64317]_ , \new_[64318]_ , \new_[64322]_ , \new_[64323]_ ,
    \new_[64326]_ , \new_[64329]_ , \new_[64330]_ , \new_[64331]_ ,
    \new_[64335]_ , \new_[64336]_ , \new_[64339]_ , \new_[64342]_ ,
    \new_[64343]_ , \new_[64344]_ , \new_[64348]_ , \new_[64349]_ ,
    \new_[64352]_ , \new_[64355]_ , \new_[64356]_ , \new_[64357]_ ,
    \new_[64361]_ , \new_[64362]_ , \new_[64365]_ , \new_[64368]_ ,
    \new_[64369]_ , \new_[64370]_ , \new_[64374]_ , \new_[64375]_ ,
    \new_[64378]_ , \new_[64381]_ , \new_[64382]_ , \new_[64383]_ ,
    \new_[64387]_ , \new_[64388]_ , \new_[64391]_ , \new_[64394]_ ,
    \new_[64395]_ , \new_[64396]_ , \new_[64400]_ , \new_[64401]_ ,
    \new_[64404]_ , \new_[64407]_ , \new_[64408]_ , \new_[64409]_ ,
    \new_[64413]_ , \new_[64414]_ , \new_[64417]_ , \new_[64420]_ ,
    \new_[64421]_ , \new_[64422]_ , \new_[64426]_ , \new_[64427]_ ,
    \new_[64430]_ , \new_[64433]_ , \new_[64434]_ , \new_[64435]_ ,
    \new_[64439]_ , \new_[64440]_ , \new_[64443]_ , \new_[64446]_ ,
    \new_[64447]_ , \new_[64448]_ , \new_[64452]_ , \new_[64453]_ ,
    \new_[64456]_ , \new_[64459]_ , \new_[64460]_ , \new_[64461]_ ,
    \new_[64465]_ , \new_[64466]_ , \new_[64469]_ , \new_[64472]_ ,
    \new_[64473]_ , \new_[64474]_ , \new_[64478]_ , \new_[64479]_ ,
    \new_[64482]_ , \new_[64485]_ , \new_[64486]_ , \new_[64487]_ ,
    \new_[64491]_ , \new_[64492]_ , \new_[64495]_ , \new_[64498]_ ,
    \new_[64499]_ , \new_[64500]_ , \new_[64504]_ , \new_[64505]_ ,
    \new_[64508]_ , \new_[64511]_ , \new_[64512]_ , \new_[64513]_ ,
    \new_[64517]_ , \new_[64518]_ , \new_[64521]_ , \new_[64524]_ ,
    \new_[64525]_ , \new_[64526]_ , \new_[64530]_ , \new_[64531]_ ,
    \new_[64534]_ , \new_[64537]_ , \new_[64538]_ , \new_[64539]_ ,
    \new_[64543]_ , \new_[64544]_ , \new_[64547]_ , \new_[64550]_ ,
    \new_[64551]_ , \new_[64552]_ , \new_[64556]_ , \new_[64557]_ ,
    \new_[64560]_ , \new_[64563]_ , \new_[64564]_ , \new_[64565]_ ,
    \new_[64569]_ , \new_[64570]_ , \new_[64573]_ , \new_[64576]_ ,
    \new_[64577]_ , \new_[64578]_ , \new_[64582]_ , \new_[64583]_ ,
    \new_[64586]_ , \new_[64589]_ , \new_[64590]_ , \new_[64591]_ ,
    \new_[64595]_ , \new_[64596]_ , \new_[64599]_ , \new_[64602]_ ,
    \new_[64603]_ , \new_[64604]_ , \new_[64608]_ , \new_[64609]_ ,
    \new_[64612]_ , \new_[64615]_ , \new_[64616]_ , \new_[64617]_ ,
    \new_[64621]_ , \new_[64622]_ , \new_[64625]_ , \new_[64628]_ ,
    \new_[64629]_ , \new_[64630]_ , \new_[64634]_ , \new_[64635]_ ,
    \new_[64638]_ , \new_[64641]_ , \new_[64642]_ , \new_[64643]_ ,
    \new_[64647]_ , \new_[64648]_ , \new_[64651]_ , \new_[64654]_ ,
    \new_[64655]_ , \new_[64656]_ , \new_[64660]_ , \new_[64661]_ ,
    \new_[64664]_ , \new_[64667]_ , \new_[64668]_ , \new_[64669]_ ,
    \new_[64673]_ , \new_[64674]_ , \new_[64677]_ , \new_[64680]_ ,
    \new_[64681]_ , \new_[64682]_ , \new_[64686]_ , \new_[64687]_ ,
    \new_[64690]_ , \new_[64693]_ , \new_[64694]_ , \new_[64695]_ ,
    \new_[64699]_ , \new_[64700]_ , \new_[64703]_ , \new_[64706]_ ,
    \new_[64707]_ , \new_[64708]_ , \new_[64712]_ , \new_[64713]_ ,
    \new_[64716]_ , \new_[64719]_ , \new_[64720]_ , \new_[64721]_ ,
    \new_[64725]_ , \new_[64726]_ , \new_[64729]_ , \new_[64732]_ ,
    \new_[64733]_ , \new_[64734]_ , \new_[64738]_ , \new_[64739]_ ,
    \new_[64742]_ , \new_[64745]_ , \new_[64746]_ , \new_[64747]_ ,
    \new_[64751]_ , \new_[64752]_ , \new_[64755]_ , \new_[64758]_ ,
    \new_[64759]_ , \new_[64760]_ , \new_[64764]_ , \new_[64765]_ ,
    \new_[64768]_ , \new_[64771]_ , \new_[64772]_ , \new_[64773]_ ,
    \new_[64777]_ , \new_[64778]_ , \new_[64781]_ , \new_[64784]_ ,
    \new_[64785]_ , \new_[64786]_ , \new_[64790]_ , \new_[64791]_ ,
    \new_[64794]_ , \new_[64797]_ , \new_[64798]_ , \new_[64799]_ ,
    \new_[64803]_ , \new_[64804]_ , \new_[64807]_ , \new_[64810]_ ,
    \new_[64811]_ , \new_[64812]_ , \new_[64816]_ , \new_[64817]_ ,
    \new_[64820]_ , \new_[64823]_ , \new_[64824]_ , \new_[64825]_ ,
    \new_[64829]_ , \new_[64830]_ , \new_[64833]_ , \new_[64836]_ ,
    \new_[64837]_ , \new_[64838]_ , \new_[64842]_ , \new_[64843]_ ,
    \new_[64846]_ , \new_[64849]_ , \new_[64850]_ , \new_[64851]_ ,
    \new_[64855]_ , \new_[64856]_ , \new_[64859]_ , \new_[64862]_ ,
    \new_[64863]_ , \new_[64864]_ , \new_[64868]_ , \new_[64869]_ ,
    \new_[64872]_ , \new_[64875]_ , \new_[64876]_ , \new_[64877]_ ,
    \new_[64881]_ , \new_[64882]_ , \new_[64885]_ , \new_[64888]_ ,
    \new_[64889]_ , \new_[64890]_ , \new_[64894]_ , \new_[64895]_ ,
    \new_[64898]_ , \new_[64901]_ , \new_[64902]_ , \new_[64903]_ ,
    \new_[64907]_ , \new_[64908]_ , \new_[64911]_ , \new_[64914]_ ,
    \new_[64915]_ , \new_[64916]_ , \new_[64920]_ , \new_[64921]_ ,
    \new_[64924]_ , \new_[64927]_ , \new_[64928]_ , \new_[64929]_ ,
    \new_[64933]_ , \new_[64934]_ , \new_[64937]_ , \new_[64940]_ ,
    \new_[64941]_ , \new_[64942]_ , \new_[64946]_ , \new_[64947]_ ,
    \new_[64950]_ , \new_[64953]_ , \new_[64954]_ , \new_[64955]_ ,
    \new_[64959]_ , \new_[64960]_ , \new_[64963]_ , \new_[64966]_ ,
    \new_[64967]_ , \new_[64968]_ , \new_[64972]_ , \new_[64973]_ ,
    \new_[64976]_ , \new_[64979]_ , \new_[64980]_ , \new_[64981]_ ,
    \new_[64985]_ , \new_[64986]_ , \new_[64989]_ , \new_[64992]_ ,
    \new_[64993]_ , \new_[64994]_ , \new_[64998]_ , \new_[64999]_ ,
    \new_[65002]_ , \new_[65005]_ , \new_[65006]_ , \new_[65007]_ ,
    \new_[65011]_ , \new_[65012]_ , \new_[65015]_ , \new_[65018]_ ,
    \new_[65019]_ , \new_[65020]_ , \new_[65024]_ , \new_[65025]_ ,
    \new_[65028]_ , \new_[65031]_ , \new_[65032]_ , \new_[65033]_ ,
    \new_[65037]_ , \new_[65038]_ , \new_[65041]_ , \new_[65044]_ ,
    \new_[65045]_ , \new_[65046]_ , \new_[65050]_ , \new_[65051]_ ,
    \new_[65054]_ , \new_[65057]_ , \new_[65058]_ , \new_[65059]_ ,
    \new_[65063]_ , \new_[65064]_ , \new_[65067]_ , \new_[65070]_ ,
    \new_[65071]_ , \new_[65072]_ , \new_[65076]_ , \new_[65077]_ ,
    \new_[65080]_ , \new_[65083]_ , \new_[65084]_ , \new_[65085]_ ,
    \new_[65089]_ , \new_[65090]_ , \new_[65093]_ , \new_[65096]_ ,
    \new_[65097]_ , \new_[65098]_ , \new_[65102]_ , \new_[65103]_ ,
    \new_[65106]_ , \new_[65109]_ , \new_[65110]_ , \new_[65111]_ ,
    \new_[65115]_ , \new_[65116]_ , \new_[65119]_ , \new_[65122]_ ,
    \new_[65123]_ , \new_[65124]_ , \new_[65128]_ , \new_[65129]_ ,
    \new_[65132]_ , \new_[65135]_ , \new_[65136]_ , \new_[65137]_ ,
    \new_[65141]_ , \new_[65142]_ , \new_[65145]_ , \new_[65148]_ ,
    \new_[65149]_ , \new_[65150]_ , \new_[65154]_ , \new_[65155]_ ,
    \new_[65158]_ , \new_[65161]_ , \new_[65162]_ , \new_[65163]_ ,
    \new_[65167]_ , \new_[65168]_ , \new_[65171]_ , \new_[65174]_ ,
    \new_[65175]_ , \new_[65176]_ , \new_[65180]_ , \new_[65181]_ ,
    \new_[65184]_ , \new_[65187]_ , \new_[65188]_ , \new_[65189]_ ,
    \new_[65193]_ , \new_[65194]_ , \new_[65197]_ , \new_[65200]_ ,
    \new_[65201]_ , \new_[65202]_ , \new_[65206]_ , \new_[65207]_ ,
    \new_[65210]_ , \new_[65213]_ , \new_[65214]_ , \new_[65215]_ ,
    \new_[65219]_ , \new_[65220]_ , \new_[65223]_ , \new_[65226]_ ,
    \new_[65227]_ , \new_[65228]_ , \new_[65232]_ , \new_[65233]_ ,
    \new_[65236]_ , \new_[65239]_ , \new_[65240]_ , \new_[65241]_ ,
    \new_[65245]_ , \new_[65246]_ , \new_[65249]_ , \new_[65252]_ ,
    \new_[65253]_ , \new_[65254]_ , \new_[65258]_ , \new_[65259]_ ,
    \new_[65262]_ , \new_[65265]_ , \new_[65266]_ , \new_[65267]_ ,
    \new_[65271]_ , \new_[65272]_ , \new_[65275]_ , \new_[65278]_ ,
    \new_[65279]_ , \new_[65280]_ , \new_[65284]_ , \new_[65285]_ ,
    \new_[65288]_ , \new_[65291]_ , \new_[65292]_ , \new_[65293]_ ,
    \new_[65297]_ , \new_[65298]_ , \new_[65301]_ , \new_[65304]_ ,
    \new_[65305]_ , \new_[65306]_ , \new_[65310]_ , \new_[65311]_ ,
    \new_[65314]_ , \new_[65317]_ , \new_[65318]_ , \new_[65319]_ ,
    \new_[65323]_ , \new_[65324]_ , \new_[65327]_ , \new_[65330]_ ,
    \new_[65331]_ , \new_[65332]_ , \new_[65336]_ , \new_[65337]_ ,
    \new_[65340]_ , \new_[65343]_ , \new_[65344]_ , \new_[65345]_ ,
    \new_[65349]_ , \new_[65350]_ , \new_[65353]_ , \new_[65356]_ ,
    \new_[65357]_ , \new_[65358]_ , \new_[65362]_ , \new_[65363]_ ,
    \new_[65366]_ , \new_[65369]_ , \new_[65370]_ , \new_[65371]_ ,
    \new_[65375]_ , \new_[65376]_ , \new_[65379]_ , \new_[65382]_ ,
    \new_[65383]_ , \new_[65384]_ , \new_[65388]_ , \new_[65389]_ ,
    \new_[65392]_ , \new_[65395]_ , \new_[65396]_ , \new_[65397]_ ,
    \new_[65401]_ , \new_[65402]_ , \new_[65405]_ , \new_[65408]_ ,
    \new_[65409]_ , \new_[65410]_ , \new_[65414]_ , \new_[65415]_ ,
    \new_[65418]_ , \new_[65421]_ , \new_[65422]_ , \new_[65423]_ ,
    \new_[65427]_ , \new_[65428]_ , \new_[65431]_ , \new_[65434]_ ,
    \new_[65435]_ , \new_[65436]_ , \new_[65440]_ , \new_[65441]_ ,
    \new_[65444]_ , \new_[65447]_ , \new_[65448]_ , \new_[65449]_ ,
    \new_[65453]_ , \new_[65454]_ , \new_[65457]_ , \new_[65460]_ ,
    \new_[65461]_ , \new_[65462]_ , \new_[65466]_ , \new_[65467]_ ,
    \new_[65470]_ , \new_[65473]_ , \new_[65474]_ , \new_[65475]_ ,
    \new_[65479]_ , \new_[65480]_ , \new_[65483]_ , \new_[65486]_ ,
    \new_[65487]_ , \new_[65488]_ , \new_[65492]_ , \new_[65493]_ ,
    \new_[65496]_ , \new_[65499]_ , \new_[65500]_ , \new_[65501]_ ,
    \new_[65505]_ , \new_[65506]_ , \new_[65509]_ , \new_[65512]_ ,
    \new_[65513]_ , \new_[65514]_ , \new_[65518]_ , \new_[65519]_ ,
    \new_[65522]_ , \new_[65525]_ , \new_[65526]_ , \new_[65527]_ ,
    \new_[65531]_ , \new_[65532]_ , \new_[65535]_ , \new_[65538]_ ,
    \new_[65539]_ , \new_[65540]_ , \new_[65544]_ , \new_[65545]_ ,
    \new_[65548]_ , \new_[65551]_ , \new_[65552]_ , \new_[65553]_ ,
    \new_[65557]_ , \new_[65558]_ , \new_[65561]_ , \new_[65564]_ ,
    \new_[65565]_ , \new_[65566]_ , \new_[65570]_ , \new_[65571]_ ,
    \new_[65574]_ , \new_[65577]_ , \new_[65578]_ , \new_[65579]_ ,
    \new_[65583]_ , \new_[65584]_ , \new_[65587]_ , \new_[65590]_ ,
    \new_[65591]_ , \new_[65592]_ , \new_[65596]_ , \new_[65597]_ ,
    \new_[65600]_ , \new_[65603]_ , \new_[65604]_ , \new_[65605]_ ,
    \new_[65609]_ , \new_[65610]_ , \new_[65613]_ , \new_[65616]_ ,
    \new_[65617]_ , \new_[65618]_ , \new_[65622]_ , \new_[65623]_ ,
    \new_[65626]_ , \new_[65629]_ , \new_[65630]_ , \new_[65631]_ ,
    \new_[65635]_ , \new_[65636]_ , \new_[65639]_ , \new_[65642]_ ,
    \new_[65643]_ , \new_[65644]_ , \new_[65648]_ , \new_[65649]_ ,
    \new_[65652]_ , \new_[65655]_ , \new_[65656]_ , \new_[65657]_ ,
    \new_[65661]_ , \new_[65662]_ , \new_[65665]_ , \new_[65668]_ ,
    \new_[65669]_ , \new_[65670]_ , \new_[65674]_ , \new_[65675]_ ,
    \new_[65678]_ , \new_[65681]_ , \new_[65682]_ , \new_[65683]_ ,
    \new_[65687]_ , \new_[65688]_ , \new_[65691]_ , \new_[65694]_ ,
    \new_[65695]_ , \new_[65696]_ , \new_[65700]_ , \new_[65701]_ ,
    \new_[65704]_ , \new_[65707]_ , \new_[65708]_ , \new_[65709]_ ,
    \new_[65713]_ , \new_[65714]_ , \new_[65717]_ , \new_[65720]_ ,
    \new_[65721]_ , \new_[65722]_ , \new_[65726]_ , \new_[65727]_ ,
    \new_[65730]_ , \new_[65733]_ , \new_[65734]_ , \new_[65735]_ ,
    \new_[65739]_ , \new_[65740]_ , \new_[65743]_ , \new_[65746]_ ,
    \new_[65747]_ , \new_[65748]_ , \new_[65752]_ , \new_[65753]_ ,
    \new_[65756]_ , \new_[65759]_ , \new_[65760]_ , \new_[65761]_ ,
    \new_[65765]_ , \new_[65766]_ , \new_[65769]_ , \new_[65772]_ ,
    \new_[65773]_ , \new_[65774]_ , \new_[65778]_ , \new_[65779]_ ,
    \new_[65782]_ , \new_[65785]_ , \new_[65786]_ , \new_[65787]_ ,
    \new_[65791]_ , \new_[65792]_ , \new_[65795]_ , \new_[65798]_ ,
    \new_[65799]_ , \new_[65800]_ , \new_[65804]_ , \new_[65805]_ ,
    \new_[65808]_ , \new_[65811]_ , \new_[65812]_ , \new_[65813]_ ,
    \new_[65817]_ , \new_[65818]_ , \new_[65821]_ , \new_[65824]_ ,
    \new_[65825]_ , \new_[65826]_ , \new_[65830]_ , \new_[65831]_ ,
    \new_[65834]_ , \new_[65837]_ , \new_[65838]_ , \new_[65839]_ ,
    \new_[65843]_ , \new_[65844]_ , \new_[65847]_ , \new_[65850]_ ,
    \new_[65851]_ , \new_[65852]_ , \new_[65856]_ , \new_[65857]_ ,
    \new_[65860]_ , \new_[65863]_ , \new_[65864]_ , \new_[65865]_ ,
    \new_[65869]_ , \new_[65870]_ , \new_[65873]_ , \new_[65876]_ ,
    \new_[65877]_ , \new_[65878]_ , \new_[65882]_ , \new_[65883]_ ,
    \new_[65886]_ , \new_[65889]_ , \new_[65890]_ , \new_[65891]_ ,
    \new_[65895]_ , \new_[65896]_ , \new_[65899]_ , \new_[65902]_ ,
    \new_[65903]_ , \new_[65904]_ , \new_[65908]_ , \new_[65909]_ ,
    \new_[65912]_ , \new_[65915]_ , \new_[65916]_ , \new_[65917]_ ,
    \new_[65921]_ , \new_[65922]_ , \new_[65925]_ , \new_[65928]_ ,
    \new_[65929]_ , \new_[65930]_ , \new_[65934]_ , \new_[65935]_ ,
    \new_[65938]_ , \new_[65941]_ , \new_[65942]_ , \new_[65943]_ ,
    \new_[65947]_ , \new_[65948]_ , \new_[65951]_ , \new_[65954]_ ,
    \new_[65955]_ , \new_[65956]_ , \new_[65960]_ , \new_[65961]_ ,
    \new_[65964]_ , \new_[65967]_ , \new_[65968]_ , \new_[65969]_ ,
    \new_[65973]_ , \new_[65974]_ , \new_[65977]_ , \new_[65980]_ ,
    \new_[65981]_ , \new_[65982]_ , \new_[65986]_ , \new_[65987]_ ,
    \new_[65990]_ , \new_[65993]_ , \new_[65994]_ , \new_[65995]_ ,
    \new_[65999]_ , \new_[66000]_ , \new_[66003]_ , \new_[66006]_ ,
    \new_[66007]_ , \new_[66008]_ , \new_[66012]_ , \new_[66013]_ ,
    \new_[66016]_ , \new_[66019]_ , \new_[66020]_ , \new_[66021]_ ,
    \new_[66025]_ , \new_[66026]_ , \new_[66029]_ , \new_[66032]_ ,
    \new_[66033]_ , \new_[66034]_ , \new_[66038]_ , \new_[66039]_ ,
    \new_[66042]_ , \new_[66045]_ , \new_[66046]_ , \new_[66047]_ ,
    \new_[66051]_ , \new_[66052]_ , \new_[66055]_ , \new_[66058]_ ,
    \new_[66059]_ , \new_[66060]_ , \new_[66064]_ , \new_[66065]_ ,
    \new_[66068]_ , \new_[66071]_ , \new_[66072]_ , \new_[66073]_ ,
    \new_[66077]_ , \new_[66078]_ , \new_[66081]_ , \new_[66084]_ ,
    \new_[66085]_ , \new_[66086]_ , \new_[66090]_ , \new_[66091]_ ,
    \new_[66094]_ , \new_[66097]_ , \new_[66098]_ , \new_[66099]_ ,
    \new_[66103]_ , \new_[66104]_ , \new_[66107]_ , \new_[66110]_ ,
    \new_[66111]_ , \new_[66112]_ , \new_[66116]_ , \new_[66117]_ ,
    \new_[66120]_ , \new_[66123]_ , \new_[66124]_ , \new_[66125]_ ,
    \new_[66129]_ , \new_[66130]_ , \new_[66133]_ , \new_[66136]_ ,
    \new_[66137]_ , \new_[66138]_ , \new_[66142]_ , \new_[66143]_ ,
    \new_[66146]_ , \new_[66149]_ , \new_[66150]_ , \new_[66151]_ ,
    \new_[66155]_ , \new_[66156]_ , \new_[66159]_ , \new_[66162]_ ,
    \new_[66163]_ , \new_[66164]_ , \new_[66168]_ , \new_[66169]_ ,
    \new_[66172]_ , \new_[66175]_ , \new_[66176]_ , \new_[66177]_ ,
    \new_[66181]_ , \new_[66182]_ , \new_[66185]_ , \new_[66188]_ ,
    \new_[66189]_ , \new_[66190]_ , \new_[66194]_ , \new_[66195]_ ,
    \new_[66198]_ , \new_[66201]_ , \new_[66202]_ , \new_[66203]_ ,
    \new_[66207]_ , \new_[66208]_ , \new_[66211]_ , \new_[66214]_ ,
    \new_[66215]_ , \new_[66216]_ , \new_[66220]_ , \new_[66221]_ ,
    \new_[66224]_ , \new_[66227]_ , \new_[66228]_ , \new_[66229]_ ,
    \new_[66233]_ , \new_[66234]_ , \new_[66237]_ , \new_[66240]_ ,
    \new_[66241]_ , \new_[66242]_ , \new_[66246]_ , \new_[66247]_ ,
    \new_[66250]_ , \new_[66253]_ , \new_[66254]_ , \new_[66255]_ ,
    \new_[66259]_ , \new_[66260]_ , \new_[66263]_ , \new_[66266]_ ,
    \new_[66267]_ , \new_[66268]_ , \new_[66272]_ , \new_[66273]_ ,
    \new_[66276]_ , \new_[66279]_ , \new_[66280]_ , \new_[66281]_ ,
    \new_[66285]_ , \new_[66286]_ , \new_[66289]_ , \new_[66292]_ ,
    \new_[66293]_ , \new_[66294]_ , \new_[66298]_ , \new_[66299]_ ,
    \new_[66302]_ , \new_[66305]_ , \new_[66306]_ , \new_[66307]_ ,
    \new_[66311]_ , \new_[66312]_ , \new_[66315]_ , \new_[66318]_ ,
    \new_[66319]_ , \new_[66320]_ , \new_[66324]_ , \new_[66325]_ ,
    \new_[66328]_ , \new_[66331]_ , \new_[66332]_ , \new_[66333]_ ,
    \new_[66337]_ , \new_[66338]_ , \new_[66341]_ , \new_[66344]_ ,
    \new_[66345]_ , \new_[66346]_ , \new_[66350]_ , \new_[66351]_ ,
    \new_[66354]_ , \new_[66357]_ , \new_[66358]_ , \new_[66359]_ ,
    \new_[66363]_ , \new_[66364]_ , \new_[66367]_ , \new_[66370]_ ,
    \new_[66371]_ , \new_[66372]_ , \new_[66376]_ , \new_[66377]_ ,
    \new_[66380]_ , \new_[66383]_ , \new_[66384]_ , \new_[66385]_ ,
    \new_[66389]_ , \new_[66390]_ , \new_[66393]_ , \new_[66396]_ ,
    \new_[66397]_ , \new_[66398]_ , \new_[66402]_ , \new_[66403]_ ,
    \new_[66406]_ , \new_[66409]_ , \new_[66410]_ , \new_[66411]_ ,
    \new_[66415]_ , \new_[66416]_ , \new_[66419]_ , \new_[66422]_ ,
    \new_[66423]_ , \new_[66424]_ , \new_[66428]_ , \new_[66429]_ ,
    \new_[66432]_ , \new_[66435]_ , \new_[66436]_ , \new_[66437]_ ,
    \new_[66441]_ , \new_[66442]_ , \new_[66445]_ , \new_[66448]_ ,
    \new_[66449]_ , \new_[66450]_ , \new_[66454]_ , \new_[66455]_ ,
    \new_[66458]_ , \new_[66461]_ , \new_[66462]_ , \new_[66463]_ ,
    \new_[66467]_ , \new_[66468]_ , \new_[66471]_ , \new_[66474]_ ,
    \new_[66475]_ , \new_[66476]_ , \new_[66480]_ , \new_[66481]_ ,
    \new_[66484]_ , \new_[66487]_ , \new_[66488]_ , \new_[66489]_ ,
    \new_[66493]_ , \new_[66494]_ , \new_[66497]_ , \new_[66500]_ ,
    \new_[66501]_ , \new_[66502]_ , \new_[66506]_ , \new_[66507]_ ,
    \new_[66510]_ , \new_[66513]_ , \new_[66514]_ , \new_[66515]_ ,
    \new_[66519]_ , \new_[66520]_ , \new_[66523]_ , \new_[66526]_ ,
    \new_[66527]_ , \new_[66528]_ , \new_[66532]_ , \new_[66533]_ ,
    \new_[66536]_ , \new_[66539]_ , \new_[66540]_ , \new_[66541]_ ,
    \new_[66545]_ , \new_[66546]_ , \new_[66549]_ , \new_[66552]_ ,
    \new_[66553]_ , \new_[66554]_ , \new_[66558]_ , \new_[66559]_ ,
    \new_[66562]_ , \new_[66565]_ , \new_[66566]_ , \new_[66567]_ ,
    \new_[66571]_ , \new_[66572]_ , \new_[66575]_ , \new_[66578]_ ,
    \new_[66579]_ , \new_[66580]_ , \new_[66584]_ , \new_[66585]_ ,
    \new_[66588]_ , \new_[66591]_ , \new_[66592]_ , \new_[66593]_ ,
    \new_[66597]_ , \new_[66598]_ , \new_[66601]_ , \new_[66604]_ ,
    \new_[66605]_ , \new_[66606]_ , \new_[66610]_ , \new_[66611]_ ,
    \new_[66614]_ , \new_[66617]_ , \new_[66618]_ , \new_[66619]_ ,
    \new_[66623]_ , \new_[66624]_ , \new_[66627]_ , \new_[66630]_ ,
    \new_[66631]_ , \new_[66632]_ , \new_[66636]_ , \new_[66637]_ ,
    \new_[66640]_ , \new_[66643]_ , \new_[66644]_ , \new_[66645]_ ,
    \new_[66649]_ , \new_[66650]_ , \new_[66653]_ , \new_[66656]_ ,
    \new_[66657]_ , \new_[66658]_ , \new_[66662]_ , \new_[66663]_ ,
    \new_[66666]_ , \new_[66669]_ , \new_[66670]_ , \new_[66671]_ ,
    \new_[66675]_ , \new_[66676]_ , \new_[66679]_ , \new_[66682]_ ,
    \new_[66683]_ , \new_[66684]_ , \new_[66688]_ , \new_[66689]_ ,
    \new_[66692]_ , \new_[66695]_ , \new_[66696]_ , \new_[66697]_ ,
    \new_[66701]_ , \new_[66702]_ , \new_[66705]_ , \new_[66708]_ ,
    \new_[66709]_ , \new_[66710]_ , \new_[66714]_ , \new_[66715]_ ,
    \new_[66718]_ , \new_[66721]_ , \new_[66722]_ , \new_[66723]_ ,
    \new_[66727]_ , \new_[66728]_ , \new_[66731]_ , \new_[66734]_ ,
    \new_[66735]_ , \new_[66736]_ , \new_[66740]_ , \new_[66741]_ ,
    \new_[66744]_ , \new_[66747]_ , \new_[66748]_ , \new_[66749]_ ,
    \new_[66753]_ , \new_[66754]_ , \new_[66757]_ , \new_[66760]_ ,
    \new_[66761]_ , \new_[66762]_ , \new_[66766]_ , \new_[66767]_ ,
    \new_[66770]_ , \new_[66773]_ , \new_[66774]_ , \new_[66775]_ ,
    \new_[66779]_ , \new_[66780]_ , \new_[66783]_ , \new_[66786]_ ,
    \new_[66787]_ , \new_[66788]_ , \new_[66792]_ , \new_[66793]_ ,
    \new_[66796]_ , \new_[66799]_ , \new_[66800]_ , \new_[66801]_ ,
    \new_[66805]_ , \new_[66806]_ , \new_[66809]_ , \new_[66812]_ ,
    \new_[66813]_ , \new_[66814]_ , \new_[66818]_ , \new_[66819]_ ,
    \new_[66822]_ , \new_[66825]_ , \new_[66826]_ , \new_[66827]_ ,
    \new_[66831]_ , \new_[66832]_ , \new_[66835]_ , \new_[66838]_ ,
    \new_[66839]_ , \new_[66840]_ , \new_[66844]_ , \new_[66845]_ ,
    \new_[66848]_ , \new_[66851]_ , \new_[66852]_ , \new_[66853]_ ,
    \new_[66857]_ , \new_[66858]_ , \new_[66861]_ , \new_[66864]_ ,
    \new_[66865]_ , \new_[66866]_ , \new_[66870]_ , \new_[66871]_ ,
    \new_[66874]_ , \new_[66877]_ , \new_[66878]_ , \new_[66879]_ ,
    \new_[66883]_ , \new_[66884]_ , \new_[66887]_ , \new_[66890]_ ,
    \new_[66891]_ , \new_[66892]_ , \new_[66896]_ , \new_[66897]_ ,
    \new_[66900]_ , \new_[66903]_ , \new_[66904]_ , \new_[66905]_ ,
    \new_[66909]_ , \new_[66910]_ , \new_[66913]_ , \new_[66916]_ ,
    \new_[66917]_ , \new_[66918]_ , \new_[66922]_ , \new_[66923]_ ,
    \new_[66926]_ , \new_[66929]_ , \new_[66930]_ , \new_[66931]_ ,
    \new_[66935]_ , \new_[66936]_ , \new_[66939]_ , \new_[66942]_ ,
    \new_[66943]_ , \new_[66944]_ , \new_[66948]_ , \new_[66949]_ ,
    \new_[66952]_ , \new_[66955]_ , \new_[66956]_ , \new_[66957]_ ,
    \new_[66961]_ , \new_[66962]_ , \new_[66965]_ , \new_[66968]_ ,
    \new_[66969]_ , \new_[66970]_ , \new_[66974]_ , \new_[66975]_ ,
    \new_[66978]_ , \new_[66981]_ , \new_[66982]_ , \new_[66983]_ ,
    \new_[66987]_ , \new_[66988]_ , \new_[66991]_ , \new_[66994]_ ,
    \new_[66995]_ , \new_[66996]_ , \new_[67000]_ , \new_[67001]_ ,
    \new_[67004]_ , \new_[67007]_ , \new_[67008]_ , \new_[67009]_ ,
    \new_[67013]_ , \new_[67014]_ , \new_[67017]_ , \new_[67020]_ ,
    \new_[67021]_ , \new_[67022]_ , \new_[67026]_ , \new_[67027]_ ,
    \new_[67030]_ , \new_[67033]_ , \new_[67034]_ , \new_[67035]_ ,
    \new_[67039]_ , \new_[67040]_ , \new_[67043]_ , \new_[67046]_ ,
    \new_[67047]_ , \new_[67048]_ , \new_[67052]_ , \new_[67053]_ ,
    \new_[67056]_ , \new_[67059]_ , \new_[67060]_ , \new_[67061]_ ,
    \new_[67065]_ , \new_[67066]_ , \new_[67069]_ , \new_[67072]_ ,
    \new_[67073]_ , \new_[67074]_ , \new_[67078]_ , \new_[67079]_ ,
    \new_[67082]_ , \new_[67085]_ , \new_[67086]_ , \new_[67087]_ ,
    \new_[67091]_ , \new_[67092]_ , \new_[67095]_ , \new_[67098]_ ,
    \new_[67099]_ , \new_[67100]_ , \new_[67104]_ , \new_[67105]_ ,
    \new_[67108]_ , \new_[67111]_ , \new_[67112]_ , \new_[67113]_ ,
    \new_[67117]_ , \new_[67118]_ , \new_[67121]_ , \new_[67124]_ ,
    \new_[67125]_ , \new_[67126]_ , \new_[67130]_ , \new_[67131]_ ,
    \new_[67134]_ , \new_[67137]_ , \new_[67138]_ , \new_[67139]_ ,
    \new_[67143]_ , \new_[67144]_ , \new_[67147]_ , \new_[67150]_ ,
    \new_[67151]_ , \new_[67152]_ , \new_[67156]_ , \new_[67157]_ ,
    \new_[67160]_ , \new_[67163]_ , \new_[67164]_ , \new_[67165]_ ,
    \new_[67169]_ , \new_[67170]_ , \new_[67173]_ , \new_[67176]_ ,
    \new_[67177]_ , \new_[67178]_ , \new_[67182]_ , \new_[67183]_ ,
    \new_[67186]_ , \new_[67189]_ , \new_[67190]_ , \new_[67191]_ ,
    \new_[67195]_ , \new_[67196]_ , \new_[67199]_ , \new_[67202]_ ,
    \new_[67203]_ , \new_[67204]_ , \new_[67208]_ , \new_[67209]_ ,
    \new_[67212]_ , \new_[67215]_ , \new_[67216]_ , \new_[67217]_ ,
    \new_[67221]_ , \new_[67222]_ , \new_[67225]_ , \new_[67228]_ ,
    \new_[67229]_ , \new_[67230]_ , \new_[67234]_ , \new_[67235]_ ,
    \new_[67238]_ , \new_[67241]_ , \new_[67242]_ , \new_[67243]_ ,
    \new_[67247]_ , \new_[67248]_ , \new_[67251]_ , \new_[67254]_ ,
    \new_[67255]_ , \new_[67256]_ , \new_[67260]_ , \new_[67261]_ ,
    \new_[67264]_ , \new_[67267]_ , \new_[67268]_ , \new_[67269]_ ,
    \new_[67273]_ , \new_[67274]_ , \new_[67277]_ , \new_[67280]_ ,
    \new_[67281]_ , \new_[67282]_ , \new_[67286]_ , \new_[67287]_ ,
    \new_[67290]_ , \new_[67293]_ , \new_[67294]_ , \new_[67295]_ ,
    \new_[67299]_ , \new_[67300]_ , \new_[67303]_ , \new_[67306]_ ,
    \new_[67307]_ , \new_[67308]_ , \new_[67312]_ , \new_[67313]_ ,
    \new_[67316]_ , \new_[67319]_ , \new_[67320]_ , \new_[67321]_ ,
    \new_[67325]_ , \new_[67326]_ , \new_[67329]_ , \new_[67332]_ ,
    \new_[67333]_ , \new_[67334]_ , \new_[67338]_ , \new_[67339]_ ,
    \new_[67342]_ , \new_[67345]_ , \new_[67346]_ , \new_[67347]_ ,
    \new_[67351]_ , \new_[67352]_ , \new_[67355]_ , \new_[67358]_ ,
    \new_[67359]_ , \new_[67360]_ , \new_[67364]_ , \new_[67365]_ ,
    \new_[67368]_ , \new_[67371]_ , \new_[67372]_ , \new_[67373]_ ,
    \new_[67377]_ , \new_[67378]_ , \new_[67381]_ , \new_[67384]_ ,
    \new_[67385]_ , \new_[67386]_ , \new_[67390]_ , \new_[67391]_ ,
    \new_[67394]_ , \new_[67397]_ , \new_[67398]_ , \new_[67399]_ ,
    \new_[67403]_ , \new_[67404]_ , \new_[67407]_ , \new_[67410]_ ,
    \new_[67411]_ , \new_[67412]_ , \new_[67416]_ , \new_[67417]_ ,
    \new_[67420]_ , \new_[67423]_ , \new_[67424]_ , \new_[67425]_ ,
    \new_[67429]_ , \new_[67430]_ , \new_[67433]_ , \new_[67436]_ ,
    \new_[67437]_ , \new_[67438]_ , \new_[67442]_ , \new_[67443]_ ,
    \new_[67446]_ , \new_[67449]_ , \new_[67450]_ , \new_[67451]_ ,
    \new_[67455]_ , \new_[67456]_ , \new_[67459]_ , \new_[67462]_ ,
    \new_[67463]_ , \new_[67464]_ , \new_[67468]_ , \new_[67469]_ ,
    \new_[67472]_ , \new_[67475]_ , \new_[67476]_ , \new_[67477]_ ,
    \new_[67481]_ , \new_[67482]_ , \new_[67485]_ , \new_[67488]_ ,
    \new_[67489]_ , \new_[67490]_ , \new_[67494]_ , \new_[67495]_ ,
    \new_[67498]_ , \new_[67501]_ , \new_[67502]_ , \new_[67503]_ ,
    \new_[67507]_ , \new_[67508]_ , \new_[67511]_ , \new_[67514]_ ,
    \new_[67515]_ , \new_[67516]_ , \new_[67520]_ , \new_[67521]_ ,
    \new_[67524]_ , \new_[67527]_ , \new_[67528]_ , \new_[67529]_ ,
    \new_[67533]_ , \new_[67534]_ , \new_[67537]_ , \new_[67540]_ ,
    \new_[67541]_ , \new_[67542]_ , \new_[67546]_ , \new_[67547]_ ,
    \new_[67550]_ , \new_[67553]_ , \new_[67554]_ , \new_[67555]_ ,
    \new_[67559]_ , \new_[67560]_ , \new_[67563]_ , \new_[67566]_ ,
    \new_[67567]_ , \new_[67568]_ , \new_[67572]_ , \new_[67573]_ ,
    \new_[67576]_ , \new_[67579]_ , \new_[67580]_ , \new_[67581]_ ,
    \new_[67585]_ , \new_[67586]_ , \new_[67589]_ , \new_[67592]_ ,
    \new_[67593]_ , \new_[67594]_ , \new_[67598]_ , \new_[67599]_ ,
    \new_[67602]_ , \new_[67605]_ , \new_[67606]_ , \new_[67607]_ ,
    \new_[67611]_ , \new_[67612]_ , \new_[67615]_ , \new_[67618]_ ,
    \new_[67619]_ , \new_[67620]_ , \new_[67624]_ , \new_[67625]_ ,
    \new_[67628]_ , \new_[67631]_ , \new_[67632]_ , \new_[67633]_ ,
    \new_[67637]_ , \new_[67638]_ , \new_[67641]_ , \new_[67644]_ ,
    \new_[67645]_ , \new_[67646]_ , \new_[67650]_ , \new_[67651]_ ,
    \new_[67654]_ , \new_[67657]_ , \new_[67658]_ , \new_[67659]_ ,
    \new_[67663]_ , \new_[67664]_ , \new_[67667]_ , \new_[67670]_ ,
    \new_[67671]_ , \new_[67672]_ , \new_[67676]_ , \new_[67677]_ ,
    \new_[67680]_ , \new_[67683]_ , \new_[67684]_ , \new_[67685]_ ,
    \new_[67689]_ , \new_[67690]_ , \new_[67693]_ , \new_[67696]_ ,
    \new_[67697]_ , \new_[67698]_ , \new_[67702]_ , \new_[67703]_ ,
    \new_[67706]_ , \new_[67709]_ , \new_[67710]_ , \new_[67711]_ ,
    \new_[67715]_ , \new_[67716]_ , \new_[67719]_ , \new_[67722]_ ,
    \new_[67723]_ , \new_[67724]_ , \new_[67728]_ , \new_[67729]_ ,
    \new_[67732]_ , \new_[67735]_ , \new_[67736]_ , \new_[67737]_ ,
    \new_[67741]_ , \new_[67742]_ , \new_[67745]_ , \new_[67748]_ ,
    \new_[67749]_ , \new_[67750]_ , \new_[67754]_ , \new_[67755]_ ,
    \new_[67758]_ , \new_[67761]_ , \new_[67762]_ , \new_[67763]_ ,
    \new_[67767]_ , \new_[67768]_ , \new_[67771]_ , \new_[67774]_ ,
    \new_[67775]_ , \new_[67776]_ , \new_[67780]_ , \new_[67781]_ ,
    \new_[67784]_ , \new_[67787]_ , \new_[67788]_ , \new_[67789]_ ,
    \new_[67793]_ , \new_[67794]_ , \new_[67797]_ , \new_[67800]_ ,
    \new_[67801]_ , \new_[67802]_ , \new_[67806]_ , \new_[67807]_ ,
    \new_[67810]_ , \new_[67813]_ , \new_[67814]_ , \new_[67815]_ ,
    \new_[67819]_ , \new_[67820]_ , \new_[67823]_ , \new_[67826]_ ,
    \new_[67827]_ , \new_[67828]_ , \new_[67832]_ , \new_[67833]_ ,
    \new_[67836]_ , \new_[67839]_ , \new_[67840]_ , \new_[67841]_ ,
    \new_[67845]_ , \new_[67846]_ , \new_[67849]_ , \new_[67852]_ ,
    \new_[67853]_ , \new_[67854]_ , \new_[67858]_ , \new_[67859]_ ,
    \new_[67862]_ , \new_[67865]_ , \new_[67866]_ , \new_[67867]_ ,
    \new_[67871]_ , \new_[67872]_ , \new_[67875]_ , \new_[67878]_ ,
    \new_[67879]_ , \new_[67880]_ , \new_[67884]_ , \new_[67885]_ ,
    \new_[67888]_ , \new_[67891]_ , \new_[67892]_ , \new_[67893]_ ,
    \new_[67897]_ , \new_[67898]_ , \new_[67901]_ , \new_[67904]_ ,
    \new_[67905]_ , \new_[67906]_ , \new_[67910]_ , \new_[67911]_ ,
    \new_[67914]_ , \new_[67917]_ , \new_[67918]_ , \new_[67919]_ ,
    \new_[67923]_ , \new_[67924]_ , \new_[67927]_ , \new_[67930]_ ,
    \new_[67931]_ , \new_[67932]_ , \new_[67936]_ , \new_[67937]_ ,
    \new_[67940]_ , \new_[67943]_ , \new_[67944]_ , \new_[67945]_ ,
    \new_[67949]_ , \new_[67950]_ , \new_[67953]_ , \new_[67956]_ ,
    \new_[67957]_ , \new_[67958]_ , \new_[67962]_ , \new_[67963]_ ,
    \new_[67966]_ , \new_[67969]_ , \new_[67970]_ , \new_[67971]_ ,
    \new_[67975]_ , \new_[67976]_ , \new_[67979]_ , \new_[67982]_ ,
    \new_[67983]_ , \new_[67984]_ , \new_[67988]_ , \new_[67989]_ ,
    \new_[67992]_ , \new_[67995]_ , \new_[67996]_ , \new_[67997]_ ,
    \new_[68001]_ , \new_[68002]_ , \new_[68005]_ , \new_[68008]_ ,
    \new_[68009]_ , \new_[68010]_ , \new_[68014]_ , \new_[68015]_ ,
    \new_[68018]_ , \new_[68021]_ , \new_[68022]_ , \new_[68023]_ ,
    \new_[68027]_ , \new_[68028]_ , \new_[68031]_ , \new_[68034]_ ,
    \new_[68035]_ , \new_[68036]_ , \new_[68040]_ , \new_[68041]_ ,
    \new_[68044]_ , \new_[68047]_ , \new_[68048]_ , \new_[68049]_ ,
    \new_[68053]_ , \new_[68054]_ , \new_[68057]_ , \new_[68060]_ ,
    \new_[68061]_ , \new_[68062]_ , \new_[68066]_ , \new_[68067]_ ,
    \new_[68070]_ , \new_[68073]_ , \new_[68074]_ , \new_[68075]_ ,
    \new_[68079]_ , \new_[68080]_ , \new_[68083]_ , \new_[68086]_ ,
    \new_[68087]_ , \new_[68088]_ , \new_[68092]_ , \new_[68093]_ ,
    \new_[68096]_ , \new_[68099]_ , \new_[68100]_ , \new_[68101]_ ,
    \new_[68105]_ , \new_[68106]_ , \new_[68109]_ , \new_[68112]_ ,
    \new_[68113]_ , \new_[68114]_ , \new_[68118]_ , \new_[68119]_ ,
    \new_[68122]_ , \new_[68125]_ , \new_[68126]_ , \new_[68127]_ ,
    \new_[68131]_ , \new_[68132]_ , \new_[68135]_ , \new_[68138]_ ,
    \new_[68139]_ , \new_[68140]_ , \new_[68144]_ , \new_[68145]_ ,
    \new_[68148]_ , \new_[68151]_ , \new_[68152]_ , \new_[68153]_ ,
    \new_[68157]_ , \new_[68158]_ , \new_[68161]_ , \new_[68164]_ ,
    \new_[68165]_ , \new_[68166]_ , \new_[68170]_ , \new_[68171]_ ,
    \new_[68174]_ , \new_[68177]_ , \new_[68178]_ , \new_[68179]_ ,
    \new_[68183]_ , \new_[68184]_ , \new_[68187]_ , \new_[68190]_ ,
    \new_[68191]_ , \new_[68192]_ , \new_[68196]_ , \new_[68197]_ ,
    \new_[68200]_ , \new_[68203]_ , \new_[68204]_ , \new_[68205]_ ,
    \new_[68209]_ , \new_[68210]_ , \new_[68213]_ , \new_[68216]_ ,
    \new_[68217]_ , \new_[68218]_ , \new_[68222]_ , \new_[68223]_ ,
    \new_[68226]_ , \new_[68229]_ , \new_[68230]_ , \new_[68231]_ ,
    \new_[68235]_ , \new_[68236]_ , \new_[68239]_ , \new_[68242]_ ,
    \new_[68243]_ , \new_[68244]_ , \new_[68248]_ , \new_[68249]_ ,
    \new_[68252]_ , \new_[68255]_ , \new_[68256]_ , \new_[68257]_ ,
    \new_[68261]_ , \new_[68262]_ , \new_[68265]_ , \new_[68268]_ ,
    \new_[68269]_ , \new_[68270]_ , \new_[68274]_ , \new_[68275]_ ,
    \new_[68278]_ , \new_[68281]_ , \new_[68282]_ , \new_[68283]_ ,
    \new_[68287]_ , \new_[68288]_ , \new_[68291]_ , \new_[68294]_ ,
    \new_[68295]_ , \new_[68296]_ , \new_[68300]_ , \new_[68301]_ ,
    \new_[68304]_ , \new_[68307]_ , \new_[68308]_ , \new_[68309]_ ,
    \new_[68313]_ , \new_[68314]_ , \new_[68317]_ , \new_[68320]_ ,
    \new_[68321]_ , \new_[68322]_ , \new_[68326]_ , \new_[68327]_ ,
    \new_[68330]_ , \new_[68333]_ , \new_[68334]_ , \new_[68335]_ ,
    \new_[68339]_ , \new_[68340]_ , \new_[68343]_ , \new_[68346]_ ,
    \new_[68347]_ , \new_[68348]_ , \new_[68352]_ , \new_[68353]_ ,
    \new_[68356]_ , \new_[68359]_ , \new_[68360]_ , \new_[68361]_ ,
    \new_[68365]_ , \new_[68366]_ , \new_[68369]_ , \new_[68372]_ ,
    \new_[68373]_ , \new_[68374]_ , \new_[68378]_ , \new_[68379]_ ,
    \new_[68382]_ , \new_[68385]_ , \new_[68386]_ , \new_[68387]_ ,
    \new_[68391]_ , \new_[68392]_ , \new_[68395]_ , \new_[68398]_ ,
    \new_[68399]_ , \new_[68400]_ , \new_[68404]_ , \new_[68405]_ ,
    \new_[68408]_ , \new_[68411]_ , \new_[68412]_ , \new_[68413]_ ,
    \new_[68417]_ , \new_[68418]_ , \new_[68421]_ , \new_[68424]_ ,
    \new_[68425]_ , \new_[68426]_ , \new_[68430]_ , \new_[68431]_ ,
    \new_[68434]_ , \new_[68437]_ , \new_[68438]_ , \new_[68439]_ ,
    \new_[68443]_ , \new_[68444]_ , \new_[68447]_ , \new_[68450]_ ,
    \new_[68451]_ , \new_[68452]_ , \new_[68456]_ , \new_[68457]_ ,
    \new_[68460]_ , \new_[68463]_ , \new_[68464]_ , \new_[68465]_ ,
    \new_[68469]_ , \new_[68470]_ , \new_[68473]_ , \new_[68476]_ ,
    \new_[68477]_ , \new_[68478]_ , \new_[68482]_ , \new_[68483]_ ,
    \new_[68486]_ , \new_[68489]_ , \new_[68490]_ , \new_[68491]_ ,
    \new_[68495]_ , \new_[68496]_ , \new_[68499]_ , \new_[68502]_ ,
    \new_[68503]_ , \new_[68504]_ , \new_[68508]_ , \new_[68509]_ ,
    \new_[68512]_ , \new_[68515]_ , \new_[68516]_ , \new_[68517]_ ,
    \new_[68521]_ , \new_[68522]_ , \new_[68525]_ , \new_[68528]_ ,
    \new_[68529]_ , \new_[68530]_ , \new_[68534]_ , \new_[68535]_ ,
    \new_[68538]_ , \new_[68541]_ , \new_[68542]_ , \new_[68543]_ ,
    \new_[68547]_ , \new_[68548]_ , \new_[68551]_ , \new_[68554]_ ,
    \new_[68555]_ , \new_[68556]_ , \new_[68560]_ , \new_[68561]_ ,
    \new_[68564]_ , \new_[68567]_ , \new_[68568]_ , \new_[68569]_ ,
    \new_[68573]_ , \new_[68574]_ , \new_[68577]_ , \new_[68580]_ ,
    \new_[68581]_ , \new_[68582]_ , \new_[68586]_ , \new_[68587]_ ,
    \new_[68590]_ , \new_[68593]_ , \new_[68594]_ , \new_[68595]_ ,
    \new_[68599]_ , \new_[68600]_ , \new_[68603]_ , \new_[68606]_ ,
    \new_[68607]_ , \new_[68608]_ , \new_[68612]_ , \new_[68613]_ ,
    \new_[68616]_ , \new_[68619]_ , \new_[68620]_ , \new_[68621]_ ,
    \new_[68625]_ , \new_[68626]_ , \new_[68629]_ , \new_[68632]_ ,
    \new_[68633]_ , \new_[68634]_ , \new_[68638]_ , \new_[68639]_ ,
    \new_[68642]_ , \new_[68645]_ , \new_[68646]_ , \new_[68647]_ ,
    \new_[68651]_ , \new_[68652]_ , \new_[68655]_ , \new_[68658]_ ,
    \new_[68659]_ , \new_[68660]_ , \new_[68664]_ , \new_[68665]_ ,
    \new_[68668]_ , \new_[68671]_ , \new_[68672]_ , \new_[68673]_ ,
    \new_[68677]_ , \new_[68678]_ , \new_[68681]_ , \new_[68684]_ ,
    \new_[68685]_ , \new_[68686]_ , \new_[68690]_ , \new_[68691]_ ,
    \new_[68694]_ , \new_[68697]_ , \new_[68698]_ , \new_[68699]_ ,
    \new_[68703]_ , \new_[68704]_ , \new_[68707]_ , \new_[68710]_ ,
    \new_[68711]_ , \new_[68712]_ , \new_[68716]_ , \new_[68717]_ ,
    \new_[68720]_ , \new_[68723]_ , \new_[68724]_ , \new_[68725]_ ,
    \new_[68729]_ , \new_[68730]_ , \new_[68733]_ , \new_[68736]_ ,
    \new_[68737]_ , \new_[68738]_ , \new_[68742]_ , \new_[68743]_ ,
    \new_[68746]_ , \new_[68749]_ , \new_[68750]_ , \new_[68751]_ ,
    \new_[68755]_ , \new_[68756]_ , \new_[68759]_ , \new_[68762]_ ,
    \new_[68763]_ , \new_[68764]_ , \new_[68768]_ , \new_[68769]_ ,
    \new_[68772]_ , \new_[68775]_ , \new_[68776]_ , \new_[68777]_ ,
    \new_[68781]_ , \new_[68782]_ , \new_[68785]_ , \new_[68788]_ ,
    \new_[68789]_ , \new_[68790]_ , \new_[68794]_ , \new_[68795]_ ,
    \new_[68798]_ , \new_[68801]_ , \new_[68802]_ , \new_[68803]_ ,
    \new_[68807]_ , \new_[68808]_ , \new_[68811]_ , \new_[68814]_ ,
    \new_[68815]_ , \new_[68816]_ , \new_[68820]_ , \new_[68821]_ ,
    \new_[68824]_ , \new_[68827]_ , \new_[68828]_ , \new_[68829]_ ,
    \new_[68833]_ , \new_[68834]_ , \new_[68837]_ , \new_[68840]_ ,
    \new_[68841]_ , \new_[68842]_ , \new_[68846]_ , \new_[68847]_ ,
    \new_[68850]_ , \new_[68853]_ , \new_[68854]_ , \new_[68855]_ ,
    \new_[68859]_ , \new_[68860]_ , \new_[68863]_ , \new_[68866]_ ,
    \new_[68867]_ , \new_[68868]_ , \new_[68872]_ , \new_[68873]_ ,
    \new_[68876]_ , \new_[68879]_ , \new_[68880]_ , \new_[68881]_ ,
    \new_[68885]_ , \new_[68886]_ , \new_[68889]_ , \new_[68892]_ ,
    \new_[68893]_ , \new_[68894]_ , \new_[68898]_ , \new_[68899]_ ,
    \new_[68902]_ , \new_[68905]_ , \new_[68906]_ , \new_[68907]_ ,
    \new_[68911]_ , \new_[68912]_ , \new_[68915]_ , \new_[68918]_ ,
    \new_[68919]_ , \new_[68920]_ , \new_[68924]_ , \new_[68925]_ ,
    \new_[68928]_ , \new_[68931]_ , \new_[68932]_ , \new_[68933]_ ,
    \new_[68937]_ , \new_[68938]_ , \new_[68941]_ , \new_[68944]_ ,
    \new_[68945]_ , \new_[68946]_ , \new_[68950]_ , \new_[68951]_ ,
    \new_[68954]_ , \new_[68957]_ , \new_[68958]_ , \new_[68959]_ ,
    \new_[68963]_ , \new_[68964]_ , \new_[68967]_ , \new_[68970]_ ,
    \new_[68971]_ , \new_[68972]_ , \new_[68976]_ , \new_[68977]_ ,
    \new_[68980]_ , \new_[68983]_ , \new_[68984]_ , \new_[68985]_ ,
    \new_[68989]_ , \new_[68990]_ , \new_[68993]_ , \new_[68996]_ ,
    \new_[68997]_ , \new_[68998]_ , \new_[69002]_ , \new_[69003]_ ,
    \new_[69006]_ , \new_[69009]_ , \new_[69010]_ , \new_[69011]_ ,
    \new_[69015]_ , \new_[69016]_ , \new_[69019]_ , \new_[69022]_ ,
    \new_[69023]_ , \new_[69024]_ , \new_[69028]_ , \new_[69029]_ ,
    \new_[69032]_ , \new_[69035]_ , \new_[69036]_ , \new_[69037]_ ,
    \new_[69041]_ , \new_[69042]_ , \new_[69045]_ , \new_[69048]_ ,
    \new_[69049]_ , \new_[69050]_ , \new_[69054]_ , \new_[69055]_ ,
    \new_[69058]_ , \new_[69061]_ , \new_[69062]_ , \new_[69063]_ ,
    \new_[69067]_ , \new_[69068]_ , \new_[69071]_ , \new_[69074]_ ,
    \new_[69075]_ , \new_[69076]_ , \new_[69080]_ , \new_[69081]_ ,
    \new_[69084]_ , \new_[69087]_ , \new_[69088]_ , \new_[69089]_ ,
    \new_[69093]_ , \new_[69094]_ , \new_[69097]_ , \new_[69100]_ ,
    \new_[69101]_ , \new_[69102]_ , \new_[69106]_ , \new_[69107]_ ,
    \new_[69110]_ , \new_[69113]_ , \new_[69114]_ , \new_[69115]_ ,
    \new_[69119]_ , \new_[69120]_ , \new_[69123]_ , \new_[69126]_ ,
    \new_[69127]_ , \new_[69128]_ , \new_[69132]_ , \new_[69133]_ ,
    \new_[69136]_ , \new_[69139]_ , \new_[69140]_ , \new_[69141]_ ,
    \new_[69145]_ , \new_[69146]_ , \new_[69149]_ , \new_[69152]_ ,
    \new_[69153]_ , \new_[69154]_ , \new_[69158]_ , \new_[69159]_ ,
    \new_[69162]_ , \new_[69165]_ , \new_[69166]_ , \new_[69167]_ ,
    \new_[69171]_ , \new_[69172]_ , \new_[69175]_ , \new_[69178]_ ,
    \new_[69179]_ , \new_[69180]_ , \new_[69184]_ , \new_[69185]_ ,
    \new_[69188]_ , \new_[69191]_ , \new_[69192]_ , \new_[69193]_ ,
    \new_[69197]_ , \new_[69198]_ , \new_[69201]_ , \new_[69204]_ ,
    \new_[69205]_ , \new_[69206]_ , \new_[69210]_ , \new_[69211]_ ,
    \new_[69214]_ , \new_[69217]_ , \new_[69218]_ , \new_[69219]_ ,
    \new_[69223]_ , \new_[69224]_ , \new_[69227]_ , \new_[69230]_ ,
    \new_[69231]_ , \new_[69232]_ , \new_[69236]_ , \new_[69237]_ ,
    \new_[69240]_ , \new_[69243]_ , \new_[69244]_ , \new_[69245]_ ,
    \new_[69249]_ , \new_[69250]_ , \new_[69253]_ , \new_[69256]_ ,
    \new_[69257]_ , \new_[69258]_ , \new_[69262]_ , \new_[69263]_ ,
    \new_[69266]_ , \new_[69269]_ , \new_[69270]_ , \new_[69271]_ ,
    \new_[69275]_ , \new_[69276]_ , \new_[69279]_ , \new_[69282]_ ,
    \new_[69283]_ , \new_[69284]_ , \new_[69288]_ , \new_[69289]_ ,
    \new_[69292]_ , \new_[69295]_ , \new_[69296]_ , \new_[69297]_ ,
    \new_[69301]_ , \new_[69302]_ , \new_[69305]_ , \new_[69308]_ ,
    \new_[69309]_ , \new_[69310]_ , \new_[69314]_ , \new_[69315]_ ,
    \new_[69318]_ , \new_[69321]_ , \new_[69322]_ , \new_[69323]_ ,
    \new_[69327]_ , \new_[69328]_ , \new_[69331]_ , \new_[69334]_ ,
    \new_[69335]_ , \new_[69336]_ , \new_[69340]_ , \new_[69341]_ ,
    \new_[69344]_ , \new_[69347]_ , \new_[69348]_ , \new_[69349]_ ,
    \new_[69353]_ , \new_[69354]_ , \new_[69357]_ , \new_[69360]_ ,
    \new_[69361]_ , \new_[69362]_ , \new_[69366]_ , \new_[69367]_ ,
    \new_[69370]_ , \new_[69373]_ , \new_[69374]_ , \new_[69375]_ ,
    \new_[69379]_ , \new_[69380]_ , \new_[69383]_ , \new_[69386]_ ,
    \new_[69387]_ , \new_[69388]_ , \new_[69392]_ , \new_[69393]_ ,
    \new_[69396]_ , \new_[69399]_ , \new_[69400]_ , \new_[69401]_ ,
    \new_[69405]_ , \new_[69406]_ , \new_[69409]_ , \new_[69412]_ ,
    \new_[69413]_ , \new_[69414]_ , \new_[69418]_ , \new_[69419]_ ,
    \new_[69422]_ , \new_[69425]_ , \new_[69426]_ , \new_[69427]_ ,
    \new_[69431]_ , \new_[69432]_ , \new_[69435]_ , \new_[69438]_ ,
    \new_[69439]_ , \new_[69440]_ , \new_[69444]_ , \new_[69445]_ ,
    \new_[69448]_ , \new_[69451]_ , \new_[69452]_ , \new_[69453]_ ,
    \new_[69457]_ , \new_[69458]_ , \new_[69461]_ , \new_[69464]_ ,
    \new_[69465]_ , \new_[69466]_ , \new_[69470]_ , \new_[69471]_ ,
    \new_[69474]_ , \new_[69477]_ , \new_[69478]_ , \new_[69479]_ ,
    \new_[69483]_ , \new_[69484]_ , \new_[69487]_ , \new_[69490]_ ,
    \new_[69491]_ , \new_[69492]_ , \new_[69496]_ , \new_[69497]_ ,
    \new_[69500]_ , \new_[69503]_ , \new_[69504]_ , \new_[69505]_ ,
    \new_[69509]_ , \new_[69510]_ , \new_[69513]_ , \new_[69516]_ ,
    \new_[69517]_ , \new_[69518]_ , \new_[69522]_ , \new_[69523]_ ,
    \new_[69526]_ , \new_[69529]_ , \new_[69530]_ , \new_[69531]_ ,
    \new_[69535]_ , \new_[69536]_ , \new_[69539]_ , \new_[69542]_ ,
    \new_[69543]_ , \new_[69544]_ , \new_[69548]_ , \new_[69549]_ ,
    \new_[69552]_ , \new_[69555]_ , \new_[69556]_ , \new_[69557]_ ,
    \new_[69561]_ , \new_[69562]_ , \new_[69565]_ , \new_[69568]_ ,
    \new_[69569]_ , \new_[69570]_ , \new_[69574]_ , \new_[69575]_ ,
    \new_[69578]_ , \new_[69581]_ , \new_[69582]_ , \new_[69583]_ ,
    \new_[69587]_ , \new_[69588]_ , \new_[69591]_ , \new_[69594]_ ,
    \new_[69595]_ , \new_[69596]_ , \new_[69600]_ , \new_[69601]_ ,
    \new_[69604]_ , \new_[69607]_ , \new_[69608]_ , \new_[69609]_ ,
    \new_[69613]_ , \new_[69614]_ , \new_[69617]_ , \new_[69620]_ ,
    \new_[69621]_ , \new_[69622]_ , \new_[69626]_ , \new_[69627]_ ,
    \new_[69630]_ , \new_[69633]_ , \new_[69634]_ , \new_[69635]_ ,
    \new_[69639]_ , \new_[69640]_ , \new_[69643]_ , \new_[69646]_ ,
    \new_[69647]_ , \new_[69648]_ , \new_[69652]_ , \new_[69653]_ ,
    \new_[69656]_ , \new_[69659]_ , \new_[69660]_ , \new_[69661]_ ,
    \new_[69665]_ , \new_[69666]_ , \new_[69669]_ , \new_[69672]_ ,
    \new_[69673]_ , \new_[69674]_ , \new_[69678]_ , \new_[69679]_ ,
    \new_[69682]_ , \new_[69685]_ , \new_[69686]_ , \new_[69687]_ ,
    \new_[69691]_ , \new_[69692]_ , \new_[69695]_ , \new_[69698]_ ,
    \new_[69699]_ , \new_[69700]_ , \new_[69704]_ , \new_[69705]_ ,
    \new_[69708]_ , \new_[69711]_ , \new_[69712]_ , \new_[69713]_ ,
    \new_[69717]_ , \new_[69718]_ , \new_[69721]_ , \new_[69724]_ ,
    \new_[69725]_ , \new_[69726]_ , \new_[69730]_ , \new_[69731]_ ,
    \new_[69734]_ , \new_[69737]_ , \new_[69738]_ , \new_[69739]_ ,
    \new_[69743]_ , \new_[69744]_ , \new_[69747]_ , \new_[69750]_ ,
    \new_[69751]_ , \new_[69752]_ , \new_[69756]_ , \new_[69757]_ ,
    \new_[69760]_ , \new_[69763]_ , \new_[69764]_ , \new_[69765]_ ,
    \new_[69769]_ , \new_[69770]_ , \new_[69773]_ , \new_[69776]_ ,
    \new_[69777]_ , \new_[69778]_ , \new_[69782]_ , \new_[69783]_ ,
    \new_[69786]_ , \new_[69789]_ , \new_[69790]_ , \new_[69791]_ ,
    \new_[69795]_ , \new_[69796]_ , \new_[69799]_ , \new_[69802]_ ,
    \new_[69803]_ , \new_[69804]_ , \new_[69808]_ , \new_[69809]_ ,
    \new_[69812]_ , \new_[69815]_ , \new_[69816]_ , \new_[69817]_ ,
    \new_[69821]_ , \new_[69822]_ , \new_[69825]_ , \new_[69828]_ ,
    \new_[69829]_ , \new_[69830]_ , \new_[69834]_ , \new_[69835]_ ,
    \new_[69838]_ , \new_[69841]_ , \new_[69842]_ , \new_[69843]_ ,
    \new_[69847]_ , \new_[69848]_ , \new_[69851]_ , \new_[69854]_ ,
    \new_[69855]_ , \new_[69856]_ , \new_[69860]_ , \new_[69861]_ ,
    \new_[69864]_ , \new_[69867]_ , \new_[69868]_ , \new_[69869]_ ,
    \new_[69873]_ , \new_[69874]_ , \new_[69877]_ , \new_[69880]_ ,
    \new_[69881]_ , \new_[69882]_ , \new_[69886]_ , \new_[69887]_ ,
    \new_[69890]_ , \new_[69893]_ , \new_[69894]_ , \new_[69895]_ ,
    \new_[69899]_ , \new_[69900]_ , \new_[69903]_ , \new_[69906]_ ,
    \new_[69907]_ , \new_[69908]_ , \new_[69912]_ , \new_[69913]_ ,
    \new_[69916]_ , \new_[69919]_ , \new_[69920]_ , \new_[69921]_ ,
    \new_[69925]_ , \new_[69926]_ , \new_[69929]_ , \new_[69932]_ ,
    \new_[69933]_ , \new_[69934]_ , \new_[69938]_ , \new_[69939]_ ,
    \new_[69942]_ , \new_[69945]_ , \new_[69946]_ , \new_[69947]_ ,
    \new_[69951]_ , \new_[69952]_ , \new_[69955]_ , \new_[69958]_ ,
    \new_[69959]_ , \new_[69960]_ , \new_[69964]_ , \new_[69965]_ ,
    \new_[69968]_ , \new_[69971]_ , \new_[69972]_ , \new_[69973]_ ,
    \new_[69977]_ , \new_[69978]_ , \new_[69981]_ , \new_[69984]_ ,
    \new_[69985]_ , \new_[69986]_ , \new_[69990]_ , \new_[69991]_ ,
    \new_[69994]_ , \new_[69997]_ , \new_[69998]_ , \new_[69999]_ ,
    \new_[70003]_ , \new_[70004]_ , \new_[70007]_ , \new_[70010]_ ,
    \new_[70011]_ , \new_[70012]_ , \new_[70016]_ , \new_[70017]_ ,
    \new_[70020]_ , \new_[70023]_ , \new_[70024]_ , \new_[70025]_ ,
    \new_[70029]_ , \new_[70030]_ , \new_[70033]_ , \new_[70036]_ ,
    \new_[70037]_ , \new_[70038]_ , \new_[70042]_ , \new_[70043]_ ,
    \new_[70046]_ , \new_[70049]_ , \new_[70050]_ , \new_[70051]_ ,
    \new_[70055]_ , \new_[70056]_ , \new_[70059]_ , \new_[70062]_ ,
    \new_[70063]_ , \new_[70064]_ , \new_[70068]_ , \new_[70069]_ ,
    \new_[70072]_ , \new_[70075]_ , \new_[70076]_ , \new_[70077]_ ,
    \new_[70081]_ , \new_[70082]_ , \new_[70085]_ , \new_[70088]_ ,
    \new_[70089]_ , \new_[70090]_ , \new_[70094]_ , \new_[70095]_ ,
    \new_[70098]_ , \new_[70101]_ , \new_[70102]_ , \new_[70103]_ ,
    \new_[70107]_ , \new_[70108]_ , \new_[70111]_ , \new_[70114]_ ,
    \new_[70115]_ , \new_[70116]_ , \new_[70120]_ , \new_[70121]_ ,
    \new_[70124]_ , \new_[70127]_ , \new_[70128]_ , \new_[70129]_ ,
    \new_[70133]_ , \new_[70134]_ , \new_[70137]_ , \new_[70140]_ ,
    \new_[70141]_ , \new_[70142]_ , \new_[70146]_ , \new_[70147]_ ,
    \new_[70150]_ , \new_[70153]_ , \new_[70154]_ , \new_[70155]_ ,
    \new_[70159]_ , \new_[70160]_ , \new_[70163]_ , \new_[70166]_ ,
    \new_[70167]_ , \new_[70168]_ , \new_[70172]_ , \new_[70173]_ ,
    \new_[70176]_ , \new_[70179]_ , \new_[70180]_ , \new_[70181]_ ,
    \new_[70185]_ , \new_[70186]_ , \new_[70189]_ , \new_[70192]_ ,
    \new_[70193]_ , \new_[70194]_ , \new_[70198]_ , \new_[70199]_ ,
    \new_[70202]_ , \new_[70205]_ , \new_[70206]_ , \new_[70207]_ ,
    \new_[70211]_ , \new_[70212]_ , \new_[70215]_ , \new_[70218]_ ,
    \new_[70219]_ , \new_[70220]_ , \new_[70224]_ , \new_[70225]_ ,
    \new_[70228]_ , \new_[70231]_ , \new_[70232]_ , \new_[70233]_ ,
    \new_[70237]_ , \new_[70238]_ , \new_[70241]_ , \new_[70244]_ ,
    \new_[70245]_ , \new_[70246]_ , \new_[70250]_ , \new_[70251]_ ,
    \new_[70254]_ , \new_[70257]_ , \new_[70258]_ , \new_[70259]_ ,
    \new_[70263]_ , \new_[70264]_ , \new_[70267]_ , \new_[70270]_ ,
    \new_[70271]_ , \new_[70272]_ , \new_[70276]_ , \new_[70277]_ ,
    \new_[70280]_ , \new_[70283]_ , \new_[70284]_ , \new_[70285]_ ,
    \new_[70289]_ , \new_[70290]_ , \new_[70293]_ , \new_[70296]_ ,
    \new_[70297]_ , \new_[70298]_ , \new_[70302]_ , \new_[70303]_ ,
    \new_[70306]_ , \new_[70309]_ , \new_[70310]_ , \new_[70311]_ ,
    \new_[70315]_ , \new_[70316]_ , \new_[70319]_ , \new_[70322]_ ,
    \new_[70323]_ , \new_[70324]_ , \new_[70328]_ , \new_[70329]_ ,
    \new_[70332]_ , \new_[70335]_ , \new_[70336]_ , \new_[70337]_ ,
    \new_[70341]_ , \new_[70342]_ , \new_[70345]_ , \new_[70348]_ ,
    \new_[70349]_ , \new_[70350]_ , \new_[70354]_ , \new_[70355]_ ,
    \new_[70358]_ , \new_[70361]_ , \new_[70362]_ , \new_[70363]_ ,
    \new_[70367]_ , \new_[70368]_ , \new_[70371]_ , \new_[70374]_ ,
    \new_[70375]_ , \new_[70376]_ , \new_[70380]_ , \new_[70381]_ ,
    \new_[70384]_ , \new_[70387]_ , \new_[70388]_ , \new_[70389]_ ,
    \new_[70393]_ , \new_[70394]_ , \new_[70397]_ , \new_[70400]_ ,
    \new_[70401]_ , \new_[70402]_ , \new_[70406]_ , \new_[70407]_ ,
    \new_[70410]_ , \new_[70413]_ , \new_[70414]_ , \new_[70415]_ ,
    \new_[70419]_ , \new_[70420]_ , \new_[70423]_ , \new_[70426]_ ,
    \new_[70427]_ , \new_[70428]_ , \new_[70432]_ , \new_[70433]_ ,
    \new_[70436]_ , \new_[70439]_ , \new_[70440]_ , \new_[70441]_ ,
    \new_[70445]_ , \new_[70446]_ , \new_[70449]_ , \new_[70452]_ ,
    \new_[70453]_ , \new_[70454]_ , \new_[70458]_ , \new_[70459]_ ,
    \new_[70462]_ , \new_[70465]_ , \new_[70466]_ , \new_[70467]_ ,
    \new_[70471]_ , \new_[70472]_ , \new_[70475]_ , \new_[70478]_ ,
    \new_[70479]_ , \new_[70480]_ , \new_[70484]_ , \new_[70485]_ ,
    \new_[70488]_ , \new_[70491]_ , \new_[70492]_ , \new_[70493]_ ,
    \new_[70497]_ , \new_[70498]_ , \new_[70501]_ , \new_[70504]_ ,
    \new_[70505]_ , \new_[70506]_ , \new_[70510]_ , \new_[70511]_ ,
    \new_[70514]_ , \new_[70517]_ , \new_[70518]_ , \new_[70519]_ ,
    \new_[70523]_ , \new_[70524]_ , \new_[70527]_ , \new_[70530]_ ,
    \new_[70531]_ , \new_[70532]_ , \new_[70536]_ , \new_[70537]_ ,
    \new_[70540]_ , \new_[70543]_ , \new_[70544]_ , \new_[70545]_ ,
    \new_[70549]_ , \new_[70550]_ , \new_[70553]_ , \new_[70556]_ ,
    \new_[70557]_ , \new_[70558]_ , \new_[70562]_ , \new_[70563]_ ,
    \new_[70566]_ , \new_[70569]_ , \new_[70570]_ , \new_[70571]_ ,
    \new_[70575]_ , \new_[70576]_ , \new_[70579]_ , \new_[70582]_ ,
    \new_[70583]_ , \new_[70584]_ , \new_[70588]_ , \new_[70589]_ ,
    \new_[70592]_ , \new_[70595]_ , \new_[70596]_ , \new_[70597]_ ,
    \new_[70601]_ , \new_[70602]_ , \new_[70605]_ , \new_[70608]_ ,
    \new_[70609]_ , \new_[70610]_ , \new_[70614]_ , \new_[70615]_ ,
    \new_[70618]_ , \new_[70621]_ , \new_[70622]_ , \new_[70623]_ ,
    \new_[70627]_ , \new_[70628]_ , \new_[70631]_ , \new_[70634]_ ,
    \new_[70635]_ , \new_[70636]_ , \new_[70640]_ , \new_[70641]_ ,
    \new_[70644]_ , \new_[70647]_ , \new_[70648]_ , \new_[70649]_ ,
    \new_[70653]_ , \new_[70654]_ , \new_[70657]_ , \new_[70660]_ ,
    \new_[70661]_ , \new_[70662]_ , \new_[70666]_ , \new_[70667]_ ,
    \new_[70670]_ , \new_[70673]_ , \new_[70674]_ , \new_[70675]_ ,
    \new_[70679]_ , \new_[70680]_ , \new_[70683]_ , \new_[70686]_ ,
    \new_[70687]_ , \new_[70688]_ , \new_[70692]_ , \new_[70693]_ ,
    \new_[70696]_ , \new_[70699]_ , \new_[70700]_ , \new_[70701]_ ,
    \new_[70705]_ , \new_[70706]_ , \new_[70709]_ , \new_[70712]_ ,
    \new_[70713]_ , \new_[70714]_ , \new_[70718]_ , \new_[70719]_ ,
    \new_[70722]_ , \new_[70725]_ , \new_[70726]_ , \new_[70727]_ ,
    \new_[70731]_ , \new_[70732]_ , \new_[70735]_ , \new_[70738]_ ,
    \new_[70739]_ , \new_[70740]_ , \new_[70744]_ , \new_[70745]_ ,
    \new_[70748]_ , \new_[70751]_ , \new_[70752]_ , \new_[70753]_ ,
    \new_[70757]_ , \new_[70758]_ , \new_[70761]_ , \new_[70764]_ ,
    \new_[70765]_ , \new_[70766]_ , \new_[70770]_ , \new_[70771]_ ,
    \new_[70774]_ , \new_[70777]_ , \new_[70778]_ , \new_[70779]_ ,
    \new_[70783]_ , \new_[70784]_ , \new_[70787]_ , \new_[70790]_ ,
    \new_[70791]_ , \new_[70792]_ , \new_[70796]_ , \new_[70797]_ ,
    \new_[70800]_ , \new_[70803]_ , \new_[70804]_ , \new_[70805]_ ,
    \new_[70809]_ , \new_[70810]_ , \new_[70813]_ , \new_[70816]_ ,
    \new_[70817]_ , \new_[70818]_ , \new_[70822]_ , \new_[70823]_ ,
    \new_[70826]_ , \new_[70829]_ , \new_[70830]_ , \new_[70831]_ ,
    \new_[70835]_ , \new_[70836]_ , \new_[70839]_ , \new_[70842]_ ,
    \new_[70843]_ , \new_[70844]_ , \new_[70848]_ , \new_[70849]_ ,
    \new_[70852]_ , \new_[70855]_ , \new_[70856]_ , \new_[70857]_ ,
    \new_[70861]_ , \new_[70862]_ , \new_[70865]_ , \new_[70868]_ ,
    \new_[70869]_ , \new_[70870]_ , \new_[70874]_ , \new_[70875]_ ,
    \new_[70878]_ , \new_[70881]_ , \new_[70882]_ , \new_[70883]_ ,
    \new_[70887]_ , \new_[70888]_ , \new_[70891]_ , \new_[70894]_ ,
    \new_[70895]_ , \new_[70896]_ , \new_[70900]_ , \new_[70901]_ ,
    \new_[70904]_ , \new_[70907]_ , \new_[70908]_ , \new_[70909]_ ,
    \new_[70913]_ , \new_[70914]_ , \new_[70917]_ , \new_[70920]_ ,
    \new_[70921]_ , \new_[70922]_ , \new_[70926]_ , \new_[70927]_ ,
    \new_[70930]_ , \new_[70933]_ , \new_[70934]_ , \new_[70935]_ ,
    \new_[70939]_ , \new_[70940]_ , \new_[70943]_ , \new_[70946]_ ,
    \new_[70947]_ , \new_[70948]_ , \new_[70952]_ , \new_[70953]_ ,
    \new_[70956]_ , \new_[70959]_ , \new_[70960]_ , \new_[70961]_ ,
    \new_[70965]_ , \new_[70966]_ , \new_[70969]_ , \new_[70972]_ ,
    \new_[70973]_ , \new_[70974]_ , \new_[70978]_ , \new_[70979]_ ,
    \new_[70982]_ , \new_[70985]_ , \new_[70986]_ , \new_[70987]_ ,
    \new_[70991]_ , \new_[70992]_ , \new_[70995]_ , \new_[70998]_ ,
    \new_[70999]_ , \new_[71000]_ , \new_[71004]_ , \new_[71005]_ ,
    \new_[71008]_ , \new_[71011]_ , \new_[71012]_ , \new_[71013]_ ,
    \new_[71017]_ , \new_[71018]_ , \new_[71021]_ , \new_[71024]_ ,
    \new_[71025]_ , \new_[71026]_ , \new_[71030]_ , \new_[71031]_ ,
    \new_[71034]_ , \new_[71037]_ , \new_[71038]_ , \new_[71039]_ ,
    \new_[71043]_ , \new_[71044]_ , \new_[71047]_ , \new_[71050]_ ,
    \new_[71051]_ , \new_[71052]_ , \new_[71056]_ , \new_[71057]_ ,
    \new_[71060]_ , \new_[71063]_ , \new_[71064]_ , \new_[71065]_ ,
    \new_[71069]_ , \new_[71070]_ , \new_[71073]_ , \new_[71076]_ ,
    \new_[71077]_ , \new_[71078]_ , \new_[71082]_ , \new_[71083]_ ,
    \new_[71086]_ , \new_[71089]_ , \new_[71090]_ , \new_[71091]_ ,
    \new_[71095]_ , \new_[71096]_ , \new_[71099]_ , \new_[71102]_ ,
    \new_[71103]_ , \new_[71104]_ , \new_[71108]_ , \new_[71109]_ ,
    \new_[71112]_ , \new_[71115]_ , \new_[71116]_ , \new_[71117]_ ,
    \new_[71121]_ , \new_[71122]_ , \new_[71125]_ , \new_[71128]_ ,
    \new_[71129]_ , \new_[71130]_ , \new_[71134]_ , \new_[71135]_ ,
    \new_[71138]_ , \new_[71141]_ , \new_[71142]_ , \new_[71143]_ ,
    \new_[71147]_ , \new_[71148]_ , \new_[71151]_ , \new_[71154]_ ,
    \new_[71155]_ , \new_[71156]_ , \new_[71160]_ , \new_[71161]_ ,
    \new_[71164]_ , \new_[71167]_ , \new_[71168]_ , \new_[71169]_ ,
    \new_[71173]_ , \new_[71174]_ , \new_[71177]_ , \new_[71180]_ ,
    \new_[71181]_ , \new_[71182]_ , \new_[71186]_ , \new_[71187]_ ,
    \new_[71190]_ , \new_[71193]_ , \new_[71194]_ , \new_[71195]_ ,
    \new_[71199]_ , \new_[71200]_ , \new_[71203]_ , \new_[71206]_ ,
    \new_[71207]_ , \new_[71208]_ , \new_[71212]_ , \new_[71213]_ ,
    \new_[71216]_ , \new_[71219]_ , \new_[71220]_ , \new_[71221]_ ,
    \new_[71225]_ , \new_[71226]_ , \new_[71229]_ , \new_[71232]_ ,
    \new_[71233]_ , \new_[71234]_ , \new_[71238]_ , \new_[71239]_ ,
    \new_[71242]_ , \new_[71245]_ , \new_[71246]_ , \new_[71247]_ ,
    \new_[71251]_ , \new_[71252]_ , \new_[71255]_ , \new_[71258]_ ,
    \new_[71259]_ , \new_[71260]_ , \new_[71264]_ , \new_[71265]_ ,
    \new_[71268]_ , \new_[71271]_ , \new_[71272]_ , \new_[71273]_ ,
    \new_[71277]_ , \new_[71278]_ , \new_[71281]_ , \new_[71284]_ ,
    \new_[71285]_ , \new_[71286]_ , \new_[71290]_ , \new_[71291]_ ,
    \new_[71294]_ , \new_[71297]_ , \new_[71298]_ , \new_[71299]_ ,
    \new_[71303]_ , \new_[71304]_ , \new_[71307]_ , \new_[71310]_ ,
    \new_[71311]_ , \new_[71312]_ , \new_[71316]_ , \new_[71317]_ ,
    \new_[71320]_ , \new_[71323]_ , \new_[71324]_ , \new_[71325]_ ,
    \new_[71329]_ , \new_[71330]_ , \new_[71333]_ , \new_[71336]_ ,
    \new_[71337]_ , \new_[71338]_ , \new_[71342]_ , \new_[71343]_ ,
    \new_[71346]_ , \new_[71349]_ , \new_[71350]_ , \new_[71351]_ ,
    \new_[71355]_ , \new_[71356]_ , \new_[71359]_ , \new_[71362]_ ,
    \new_[71363]_ , \new_[71364]_ , \new_[71368]_ , \new_[71369]_ ,
    \new_[71372]_ , \new_[71375]_ , \new_[71376]_ , \new_[71377]_ ,
    \new_[71381]_ , \new_[71382]_ , \new_[71385]_ , \new_[71388]_ ,
    \new_[71389]_ , \new_[71390]_ , \new_[71394]_ , \new_[71395]_ ,
    \new_[71398]_ , \new_[71401]_ , \new_[71402]_ , \new_[71403]_ ,
    \new_[71407]_ , \new_[71408]_ , \new_[71411]_ , \new_[71414]_ ,
    \new_[71415]_ , \new_[71416]_ , \new_[71420]_ , \new_[71421]_ ,
    \new_[71424]_ , \new_[71427]_ , \new_[71428]_ , \new_[71429]_ ,
    \new_[71433]_ , \new_[71434]_ , \new_[71437]_ , \new_[71440]_ ,
    \new_[71441]_ , \new_[71442]_ , \new_[71446]_ , \new_[71447]_ ,
    \new_[71450]_ , \new_[71453]_ , \new_[71454]_ , \new_[71455]_ ,
    \new_[71459]_ , \new_[71460]_ , \new_[71463]_ , \new_[71466]_ ,
    \new_[71467]_ , \new_[71468]_ , \new_[71472]_ , \new_[71473]_ ,
    \new_[71476]_ , \new_[71479]_ , \new_[71480]_ , \new_[71481]_ ,
    \new_[71485]_ , \new_[71486]_ , \new_[71489]_ , \new_[71492]_ ,
    \new_[71493]_ , \new_[71494]_ , \new_[71498]_ , \new_[71499]_ ,
    \new_[71502]_ , \new_[71505]_ , \new_[71506]_ , \new_[71507]_ ,
    \new_[71511]_ , \new_[71512]_ , \new_[71515]_ , \new_[71518]_ ,
    \new_[71519]_ , \new_[71520]_ , \new_[71524]_ , \new_[71525]_ ,
    \new_[71528]_ , \new_[71531]_ , \new_[71532]_ , \new_[71533]_ ,
    \new_[71537]_ , \new_[71538]_ , \new_[71541]_ , \new_[71544]_ ,
    \new_[71545]_ , \new_[71546]_ , \new_[71550]_ , \new_[71551]_ ,
    \new_[71554]_ , \new_[71557]_ , \new_[71558]_ , \new_[71559]_ ,
    \new_[71563]_ , \new_[71564]_ , \new_[71567]_ , \new_[71570]_ ,
    \new_[71571]_ , \new_[71572]_ , \new_[71576]_ , \new_[71577]_ ,
    \new_[71580]_ , \new_[71583]_ , \new_[71584]_ , \new_[71585]_ ,
    \new_[71589]_ , \new_[71590]_ , \new_[71593]_ , \new_[71596]_ ,
    \new_[71597]_ , \new_[71598]_ , \new_[71602]_ , \new_[71603]_ ,
    \new_[71606]_ , \new_[71609]_ , \new_[71610]_ , \new_[71611]_ ,
    \new_[71615]_ , \new_[71616]_ , \new_[71619]_ , \new_[71622]_ ,
    \new_[71623]_ , \new_[71624]_ , \new_[71628]_ , \new_[71629]_ ,
    \new_[71632]_ , \new_[71635]_ , \new_[71636]_ , \new_[71637]_ ,
    \new_[71641]_ , \new_[71642]_ , \new_[71645]_ , \new_[71648]_ ,
    \new_[71649]_ , \new_[71650]_ , \new_[71654]_ , \new_[71655]_ ,
    \new_[71658]_ , \new_[71661]_ , \new_[71662]_ , \new_[71663]_ ,
    \new_[71667]_ , \new_[71668]_ , \new_[71671]_ , \new_[71674]_ ,
    \new_[71675]_ , \new_[71676]_ , \new_[71680]_ , \new_[71681]_ ,
    \new_[71684]_ , \new_[71687]_ , \new_[71688]_ , \new_[71689]_ ,
    \new_[71693]_ , \new_[71694]_ , \new_[71697]_ , \new_[71700]_ ,
    \new_[71701]_ , \new_[71702]_ , \new_[71706]_ , \new_[71707]_ ,
    \new_[71710]_ , \new_[71713]_ , \new_[71714]_ , \new_[71715]_ ,
    \new_[71719]_ , \new_[71720]_ , \new_[71723]_ , \new_[71726]_ ,
    \new_[71727]_ , \new_[71728]_ , \new_[71732]_ , \new_[71733]_ ,
    \new_[71736]_ , \new_[71739]_ , \new_[71740]_ , \new_[71741]_ ,
    \new_[71745]_ , \new_[71746]_ , \new_[71749]_ , \new_[71752]_ ,
    \new_[71753]_ , \new_[71754]_ , \new_[71758]_ , \new_[71759]_ ,
    \new_[71762]_ , \new_[71765]_ , \new_[71766]_ , \new_[71767]_ ,
    \new_[71771]_ , \new_[71772]_ , \new_[71775]_ , \new_[71778]_ ,
    \new_[71779]_ , \new_[71780]_ , \new_[71784]_ , \new_[71785]_ ,
    \new_[71788]_ , \new_[71791]_ , \new_[71792]_ , \new_[71793]_ ,
    \new_[71797]_ , \new_[71798]_ , \new_[71801]_ , \new_[71804]_ ,
    \new_[71805]_ , \new_[71806]_ , \new_[71810]_ , \new_[71811]_ ,
    \new_[71814]_ , \new_[71817]_ , \new_[71818]_ , \new_[71819]_ ,
    \new_[71823]_ , \new_[71824]_ , \new_[71827]_ , \new_[71830]_ ,
    \new_[71831]_ , \new_[71832]_ , \new_[71836]_ , \new_[71837]_ ,
    \new_[71840]_ , \new_[71843]_ , \new_[71844]_ , \new_[71845]_ ,
    \new_[71849]_ , \new_[71850]_ , \new_[71853]_ , \new_[71856]_ ,
    \new_[71857]_ , \new_[71858]_ , \new_[71862]_ , \new_[71863]_ ,
    \new_[71866]_ , \new_[71869]_ , \new_[71870]_ , \new_[71871]_ ,
    \new_[71875]_ , \new_[71876]_ , \new_[71879]_ , \new_[71882]_ ,
    \new_[71883]_ , \new_[71884]_ , \new_[71888]_ , \new_[71889]_ ,
    \new_[71892]_ , \new_[71895]_ , \new_[71896]_ , \new_[71897]_ ,
    \new_[71901]_ , \new_[71902]_ , \new_[71905]_ , \new_[71908]_ ,
    \new_[71909]_ , \new_[71910]_ , \new_[71914]_ , \new_[71915]_ ,
    \new_[71918]_ , \new_[71921]_ , \new_[71922]_ , \new_[71923]_ ,
    \new_[71927]_ , \new_[71928]_ , \new_[71931]_ , \new_[71934]_ ,
    \new_[71935]_ , \new_[71936]_ , \new_[71940]_ , \new_[71941]_ ,
    \new_[71944]_ , \new_[71947]_ , \new_[71948]_ , \new_[71949]_ ,
    \new_[71953]_ , \new_[71954]_ , \new_[71957]_ , \new_[71960]_ ,
    \new_[71961]_ , \new_[71962]_ , \new_[71966]_ , \new_[71967]_ ,
    \new_[71970]_ , \new_[71973]_ , \new_[71974]_ , \new_[71975]_ ,
    \new_[71979]_ , \new_[71980]_ , \new_[71983]_ , \new_[71986]_ ,
    \new_[71987]_ , \new_[71988]_ , \new_[71992]_ , \new_[71993]_ ,
    \new_[71996]_ , \new_[71999]_ , \new_[72000]_ , \new_[72001]_ ,
    \new_[72005]_ , \new_[72006]_ , \new_[72009]_ , \new_[72012]_ ,
    \new_[72013]_ , \new_[72014]_ , \new_[72018]_ , \new_[72019]_ ,
    \new_[72022]_ , \new_[72025]_ , \new_[72026]_ , \new_[72027]_ ,
    \new_[72031]_ , \new_[72032]_ , \new_[72035]_ , \new_[72038]_ ,
    \new_[72039]_ , \new_[72040]_ , \new_[72044]_ , \new_[72045]_ ,
    \new_[72048]_ , \new_[72051]_ , \new_[72052]_ , \new_[72053]_ ,
    \new_[72057]_ , \new_[72058]_ , \new_[72061]_ , \new_[72064]_ ,
    \new_[72065]_ , \new_[72066]_ , \new_[72070]_ , \new_[72071]_ ,
    \new_[72074]_ , \new_[72077]_ , \new_[72078]_ , \new_[72079]_ ,
    \new_[72083]_ , \new_[72084]_ , \new_[72087]_ , \new_[72090]_ ,
    \new_[72091]_ , \new_[72092]_ , \new_[72096]_ , \new_[72097]_ ,
    \new_[72100]_ , \new_[72103]_ , \new_[72104]_ , \new_[72105]_ ,
    \new_[72109]_ , \new_[72110]_ , \new_[72113]_ , \new_[72116]_ ,
    \new_[72117]_ , \new_[72118]_ , \new_[72122]_ , \new_[72123]_ ,
    \new_[72126]_ , \new_[72129]_ , \new_[72130]_ , \new_[72131]_ ,
    \new_[72135]_ , \new_[72136]_ , \new_[72139]_ , \new_[72142]_ ,
    \new_[72143]_ , \new_[72144]_ , \new_[72148]_ , \new_[72149]_ ,
    \new_[72152]_ , \new_[72155]_ , \new_[72156]_ , \new_[72157]_ ,
    \new_[72161]_ , \new_[72162]_ , \new_[72165]_ , \new_[72168]_ ,
    \new_[72169]_ , \new_[72170]_ , \new_[72174]_ , \new_[72175]_ ,
    \new_[72178]_ , \new_[72181]_ , \new_[72182]_ , \new_[72183]_ ,
    \new_[72187]_ , \new_[72188]_ , \new_[72191]_ , \new_[72194]_ ,
    \new_[72195]_ , \new_[72196]_ , \new_[72200]_ , \new_[72201]_ ,
    \new_[72204]_ , \new_[72207]_ , \new_[72208]_ , \new_[72209]_ ,
    \new_[72213]_ , \new_[72214]_ , \new_[72217]_ , \new_[72220]_ ,
    \new_[72221]_ , \new_[72222]_ , \new_[72226]_ , \new_[72227]_ ,
    \new_[72230]_ , \new_[72233]_ , \new_[72234]_ , \new_[72235]_ ,
    \new_[72239]_ , \new_[72240]_ , \new_[72243]_ , \new_[72246]_ ,
    \new_[72247]_ , \new_[72248]_ , \new_[72252]_ , \new_[72253]_ ,
    \new_[72256]_ , \new_[72259]_ , \new_[72260]_ , \new_[72261]_ ,
    \new_[72265]_ , \new_[72266]_ , \new_[72269]_ , \new_[72272]_ ,
    \new_[72273]_ , \new_[72274]_ , \new_[72278]_ , \new_[72279]_ ,
    \new_[72282]_ , \new_[72285]_ , \new_[72286]_ , \new_[72287]_ ,
    \new_[72291]_ , \new_[72292]_ , \new_[72295]_ , \new_[72298]_ ,
    \new_[72299]_ , \new_[72300]_ , \new_[72304]_ , \new_[72305]_ ,
    \new_[72308]_ , \new_[72311]_ , \new_[72312]_ , \new_[72313]_ ,
    \new_[72317]_ , \new_[72318]_ , \new_[72321]_ , \new_[72324]_ ,
    \new_[72325]_ , \new_[72326]_ , \new_[72330]_ , \new_[72331]_ ,
    \new_[72334]_ , \new_[72337]_ , \new_[72338]_ , \new_[72339]_ ,
    \new_[72343]_ , \new_[72344]_ , \new_[72347]_ , \new_[72350]_ ,
    \new_[72351]_ , \new_[72352]_ , \new_[72356]_ , \new_[72357]_ ,
    \new_[72360]_ , \new_[72363]_ , \new_[72364]_ , \new_[72365]_ ,
    \new_[72369]_ , \new_[72370]_ , \new_[72373]_ , \new_[72376]_ ,
    \new_[72377]_ , \new_[72378]_ , \new_[72382]_ , \new_[72383]_ ,
    \new_[72386]_ , \new_[72389]_ , \new_[72390]_ , \new_[72391]_ ,
    \new_[72395]_ , \new_[72396]_ , \new_[72399]_ , \new_[72402]_ ,
    \new_[72403]_ , \new_[72404]_ , \new_[72408]_ , \new_[72409]_ ,
    \new_[72412]_ , \new_[72415]_ , \new_[72416]_ , \new_[72417]_ ,
    \new_[72421]_ , \new_[72422]_ , \new_[72425]_ , \new_[72428]_ ,
    \new_[72429]_ , \new_[72430]_ , \new_[72434]_ , \new_[72435]_ ,
    \new_[72438]_ , \new_[72441]_ , \new_[72442]_ , \new_[72443]_ ,
    \new_[72447]_ , \new_[72448]_ , \new_[72451]_ , \new_[72454]_ ,
    \new_[72455]_ , \new_[72456]_ , \new_[72460]_ , \new_[72461]_ ,
    \new_[72464]_ , \new_[72467]_ , \new_[72468]_ , \new_[72469]_ ,
    \new_[72473]_ , \new_[72474]_ , \new_[72477]_ , \new_[72480]_ ,
    \new_[72481]_ , \new_[72482]_ , \new_[72486]_ , \new_[72487]_ ,
    \new_[72490]_ , \new_[72493]_ , \new_[72494]_ , \new_[72495]_ ,
    \new_[72499]_ , \new_[72500]_ , \new_[72503]_ , \new_[72506]_ ,
    \new_[72507]_ , \new_[72508]_ , \new_[72512]_ , \new_[72513]_ ,
    \new_[72516]_ , \new_[72519]_ , \new_[72520]_ , \new_[72521]_ ,
    \new_[72525]_ , \new_[72526]_ , \new_[72529]_ , \new_[72532]_ ,
    \new_[72533]_ , \new_[72534]_ , \new_[72538]_ , \new_[72539]_ ,
    \new_[72542]_ , \new_[72545]_ , \new_[72546]_ , \new_[72547]_ ,
    \new_[72551]_ , \new_[72552]_ , \new_[72555]_ , \new_[72558]_ ,
    \new_[72559]_ , \new_[72560]_ , \new_[72564]_ , \new_[72565]_ ,
    \new_[72568]_ , \new_[72571]_ , \new_[72572]_ , \new_[72573]_ ,
    \new_[72577]_ , \new_[72578]_ , \new_[72581]_ , \new_[72584]_ ,
    \new_[72585]_ , \new_[72586]_ , \new_[72590]_ , \new_[72591]_ ,
    \new_[72594]_ , \new_[72597]_ , \new_[72598]_ , \new_[72599]_ ,
    \new_[72603]_ , \new_[72604]_ , \new_[72607]_ , \new_[72610]_ ,
    \new_[72611]_ , \new_[72612]_ , \new_[72616]_ , \new_[72617]_ ,
    \new_[72620]_ , \new_[72623]_ , \new_[72624]_ , \new_[72625]_ ,
    \new_[72629]_ , \new_[72630]_ , \new_[72633]_ , \new_[72636]_ ,
    \new_[72637]_ , \new_[72638]_ , \new_[72642]_ , \new_[72643]_ ,
    \new_[72646]_ , \new_[72649]_ , \new_[72650]_ , \new_[72651]_ ,
    \new_[72655]_ , \new_[72656]_ , \new_[72659]_ , \new_[72662]_ ,
    \new_[72663]_ , \new_[72664]_ , \new_[72668]_ , \new_[72669]_ ,
    \new_[72672]_ , \new_[72675]_ , \new_[72676]_ , \new_[72677]_ ,
    \new_[72681]_ , \new_[72682]_ , \new_[72685]_ , \new_[72688]_ ,
    \new_[72689]_ , \new_[72690]_ , \new_[72694]_ , \new_[72695]_ ,
    \new_[72698]_ , \new_[72701]_ , \new_[72702]_ , \new_[72703]_ ,
    \new_[72707]_ , \new_[72708]_ , \new_[72711]_ , \new_[72714]_ ,
    \new_[72715]_ , \new_[72716]_ , \new_[72720]_ , \new_[72721]_ ,
    \new_[72724]_ , \new_[72727]_ , \new_[72728]_ , \new_[72729]_ ,
    \new_[72733]_ , \new_[72734]_ , \new_[72737]_ , \new_[72740]_ ,
    \new_[72741]_ , \new_[72742]_ , \new_[72746]_ , \new_[72747]_ ,
    \new_[72750]_ , \new_[72753]_ , \new_[72754]_ , \new_[72755]_ ,
    \new_[72759]_ , \new_[72760]_ , \new_[72763]_ , \new_[72766]_ ,
    \new_[72767]_ , \new_[72768]_ , \new_[72772]_ , \new_[72773]_ ,
    \new_[72776]_ , \new_[72779]_ , \new_[72780]_ , \new_[72781]_ ,
    \new_[72785]_ , \new_[72786]_ , \new_[72789]_ , \new_[72792]_ ,
    \new_[72793]_ , \new_[72794]_ , \new_[72798]_ , \new_[72799]_ ,
    \new_[72802]_ , \new_[72805]_ , \new_[72806]_ , \new_[72807]_ ,
    \new_[72811]_ , \new_[72812]_ , \new_[72815]_ , \new_[72818]_ ,
    \new_[72819]_ , \new_[72820]_ , \new_[72824]_ , \new_[72825]_ ,
    \new_[72828]_ , \new_[72831]_ , \new_[72832]_ , \new_[72833]_ ,
    \new_[72837]_ , \new_[72838]_ , \new_[72841]_ , \new_[72844]_ ,
    \new_[72845]_ , \new_[72846]_ , \new_[72850]_ , \new_[72851]_ ,
    \new_[72854]_ , \new_[72857]_ , \new_[72858]_ , \new_[72859]_ ,
    \new_[72863]_ , \new_[72864]_ , \new_[72867]_ , \new_[72870]_ ,
    \new_[72871]_ , \new_[72872]_ , \new_[72876]_ , \new_[72877]_ ,
    \new_[72880]_ , \new_[72883]_ , \new_[72884]_ , \new_[72885]_ ,
    \new_[72889]_ , \new_[72890]_ , \new_[72893]_ , \new_[72896]_ ,
    \new_[72897]_ , \new_[72898]_ , \new_[72902]_ , \new_[72903]_ ,
    \new_[72906]_ , \new_[72909]_ , \new_[72910]_ , \new_[72911]_ ,
    \new_[72915]_ , \new_[72916]_ , \new_[72919]_ , \new_[72922]_ ,
    \new_[72923]_ , \new_[72924]_ , \new_[72928]_ , \new_[72929]_ ,
    \new_[72932]_ , \new_[72935]_ , \new_[72936]_ , \new_[72937]_ ,
    \new_[72941]_ , \new_[72942]_ , \new_[72945]_ , \new_[72948]_ ,
    \new_[72949]_ , \new_[72950]_ , \new_[72954]_ , \new_[72955]_ ,
    \new_[72958]_ , \new_[72961]_ , \new_[72962]_ , \new_[72963]_ ,
    \new_[72967]_ , \new_[72968]_ , \new_[72971]_ , \new_[72974]_ ,
    \new_[72975]_ , \new_[72976]_ , \new_[72980]_ , \new_[72981]_ ,
    \new_[72984]_ , \new_[72987]_ , \new_[72988]_ , \new_[72989]_ ,
    \new_[72993]_ , \new_[72994]_ , \new_[72997]_ , \new_[73000]_ ,
    \new_[73001]_ , \new_[73002]_ , \new_[73006]_ , \new_[73007]_ ,
    \new_[73010]_ , \new_[73013]_ , \new_[73014]_ , \new_[73015]_ ,
    \new_[73019]_ , \new_[73020]_ , \new_[73023]_ , \new_[73026]_ ,
    \new_[73027]_ , \new_[73028]_ , \new_[73032]_ , \new_[73033]_ ,
    \new_[73036]_ , \new_[73039]_ , \new_[73040]_ , \new_[73041]_ ,
    \new_[73045]_ , \new_[73046]_ , \new_[73049]_ , \new_[73052]_ ,
    \new_[73053]_ , \new_[73054]_ , \new_[73058]_ , \new_[73059]_ ,
    \new_[73062]_ , \new_[73065]_ , \new_[73066]_ , \new_[73067]_ ,
    \new_[73071]_ , \new_[73072]_ , \new_[73075]_ , \new_[73078]_ ,
    \new_[73079]_ , \new_[73080]_ , \new_[73084]_ , \new_[73085]_ ,
    \new_[73088]_ , \new_[73091]_ , \new_[73092]_ , \new_[73093]_ ,
    \new_[73097]_ , \new_[73098]_ , \new_[73101]_ , \new_[73104]_ ,
    \new_[73105]_ , \new_[73106]_ , \new_[73110]_ , \new_[73111]_ ,
    \new_[73114]_ , \new_[73117]_ , \new_[73118]_ , \new_[73119]_ ,
    \new_[73123]_ , \new_[73124]_ , \new_[73127]_ , \new_[73130]_ ,
    \new_[73131]_ , \new_[73132]_ , \new_[73136]_ , \new_[73137]_ ,
    \new_[73140]_ , \new_[73143]_ , \new_[73144]_ , \new_[73145]_ ,
    \new_[73149]_ , \new_[73150]_ , \new_[73153]_ , \new_[73156]_ ,
    \new_[73157]_ , \new_[73158]_ , \new_[73162]_ , \new_[73163]_ ,
    \new_[73166]_ , \new_[73169]_ , \new_[73170]_ , \new_[73171]_ ,
    \new_[73175]_ , \new_[73176]_ , \new_[73179]_ , \new_[73182]_ ,
    \new_[73183]_ , \new_[73184]_ , \new_[73188]_ , \new_[73189]_ ,
    \new_[73192]_ , \new_[73195]_ , \new_[73196]_ , \new_[73197]_ ,
    \new_[73201]_ , \new_[73202]_ , \new_[73205]_ , \new_[73208]_ ,
    \new_[73209]_ , \new_[73210]_ , \new_[73214]_ , \new_[73215]_ ,
    \new_[73218]_ , \new_[73221]_ , \new_[73222]_ , \new_[73223]_ ,
    \new_[73227]_ , \new_[73228]_ , \new_[73231]_ , \new_[73234]_ ,
    \new_[73235]_ , \new_[73236]_ , \new_[73240]_ , \new_[73241]_ ,
    \new_[73244]_ , \new_[73247]_ , \new_[73248]_ , \new_[73249]_ ,
    \new_[73253]_ , \new_[73254]_ , \new_[73257]_ , \new_[73260]_ ,
    \new_[73261]_ , \new_[73262]_ , \new_[73266]_ , \new_[73267]_ ,
    \new_[73270]_ , \new_[73273]_ , \new_[73274]_ , \new_[73275]_ ,
    \new_[73279]_ , \new_[73280]_ , \new_[73283]_ , \new_[73286]_ ,
    \new_[73287]_ , \new_[73288]_ , \new_[73292]_ , \new_[73293]_ ,
    \new_[73296]_ , \new_[73299]_ , \new_[73300]_ , \new_[73301]_ ,
    \new_[73305]_ , \new_[73306]_ , \new_[73309]_ , \new_[73312]_ ,
    \new_[73313]_ , \new_[73314]_ , \new_[73318]_ , \new_[73319]_ ,
    \new_[73322]_ , \new_[73325]_ , \new_[73326]_ , \new_[73327]_ ,
    \new_[73331]_ , \new_[73332]_ , \new_[73335]_ , \new_[73338]_ ,
    \new_[73339]_ , \new_[73340]_ , \new_[73344]_ , \new_[73345]_ ,
    \new_[73348]_ , \new_[73351]_ , \new_[73352]_ , \new_[73353]_ ,
    \new_[73357]_ , \new_[73358]_ , \new_[73361]_ , \new_[73364]_ ,
    \new_[73365]_ , \new_[73366]_ , \new_[73370]_ , \new_[73371]_ ,
    \new_[73374]_ , \new_[73377]_ , \new_[73378]_ , \new_[73379]_ ,
    \new_[73383]_ , \new_[73384]_ , \new_[73387]_ , \new_[73390]_ ,
    \new_[73391]_ , \new_[73392]_ , \new_[73396]_ , \new_[73397]_ ,
    \new_[73400]_ , \new_[73403]_ , \new_[73404]_ , \new_[73405]_ ,
    \new_[73409]_ , \new_[73410]_ , \new_[73413]_ , \new_[73416]_ ,
    \new_[73417]_ , \new_[73418]_ , \new_[73422]_ , \new_[73423]_ ,
    \new_[73426]_ , \new_[73429]_ , \new_[73430]_ , \new_[73431]_ ,
    \new_[73435]_ , \new_[73436]_ , \new_[73439]_ , \new_[73442]_ ,
    \new_[73443]_ , \new_[73444]_ , \new_[73448]_ , \new_[73449]_ ,
    \new_[73452]_ , \new_[73455]_ , \new_[73456]_ , \new_[73457]_ ,
    \new_[73461]_ , \new_[73462]_ , \new_[73465]_ , \new_[73468]_ ,
    \new_[73469]_ , \new_[73470]_ , \new_[73474]_ , \new_[73475]_ ,
    \new_[73478]_ , \new_[73481]_ , \new_[73482]_ , \new_[73483]_ ,
    \new_[73487]_ , \new_[73488]_ , \new_[73491]_ , \new_[73494]_ ,
    \new_[73495]_ , \new_[73496]_ , \new_[73500]_ , \new_[73501]_ ,
    \new_[73504]_ , \new_[73507]_ , \new_[73508]_ , \new_[73509]_ ,
    \new_[73513]_ , \new_[73514]_ , \new_[73517]_ , \new_[73520]_ ,
    \new_[73521]_ , \new_[73522]_ , \new_[73526]_ , \new_[73527]_ ,
    \new_[73530]_ , \new_[73533]_ , \new_[73534]_ , \new_[73535]_ ,
    \new_[73539]_ , \new_[73540]_ , \new_[73543]_ , \new_[73546]_ ,
    \new_[73547]_ , \new_[73548]_ , \new_[73552]_ , \new_[73553]_ ,
    \new_[73556]_ , \new_[73559]_ , \new_[73560]_ , \new_[73561]_ ,
    \new_[73565]_ , \new_[73566]_ , \new_[73569]_ , \new_[73572]_ ,
    \new_[73573]_ , \new_[73574]_ , \new_[73578]_ , \new_[73579]_ ,
    \new_[73582]_ , \new_[73585]_ , \new_[73586]_ , \new_[73587]_ ,
    \new_[73591]_ , \new_[73592]_ , \new_[73595]_ , \new_[73598]_ ,
    \new_[73599]_ , \new_[73600]_ , \new_[73604]_ , \new_[73605]_ ,
    \new_[73608]_ , \new_[73611]_ , \new_[73612]_ , \new_[73613]_ ,
    \new_[73617]_ , \new_[73618]_ , \new_[73621]_ , \new_[73624]_ ,
    \new_[73625]_ , \new_[73626]_ , \new_[73630]_ , \new_[73631]_ ,
    \new_[73634]_ , \new_[73637]_ , \new_[73638]_ , \new_[73639]_ ,
    \new_[73643]_ , \new_[73644]_ , \new_[73647]_ , \new_[73650]_ ,
    \new_[73651]_ , \new_[73652]_ , \new_[73656]_ , \new_[73657]_ ,
    \new_[73660]_ , \new_[73663]_ , \new_[73664]_ , \new_[73665]_ ,
    \new_[73669]_ , \new_[73670]_ , \new_[73673]_ , \new_[73676]_ ,
    \new_[73677]_ , \new_[73678]_ , \new_[73682]_ , \new_[73683]_ ,
    \new_[73686]_ , \new_[73689]_ , \new_[73690]_ , \new_[73691]_ ,
    \new_[73695]_ , \new_[73696]_ , \new_[73699]_ , \new_[73702]_ ,
    \new_[73703]_ , \new_[73704]_ , \new_[73708]_ , \new_[73709]_ ,
    \new_[73712]_ , \new_[73715]_ , \new_[73716]_ , \new_[73717]_ ,
    \new_[73721]_ , \new_[73722]_ , \new_[73725]_ , \new_[73728]_ ,
    \new_[73729]_ , \new_[73730]_ , \new_[73734]_ , \new_[73735]_ ,
    \new_[73738]_ , \new_[73741]_ , \new_[73742]_ , \new_[73743]_ ,
    \new_[73747]_ , \new_[73748]_ , \new_[73751]_ , \new_[73754]_ ,
    \new_[73755]_ , \new_[73756]_ , \new_[73760]_ , \new_[73761]_ ,
    \new_[73764]_ , \new_[73767]_ , \new_[73768]_ , \new_[73769]_ ,
    \new_[73773]_ , \new_[73774]_ , \new_[73777]_ , \new_[73780]_ ,
    \new_[73781]_ , \new_[73782]_ , \new_[73786]_ , \new_[73787]_ ,
    \new_[73790]_ , \new_[73793]_ , \new_[73794]_ , \new_[73795]_ ,
    \new_[73799]_ , \new_[73800]_ , \new_[73803]_ , \new_[73806]_ ,
    \new_[73807]_ , \new_[73808]_ , \new_[73812]_ , \new_[73813]_ ,
    \new_[73816]_ , \new_[73819]_ , \new_[73820]_ , \new_[73821]_ ,
    \new_[73825]_ , \new_[73826]_ , \new_[73829]_ , \new_[73832]_ ,
    \new_[73833]_ , \new_[73834]_ , \new_[73838]_ , \new_[73839]_ ,
    \new_[73842]_ , \new_[73845]_ , \new_[73846]_ , \new_[73847]_ ,
    \new_[73851]_ , \new_[73852]_ , \new_[73855]_ , \new_[73858]_ ,
    \new_[73859]_ , \new_[73860]_ , \new_[73864]_ , \new_[73865]_ ,
    \new_[73868]_ , \new_[73871]_ , \new_[73872]_ , \new_[73873]_ ,
    \new_[73877]_ , \new_[73878]_ , \new_[73881]_ , \new_[73884]_ ,
    \new_[73885]_ , \new_[73886]_ , \new_[73890]_ , \new_[73891]_ ,
    \new_[73894]_ , \new_[73897]_ , \new_[73898]_ , \new_[73899]_ ,
    \new_[73903]_ , \new_[73904]_ , \new_[73907]_ , \new_[73910]_ ,
    \new_[73911]_ , \new_[73912]_ , \new_[73916]_ , \new_[73917]_ ,
    \new_[73920]_ , \new_[73923]_ , \new_[73924]_ , \new_[73925]_ ,
    \new_[73929]_ , \new_[73930]_ , \new_[73933]_ , \new_[73936]_ ,
    \new_[73937]_ , \new_[73938]_ , \new_[73942]_ , \new_[73943]_ ,
    \new_[73946]_ , \new_[73949]_ , \new_[73950]_ , \new_[73951]_ ,
    \new_[73955]_ , \new_[73956]_ , \new_[73959]_ , \new_[73962]_ ,
    \new_[73963]_ , \new_[73964]_ , \new_[73968]_ , \new_[73969]_ ,
    \new_[73972]_ , \new_[73975]_ , \new_[73976]_ , \new_[73977]_ ,
    \new_[73981]_ , \new_[73982]_ , \new_[73985]_ , \new_[73988]_ ,
    \new_[73989]_ , \new_[73990]_ , \new_[73994]_ , \new_[73995]_ ,
    \new_[73998]_ , \new_[74001]_ , \new_[74002]_ , \new_[74003]_ ,
    \new_[74007]_ , \new_[74008]_ , \new_[74011]_ , \new_[74014]_ ,
    \new_[74015]_ , \new_[74016]_ , \new_[74020]_ , \new_[74021]_ ,
    \new_[74024]_ , \new_[74027]_ , \new_[74028]_ , \new_[74029]_ ,
    \new_[74033]_ , \new_[74034]_ , \new_[74037]_ , \new_[74040]_ ,
    \new_[74041]_ , \new_[74042]_ , \new_[74046]_ , \new_[74047]_ ,
    \new_[74050]_ , \new_[74053]_ , \new_[74054]_ , \new_[74055]_ ,
    \new_[74059]_ , \new_[74060]_ , \new_[74063]_ , \new_[74066]_ ,
    \new_[74067]_ , \new_[74068]_ , \new_[74072]_ , \new_[74073]_ ,
    \new_[74076]_ , \new_[74079]_ , \new_[74080]_ , \new_[74081]_ ,
    \new_[74085]_ , \new_[74086]_ , \new_[74089]_ , \new_[74092]_ ,
    \new_[74093]_ , \new_[74094]_ , \new_[74098]_ , \new_[74099]_ ,
    \new_[74102]_ , \new_[74105]_ , \new_[74106]_ , \new_[74107]_ ,
    \new_[74111]_ , \new_[74112]_ , \new_[74115]_ , \new_[74118]_ ,
    \new_[74119]_ , \new_[74120]_ , \new_[74124]_ , \new_[74125]_ ,
    \new_[74128]_ , \new_[74131]_ , \new_[74132]_ , \new_[74133]_ ,
    \new_[74137]_ , \new_[74138]_ , \new_[74141]_ , \new_[74144]_ ,
    \new_[74145]_ , \new_[74146]_ , \new_[74150]_ , \new_[74151]_ ,
    \new_[74154]_ , \new_[74157]_ , \new_[74158]_ , \new_[74159]_ ,
    \new_[74163]_ , \new_[74164]_ , \new_[74167]_ , \new_[74170]_ ,
    \new_[74171]_ , \new_[74172]_ , \new_[74176]_ , \new_[74177]_ ,
    \new_[74180]_ , \new_[74183]_ , \new_[74184]_ , \new_[74185]_ ,
    \new_[74189]_ , \new_[74190]_ , \new_[74193]_ , \new_[74196]_ ,
    \new_[74197]_ , \new_[74198]_ , \new_[74202]_ , \new_[74203]_ ,
    \new_[74206]_ , \new_[74209]_ , \new_[74210]_ , \new_[74211]_ ,
    \new_[74215]_ , \new_[74216]_ , \new_[74219]_ , \new_[74222]_ ,
    \new_[74223]_ , \new_[74224]_ , \new_[74228]_ , \new_[74229]_ ,
    \new_[74232]_ , \new_[74235]_ , \new_[74236]_ , \new_[74237]_ ,
    \new_[74241]_ , \new_[74242]_ , \new_[74245]_ , \new_[74248]_ ,
    \new_[74249]_ , \new_[74250]_ , \new_[74254]_ , \new_[74255]_ ,
    \new_[74258]_ , \new_[74261]_ , \new_[74262]_ , \new_[74263]_ ,
    \new_[74267]_ , \new_[74268]_ , \new_[74271]_ , \new_[74274]_ ,
    \new_[74275]_ , \new_[74276]_ , \new_[74280]_ , \new_[74281]_ ,
    \new_[74284]_ , \new_[74287]_ , \new_[74288]_ , \new_[74289]_ ,
    \new_[74292]_ , \new_[74295]_ , \new_[74296]_ , \new_[74299]_ ,
    \new_[74302]_ , \new_[74303]_ , \new_[74304]_ , \new_[74308]_ ,
    \new_[74309]_ , \new_[74312]_ , \new_[74315]_ , \new_[74316]_ ,
    \new_[74317]_ , \new_[74320]_ , \new_[74323]_ , \new_[74324]_ ,
    \new_[74327]_ , \new_[74330]_ , \new_[74331]_ , \new_[74332]_ ,
    \new_[74336]_ , \new_[74337]_ , \new_[74340]_ , \new_[74343]_ ,
    \new_[74344]_ , \new_[74345]_ , \new_[74348]_ , \new_[74351]_ ,
    \new_[74352]_ , \new_[74355]_ , \new_[74358]_ , \new_[74359]_ ,
    \new_[74360]_ , \new_[74364]_ , \new_[74365]_ , \new_[74368]_ ,
    \new_[74371]_ , \new_[74372]_ , \new_[74373]_ , \new_[74376]_ ,
    \new_[74379]_ , \new_[74380]_ , \new_[74383]_ , \new_[74386]_ ,
    \new_[74387]_ , \new_[74388]_ , \new_[74392]_ , \new_[74393]_ ,
    \new_[74396]_ , \new_[74399]_ , \new_[74400]_ , \new_[74401]_ ,
    \new_[74404]_ , \new_[74407]_ , \new_[74408]_ , \new_[74411]_ ,
    \new_[74414]_ , \new_[74415]_ , \new_[74416]_ , \new_[74420]_ ,
    \new_[74421]_ , \new_[74424]_ , \new_[74427]_ , \new_[74428]_ ,
    \new_[74429]_ , \new_[74432]_ , \new_[74435]_ , \new_[74436]_ ,
    \new_[74439]_ , \new_[74442]_ , \new_[74443]_ , \new_[74444]_ ,
    \new_[74448]_ , \new_[74449]_ , \new_[74452]_ , \new_[74455]_ ,
    \new_[74456]_ , \new_[74457]_ , \new_[74460]_ , \new_[74463]_ ,
    \new_[74464]_ , \new_[74467]_ , \new_[74470]_ , \new_[74471]_ ,
    \new_[74472]_ , \new_[74476]_ , \new_[74477]_ , \new_[74480]_ ,
    \new_[74483]_ , \new_[74484]_ , \new_[74485]_ , \new_[74488]_ ,
    \new_[74491]_ , \new_[74492]_ , \new_[74495]_ , \new_[74498]_ ,
    \new_[74499]_ , \new_[74500]_ , \new_[74504]_ , \new_[74505]_ ,
    \new_[74508]_ , \new_[74511]_ , \new_[74512]_ , \new_[74513]_ ,
    \new_[74516]_ , \new_[74519]_ , \new_[74520]_ , \new_[74523]_ ,
    \new_[74526]_ , \new_[74527]_ , \new_[74528]_ , \new_[74532]_ ,
    \new_[74533]_ , \new_[74536]_ , \new_[74539]_ , \new_[74540]_ ,
    \new_[74541]_ , \new_[74544]_ , \new_[74547]_ , \new_[74548]_ ,
    \new_[74551]_ , \new_[74554]_ , \new_[74555]_ , \new_[74556]_ ,
    \new_[74560]_ , \new_[74561]_ , \new_[74564]_ , \new_[74567]_ ,
    \new_[74568]_ , \new_[74569]_ , \new_[74572]_ , \new_[74575]_ ,
    \new_[74576]_ , \new_[74579]_ , \new_[74582]_ , \new_[74583]_ ,
    \new_[74584]_ , \new_[74588]_ , \new_[74589]_ , \new_[74592]_ ,
    \new_[74595]_ , \new_[74596]_ , \new_[74597]_ , \new_[74600]_ ,
    \new_[74603]_ , \new_[74604]_ , \new_[74607]_ , \new_[74610]_ ,
    \new_[74611]_ , \new_[74612]_ , \new_[74616]_ , \new_[74617]_ ,
    \new_[74620]_ , \new_[74623]_ , \new_[74624]_ , \new_[74625]_ ,
    \new_[74628]_ , \new_[74631]_ , \new_[74632]_ , \new_[74635]_ ,
    \new_[74638]_ , \new_[74639]_ , \new_[74640]_ , \new_[74644]_ ,
    \new_[74645]_ , \new_[74648]_ , \new_[74651]_ , \new_[74652]_ ,
    \new_[74653]_ , \new_[74656]_ , \new_[74659]_ , \new_[74660]_ ,
    \new_[74663]_ , \new_[74666]_ , \new_[74667]_ , \new_[74668]_ ,
    \new_[74672]_ , \new_[74673]_ , \new_[74676]_ , \new_[74679]_ ,
    \new_[74680]_ , \new_[74681]_ , \new_[74684]_ , \new_[74687]_ ,
    \new_[74688]_ , \new_[74691]_ , \new_[74694]_ , \new_[74695]_ ,
    \new_[74696]_ , \new_[74700]_ , \new_[74701]_ , \new_[74704]_ ,
    \new_[74707]_ , \new_[74708]_ , \new_[74709]_ , \new_[74712]_ ,
    \new_[74715]_ , \new_[74716]_ , \new_[74719]_ , \new_[74722]_ ,
    \new_[74723]_ , \new_[74724]_ , \new_[74728]_ , \new_[74729]_ ,
    \new_[74732]_ , \new_[74735]_ , \new_[74736]_ , \new_[74737]_ ,
    \new_[74740]_ , \new_[74743]_ , \new_[74744]_ , \new_[74747]_ ,
    \new_[74750]_ , \new_[74751]_ , \new_[74752]_ , \new_[74756]_ ,
    \new_[74757]_ , \new_[74760]_ , \new_[74763]_ , \new_[74764]_ ,
    \new_[74765]_ , \new_[74768]_ , \new_[74771]_ , \new_[74772]_ ,
    \new_[74775]_ , \new_[74778]_ , \new_[74779]_ , \new_[74780]_ ,
    \new_[74784]_ , \new_[74785]_ , \new_[74788]_ , \new_[74791]_ ,
    \new_[74792]_ , \new_[74793]_ , \new_[74796]_ , \new_[74799]_ ,
    \new_[74800]_ , \new_[74803]_ , \new_[74806]_ , \new_[74807]_ ,
    \new_[74808]_ , \new_[74812]_ , \new_[74813]_ , \new_[74816]_ ,
    \new_[74819]_ , \new_[74820]_ , \new_[74821]_ , \new_[74824]_ ,
    \new_[74827]_ , \new_[74828]_ , \new_[74831]_ , \new_[74834]_ ,
    \new_[74835]_ , \new_[74836]_ , \new_[74840]_ , \new_[74841]_ ,
    \new_[74844]_ , \new_[74847]_ , \new_[74848]_ , \new_[74849]_ ,
    \new_[74852]_ , \new_[74855]_ , \new_[74856]_ , \new_[74859]_ ,
    \new_[74862]_ , \new_[74863]_ , \new_[74864]_ , \new_[74868]_ ,
    \new_[74869]_ , \new_[74872]_ , \new_[74875]_ , \new_[74876]_ ,
    \new_[74877]_ , \new_[74880]_ , \new_[74883]_ , \new_[74884]_ ,
    \new_[74887]_ , \new_[74890]_ , \new_[74891]_ , \new_[74892]_ ,
    \new_[74896]_ , \new_[74897]_ , \new_[74900]_ , \new_[74903]_ ,
    \new_[74904]_ , \new_[74905]_ , \new_[74908]_ , \new_[74911]_ ,
    \new_[74912]_ , \new_[74915]_ , \new_[74918]_ , \new_[74919]_ ,
    \new_[74920]_ , \new_[74924]_ , \new_[74925]_ , \new_[74928]_ ,
    \new_[74931]_ , \new_[74932]_ , \new_[74933]_ , \new_[74936]_ ,
    \new_[74939]_ , \new_[74940]_ , \new_[74943]_ , \new_[74946]_ ,
    \new_[74947]_ , \new_[74948]_ , \new_[74952]_ , \new_[74953]_ ,
    \new_[74956]_ , \new_[74959]_ , \new_[74960]_ , \new_[74961]_ ,
    \new_[74964]_ , \new_[74967]_ , \new_[74968]_ , \new_[74971]_ ,
    \new_[74974]_ , \new_[74975]_ , \new_[74976]_ , \new_[74980]_ ,
    \new_[74981]_ , \new_[74984]_ , \new_[74987]_ , \new_[74988]_ ,
    \new_[74989]_ , \new_[74992]_ , \new_[74995]_ , \new_[74996]_ ,
    \new_[74999]_ , \new_[75002]_ , \new_[75003]_ , \new_[75004]_ ,
    \new_[75008]_ , \new_[75009]_ , \new_[75012]_ , \new_[75015]_ ,
    \new_[75016]_ , \new_[75017]_ , \new_[75020]_ , \new_[75023]_ ,
    \new_[75024]_ , \new_[75027]_ , \new_[75030]_ , \new_[75031]_ ,
    \new_[75032]_ , \new_[75036]_ , \new_[75037]_ , \new_[75040]_ ,
    \new_[75043]_ , \new_[75044]_ , \new_[75045]_ , \new_[75048]_ ,
    \new_[75051]_ , \new_[75052]_ , \new_[75055]_ , \new_[75058]_ ,
    \new_[75059]_ , \new_[75060]_ , \new_[75064]_ , \new_[75065]_ ,
    \new_[75068]_ , \new_[75071]_ , \new_[75072]_ , \new_[75073]_ ,
    \new_[75076]_ , \new_[75079]_ , \new_[75080]_ , \new_[75083]_ ,
    \new_[75086]_ , \new_[75087]_ , \new_[75088]_ , \new_[75092]_ ,
    \new_[75093]_ , \new_[75096]_ , \new_[75099]_ , \new_[75100]_ ,
    \new_[75101]_ , \new_[75104]_ , \new_[75107]_ , \new_[75108]_ ,
    \new_[75111]_ , \new_[75114]_ , \new_[75115]_ , \new_[75116]_ ,
    \new_[75120]_ , \new_[75121]_ , \new_[75124]_ , \new_[75127]_ ,
    \new_[75128]_ , \new_[75129]_ , \new_[75132]_ , \new_[75135]_ ,
    \new_[75136]_ , \new_[75139]_ , \new_[75142]_ , \new_[75143]_ ,
    \new_[75144]_ , \new_[75148]_ , \new_[75149]_ , \new_[75152]_ ,
    \new_[75155]_ , \new_[75156]_ , \new_[75157]_ , \new_[75160]_ ,
    \new_[75163]_ , \new_[75164]_ , \new_[75167]_ , \new_[75170]_ ,
    \new_[75171]_ , \new_[75172]_ , \new_[75176]_ , \new_[75177]_ ,
    \new_[75180]_ , \new_[75183]_ , \new_[75184]_ , \new_[75185]_ ,
    \new_[75188]_ , \new_[75191]_ , \new_[75192]_ , \new_[75195]_ ,
    \new_[75198]_ , \new_[75199]_ , \new_[75200]_ , \new_[75204]_ ,
    \new_[75205]_ , \new_[75208]_ , \new_[75211]_ , \new_[75212]_ ,
    \new_[75213]_ , \new_[75216]_ , \new_[75219]_ , \new_[75220]_ ,
    \new_[75223]_ , \new_[75226]_ , \new_[75227]_ , \new_[75228]_ ,
    \new_[75232]_ , \new_[75233]_ , \new_[75236]_ , \new_[75239]_ ,
    \new_[75240]_ , \new_[75241]_ , \new_[75244]_ , \new_[75247]_ ,
    \new_[75248]_ , \new_[75251]_ , \new_[75254]_ , \new_[75255]_ ,
    \new_[75256]_ , \new_[75260]_ , \new_[75261]_ , \new_[75264]_ ,
    \new_[75267]_ , \new_[75268]_ , \new_[75269]_ , \new_[75272]_ ,
    \new_[75275]_ , \new_[75276]_ , \new_[75279]_ , \new_[75282]_ ,
    \new_[75283]_ , \new_[75284]_ , \new_[75288]_ , \new_[75289]_ ,
    \new_[75292]_ , \new_[75295]_ , \new_[75296]_ , \new_[75297]_ ,
    \new_[75300]_ , \new_[75303]_ , \new_[75304]_ , \new_[75307]_ ,
    \new_[75310]_ , \new_[75311]_ , \new_[75312]_ , \new_[75316]_ ,
    \new_[75317]_ , \new_[75320]_ , \new_[75323]_ , \new_[75324]_ ,
    \new_[75325]_ , \new_[75328]_ , \new_[75331]_ , \new_[75332]_ ,
    \new_[75335]_ , \new_[75338]_ , \new_[75339]_ , \new_[75340]_ ,
    \new_[75344]_ , \new_[75345]_ , \new_[75348]_ , \new_[75351]_ ,
    \new_[75352]_ , \new_[75353]_ , \new_[75356]_ , \new_[75359]_ ,
    \new_[75360]_ , \new_[75363]_ , \new_[75366]_ , \new_[75367]_ ,
    \new_[75368]_ , \new_[75372]_ , \new_[75373]_ , \new_[75376]_ ,
    \new_[75379]_ , \new_[75380]_ , \new_[75381]_ , \new_[75384]_ ,
    \new_[75387]_ , \new_[75388]_ , \new_[75391]_ , \new_[75394]_ ,
    \new_[75395]_ , \new_[75396]_ , \new_[75400]_ , \new_[75401]_ ,
    \new_[75404]_ , \new_[75407]_ , \new_[75408]_ , \new_[75409]_ ,
    \new_[75412]_ , \new_[75415]_ , \new_[75416]_ , \new_[75419]_ ,
    \new_[75422]_ , \new_[75423]_ , \new_[75424]_ , \new_[75428]_ ,
    \new_[75429]_ , \new_[75432]_ , \new_[75435]_ , \new_[75436]_ ,
    \new_[75437]_ , \new_[75440]_ , \new_[75443]_ , \new_[75444]_ ,
    \new_[75447]_ , \new_[75450]_ , \new_[75451]_ , \new_[75452]_ ,
    \new_[75456]_ , \new_[75457]_ , \new_[75460]_ , \new_[75463]_ ,
    \new_[75464]_ , \new_[75465]_ , \new_[75468]_ , \new_[75471]_ ,
    \new_[75472]_ , \new_[75475]_ , \new_[75478]_ , \new_[75479]_ ,
    \new_[75480]_ , \new_[75484]_ , \new_[75485]_ , \new_[75488]_ ,
    \new_[75491]_ , \new_[75492]_ , \new_[75493]_ , \new_[75496]_ ,
    \new_[75499]_ , \new_[75500]_ , \new_[75503]_ , \new_[75506]_ ,
    \new_[75507]_ , \new_[75508]_ , \new_[75512]_ , \new_[75513]_ ,
    \new_[75516]_ , \new_[75519]_ , \new_[75520]_ , \new_[75521]_ ,
    \new_[75524]_ , \new_[75527]_ , \new_[75528]_ , \new_[75531]_ ,
    \new_[75534]_ , \new_[75535]_ , \new_[75536]_ , \new_[75540]_ ,
    \new_[75541]_ , \new_[75544]_ , \new_[75547]_ , \new_[75548]_ ,
    \new_[75549]_ , \new_[75552]_ , \new_[75555]_ , \new_[75556]_ ,
    \new_[75559]_ , \new_[75562]_ , \new_[75563]_ , \new_[75564]_ ,
    \new_[75568]_ , \new_[75569]_ , \new_[75572]_ , \new_[75575]_ ,
    \new_[75576]_ , \new_[75577]_ , \new_[75580]_ , \new_[75583]_ ,
    \new_[75584]_ , \new_[75587]_ , \new_[75590]_ , \new_[75591]_ ,
    \new_[75592]_ , \new_[75596]_ , \new_[75597]_ , \new_[75600]_ ,
    \new_[75603]_ , \new_[75604]_ , \new_[75605]_ , \new_[75608]_ ,
    \new_[75611]_ , \new_[75612]_ , \new_[75615]_ , \new_[75618]_ ,
    \new_[75619]_ , \new_[75620]_ , \new_[75624]_ , \new_[75625]_ ,
    \new_[75628]_ , \new_[75631]_ , \new_[75632]_ , \new_[75633]_ ,
    \new_[75636]_ , \new_[75639]_ , \new_[75640]_ , \new_[75643]_ ,
    \new_[75646]_ , \new_[75647]_ , \new_[75648]_ , \new_[75652]_ ,
    \new_[75653]_ , \new_[75656]_ , \new_[75659]_ , \new_[75660]_ ,
    \new_[75661]_ , \new_[75664]_ , \new_[75667]_ , \new_[75668]_ ,
    \new_[75671]_ , \new_[75674]_ , \new_[75675]_ , \new_[75676]_ ,
    \new_[75680]_ , \new_[75681]_ , \new_[75684]_ , \new_[75687]_ ,
    \new_[75688]_ , \new_[75689]_ , \new_[75692]_ , \new_[75695]_ ,
    \new_[75696]_ , \new_[75699]_ , \new_[75702]_ , \new_[75703]_ ,
    \new_[75704]_ , \new_[75708]_ , \new_[75709]_ , \new_[75712]_ ,
    \new_[75715]_ , \new_[75716]_ , \new_[75717]_ , \new_[75720]_ ,
    \new_[75723]_ , \new_[75724]_ , \new_[75727]_ , \new_[75730]_ ,
    \new_[75731]_ , \new_[75732]_ , \new_[75736]_ , \new_[75737]_ ,
    \new_[75740]_ , \new_[75743]_ , \new_[75744]_ , \new_[75745]_ ,
    \new_[75748]_ , \new_[75751]_ , \new_[75752]_ , \new_[75755]_ ,
    \new_[75758]_ , \new_[75759]_ , \new_[75760]_ , \new_[75764]_ ,
    \new_[75765]_ , \new_[75768]_ , \new_[75771]_ , \new_[75772]_ ,
    \new_[75773]_ , \new_[75776]_ , \new_[75779]_ , \new_[75780]_ ,
    \new_[75783]_ , \new_[75786]_ , \new_[75787]_ , \new_[75788]_ ,
    \new_[75792]_ , \new_[75793]_ , \new_[75796]_ , \new_[75799]_ ,
    \new_[75800]_ , \new_[75801]_ , \new_[75804]_ , \new_[75807]_ ,
    \new_[75808]_ , \new_[75811]_ , \new_[75814]_ , \new_[75815]_ ,
    \new_[75816]_ , \new_[75820]_ , \new_[75821]_ , \new_[75824]_ ,
    \new_[75827]_ , \new_[75828]_ , \new_[75829]_ , \new_[75832]_ ,
    \new_[75835]_ , \new_[75836]_ , \new_[75839]_ , \new_[75842]_ ,
    \new_[75843]_ , \new_[75844]_ , \new_[75848]_ , \new_[75849]_ ,
    \new_[75852]_ , \new_[75855]_ , \new_[75856]_ , \new_[75857]_ ,
    \new_[75860]_ , \new_[75863]_ , \new_[75864]_ , \new_[75867]_ ,
    \new_[75870]_ , \new_[75871]_ , \new_[75872]_ , \new_[75876]_ ,
    \new_[75877]_ , \new_[75880]_ , \new_[75883]_ , \new_[75884]_ ,
    \new_[75885]_ , \new_[75888]_ , \new_[75891]_ , \new_[75892]_ ,
    \new_[75895]_ , \new_[75898]_ , \new_[75899]_ , \new_[75900]_ ,
    \new_[75904]_ , \new_[75905]_ , \new_[75908]_ , \new_[75911]_ ,
    \new_[75912]_ , \new_[75913]_ , \new_[75916]_ , \new_[75919]_ ,
    \new_[75920]_ , \new_[75923]_ , \new_[75926]_ , \new_[75927]_ ,
    \new_[75928]_ , \new_[75932]_ , \new_[75933]_ , \new_[75936]_ ,
    \new_[75939]_ , \new_[75940]_ , \new_[75941]_ , \new_[75944]_ ,
    \new_[75947]_ , \new_[75948]_ , \new_[75951]_ , \new_[75954]_ ,
    \new_[75955]_ , \new_[75956]_ , \new_[75960]_ , \new_[75961]_ ,
    \new_[75964]_ , \new_[75967]_ , \new_[75968]_ , \new_[75969]_ ,
    \new_[75972]_ , \new_[75975]_ , \new_[75976]_ , \new_[75979]_ ,
    \new_[75982]_ , \new_[75983]_ , \new_[75984]_ , \new_[75988]_ ,
    \new_[75989]_ , \new_[75992]_ , \new_[75995]_ , \new_[75996]_ ,
    \new_[75997]_ , \new_[76000]_ , \new_[76003]_ , \new_[76004]_ ,
    \new_[76007]_ , \new_[76010]_ , \new_[76011]_ , \new_[76012]_ ,
    \new_[76016]_ , \new_[76017]_ , \new_[76020]_ , \new_[76023]_ ,
    \new_[76024]_ , \new_[76025]_ , \new_[76028]_ , \new_[76031]_ ,
    \new_[76032]_ , \new_[76035]_ , \new_[76038]_ , \new_[76039]_ ,
    \new_[76040]_ , \new_[76044]_ , \new_[76045]_ , \new_[76048]_ ,
    \new_[76051]_ , \new_[76052]_ , \new_[76053]_ , \new_[76056]_ ,
    \new_[76059]_ , \new_[76060]_ , \new_[76063]_ , \new_[76066]_ ,
    \new_[76067]_ , \new_[76068]_ , \new_[76072]_ , \new_[76073]_ ,
    \new_[76076]_ , \new_[76079]_ , \new_[76080]_ , \new_[76081]_ ,
    \new_[76084]_ , \new_[76087]_ , \new_[76088]_ , \new_[76091]_ ,
    \new_[76094]_ , \new_[76095]_ , \new_[76096]_ , \new_[76100]_ ,
    \new_[76101]_ , \new_[76104]_ , \new_[76107]_ , \new_[76108]_ ,
    \new_[76109]_ , \new_[76112]_ , \new_[76115]_ , \new_[76116]_ ,
    \new_[76119]_ , \new_[76122]_ , \new_[76123]_ , \new_[76124]_ ,
    \new_[76128]_ , \new_[76129]_ , \new_[76132]_ , \new_[76135]_ ,
    \new_[76136]_ , \new_[76137]_ , \new_[76140]_ , \new_[76143]_ ,
    \new_[76144]_ , \new_[76147]_ , \new_[76150]_ , \new_[76151]_ ,
    \new_[76152]_ , \new_[76156]_ , \new_[76157]_ , \new_[76160]_ ,
    \new_[76163]_ , \new_[76164]_ , \new_[76165]_ , \new_[76168]_ ,
    \new_[76171]_ , \new_[76172]_ , \new_[76175]_ , \new_[76178]_ ,
    \new_[76179]_ , \new_[76180]_ , \new_[76184]_ , \new_[76185]_ ,
    \new_[76188]_ , \new_[76191]_ , \new_[76192]_ , \new_[76193]_ ,
    \new_[76196]_ , \new_[76199]_ , \new_[76200]_ , \new_[76203]_ ,
    \new_[76206]_ , \new_[76207]_ , \new_[76208]_ , \new_[76212]_ ,
    \new_[76213]_ , \new_[76216]_ , \new_[76219]_ , \new_[76220]_ ,
    \new_[76221]_ , \new_[76224]_ , \new_[76227]_ , \new_[76228]_ ,
    \new_[76231]_ , \new_[76234]_ , \new_[76235]_ , \new_[76236]_ ,
    \new_[76240]_ , \new_[76241]_ , \new_[76244]_ , \new_[76247]_ ,
    \new_[76248]_ , \new_[76249]_ , \new_[76252]_ , \new_[76255]_ ,
    \new_[76256]_ , \new_[76259]_ , \new_[76262]_ , \new_[76263]_ ,
    \new_[76264]_ , \new_[76268]_ , \new_[76269]_ , \new_[76272]_ ,
    \new_[76275]_ , \new_[76276]_ , \new_[76277]_ , \new_[76280]_ ,
    \new_[76283]_ , \new_[76284]_ , \new_[76287]_ , \new_[76290]_ ,
    \new_[76291]_ , \new_[76292]_ , \new_[76296]_ , \new_[76297]_ ,
    \new_[76300]_ , \new_[76303]_ , \new_[76304]_ , \new_[76305]_ ,
    \new_[76308]_ , \new_[76311]_ , \new_[76312]_ , \new_[76315]_ ,
    \new_[76318]_ , \new_[76319]_ , \new_[76320]_ , \new_[76324]_ ,
    \new_[76325]_ , \new_[76328]_ , \new_[76331]_ , \new_[76332]_ ,
    \new_[76333]_ , \new_[76336]_ , \new_[76339]_ , \new_[76340]_ ,
    \new_[76343]_ , \new_[76346]_ , \new_[76347]_ , \new_[76348]_ ,
    \new_[76352]_ , \new_[76353]_ , \new_[76356]_ , \new_[76359]_ ,
    \new_[76360]_ , \new_[76361]_ , \new_[76364]_ , \new_[76367]_ ,
    \new_[76368]_ , \new_[76371]_ , \new_[76374]_ , \new_[76375]_ ,
    \new_[76376]_ , \new_[76380]_ , \new_[76381]_ , \new_[76384]_ ,
    \new_[76387]_ , \new_[76388]_ , \new_[76389]_ , \new_[76392]_ ,
    \new_[76395]_ , \new_[76396]_ , \new_[76399]_ , \new_[76402]_ ,
    \new_[76403]_ , \new_[76404]_ , \new_[76408]_ , \new_[76409]_ ,
    \new_[76412]_ , \new_[76415]_ , \new_[76416]_ , \new_[76417]_ ,
    \new_[76420]_ , \new_[76423]_ , \new_[76424]_ , \new_[76427]_ ,
    \new_[76430]_ , \new_[76431]_ , \new_[76432]_ , \new_[76436]_ ,
    \new_[76437]_ , \new_[76440]_ , \new_[76443]_ , \new_[76444]_ ,
    \new_[76445]_ , \new_[76448]_ , \new_[76451]_ , \new_[76452]_ ,
    \new_[76455]_ , \new_[76458]_ , \new_[76459]_ , \new_[76460]_ ,
    \new_[76464]_ , \new_[76465]_ , \new_[76468]_ , \new_[76471]_ ,
    \new_[76472]_ , \new_[76473]_ , \new_[76476]_ , \new_[76479]_ ,
    \new_[76480]_ , \new_[76483]_ , \new_[76486]_ , \new_[76487]_ ,
    \new_[76488]_ , \new_[76492]_ , \new_[76493]_ , \new_[76496]_ ,
    \new_[76499]_ , \new_[76500]_ , \new_[76501]_ , \new_[76504]_ ,
    \new_[76507]_ , \new_[76508]_ , \new_[76511]_ , \new_[76514]_ ,
    \new_[76515]_ , \new_[76516]_ , \new_[76520]_ , \new_[76521]_ ,
    \new_[76524]_ , \new_[76527]_ , \new_[76528]_ , \new_[76529]_ ,
    \new_[76532]_ , \new_[76535]_ , \new_[76536]_ , \new_[76539]_ ,
    \new_[76542]_ , \new_[76543]_ , \new_[76544]_ , \new_[76548]_ ,
    \new_[76549]_ , \new_[76552]_ , \new_[76555]_ , \new_[76556]_ ,
    \new_[76557]_ , \new_[76560]_ , \new_[76563]_ , \new_[76564]_ ,
    \new_[76567]_ , \new_[76570]_ , \new_[76571]_ , \new_[76572]_ ,
    \new_[76576]_ , \new_[76577]_ , \new_[76580]_ , \new_[76583]_ ,
    \new_[76584]_ , \new_[76585]_ , \new_[76588]_ , \new_[76591]_ ,
    \new_[76592]_ , \new_[76595]_ , \new_[76598]_ , \new_[76599]_ ,
    \new_[76600]_ , \new_[76604]_ , \new_[76605]_ , \new_[76608]_ ,
    \new_[76611]_ , \new_[76612]_ , \new_[76613]_ , \new_[76616]_ ,
    \new_[76619]_ , \new_[76620]_ , \new_[76623]_ , \new_[76626]_ ,
    \new_[76627]_ , \new_[76628]_ , \new_[76632]_ , \new_[76633]_ ,
    \new_[76636]_ , \new_[76639]_ , \new_[76640]_ , \new_[76641]_ ,
    \new_[76644]_ , \new_[76647]_ , \new_[76648]_ , \new_[76651]_ ,
    \new_[76654]_ , \new_[76655]_ , \new_[76656]_ , \new_[76660]_ ,
    \new_[76661]_ , \new_[76664]_ , \new_[76667]_ , \new_[76668]_ ,
    \new_[76669]_ , \new_[76672]_ , \new_[76675]_ , \new_[76676]_ ,
    \new_[76679]_ , \new_[76682]_ , \new_[76683]_ , \new_[76684]_ ,
    \new_[76688]_ , \new_[76689]_ , \new_[76692]_ , \new_[76695]_ ,
    \new_[76696]_ , \new_[76697]_ , \new_[76700]_ , \new_[76703]_ ,
    \new_[76704]_ , \new_[76707]_ , \new_[76710]_ , \new_[76711]_ ,
    \new_[76712]_ , \new_[76716]_ , \new_[76717]_ , \new_[76720]_ ,
    \new_[76723]_ , \new_[76724]_ , \new_[76725]_ , \new_[76728]_ ,
    \new_[76731]_ , \new_[76732]_ , \new_[76735]_ , \new_[76738]_ ,
    \new_[76739]_ , \new_[76740]_ , \new_[76744]_ , \new_[76745]_ ,
    \new_[76748]_ , \new_[76751]_ , \new_[76752]_ , \new_[76753]_ ,
    \new_[76756]_ , \new_[76759]_ , \new_[76760]_ , \new_[76763]_ ,
    \new_[76766]_ , \new_[76767]_ , \new_[76768]_ , \new_[76772]_ ,
    \new_[76773]_ , \new_[76776]_ , \new_[76779]_ , \new_[76780]_ ,
    \new_[76781]_ , \new_[76784]_ , \new_[76787]_ , \new_[76788]_ ,
    \new_[76791]_ , \new_[76794]_ , \new_[76795]_ , \new_[76796]_ ,
    \new_[76800]_ , \new_[76801]_ , \new_[76804]_ , \new_[76807]_ ,
    \new_[76808]_ , \new_[76809]_ , \new_[76812]_ , \new_[76815]_ ,
    \new_[76816]_ , \new_[76819]_ , \new_[76822]_ , \new_[76823]_ ,
    \new_[76824]_ , \new_[76828]_ , \new_[76829]_ , \new_[76832]_ ,
    \new_[76835]_ , \new_[76836]_ , \new_[76837]_ , \new_[76840]_ ,
    \new_[76843]_ , \new_[76844]_ , \new_[76847]_ , \new_[76850]_ ,
    \new_[76851]_ , \new_[76852]_ , \new_[76856]_ , \new_[76857]_ ,
    \new_[76860]_ , \new_[76863]_ , \new_[76864]_ , \new_[76865]_ ,
    \new_[76868]_ , \new_[76871]_ , \new_[76872]_ , \new_[76875]_ ,
    \new_[76878]_ , \new_[76879]_ , \new_[76880]_ , \new_[76884]_ ,
    \new_[76885]_ , \new_[76888]_ , \new_[76891]_ , \new_[76892]_ ,
    \new_[76893]_ , \new_[76896]_ , \new_[76899]_ , \new_[76900]_ ,
    \new_[76903]_ , \new_[76906]_ , \new_[76907]_ , \new_[76908]_ ,
    \new_[76912]_ , \new_[76913]_ , \new_[76916]_ , \new_[76919]_ ,
    \new_[76920]_ , \new_[76921]_ , \new_[76924]_ , \new_[76927]_ ,
    \new_[76928]_ , \new_[76931]_ , \new_[76934]_ , \new_[76935]_ ,
    \new_[76936]_ , \new_[76940]_ , \new_[76941]_ , \new_[76944]_ ,
    \new_[76947]_ , \new_[76948]_ , \new_[76949]_ , \new_[76952]_ ,
    \new_[76955]_ , \new_[76956]_ , \new_[76959]_ , \new_[76962]_ ,
    \new_[76963]_ , \new_[76964]_ , \new_[76968]_ , \new_[76969]_ ,
    \new_[76972]_ , \new_[76975]_ , \new_[76976]_ , \new_[76977]_ ,
    \new_[76980]_ , \new_[76983]_ , \new_[76984]_ , \new_[76987]_ ,
    \new_[76990]_ , \new_[76991]_ , \new_[76992]_ , \new_[76996]_ ,
    \new_[76997]_ , \new_[77000]_ , \new_[77003]_ , \new_[77004]_ ,
    \new_[77005]_ , \new_[77008]_ , \new_[77011]_ , \new_[77012]_ ,
    \new_[77015]_ , \new_[77018]_ , \new_[77019]_ , \new_[77020]_ ,
    \new_[77024]_ , \new_[77025]_ , \new_[77028]_ , \new_[77031]_ ,
    \new_[77032]_ , \new_[77033]_ , \new_[77036]_ , \new_[77039]_ ,
    \new_[77040]_ , \new_[77043]_ , \new_[77046]_ , \new_[77047]_ ,
    \new_[77048]_ , \new_[77052]_ , \new_[77053]_ , \new_[77056]_ ,
    \new_[77059]_ , \new_[77060]_ , \new_[77061]_ , \new_[77064]_ ,
    \new_[77067]_ , \new_[77068]_ , \new_[77071]_ , \new_[77074]_ ,
    \new_[77075]_ , \new_[77076]_ , \new_[77080]_ , \new_[77081]_ ,
    \new_[77084]_ , \new_[77087]_ , \new_[77088]_ , \new_[77089]_ ,
    \new_[77092]_ , \new_[77095]_ , \new_[77096]_ , \new_[77099]_ ,
    \new_[77102]_ , \new_[77103]_ , \new_[77104]_ , \new_[77108]_ ,
    \new_[77109]_ , \new_[77112]_ , \new_[77115]_ , \new_[77116]_ ,
    \new_[77117]_ , \new_[77120]_ , \new_[77123]_ , \new_[77124]_ ,
    \new_[77127]_ , \new_[77130]_ , \new_[77131]_ , \new_[77132]_ ,
    \new_[77136]_ , \new_[77137]_ , \new_[77140]_ , \new_[77143]_ ,
    \new_[77144]_ , \new_[77145]_ , \new_[77148]_ , \new_[77151]_ ,
    \new_[77152]_ , \new_[77155]_ , \new_[77158]_ , \new_[77159]_ ,
    \new_[77160]_ , \new_[77164]_ , \new_[77165]_ , \new_[77168]_ ,
    \new_[77171]_ , \new_[77172]_ , \new_[77173]_ , \new_[77176]_ ,
    \new_[77179]_ , \new_[77180]_ , \new_[77183]_ , \new_[77186]_ ,
    \new_[77187]_ , \new_[77188]_ , \new_[77192]_ , \new_[77193]_ ,
    \new_[77196]_ , \new_[77199]_ , \new_[77200]_ , \new_[77201]_ ,
    \new_[77204]_ , \new_[77207]_ , \new_[77208]_ , \new_[77211]_ ,
    \new_[77214]_ , \new_[77215]_ , \new_[77216]_ , \new_[77220]_ ,
    \new_[77221]_ , \new_[77224]_ , \new_[77227]_ , \new_[77228]_ ,
    \new_[77229]_ , \new_[77232]_ , \new_[77235]_ , \new_[77236]_ ,
    \new_[77239]_ , \new_[77242]_ , \new_[77243]_ , \new_[77244]_ ,
    \new_[77248]_ , \new_[77249]_ , \new_[77252]_ , \new_[77255]_ ,
    \new_[77256]_ , \new_[77257]_ , \new_[77260]_ , \new_[77263]_ ,
    \new_[77264]_ , \new_[77267]_ , \new_[77270]_ , \new_[77271]_ ,
    \new_[77272]_ , \new_[77276]_ , \new_[77277]_ , \new_[77280]_ ,
    \new_[77283]_ , \new_[77284]_ , \new_[77285]_ , \new_[77288]_ ,
    \new_[77291]_ , \new_[77292]_ , \new_[77295]_ , \new_[77298]_ ,
    \new_[77299]_ , \new_[77300]_ , \new_[77304]_ , \new_[77305]_ ,
    \new_[77308]_ , \new_[77311]_ , \new_[77312]_ , \new_[77313]_ ,
    \new_[77316]_ , \new_[77319]_ , \new_[77320]_ , \new_[77323]_ ,
    \new_[77326]_ , \new_[77327]_ , \new_[77328]_ , \new_[77332]_ ,
    \new_[77333]_ , \new_[77336]_ , \new_[77339]_ , \new_[77340]_ ,
    \new_[77341]_ , \new_[77344]_ , \new_[77347]_ , \new_[77348]_ ,
    \new_[77351]_ , \new_[77354]_ , \new_[77355]_ , \new_[77356]_ ,
    \new_[77360]_ , \new_[77361]_ , \new_[77364]_ , \new_[77367]_ ,
    \new_[77368]_ , \new_[77369]_ , \new_[77372]_ , \new_[77375]_ ,
    \new_[77376]_ , \new_[77379]_ , \new_[77382]_ , \new_[77383]_ ,
    \new_[77384]_ , \new_[77388]_ , \new_[77389]_ , \new_[77392]_ ,
    \new_[77395]_ , \new_[77396]_ , \new_[77397]_ , \new_[77400]_ ,
    \new_[77403]_ , \new_[77404]_ , \new_[77407]_ , \new_[77410]_ ,
    \new_[77411]_ , \new_[77412]_ , \new_[77416]_ , \new_[77417]_ ,
    \new_[77420]_ , \new_[77423]_ , \new_[77424]_ , \new_[77425]_ ,
    \new_[77428]_ , \new_[77431]_ , \new_[77432]_ , \new_[77435]_ ,
    \new_[77438]_ , \new_[77439]_ , \new_[77440]_ , \new_[77444]_ ,
    \new_[77445]_ , \new_[77448]_ , \new_[77451]_ , \new_[77452]_ ,
    \new_[77453]_ , \new_[77456]_ , \new_[77459]_ , \new_[77460]_ ,
    \new_[77463]_ , \new_[77466]_ , \new_[77467]_ , \new_[77468]_ ,
    \new_[77472]_ , \new_[77473]_ , \new_[77476]_ , \new_[77479]_ ,
    \new_[77480]_ , \new_[77481]_ , \new_[77484]_ , \new_[77487]_ ,
    \new_[77488]_ , \new_[77491]_ , \new_[77494]_ , \new_[77495]_ ,
    \new_[77496]_ , \new_[77500]_ , \new_[77501]_ , \new_[77504]_ ,
    \new_[77507]_ , \new_[77508]_ , \new_[77509]_ , \new_[77512]_ ,
    \new_[77515]_ , \new_[77516]_ , \new_[77519]_ , \new_[77522]_ ,
    \new_[77523]_ , \new_[77524]_ , \new_[77528]_ , \new_[77529]_ ,
    \new_[77532]_ , \new_[77535]_ , \new_[77536]_ , \new_[77537]_ ,
    \new_[77540]_ , \new_[77543]_ , \new_[77544]_ , \new_[77547]_ ,
    \new_[77550]_ , \new_[77551]_ , \new_[77552]_ , \new_[77556]_ ,
    \new_[77557]_ , \new_[77560]_ , \new_[77563]_ , \new_[77564]_ ,
    \new_[77565]_ , \new_[77568]_ , \new_[77571]_ , \new_[77572]_ ,
    \new_[77575]_ , \new_[77578]_ , \new_[77579]_ , \new_[77580]_ ,
    \new_[77584]_ , \new_[77585]_ , \new_[77588]_ , \new_[77591]_ ,
    \new_[77592]_ , \new_[77593]_ , \new_[77596]_ , \new_[77599]_ ,
    \new_[77600]_ , \new_[77603]_ , \new_[77606]_ , \new_[77607]_ ,
    \new_[77608]_ , \new_[77612]_ , \new_[77613]_ , \new_[77616]_ ,
    \new_[77619]_ , \new_[77620]_ , \new_[77621]_ , \new_[77624]_ ,
    \new_[77627]_ , \new_[77628]_ , \new_[77631]_ , \new_[77634]_ ,
    \new_[77635]_ , \new_[77636]_ , \new_[77640]_ , \new_[77641]_ ,
    \new_[77644]_ , \new_[77647]_ , \new_[77648]_ , \new_[77649]_ ,
    \new_[77652]_ , \new_[77655]_ , \new_[77656]_ , \new_[77659]_ ,
    \new_[77662]_ , \new_[77663]_ , \new_[77664]_ , \new_[77668]_ ,
    \new_[77669]_ , \new_[77672]_ , \new_[77675]_ , \new_[77676]_ ,
    \new_[77677]_ , \new_[77680]_ , \new_[77683]_ , \new_[77684]_ ,
    \new_[77687]_ , \new_[77690]_ , \new_[77691]_ , \new_[77692]_ ,
    \new_[77696]_ , \new_[77697]_ , \new_[77700]_ , \new_[77703]_ ,
    \new_[77704]_ , \new_[77705]_ , \new_[77708]_ , \new_[77711]_ ,
    \new_[77712]_ , \new_[77715]_ , \new_[77718]_ , \new_[77719]_ ,
    \new_[77720]_ , \new_[77724]_ , \new_[77725]_ , \new_[77728]_ ,
    \new_[77731]_ , \new_[77732]_ , \new_[77733]_ , \new_[77736]_ ,
    \new_[77739]_ , \new_[77740]_ , \new_[77743]_ , \new_[77746]_ ,
    \new_[77747]_ , \new_[77748]_ , \new_[77752]_ , \new_[77753]_ ,
    \new_[77756]_ , \new_[77759]_ , \new_[77760]_ , \new_[77761]_ ,
    \new_[77764]_ , \new_[77767]_ , \new_[77768]_ , \new_[77771]_ ,
    \new_[77774]_ , \new_[77775]_ , \new_[77776]_ , \new_[77780]_ ,
    \new_[77781]_ , \new_[77784]_ , \new_[77787]_ , \new_[77788]_ ,
    \new_[77789]_ , \new_[77792]_ , \new_[77795]_ , \new_[77796]_ ,
    \new_[77799]_ , \new_[77802]_ , \new_[77803]_ , \new_[77804]_ ,
    \new_[77808]_ , \new_[77809]_ , \new_[77812]_ , \new_[77815]_ ,
    \new_[77816]_ , \new_[77817]_ , \new_[77820]_ , \new_[77823]_ ,
    \new_[77824]_ , \new_[77827]_ , \new_[77830]_ , \new_[77831]_ ,
    \new_[77832]_ , \new_[77836]_ , \new_[77837]_ , \new_[77840]_ ,
    \new_[77843]_ , \new_[77844]_ , \new_[77845]_ , \new_[77848]_ ,
    \new_[77851]_ , \new_[77852]_ , \new_[77855]_ , \new_[77858]_ ,
    \new_[77859]_ , \new_[77860]_ , \new_[77864]_ , \new_[77865]_ ,
    \new_[77868]_ , \new_[77871]_ , \new_[77872]_ , \new_[77873]_ ,
    \new_[77876]_ , \new_[77879]_ , \new_[77880]_ , \new_[77883]_ ,
    \new_[77886]_ , \new_[77887]_ , \new_[77888]_ , \new_[77892]_ ,
    \new_[77893]_ , \new_[77896]_ , \new_[77899]_ , \new_[77900]_ ,
    \new_[77901]_ , \new_[77904]_ , \new_[77907]_ , \new_[77908]_ ,
    \new_[77911]_ , \new_[77914]_ , \new_[77915]_ , \new_[77916]_ ,
    \new_[77920]_ , \new_[77921]_ , \new_[77924]_ , \new_[77927]_ ,
    \new_[77928]_ , \new_[77929]_ , \new_[77932]_ , \new_[77935]_ ,
    \new_[77936]_ , \new_[77939]_ , \new_[77942]_ , \new_[77943]_ ,
    \new_[77944]_ , \new_[77948]_ , \new_[77949]_ , \new_[77952]_ ,
    \new_[77955]_ , \new_[77956]_ , \new_[77957]_ , \new_[77960]_ ,
    \new_[77963]_ , \new_[77964]_ , \new_[77967]_ , \new_[77970]_ ,
    \new_[77971]_ , \new_[77972]_ , \new_[77976]_ , \new_[77977]_ ,
    \new_[77980]_ , \new_[77983]_ , \new_[77984]_ , \new_[77985]_ ,
    \new_[77988]_ , \new_[77991]_ , \new_[77992]_ , \new_[77995]_ ,
    \new_[77998]_ , \new_[77999]_ , \new_[78000]_ , \new_[78004]_ ,
    \new_[78005]_ , \new_[78008]_ , \new_[78011]_ , \new_[78012]_ ,
    \new_[78013]_ , \new_[78016]_ , \new_[78019]_ , \new_[78020]_ ,
    \new_[78023]_ , \new_[78026]_ , \new_[78027]_ , \new_[78028]_ ,
    \new_[78032]_ , \new_[78033]_ , \new_[78036]_ , \new_[78039]_ ,
    \new_[78040]_ , \new_[78041]_ , \new_[78044]_ , \new_[78047]_ ,
    \new_[78048]_ , \new_[78051]_ , \new_[78054]_ , \new_[78055]_ ,
    \new_[78056]_ , \new_[78060]_ , \new_[78061]_ , \new_[78064]_ ,
    \new_[78067]_ , \new_[78068]_ , \new_[78069]_ , \new_[78072]_ ,
    \new_[78075]_ , \new_[78076]_ , \new_[78079]_ , \new_[78082]_ ,
    \new_[78083]_ , \new_[78084]_ , \new_[78088]_ , \new_[78089]_ ,
    \new_[78092]_ , \new_[78095]_ , \new_[78096]_ , \new_[78097]_ ,
    \new_[78100]_ , \new_[78103]_ , \new_[78104]_ , \new_[78107]_ ,
    \new_[78110]_ , \new_[78111]_ , \new_[78112]_ , \new_[78116]_ ,
    \new_[78117]_ , \new_[78120]_ , \new_[78123]_ , \new_[78124]_ ,
    \new_[78125]_ , \new_[78128]_ , \new_[78131]_ , \new_[78132]_ ,
    \new_[78135]_ , \new_[78138]_ , \new_[78139]_ , \new_[78140]_ ,
    \new_[78144]_ , \new_[78145]_ , \new_[78148]_ , \new_[78151]_ ,
    \new_[78152]_ , \new_[78153]_ , \new_[78156]_ , \new_[78159]_ ,
    \new_[78160]_ , \new_[78163]_ , \new_[78166]_ , \new_[78167]_ ,
    \new_[78168]_ , \new_[78172]_ , \new_[78173]_ , \new_[78176]_ ,
    \new_[78179]_ , \new_[78180]_ , \new_[78181]_ , \new_[78184]_ ,
    \new_[78187]_ , \new_[78188]_ , \new_[78191]_ , \new_[78194]_ ,
    \new_[78195]_ , \new_[78196]_ , \new_[78200]_ , \new_[78201]_ ,
    \new_[78204]_ , \new_[78207]_ , \new_[78208]_ , \new_[78209]_ ,
    \new_[78212]_ , \new_[78215]_ , \new_[78216]_ , \new_[78219]_ ,
    \new_[78222]_ , \new_[78223]_ , \new_[78224]_ , \new_[78228]_ ,
    \new_[78229]_ , \new_[78232]_ , \new_[78235]_ , \new_[78236]_ ,
    \new_[78237]_ , \new_[78240]_ , \new_[78243]_ , \new_[78244]_ ,
    \new_[78247]_ , \new_[78250]_ , \new_[78251]_ , \new_[78252]_ ,
    \new_[78256]_ , \new_[78257]_ , \new_[78260]_ , \new_[78263]_ ,
    \new_[78264]_ , \new_[78265]_ , \new_[78268]_ , \new_[78271]_ ,
    \new_[78272]_ , \new_[78275]_ , \new_[78278]_ , \new_[78279]_ ,
    \new_[78280]_ , \new_[78284]_ , \new_[78285]_ , \new_[78288]_ ,
    \new_[78291]_ , \new_[78292]_ , \new_[78293]_ , \new_[78296]_ ,
    \new_[78299]_ , \new_[78300]_ , \new_[78303]_ , \new_[78306]_ ,
    \new_[78307]_ , \new_[78308]_ , \new_[78312]_ , \new_[78313]_ ,
    \new_[78316]_ , \new_[78319]_ , \new_[78320]_ , \new_[78321]_ ,
    \new_[78324]_ , \new_[78327]_ , \new_[78328]_ , \new_[78331]_ ,
    \new_[78334]_ , \new_[78335]_ , \new_[78336]_ , \new_[78340]_ ,
    \new_[78341]_ , \new_[78344]_ , \new_[78347]_ , \new_[78348]_ ,
    \new_[78349]_ , \new_[78352]_ , \new_[78355]_ , \new_[78356]_ ,
    \new_[78359]_ , \new_[78362]_ , \new_[78363]_ , \new_[78364]_ ,
    \new_[78368]_ , \new_[78369]_ , \new_[78372]_ , \new_[78375]_ ,
    \new_[78376]_ , \new_[78377]_ , \new_[78380]_ , \new_[78383]_ ,
    \new_[78384]_ , \new_[78387]_ , \new_[78390]_ , \new_[78391]_ ,
    \new_[78392]_ , \new_[78396]_ , \new_[78397]_ , \new_[78400]_ ,
    \new_[78403]_ , \new_[78404]_ , \new_[78405]_ , \new_[78408]_ ,
    \new_[78411]_ , \new_[78412]_ , \new_[78415]_ , \new_[78418]_ ,
    \new_[78419]_ , \new_[78420]_ , \new_[78424]_ , \new_[78425]_ ,
    \new_[78428]_ , \new_[78431]_ , \new_[78432]_ , \new_[78433]_ ,
    \new_[78436]_ , \new_[78439]_ , \new_[78440]_ , \new_[78443]_ ,
    \new_[78446]_ , \new_[78447]_ , \new_[78448]_ , \new_[78452]_ ,
    \new_[78453]_ , \new_[78456]_ , \new_[78459]_ , \new_[78460]_ ,
    \new_[78461]_ , \new_[78464]_ , \new_[78467]_ , \new_[78468]_ ,
    \new_[78471]_ , \new_[78474]_ , \new_[78475]_ , \new_[78476]_ ,
    \new_[78480]_ , \new_[78481]_ , \new_[78484]_ , \new_[78487]_ ,
    \new_[78488]_ , \new_[78489]_ , \new_[78492]_ , \new_[78495]_ ,
    \new_[78496]_ , \new_[78499]_ , \new_[78502]_ , \new_[78503]_ ,
    \new_[78504]_ , \new_[78508]_ , \new_[78509]_ , \new_[78512]_ ,
    \new_[78515]_ , \new_[78516]_ , \new_[78517]_ , \new_[78520]_ ,
    \new_[78523]_ , \new_[78524]_ , \new_[78527]_ , \new_[78530]_ ,
    \new_[78531]_ , \new_[78532]_ , \new_[78536]_ , \new_[78537]_ ,
    \new_[78540]_ , \new_[78543]_ , \new_[78544]_ , \new_[78545]_ ,
    \new_[78548]_ , \new_[78551]_ , \new_[78552]_ , \new_[78555]_ ,
    \new_[78558]_ , \new_[78559]_ , \new_[78560]_ , \new_[78564]_ ,
    \new_[78565]_ , \new_[78568]_ , \new_[78571]_ , \new_[78572]_ ,
    \new_[78573]_ , \new_[78576]_ , \new_[78579]_ , \new_[78580]_ ,
    \new_[78583]_ , \new_[78586]_ , \new_[78587]_ , \new_[78588]_ ,
    \new_[78592]_ , \new_[78593]_ , \new_[78596]_ , \new_[78599]_ ,
    \new_[78600]_ , \new_[78601]_ , \new_[78604]_ , \new_[78607]_ ,
    \new_[78608]_ , \new_[78611]_ , \new_[78614]_ , \new_[78615]_ ,
    \new_[78616]_ , \new_[78620]_ , \new_[78621]_ , \new_[78624]_ ,
    \new_[78627]_ , \new_[78628]_ , \new_[78629]_ , \new_[78632]_ ,
    \new_[78635]_ , \new_[78636]_ , \new_[78639]_ , \new_[78642]_ ,
    \new_[78643]_ , \new_[78644]_ , \new_[78648]_ , \new_[78649]_ ,
    \new_[78652]_ , \new_[78655]_ , \new_[78656]_ , \new_[78657]_ ,
    \new_[78660]_ , \new_[78663]_ , \new_[78664]_ , \new_[78667]_ ,
    \new_[78670]_ , \new_[78671]_ , \new_[78672]_ , \new_[78676]_ ,
    \new_[78677]_ , \new_[78680]_ , \new_[78683]_ , \new_[78684]_ ,
    \new_[78685]_ , \new_[78688]_ , \new_[78691]_ , \new_[78692]_ ,
    \new_[78695]_ , \new_[78698]_ , \new_[78699]_ , \new_[78700]_ ,
    \new_[78704]_ , \new_[78705]_ , \new_[78708]_ , \new_[78711]_ ,
    \new_[78712]_ , \new_[78713]_ , \new_[78716]_ , \new_[78719]_ ,
    \new_[78720]_ , \new_[78723]_ , \new_[78726]_ , \new_[78727]_ ,
    \new_[78728]_ , \new_[78732]_ , \new_[78733]_ , \new_[78736]_ ,
    \new_[78739]_ , \new_[78740]_ , \new_[78741]_ , \new_[78744]_ ,
    \new_[78747]_ , \new_[78748]_ , \new_[78751]_ , \new_[78754]_ ,
    \new_[78755]_ , \new_[78756]_ , \new_[78760]_ , \new_[78761]_ ,
    \new_[78764]_ , \new_[78767]_ , \new_[78768]_ , \new_[78769]_ ,
    \new_[78772]_ , \new_[78775]_ , \new_[78776]_ , \new_[78779]_ ,
    \new_[78782]_ , \new_[78783]_ , \new_[78784]_ , \new_[78788]_ ,
    \new_[78789]_ , \new_[78792]_ , \new_[78795]_ , \new_[78796]_ ,
    \new_[78797]_ , \new_[78800]_ , \new_[78803]_ , \new_[78804]_ ,
    \new_[78807]_ , \new_[78810]_ , \new_[78811]_ , \new_[78812]_ ,
    \new_[78816]_ , \new_[78817]_ , \new_[78820]_ , \new_[78823]_ ,
    \new_[78824]_ , \new_[78825]_ , \new_[78828]_ , \new_[78831]_ ,
    \new_[78832]_ , \new_[78835]_ , \new_[78838]_ , \new_[78839]_ ,
    \new_[78840]_ , \new_[78844]_ , \new_[78845]_ , \new_[78848]_ ,
    \new_[78851]_ , \new_[78852]_ , \new_[78853]_ , \new_[78856]_ ,
    \new_[78859]_ , \new_[78860]_ , \new_[78863]_ , \new_[78866]_ ,
    \new_[78867]_ , \new_[78868]_ , \new_[78872]_ , \new_[78873]_ ,
    \new_[78876]_ , \new_[78879]_ , \new_[78880]_ , \new_[78881]_ ,
    \new_[78884]_ , \new_[78887]_ , \new_[78888]_ , \new_[78891]_ ,
    \new_[78894]_ , \new_[78895]_ , \new_[78896]_ , \new_[78900]_ ,
    \new_[78901]_ , \new_[78904]_ , \new_[78907]_ , \new_[78908]_ ,
    \new_[78909]_ , \new_[78912]_ , \new_[78915]_ , \new_[78916]_ ,
    \new_[78919]_ , \new_[78922]_ , \new_[78923]_ , \new_[78924]_ ,
    \new_[78928]_ , \new_[78929]_ , \new_[78932]_ , \new_[78935]_ ,
    \new_[78936]_ , \new_[78937]_ , \new_[78940]_ , \new_[78943]_ ,
    \new_[78944]_ , \new_[78947]_ , \new_[78950]_ , \new_[78951]_ ,
    \new_[78952]_ , \new_[78956]_ , \new_[78957]_ , \new_[78960]_ ,
    \new_[78963]_ , \new_[78964]_ , \new_[78965]_ , \new_[78968]_ ,
    \new_[78971]_ , \new_[78972]_ , \new_[78975]_ , \new_[78978]_ ,
    \new_[78979]_ , \new_[78980]_ , \new_[78984]_ , \new_[78985]_ ,
    \new_[78988]_ , \new_[78991]_ , \new_[78992]_ , \new_[78993]_ ,
    \new_[78996]_ , \new_[78999]_ , \new_[79000]_ , \new_[79003]_ ,
    \new_[79006]_ , \new_[79007]_ , \new_[79008]_ , \new_[79012]_ ,
    \new_[79013]_ , \new_[79016]_ , \new_[79019]_ , \new_[79020]_ ,
    \new_[79021]_ , \new_[79024]_ , \new_[79027]_ , \new_[79028]_ ,
    \new_[79031]_ , \new_[79034]_ , \new_[79035]_ , \new_[79036]_ ,
    \new_[79040]_ , \new_[79041]_ , \new_[79044]_ , \new_[79047]_ ,
    \new_[79048]_ , \new_[79049]_ , \new_[79052]_ , \new_[79055]_ ,
    \new_[79056]_ , \new_[79059]_ , \new_[79062]_ , \new_[79063]_ ,
    \new_[79064]_ , \new_[79068]_ , \new_[79069]_ , \new_[79072]_ ,
    \new_[79075]_ , \new_[79076]_ , \new_[79077]_ , \new_[79080]_ ,
    \new_[79083]_ , \new_[79084]_ , \new_[79087]_ , \new_[79090]_ ,
    \new_[79091]_ , \new_[79092]_ , \new_[79096]_ , \new_[79097]_ ,
    \new_[79100]_ , \new_[79103]_ , \new_[79104]_ , \new_[79105]_ ,
    \new_[79108]_ , \new_[79111]_ , \new_[79112]_ , \new_[79115]_ ,
    \new_[79118]_ , \new_[79119]_ , \new_[79120]_ , \new_[79124]_ ,
    \new_[79125]_ , \new_[79128]_ , \new_[79131]_ , \new_[79132]_ ,
    \new_[79133]_ , \new_[79136]_ , \new_[79139]_ , \new_[79140]_ ,
    \new_[79143]_ , \new_[79146]_ , \new_[79147]_ , \new_[79148]_ ,
    \new_[79152]_ , \new_[79153]_ , \new_[79156]_ , \new_[79159]_ ,
    \new_[79160]_ , \new_[79161]_ , \new_[79164]_ , \new_[79167]_ ,
    \new_[79168]_ , \new_[79171]_ , \new_[79174]_ , \new_[79175]_ ,
    \new_[79176]_ , \new_[79180]_ , \new_[79181]_ , \new_[79184]_ ,
    \new_[79187]_ , \new_[79188]_ , \new_[79189]_ , \new_[79192]_ ,
    \new_[79195]_ , \new_[79196]_ , \new_[79199]_ , \new_[79202]_ ,
    \new_[79203]_ , \new_[79204]_ , \new_[79208]_ , \new_[79209]_ ,
    \new_[79212]_ , \new_[79215]_ , \new_[79216]_ , \new_[79217]_ ,
    \new_[79220]_ , \new_[79223]_ , \new_[79224]_ , \new_[79227]_ ,
    \new_[79230]_ , \new_[79231]_ , \new_[79232]_ , \new_[79236]_ ,
    \new_[79237]_ , \new_[79240]_ , \new_[79243]_ , \new_[79244]_ ,
    \new_[79245]_ , \new_[79248]_ , \new_[79251]_ , \new_[79252]_ ,
    \new_[79255]_ , \new_[79258]_ , \new_[79259]_ , \new_[79260]_ ,
    \new_[79264]_ , \new_[79265]_ , \new_[79268]_ , \new_[79271]_ ,
    \new_[79272]_ , \new_[79273]_ , \new_[79276]_ , \new_[79279]_ ,
    \new_[79280]_ , \new_[79283]_ , \new_[79286]_ , \new_[79287]_ ,
    \new_[79288]_ , \new_[79292]_ , \new_[79293]_ , \new_[79296]_ ,
    \new_[79299]_ , \new_[79300]_ , \new_[79301]_ , \new_[79304]_ ,
    \new_[79307]_ , \new_[79308]_ , \new_[79311]_ , \new_[79314]_ ,
    \new_[79315]_ , \new_[79316]_ , \new_[79320]_ , \new_[79321]_ ,
    \new_[79324]_ , \new_[79327]_ , \new_[79328]_ , \new_[79329]_ ,
    \new_[79332]_ , \new_[79335]_ , \new_[79336]_ , \new_[79339]_ ,
    \new_[79342]_ , \new_[79343]_ , \new_[79344]_ , \new_[79348]_ ,
    \new_[79349]_ , \new_[79352]_ , \new_[79355]_ , \new_[79356]_ ,
    \new_[79357]_ , \new_[79360]_ , \new_[79363]_ , \new_[79364]_ ,
    \new_[79367]_ , \new_[79370]_ , \new_[79371]_ , \new_[79372]_ ,
    \new_[79376]_ , \new_[79377]_ , \new_[79380]_ , \new_[79383]_ ,
    \new_[79384]_ , \new_[79385]_ , \new_[79388]_ , \new_[79391]_ ,
    \new_[79392]_ , \new_[79395]_ , \new_[79398]_ , \new_[79399]_ ,
    \new_[79400]_ , \new_[79404]_ , \new_[79405]_ , \new_[79408]_ ,
    \new_[79411]_ , \new_[79412]_ , \new_[79413]_ , \new_[79416]_ ,
    \new_[79419]_ , \new_[79420]_ , \new_[79423]_ , \new_[79426]_ ,
    \new_[79427]_ , \new_[79428]_ , \new_[79432]_ , \new_[79433]_ ,
    \new_[79436]_ , \new_[79439]_ , \new_[79440]_ , \new_[79441]_ ,
    \new_[79444]_ , \new_[79447]_ , \new_[79448]_ , \new_[79451]_ ,
    \new_[79454]_ , \new_[79455]_ , \new_[79456]_ , \new_[79460]_ ,
    \new_[79461]_ , \new_[79464]_ , \new_[79467]_ , \new_[79468]_ ,
    \new_[79469]_ , \new_[79472]_ , \new_[79475]_ , \new_[79476]_ ,
    \new_[79479]_ , \new_[79482]_ , \new_[79483]_ , \new_[79484]_ ,
    \new_[79488]_ , \new_[79489]_ , \new_[79492]_ , \new_[79495]_ ,
    \new_[79496]_ , \new_[79497]_ , \new_[79500]_ , \new_[79503]_ ,
    \new_[79504]_ , \new_[79507]_ , \new_[79510]_ , \new_[79511]_ ,
    \new_[79512]_ , \new_[79516]_ , \new_[79517]_ , \new_[79520]_ ,
    \new_[79523]_ , \new_[79524]_ , \new_[79525]_ , \new_[79528]_ ,
    \new_[79531]_ , \new_[79532]_ , \new_[79535]_ , \new_[79538]_ ,
    \new_[79539]_ , \new_[79540]_ , \new_[79544]_ , \new_[79545]_ ,
    \new_[79548]_ , \new_[79551]_ , \new_[79552]_ , \new_[79553]_ ,
    \new_[79556]_ , \new_[79559]_ , \new_[79560]_ , \new_[79563]_ ,
    \new_[79566]_ , \new_[79567]_ , \new_[79568]_ , \new_[79572]_ ,
    \new_[79573]_ , \new_[79576]_ , \new_[79579]_ , \new_[79580]_ ,
    \new_[79581]_ , \new_[79584]_ , \new_[79587]_ , \new_[79588]_ ,
    \new_[79591]_ , \new_[79594]_ , \new_[79595]_ , \new_[79596]_ ,
    \new_[79600]_ , \new_[79601]_ , \new_[79604]_ , \new_[79607]_ ,
    \new_[79608]_ , \new_[79609]_ , \new_[79612]_ , \new_[79615]_ ,
    \new_[79616]_ , \new_[79619]_ , \new_[79622]_ , \new_[79623]_ ,
    \new_[79624]_ , \new_[79628]_ , \new_[79629]_ , \new_[79632]_ ,
    \new_[79635]_ , \new_[79636]_ , \new_[79637]_ , \new_[79640]_ ,
    \new_[79643]_ , \new_[79644]_ , \new_[79647]_ , \new_[79650]_ ,
    \new_[79651]_ , \new_[79652]_ , \new_[79656]_ , \new_[79657]_ ,
    \new_[79660]_ , \new_[79663]_ , \new_[79664]_ , \new_[79665]_ ,
    \new_[79668]_ , \new_[79671]_ , \new_[79672]_ , \new_[79675]_ ,
    \new_[79678]_ , \new_[79679]_ , \new_[79680]_ , \new_[79684]_ ,
    \new_[79685]_ , \new_[79688]_ , \new_[79691]_ , \new_[79692]_ ,
    \new_[79693]_ , \new_[79696]_ , \new_[79699]_ , \new_[79700]_ ,
    \new_[79703]_ , \new_[79706]_ , \new_[79707]_ , \new_[79708]_ ,
    \new_[79712]_ , \new_[79713]_ , \new_[79716]_ , \new_[79719]_ ,
    \new_[79720]_ , \new_[79721]_ , \new_[79724]_ , \new_[79727]_ ,
    \new_[79728]_ , \new_[79731]_ , \new_[79734]_ , \new_[79735]_ ,
    \new_[79736]_ , \new_[79740]_ , \new_[79741]_ , \new_[79744]_ ,
    \new_[79747]_ , \new_[79748]_ , \new_[79749]_ , \new_[79752]_ ,
    \new_[79755]_ , \new_[79756]_ , \new_[79759]_ , \new_[79762]_ ,
    \new_[79763]_ , \new_[79764]_ , \new_[79768]_ , \new_[79769]_ ,
    \new_[79772]_ , \new_[79775]_ , \new_[79776]_ , \new_[79777]_ ,
    \new_[79780]_ , \new_[79783]_ , \new_[79784]_ , \new_[79787]_ ,
    \new_[79790]_ , \new_[79791]_ , \new_[79792]_ , \new_[79796]_ ,
    \new_[79797]_ , \new_[79800]_ , \new_[79803]_ , \new_[79804]_ ,
    \new_[79805]_ , \new_[79808]_ , \new_[79811]_ , \new_[79812]_ ,
    \new_[79815]_ , \new_[79818]_ , \new_[79819]_ , \new_[79820]_ ,
    \new_[79824]_ , \new_[79825]_ , \new_[79828]_ , \new_[79831]_ ,
    \new_[79832]_ , \new_[79833]_ , \new_[79836]_ , \new_[79839]_ ,
    \new_[79840]_ , \new_[79843]_ , \new_[79846]_ , \new_[79847]_ ,
    \new_[79848]_ , \new_[79852]_ , \new_[79853]_ , \new_[79856]_ ,
    \new_[79859]_ , \new_[79860]_ , \new_[79861]_ , \new_[79864]_ ,
    \new_[79867]_ , \new_[79868]_ , \new_[79871]_ , \new_[79874]_ ,
    \new_[79875]_ , \new_[79876]_ , \new_[79880]_ , \new_[79881]_ ,
    \new_[79884]_ , \new_[79887]_ , \new_[79888]_ , \new_[79889]_ ,
    \new_[79892]_ , \new_[79895]_ , \new_[79896]_ , \new_[79899]_ ,
    \new_[79902]_ , \new_[79903]_ , \new_[79904]_ , \new_[79908]_ ,
    \new_[79909]_ , \new_[79912]_ , \new_[79915]_ , \new_[79916]_ ,
    \new_[79917]_ , \new_[79920]_ , \new_[79923]_ , \new_[79924]_ ,
    \new_[79927]_ , \new_[79930]_ , \new_[79931]_ , \new_[79932]_ ,
    \new_[79936]_ , \new_[79937]_ , \new_[79940]_ , \new_[79943]_ ,
    \new_[79944]_ , \new_[79945]_ , \new_[79948]_ , \new_[79951]_ ,
    \new_[79952]_ , \new_[79955]_ , \new_[79958]_ , \new_[79959]_ ,
    \new_[79960]_ , \new_[79964]_ , \new_[79965]_ , \new_[79968]_ ,
    \new_[79971]_ , \new_[79972]_ , \new_[79973]_ , \new_[79976]_ ,
    \new_[79979]_ , \new_[79980]_ , \new_[79983]_ , \new_[79986]_ ,
    \new_[79987]_ , \new_[79988]_ , \new_[79992]_ , \new_[79993]_ ,
    \new_[79996]_ , \new_[79999]_ , \new_[80000]_ , \new_[80001]_ ,
    \new_[80004]_ , \new_[80007]_ , \new_[80008]_ , \new_[80011]_ ,
    \new_[80014]_ , \new_[80015]_ , \new_[80016]_ , \new_[80020]_ ,
    \new_[80021]_ , \new_[80024]_ , \new_[80027]_ , \new_[80028]_ ,
    \new_[80029]_ , \new_[80032]_ , \new_[80035]_ , \new_[80036]_ ,
    \new_[80039]_ , \new_[80042]_ , \new_[80043]_ , \new_[80044]_ ,
    \new_[80048]_ , \new_[80049]_ , \new_[80052]_ , \new_[80055]_ ,
    \new_[80056]_ , \new_[80057]_ , \new_[80060]_ , \new_[80063]_ ,
    \new_[80064]_ , \new_[80067]_ , \new_[80070]_ , \new_[80071]_ ,
    \new_[80072]_ , \new_[80076]_ , \new_[80077]_ , \new_[80080]_ ,
    \new_[80083]_ , \new_[80084]_ , \new_[80085]_ , \new_[80088]_ ,
    \new_[80091]_ , \new_[80092]_ , \new_[80095]_ , \new_[80098]_ ,
    \new_[80099]_ , \new_[80100]_ , \new_[80104]_ , \new_[80105]_ ,
    \new_[80108]_ , \new_[80111]_ , \new_[80112]_ , \new_[80113]_ ,
    \new_[80116]_ , \new_[80119]_ , \new_[80120]_ , \new_[80123]_ ,
    \new_[80126]_ , \new_[80127]_ , \new_[80128]_ , \new_[80132]_ ,
    \new_[80133]_ , \new_[80136]_ , \new_[80139]_ , \new_[80140]_ ,
    \new_[80141]_ , \new_[80144]_ , \new_[80147]_ , \new_[80148]_ ,
    \new_[80151]_ , \new_[80154]_ , \new_[80155]_ , \new_[80156]_ ,
    \new_[80160]_ , \new_[80161]_ , \new_[80164]_ , \new_[80167]_ ,
    \new_[80168]_ , \new_[80169]_ , \new_[80172]_ , \new_[80175]_ ,
    \new_[80176]_ , \new_[80179]_ , \new_[80182]_ , \new_[80183]_ ,
    \new_[80184]_ , \new_[80188]_ , \new_[80189]_ , \new_[80192]_ ,
    \new_[80195]_ , \new_[80196]_ , \new_[80197]_ , \new_[80200]_ ,
    \new_[80203]_ , \new_[80204]_ , \new_[80207]_ , \new_[80210]_ ,
    \new_[80211]_ , \new_[80212]_ , \new_[80216]_ , \new_[80217]_ ,
    \new_[80220]_ , \new_[80223]_ , \new_[80224]_ , \new_[80225]_ ,
    \new_[80228]_ , \new_[80231]_ , \new_[80232]_ , \new_[80235]_ ,
    \new_[80238]_ , \new_[80239]_ , \new_[80240]_ , \new_[80244]_ ,
    \new_[80245]_ , \new_[80248]_ , \new_[80251]_ , \new_[80252]_ ,
    \new_[80253]_ , \new_[80256]_ , \new_[80259]_ , \new_[80260]_ ,
    \new_[80263]_ , \new_[80266]_ , \new_[80267]_ , \new_[80268]_ ,
    \new_[80272]_ , \new_[80273]_ , \new_[80276]_ , \new_[80279]_ ,
    \new_[80280]_ , \new_[80281]_ , \new_[80284]_ , \new_[80287]_ ,
    \new_[80288]_ , \new_[80291]_ , \new_[80294]_ , \new_[80295]_ ,
    \new_[80296]_ , \new_[80300]_ , \new_[80301]_ , \new_[80304]_ ,
    \new_[80307]_ , \new_[80308]_ , \new_[80309]_ , \new_[80312]_ ,
    \new_[80315]_ , \new_[80316]_ , \new_[80319]_ , \new_[80322]_ ,
    \new_[80323]_ , \new_[80324]_ , \new_[80328]_ , \new_[80329]_ ,
    \new_[80332]_ , \new_[80335]_ , \new_[80336]_ , \new_[80337]_ ,
    \new_[80340]_ , \new_[80343]_ , \new_[80344]_ , \new_[80347]_ ,
    \new_[80350]_ , \new_[80351]_ , \new_[80352]_ , \new_[80356]_ ,
    \new_[80357]_ , \new_[80360]_ , \new_[80363]_ , \new_[80364]_ ,
    \new_[80365]_ , \new_[80368]_ , \new_[80371]_ , \new_[80372]_ ,
    \new_[80375]_ , \new_[80378]_ , \new_[80379]_ , \new_[80380]_ ,
    \new_[80384]_ , \new_[80385]_ , \new_[80388]_ , \new_[80391]_ ,
    \new_[80392]_ , \new_[80393]_ , \new_[80396]_ , \new_[80399]_ ,
    \new_[80400]_ , \new_[80403]_ , \new_[80406]_ , \new_[80407]_ ,
    \new_[80408]_ , \new_[80412]_ , \new_[80413]_ , \new_[80416]_ ,
    \new_[80419]_ , \new_[80420]_ , \new_[80421]_ , \new_[80424]_ ,
    \new_[80427]_ , \new_[80428]_ , \new_[80431]_ , \new_[80434]_ ,
    \new_[80435]_ , \new_[80436]_ , \new_[80440]_ , \new_[80441]_ ,
    \new_[80444]_ , \new_[80447]_ , \new_[80448]_ , \new_[80449]_ ,
    \new_[80452]_ , \new_[80455]_ , \new_[80456]_ , \new_[80459]_ ,
    \new_[80462]_ , \new_[80463]_ , \new_[80464]_ , \new_[80468]_ ,
    \new_[80469]_ , \new_[80472]_ , \new_[80475]_ , \new_[80476]_ ,
    \new_[80477]_ , \new_[80480]_ , \new_[80483]_ , \new_[80484]_ ,
    \new_[80487]_ , \new_[80490]_ , \new_[80491]_ , \new_[80492]_ ,
    \new_[80496]_ , \new_[80497]_ , \new_[80500]_ , \new_[80503]_ ,
    \new_[80504]_ , \new_[80505]_ , \new_[80508]_ , \new_[80511]_ ,
    \new_[80512]_ , \new_[80515]_ , \new_[80518]_ , \new_[80519]_ ,
    \new_[80520]_ , \new_[80524]_ , \new_[80525]_ , \new_[80528]_ ,
    \new_[80531]_ , \new_[80532]_ , \new_[80533]_ , \new_[80536]_ ,
    \new_[80539]_ , \new_[80540]_ , \new_[80543]_ , \new_[80546]_ ,
    \new_[80547]_ , \new_[80548]_ , \new_[80552]_ , \new_[80553]_ ,
    \new_[80556]_ , \new_[80559]_ , \new_[80560]_ , \new_[80561]_ ,
    \new_[80564]_ , \new_[80567]_ , \new_[80568]_ , \new_[80571]_ ,
    \new_[80574]_ , \new_[80575]_ , \new_[80576]_ , \new_[80580]_ ,
    \new_[80581]_ , \new_[80584]_ , \new_[80587]_ , \new_[80588]_ ,
    \new_[80589]_ , \new_[80592]_ , \new_[80595]_ , \new_[80596]_ ,
    \new_[80599]_ , \new_[80602]_ , \new_[80603]_ , \new_[80604]_ ,
    \new_[80608]_ , \new_[80609]_ , \new_[80612]_ , \new_[80615]_ ,
    \new_[80616]_ , \new_[80617]_ , \new_[80620]_ , \new_[80623]_ ,
    \new_[80624]_ , \new_[80627]_ , \new_[80630]_ , \new_[80631]_ ,
    \new_[80632]_ , \new_[80636]_ , \new_[80637]_ , \new_[80640]_ ,
    \new_[80643]_ , \new_[80644]_ , \new_[80645]_ , \new_[80648]_ ,
    \new_[80651]_ , \new_[80652]_ , \new_[80655]_ , \new_[80658]_ ,
    \new_[80659]_ , \new_[80660]_ , \new_[80664]_ , \new_[80665]_ ,
    \new_[80668]_ , \new_[80671]_ , \new_[80672]_ , \new_[80673]_ ,
    \new_[80676]_ , \new_[80679]_ , \new_[80680]_ , \new_[80683]_ ,
    \new_[80686]_ , \new_[80687]_ , \new_[80688]_ , \new_[80692]_ ,
    \new_[80693]_ , \new_[80696]_ , \new_[80699]_ , \new_[80700]_ ,
    \new_[80701]_ , \new_[80704]_ , \new_[80707]_ , \new_[80708]_ ,
    \new_[80711]_ , \new_[80714]_ , \new_[80715]_ , \new_[80716]_ ,
    \new_[80720]_ , \new_[80721]_ , \new_[80724]_ , \new_[80727]_ ,
    \new_[80728]_ , \new_[80729]_ , \new_[80732]_ , \new_[80735]_ ,
    \new_[80736]_ , \new_[80739]_ , \new_[80742]_ , \new_[80743]_ ,
    \new_[80744]_ , \new_[80748]_ , \new_[80749]_ , \new_[80752]_ ,
    \new_[80755]_ , \new_[80756]_ , \new_[80757]_ , \new_[80760]_ ,
    \new_[80763]_ , \new_[80764]_ , \new_[80767]_ , \new_[80770]_ ,
    \new_[80771]_ , \new_[80772]_ , \new_[80776]_ , \new_[80777]_ ,
    \new_[80780]_ , \new_[80783]_ , \new_[80784]_ , \new_[80785]_ ,
    \new_[80788]_ , \new_[80791]_ , \new_[80792]_ , \new_[80795]_ ,
    \new_[80798]_ , \new_[80799]_ , \new_[80800]_ , \new_[80804]_ ,
    \new_[80805]_ , \new_[80808]_ , \new_[80811]_ , \new_[80812]_ ,
    \new_[80813]_ , \new_[80816]_ , \new_[80819]_ , \new_[80820]_ ,
    \new_[80823]_ , \new_[80826]_ , \new_[80827]_ , \new_[80828]_ ,
    \new_[80832]_ , \new_[80833]_ , \new_[80836]_ , \new_[80839]_ ,
    \new_[80840]_ , \new_[80841]_ , \new_[80844]_ , \new_[80847]_ ,
    \new_[80848]_ , \new_[80851]_ , \new_[80854]_ , \new_[80855]_ ,
    \new_[80856]_ , \new_[80860]_ , \new_[80861]_ , \new_[80864]_ ,
    \new_[80867]_ , \new_[80868]_ , \new_[80869]_ , \new_[80872]_ ,
    \new_[80875]_ , \new_[80876]_ , \new_[80879]_ , \new_[80882]_ ,
    \new_[80883]_ , \new_[80884]_ , \new_[80888]_ , \new_[80889]_ ,
    \new_[80892]_ , \new_[80895]_ , \new_[80896]_ , \new_[80897]_ ,
    \new_[80900]_ , \new_[80903]_ , \new_[80904]_ , \new_[80907]_ ,
    \new_[80910]_ , \new_[80911]_ , \new_[80912]_ , \new_[80916]_ ,
    \new_[80917]_ , \new_[80920]_ , \new_[80923]_ , \new_[80924]_ ,
    \new_[80925]_ , \new_[80928]_ , \new_[80931]_ , \new_[80932]_ ,
    \new_[80935]_ , \new_[80938]_ , \new_[80939]_ , \new_[80940]_ ,
    \new_[80944]_ , \new_[80945]_ , \new_[80948]_ , \new_[80951]_ ,
    \new_[80952]_ , \new_[80953]_ , \new_[80956]_ , \new_[80959]_ ,
    \new_[80960]_ , \new_[80963]_ , \new_[80966]_ , \new_[80967]_ ,
    \new_[80968]_ , \new_[80972]_ , \new_[80973]_ , \new_[80976]_ ,
    \new_[80979]_ , \new_[80980]_ , \new_[80981]_ , \new_[80984]_ ,
    \new_[80987]_ , \new_[80988]_ , \new_[80991]_ , \new_[80994]_ ,
    \new_[80995]_ , \new_[80996]_ , \new_[81000]_ , \new_[81001]_ ,
    \new_[81004]_ , \new_[81007]_ , \new_[81008]_ , \new_[81009]_ ,
    \new_[81012]_ , \new_[81015]_ , \new_[81016]_ , \new_[81019]_ ,
    \new_[81022]_ , \new_[81023]_ , \new_[81024]_ , \new_[81028]_ ,
    \new_[81029]_ , \new_[81032]_ , \new_[81035]_ , \new_[81036]_ ,
    \new_[81037]_ , \new_[81040]_ , \new_[81043]_ , \new_[81044]_ ,
    \new_[81047]_ , \new_[81050]_ , \new_[81051]_ , \new_[81052]_ ,
    \new_[81056]_ , \new_[81057]_ , \new_[81060]_ , \new_[81063]_ ,
    \new_[81064]_ , \new_[81065]_ , \new_[81068]_ , \new_[81071]_ ,
    \new_[81072]_ , \new_[81075]_ , \new_[81078]_ , \new_[81079]_ ,
    \new_[81080]_ , \new_[81084]_ , \new_[81085]_ , \new_[81088]_ ,
    \new_[81091]_ , \new_[81092]_ , \new_[81093]_ , \new_[81096]_ ,
    \new_[81099]_ , \new_[81100]_ , \new_[81103]_ , \new_[81106]_ ,
    \new_[81107]_ , \new_[81108]_ , \new_[81112]_ , \new_[81113]_ ,
    \new_[81116]_ , \new_[81119]_ , \new_[81120]_ , \new_[81121]_ ,
    \new_[81124]_ , \new_[81127]_ , \new_[81128]_ , \new_[81131]_ ,
    \new_[81134]_ , \new_[81135]_ , \new_[81136]_ , \new_[81140]_ ,
    \new_[81141]_ , \new_[81144]_ , \new_[81147]_ , \new_[81148]_ ,
    \new_[81149]_ , \new_[81152]_ , \new_[81155]_ , \new_[81156]_ ,
    \new_[81159]_ , \new_[81162]_ , \new_[81163]_ , \new_[81164]_ ,
    \new_[81168]_ , \new_[81169]_ , \new_[81172]_ , \new_[81175]_ ,
    \new_[81176]_ , \new_[81177]_ , \new_[81180]_ , \new_[81183]_ ,
    \new_[81184]_ , \new_[81187]_ , \new_[81190]_ , \new_[81191]_ ,
    \new_[81192]_ , \new_[81196]_ , \new_[81197]_ , \new_[81200]_ ,
    \new_[81203]_ , \new_[81204]_ , \new_[81205]_ , \new_[81208]_ ,
    \new_[81211]_ , \new_[81212]_ , \new_[81215]_ , \new_[81218]_ ,
    \new_[81219]_ , \new_[81220]_ , \new_[81224]_ , \new_[81225]_ ,
    \new_[81228]_ , \new_[81231]_ , \new_[81232]_ , \new_[81233]_ ,
    \new_[81236]_ , \new_[81239]_ , \new_[81240]_ , \new_[81243]_ ,
    \new_[81246]_ , \new_[81247]_ , \new_[81248]_ , \new_[81252]_ ,
    \new_[81253]_ , \new_[81256]_ , \new_[81259]_ , \new_[81260]_ ,
    \new_[81261]_ , \new_[81264]_ , \new_[81267]_ , \new_[81268]_ ,
    \new_[81271]_ , \new_[81274]_ , \new_[81275]_ , \new_[81276]_ ,
    \new_[81280]_ , \new_[81281]_ , \new_[81284]_ , \new_[81287]_ ,
    \new_[81288]_ , \new_[81289]_ , \new_[81292]_ , \new_[81295]_ ,
    \new_[81296]_ , \new_[81299]_ , \new_[81302]_ , \new_[81303]_ ,
    \new_[81304]_ , \new_[81308]_ , \new_[81309]_ , \new_[81312]_ ,
    \new_[81315]_ , \new_[81316]_ , \new_[81317]_ , \new_[81320]_ ,
    \new_[81323]_ , \new_[81324]_ , \new_[81327]_ , \new_[81330]_ ,
    \new_[81331]_ , \new_[81332]_ , \new_[81336]_ , \new_[81337]_ ,
    \new_[81340]_ , \new_[81343]_ , \new_[81344]_ , \new_[81345]_ ,
    \new_[81348]_ , \new_[81351]_ , \new_[81352]_ , \new_[81355]_ ,
    \new_[81358]_ , \new_[81359]_ , \new_[81360]_ , \new_[81364]_ ,
    \new_[81365]_ , \new_[81368]_ , \new_[81371]_ , \new_[81372]_ ,
    \new_[81373]_ , \new_[81376]_ , \new_[81379]_ , \new_[81380]_ ,
    \new_[81383]_ , \new_[81386]_ , \new_[81387]_ , \new_[81388]_ ,
    \new_[81392]_ , \new_[81393]_ , \new_[81396]_ , \new_[81399]_ ,
    \new_[81400]_ , \new_[81401]_ , \new_[81404]_ , \new_[81407]_ ,
    \new_[81408]_ , \new_[81411]_ , \new_[81414]_ , \new_[81415]_ ,
    \new_[81416]_ , \new_[81420]_ , \new_[81421]_ , \new_[81424]_ ,
    \new_[81427]_ , \new_[81428]_ , \new_[81429]_ , \new_[81432]_ ,
    \new_[81435]_ , \new_[81436]_ , \new_[81439]_ , \new_[81442]_ ,
    \new_[81443]_ , \new_[81444]_ , \new_[81448]_ , \new_[81449]_ ,
    \new_[81452]_ , \new_[81455]_ , \new_[81456]_ , \new_[81457]_ ,
    \new_[81460]_ , \new_[81463]_ , \new_[81464]_ , \new_[81467]_ ,
    \new_[81470]_ , \new_[81471]_ , \new_[81472]_ , \new_[81476]_ ,
    \new_[81477]_ , \new_[81480]_ , \new_[81483]_ , \new_[81484]_ ,
    \new_[81485]_ , \new_[81488]_ , \new_[81491]_ , \new_[81492]_ ,
    \new_[81495]_ , \new_[81498]_ , \new_[81499]_ , \new_[81500]_ ,
    \new_[81504]_ , \new_[81505]_ , \new_[81508]_ , \new_[81511]_ ,
    \new_[81512]_ , \new_[81513]_ , \new_[81516]_ , \new_[81519]_ ,
    \new_[81520]_ , \new_[81523]_ , \new_[81526]_ , \new_[81527]_ ,
    \new_[81528]_ , \new_[81532]_ , \new_[81533]_ , \new_[81536]_ ,
    \new_[81539]_ , \new_[81540]_ , \new_[81541]_ , \new_[81544]_ ,
    \new_[81547]_ , \new_[81548]_ , \new_[81551]_ , \new_[81554]_ ,
    \new_[81555]_ , \new_[81556]_ , \new_[81560]_ , \new_[81561]_ ,
    \new_[81564]_ , \new_[81567]_ , \new_[81568]_ , \new_[81569]_ ,
    \new_[81572]_ , \new_[81575]_ , \new_[81576]_ , \new_[81579]_ ,
    \new_[81582]_ , \new_[81583]_ , \new_[81584]_ , \new_[81588]_ ,
    \new_[81589]_ , \new_[81592]_ , \new_[81595]_ , \new_[81596]_ ,
    \new_[81597]_ , \new_[81600]_ , \new_[81603]_ , \new_[81604]_ ,
    \new_[81607]_ , \new_[81610]_ , \new_[81611]_ , \new_[81612]_ ,
    \new_[81616]_ , \new_[81617]_ , \new_[81620]_ , \new_[81623]_ ,
    \new_[81624]_ , \new_[81625]_ , \new_[81628]_ , \new_[81631]_ ,
    \new_[81632]_ , \new_[81635]_ , \new_[81638]_ , \new_[81639]_ ,
    \new_[81640]_ , \new_[81644]_ , \new_[81645]_ , \new_[81648]_ ,
    \new_[81651]_ , \new_[81652]_ , \new_[81653]_ , \new_[81656]_ ,
    \new_[81659]_ , \new_[81660]_ , \new_[81663]_ , \new_[81666]_ ,
    \new_[81667]_ , \new_[81668]_ , \new_[81672]_ , \new_[81673]_ ,
    \new_[81676]_ , \new_[81679]_ , \new_[81680]_ , \new_[81681]_ ,
    \new_[81684]_ , \new_[81687]_ , \new_[81688]_ , \new_[81691]_ ,
    \new_[81694]_ , \new_[81695]_ , \new_[81696]_ , \new_[81700]_ ,
    \new_[81701]_ , \new_[81704]_ , \new_[81707]_ , \new_[81708]_ ,
    \new_[81709]_ , \new_[81712]_ , \new_[81715]_ , \new_[81716]_ ,
    \new_[81719]_ , \new_[81722]_ , \new_[81723]_ , \new_[81724]_ ,
    \new_[81728]_ , \new_[81729]_ , \new_[81732]_ , \new_[81735]_ ,
    \new_[81736]_ , \new_[81737]_ , \new_[81740]_ , \new_[81743]_ ,
    \new_[81744]_ , \new_[81747]_ , \new_[81750]_ , \new_[81751]_ ,
    \new_[81752]_ , \new_[81756]_ , \new_[81757]_ , \new_[81760]_ ,
    \new_[81763]_ , \new_[81764]_ , \new_[81765]_ , \new_[81768]_ ,
    \new_[81771]_ , \new_[81772]_ , \new_[81775]_ , \new_[81778]_ ,
    \new_[81779]_ , \new_[81780]_ , \new_[81784]_ , \new_[81785]_ ,
    \new_[81788]_ , \new_[81791]_ , \new_[81792]_ , \new_[81793]_ ,
    \new_[81796]_ , \new_[81799]_ , \new_[81800]_ , \new_[81803]_ ,
    \new_[81806]_ , \new_[81807]_ , \new_[81808]_ , \new_[81812]_ ,
    \new_[81813]_ , \new_[81816]_ , \new_[81819]_ , \new_[81820]_ ,
    \new_[81821]_ , \new_[81824]_ , \new_[81827]_ , \new_[81828]_ ,
    \new_[81831]_ , \new_[81834]_ , \new_[81835]_ , \new_[81836]_ ,
    \new_[81840]_ , \new_[81841]_ , \new_[81844]_ , \new_[81847]_ ,
    \new_[81848]_ , \new_[81849]_ , \new_[81852]_ , \new_[81855]_ ,
    \new_[81856]_ , \new_[81859]_ , \new_[81862]_ , \new_[81863]_ ,
    \new_[81864]_ , \new_[81868]_ , \new_[81869]_ , \new_[81872]_ ,
    \new_[81875]_ , \new_[81876]_ , \new_[81877]_ , \new_[81880]_ ,
    \new_[81883]_ , \new_[81884]_ , \new_[81887]_ , \new_[81890]_ ,
    \new_[81891]_ , \new_[81892]_ , \new_[81896]_ , \new_[81897]_ ,
    \new_[81900]_ , \new_[81903]_ , \new_[81904]_ , \new_[81905]_ ,
    \new_[81908]_ , \new_[81911]_ , \new_[81912]_ , \new_[81915]_ ,
    \new_[81918]_ , \new_[81919]_ , \new_[81920]_ , \new_[81924]_ ,
    \new_[81925]_ , \new_[81928]_ , \new_[81931]_ , \new_[81932]_ ,
    \new_[81933]_ , \new_[81936]_ , \new_[81939]_ , \new_[81940]_ ,
    \new_[81943]_ , \new_[81946]_ , \new_[81947]_ , \new_[81948]_ ,
    \new_[81952]_ , \new_[81953]_ , \new_[81956]_ , \new_[81959]_ ,
    \new_[81960]_ , \new_[81961]_ , \new_[81964]_ , \new_[81967]_ ,
    \new_[81968]_ , \new_[81971]_ , \new_[81974]_ , \new_[81975]_ ,
    \new_[81976]_ , \new_[81980]_ , \new_[81981]_ , \new_[81984]_ ,
    \new_[81987]_ , \new_[81988]_ , \new_[81989]_ , \new_[81992]_ ,
    \new_[81995]_ , \new_[81996]_ , \new_[81999]_ , \new_[82002]_ ,
    \new_[82003]_ , \new_[82004]_ , \new_[82008]_ , \new_[82009]_ ,
    \new_[82012]_ , \new_[82015]_ , \new_[82016]_ , \new_[82017]_ ,
    \new_[82020]_ , \new_[82023]_ , \new_[82024]_ , \new_[82027]_ ,
    \new_[82030]_ , \new_[82031]_ , \new_[82032]_ , \new_[82036]_ ,
    \new_[82037]_ , \new_[82040]_ , \new_[82043]_ , \new_[82044]_ ,
    \new_[82045]_ , \new_[82048]_ , \new_[82051]_ , \new_[82052]_ ,
    \new_[82055]_ , \new_[82058]_ , \new_[82059]_ , \new_[82060]_ ,
    \new_[82064]_ , \new_[82065]_ , \new_[82068]_ , \new_[82071]_ ,
    \new_[82072]_ , \new_[82073]_ , \new_[82076]_ , \new_[82079]_ ,
    \new_[82080]_ , \new_[82083]_ , \new_[82086]_ , \new_[82087]_ ,
    \new_[82088]_ , \new_[82092]_ , \new_[82093]_ , \new_[82096]_ ,
    \new_[82099]_ , \new_[82100]_ , \new_[82101]_ , \new_[82104]_ ,
    \new_[82107]_ , \new_[82108]_ , \new_[82111]_ , \new_[82114]_ ,
    \new_[82115]_ , \new_[82116]_ , \new_[82120]_ , \new_[82121]_ ,
    \new_[82124]_ , \new_[82127]_ , \new_[82128]_ , \new_[82129]_ ,
    \new_[82132]_ , \new_[82135]_ , \new_[82136]_ , \new_[82139]_ ,
    \new_[82142]_ , \new_[82143]_ , \new_[82144]_ , \new_[82148]_ ,
    \new_[82149]_ , \new_[82152]_ , \new_[82155]_ , \new_[82156]_ ,
    \new_[82157]_ , \new_[82160]_ , \new_[82163]_ , \new_[82164]_ ,
    \new_[82167]_ , \new_[82170]_ , \new_[82171]_ , \new_[82172]_ ,
    \new_[82176]_ , \new_[82177]_ , \new_[82180]_ , \new_[82183]_ ,
    \new_[82184]_ , \new_[82185]_ , \new_[82188]_ , \new_[82191]_ ,
    \new_[82192]_ , \new_[82195]_ , \new_[82198]_ , \new_[82199]_ ,
    \new_[82200]_ , \new_[82204]_ , \new_[82205]_ , \new_[82208]_ ,
    \new_[82211]_ , \new_[82212]_ , \new_[82213]_ , \new_[82216]_ ,
    \new_[82219]_ , \new_[82220]_ , \new_[82223]_ , \new_[82226]_ ,
    \new_[82227]_ , \new_[82228]_ , \new_[82232]_ , \new_[82233]_ ,
    \new_[82236]_ , \new_[82239]_ , \new_[82240]_ , \new_[82241]_ ,
    \new_[82244]_ , \new_[82247]_ , \new_[82248]_ , \new_[82251]_ ,
    \new_[82254]_ , \new_[82255]_ , \new_[82256]_ , \new_[82260]_ ,
    \new_[82261]_ , \new_[82264]_ , \new_[82267]_ , \new_[82268]_ ,
    \new_[82269]_ , \new_[82272]_ , \new_[82275]_ , \new_[82276]_ ,
    \new_[82279]_ , \new_[82282]_ , \new_[82283]_ , \new_[82284]_ ,
    \new_[82288]_ , \new_[82289]_ , \new_[82292]_ , \new_[82295]_ ,
    \new_[82296]_ , \new_[82297]_ , \new_[82300]_ , \new_[82303]_ ,
    \new_[82304]_ , \new_[82307]_ , \new_[82310]_ , \new_[82311]_ ,
    \new_[82312]_ , \new_[82316]_ , \new_[82317]_ , \new_[82320]_ ,
    \new_[82323]_ , \new_[82324]_ , \new_[82325]_ , \new_[82328]_ ,
    \new_[82331]_ , \new_[82332]_ , \new_[82335]_ , \new_[82338]_ ,
    \new_[82339]_ , \new_[82340]_ , \new_[82344]_ , \new_[82345]_ ,
    \new_[82348]_ , \new_[82351]_ , \new_[82352]_ , \new_[82353]_ ,
    \new_[82356]_ , \new_[82359]_ , \new_[82360]_ , \new_[82363]_ ,
    \new_[82366]_ , \new_[82367]_ , \new_[82368]_ , \new_[82372]_ ,
    \new_[82373]_ , \new_[82376]_ , \new_[82379]_ , \new_[82380]_ ,
    \new_[82381]_ , \new_[82384]_ , \new_[82387]_ , \new_[82388]_ ,
    \new_[82391]_ , \new_[82394]_ , \new_[82395]_ , \new_[82396]_ ,
    \new_[82400]_ , \new_[82401]_ , \new_[82404]_ , \new_[82407]_ ,
    \new_[82408]_ , \new_[82409]_ , \new_[82412]_ , \new_[82415]_ ,
    \new_[82416]_ , \new_[82419]_ , \new_[82422]_ , \new_[82423]_ ,
    \new_[82424]_ , \new_[82428]_ , \new_[82429]_ , \new_[82432]_ ,
    \new_[82435]_ , \new_[82436]_ , \new_[82437]_ , \new_[82440]_ ,
    \new_[82443]_ , \new_[82444]_ , \new_[82447]_ , \new_[82450]_ ,
    \new_[82451]_ , \new_[82452]_ , \new_[82456]_ , \new_[82457]_ ,
    \new_[82460]_ , \new_[82463]_ , \new_[82464]_ , \new_[82465]_ ,
    \new_[82468]_ , \new_[82471]_ , \new_[82472]_ , \new_[82475]_ ,
    \new_[82478]_ , \new_[82479]_ , \new_[82480]_ , \new_[82484]_ ,
    \new_[82485]_ , \new_[82488]_ , \new_[82491]_ , \new_[82492]_ ,
    \new_[82493]_ , \new_[82496]_ , \new_[82499]_ , \new_[82500]_ ,
    \new_[82503]_ , \new_[82506]_ , \new_[82507]_ , \new_[82508]_ ,
    \new_[82512]_ , \new_[82513]_ , \new_[82516]_ , \new_[82519]_ ,
    \new_[82520]_ , \new_[82521]_ , \new_[82524]_ , \new_[82527]_ ,
    \new_[82528]_ , \new_[82531]_ , \new_[82534]_ , \new_[82535]_ ,
    \new_[82536]_ , \new_[82540]_ , \new_[82541]_ , \new_[82544]_ ,
    \new_[82547]_ , \new_[82548]_ , \new_[82549]_ , \new_[82552]_ ,
    \new_[82555]_ , \new_[82556]_ , \new_[82559]_ , \new_[82562]_ ,
    \new_[82563]_ , \new_[82564]_ , \new_[82568]_ , \new_[82569]_ ,
    \new_[82572]_ , \new_[82575]_ , \new_[82576]_ , \new_[82577]_ ,
    \new_[82580]_ , \new_[82583]_ , \new_[82584]_ , \new_[82587]_ ,
    \new_[82590]_ , \new_[82591]_ , \new_[82592]_ , \new_[82596]_ ,
    \new_[82597]_ , \new_[82600]_ , \new_[82603]_ , \new_[82604]_ ,
    \new_[82605]_ , \new_[82608]_ , \new_[82611]_ , \new_[82612]_ ,
    \new_[82615]_ , \new_[82618]_ , \new_[82619]_ , \new_[82620]_ ,
    \new_[82624]_ , \new_[82625]_ , \new_[82628]_ , \new_[82631]_ ,
    \new_[82632]_ , \new_[82633]_ , \new_[82636]_ , \new_[82639]_ ,
    \new_[82640]_ , \new_[82643]_ , \new_[82646]_ , \new_[82647]_ ,
    \new_[82648]_ , \new_[82652]_ , \new_[82653]_ , \new_[82656]_ ,
    \new_[82659]_ , \new_[82660]_ , \new_[82661]_ , \new_[82664]_ ,
    \new_[82667]_ , \new_[82668]_ , \new_[82671]_ , \new_[82674]_ ,
    \new_[82675]_ , \new_[82676]_ , \new_[82680]_ , \new_[82681]_ ,
    \new_[82684]_ , \new_[82687]_ , \new_[82688]_ , \new_[82689]_ ,
    \new_[82692]_ , \new_[82695]_ , \new_[82696]_ , \new_[82699]_ ,
    \new_[82702]_ , \new_[82703]_ , \new_[82704]_ , \new_[82708]_ ,
    \new_[82709]_ , \new_[82712]_ , \new_[82715]_ , \new_[82716]_ ,
    \new_[82717]_ , \new_[82720]_ , \new_[82723]_ , \new_[82724]_ ,
    \new_[82727]_ , \new_[82730]_ , \new_[82731]_ , \new_[82732]_ ,
    \new_[82736]_ , \new_[82737]_ , \new_[82740]_ , \new_[82743]_ ,
    \new_[82744]_ , \new_[82745]_ , \new_[82748]_ , \new_[82751]_ ,
    \new_[82752]_ , \new_[82755]_ , \new_[82758]_ , \new_[82759]_ ,
    \new_[82760]_ , \new_[82764]_ , \new_[82765]_ , \new_[82768]_ ,
    \new_[82771]_ , \new_[82772]_ , \new_[82773]_ , \new_[82776]_ ,
    \new_[82779]_ , \new_[82780]_ , \new_[82783]_ , \new_[82786]_ ,
    \new_[82787]_ , \new_[82788]_ , \new_[82792]_ , \new_[82793]_ ,
    \new_[82796]_ , \new_[82799]_ , \new_[82800]_ , \new_[82801]_ ,
    \new_[82804]_ , \new_[82807]_ , \new_[82808]_ , \new_[82811]_ ,
    \new_[82814]_ , \new_[82815]_ , \new_[82816]_ , \new_[82820]_ ,
    \new_[82821]_ , \new_[82824]_ , \new_[82827]_ , \new_[82828]_ ,
    \new_[82829]_ , \new_[82832]_ , \new_[82835]_ , \new_[82836]_ ,
    \new_[82839]_ , \new_[82842]_ , \new_[82843]_ , \new_[82844]_ ,
    \new_[82848]_ , \new_[82849]_ , \new_[82852]_ , \new_[82855]_ ,
    \new_[82856]_ , \new_[82857]_ , \new_[82860]_ , \new_[82863]_ ,
    \new_[82864]_ , \new_[82867]_ , \new_[82870]_ , \new_[82871]_ ,
    \new_[82872]_ , \new_[82876]_ , \new_[82877]_ , \new_[82880]_ ,
    \new_[82883]_ , \new_[82884]_ , \new_[82885]_ , \new_[82888]_ ,
    \new_[82891]_ , \new_[82892]_ , \new_[82895]_ , \new_[82898]_ ,
    \new_[82899]_ , \new_[82900]_ , \new_[82904]_ , \new_[82905]_ ,
    \new_[82908]_ , \new_[82911]_ , \new_[82912]_ , \new_[82913]_ ,
    \new_[82916]_ , \new_[82919]_ , \new_[82920]_ , \new_[82923]_ ,
    \new_[82926]_ , \new_[82927]_ , \new_[82928]_ , \new_[82932]_ ,
    \new_[82933]_ , \new_[82936]_ , \new_[82939]_ , \new_[82940]_ ,
    \new_[82941]_ , \new_[82944]_ , \new_[82947]_ , \new_[82948]_ ,
    \new_[82951]_ , \new_[82954]_ , \new_[82955]_ , \new_[82956]_ ,
    \new_[82960]_ , \new_[82961]_ , \new_[82964]_ , \new_[82967]_ ,
    \new_[82968]_ , \new_[82969]_ , \new_[82972]_ , \new_[82975]_ ,
    \new_[82976]_ , \new_[82979]_ , \new_[82982]_ , \new_[82983]_ ,
    \new_[82984]_ , \new_[82988]_ , \new_[82989]_ , \new_[82992]_ ,
    \new_[82995]_ , \new_[82996]_ , \new_[82997]_ , \new_[83000]_ ,
    \new_[83003]_ , \new_[83004]_ , \new_[83007]_ , \new_[83010]_ ,
    \new_[83011]_ , \new_[83012]_ , \new_[83016]_ , \new_[83017]_ ,
    \new_[83020]_ , \new_[83023]_ , \new_[83024]_ , \new_[83025]_ ,
    \new_[83028]_ , \new_[83031]_ , \new_[83032]_ , \new_[83035]_ ,
    \new_[83038]_ , \new_[83039]_ , \new_[83040]_ , \new_[83044]_ ,
    \new_[83045]_ , \new_[83048]_ , \new_[83051]_ , \new_[83052]_ ,
    \new_[83053]_ , \new_[83056]_ , \new_[83059]_ , \new_[83060]_ ,
    \new_[83063]_ , \new_[83066]_ , \new_[83067]_ , \new_[83068]_ ,
    \new_[83072]_ , \new_[83073]_ , \new_[83076]_ , \new_[83079]_ ,
    \new_[83080]_ , \new_[83081]_ , \new_[83084]_ , \new_[83087]_ ,
    \new_[83088]_ , \new_[83091]_ , \new_[83094]_ , \new_[83095]_ ,
    \new_[83096]_ , \new_[83100]_ , \new_[83101]_ , \new_[83104]_ ,
    \new_[83107]_ , \new_[83108]_ , \new_[83109]_ , \new_[83112]_ ,
    \new_[83115]_ , \new_[83116]_ , \new_[83119]_ , \new_[83122]_ ,
    \new_[83123]_ , \new_[83124]_ , \new_[83128]_ , \new_[83129]_ ,
    \new_[83132]_ , \new_[83135]_ , \new_[83136]_ , \new_[83137]_ ,
    \new_[83140]_ , \new_[83143]_ , \new_[83144]_ , \new_[83147]_ ,
    \new_[83150]_ , \new_[83151]_ , \new_[83152]_ , \new_[83156]_ ,
    \new_[83157]_ , \new_[83160]_ , \new_[83163]_ , \new_[83164]_ ,
    \new_[83165]_ , \new_[83168]_ , \new_[83171]_ , \new_[83172]_ ,
    \new_[83175]_ , \new_[83178]_ , \new_[83179]_ , \new_[83180]_ ,
    \new_[83184]_ , \new_[83185]_ , \new_[83188]_ , \new_[83191]_ ,
    \new_[83192]_ , \new_[83193]_ , \new_[83196]_ , \new_[83199]_ ,
    \new_[83200]_ , \new_[83203]_ , \new_[83206]_ , \new_[83207]_ ,
    \new_[83208]_ , \new_[83212]_ , \new_[83213]_ , \new_[83216]_ ,
    \new_[83219]_ , \new_[83220]_ , \new_[83221]_ , \new_[83224]_ ,
    \new_[83227]_ , \new_[83228]_ , \new_[83231]_ , \new_[83234]_ ,
    \new_[83235]_ , \new_[83236]_ , \new_[83240]_ , \new_[83241]_ ,
    \new_[83244]_ , \new_[83247]_ , \new_[83248]_ , \new_[83249]_ ,
    \new_[83252]_ , \new_[83255]_ , \new_[83256]_ , \new_[83259]_ ,
    \new_[83262]_ , \new_[83263]_ , \new_[83264]_ , \new_[83268]_ ,
    \new_[83269]_ , \new_[83272]_ , \new_[83275]_ , \new_[83276]_ ,
    \new_[83277]_ , \new_[83280]_ , \new_[83283]_ , \new_[83284]_ ,
    \new_[83287]_ , \new_[83290]_ , \new_[83291]_ , \new_[83292]_ ,
    \new_[83296]_ , \new_[83297]_ , \new_[83300]_ , \new_[83303]_ ,
    \new_[83304]_ , \new_[83305]_ , \new_[83308]_ , \new_[83311]_ ,
    \new_[83312]_ , \new_[83315]_ , \new_[83318]_ , \new_[83319]_ ,
    \new_[83320]_ , \new_[83324]_ , \new_[83325]_ , \new_[83328]_ ,
    \new_[83331]_ , \new_[83332]_ , \new_[83333]_ , \new_[83336]_ ,
    \new_[83339]_ , \new_[83340]_ , \new_[83343]_ , \new_[83346]_ ,
    \new_[83347]_ , \new_[83348]_ , \new_[83352]_ , \new_[83353]_ ,
    \new_[83356]_ , \new_[83359]_ , \new_[83360]_ , \new_[83361]_ ,
    \new_[83364]_ , \new_[83367]_ , \new_[83368]_ , \new_[83371]_ ,
    \new_[83374]_ , \new_[83375]_ , \new_[83376]_ , \new_[83380]_ ,
    \new_[83381]_ , \new_[83384]_ , \new_[83387]_ , \new_[83388]_ ,
    \new_[83389]_ , \new_[83392]_ , \new_[83395]_ , \new_[83396]_ ,
    \new_[83399]_ , \new_[83402]_ , \new_[83403]_ , \new_[83404]_ ,
    \new_[83408]_ , \new_[83409]_ , \new_[83412]_ , \new_[83415]_ ,
    \new_[83416]_ , \new_[83417]_ , \new_[83420]_ , \new_[83423]_ ,
    \new_[83424]_ , \new_[83427]_ , \new_[83430]_ , \new_[83431]_ ,
    \new_[83432]_ , \new_[83436]_ , \new_[83437]_ , \new_[83440]_ ,
    \new_[83443]_ , \new_[83444]_ , \new_[83445]_ , \new_[83448]_ ,
    \new_[83451]_ , \new_[83452]_ , \new_[83455]_ , \new_[83458]_ ,
    \new_[83459]_ , \new_[83460]_ , \new_[83464]_ , \new_[83465]_ ,
    \new_[83468]_ , \new_[83471]_ , \new_[83472]_ , \new_[83473]_ ,
    \new_[83476]_ , \new_[83479]_ , \new_[83480]_ , \new_[83483]_ ,
    \new_[83486]_ , \new_[83487]_ , \new_[83488]_ , \new_[83492]_ ,
    \new_[83493]_ , \new_[83496]_ , \new_[83499]_ , \new_[83500]_ ,
    \new_[83501]_ , \new_[83504]_ , \new_[83507]_ , \new_[83508]_ ,
    \new_[83511]_ , \new_[83514]_ , \new_[83515]_ , \new_[83516]_ ,
    \new_[83520]_ , \new_[83521]_ , \new_[83524]_ , \new_[83527]_ ,
    \new_[83528]_ , \new_[83529]_ , \new_[83532]_ , \new_[83535]_ ,
    \new_[83536]_ , \new_[83539]_ , \new_[83542]_ , \new_[83543]_ ,
    \new_[83544]_ , \new_[83548]_ , \new_[83549]_ , \new_[83552]_ ,
    \new_[83555]_ , \new_[83556]_ , \new_[83557]_ , \new_[83560]_ ,
    \new_[83563]_ , \new_[83564]_ , \new_[83567]_ , \new_[83570]_ ,
    \new_[83571]_ , \new_[83572]_ , \new_[83576]_ , \new_[83577]_ ,
    \new_[83580]_ , \new_[83583]_ , \new_[83584]_ , \new_[83585]_ ,
    \new_[83588]_ , \new_[83591]_ , \new_[83592]_ , \new_[83595]_ ,
    \new_[83598]_ , \new_[83599]_ , \new_[83600]_ , \new_[83604]_ ,
    \new_[83605]_ , \new_[83608]_ , \new_[83611]_ , \new_[83612]_ ,
    \new_[83613]_ , \new_[83616]_ , \new_[83619]_ , \new_[83620]_ ,
    \new_[83623]_ , \new_[83626]_ , \new_[83627]_ , \new_[83628]_ ,
    \new_[83632]_ , \new_[83633]_ , \new_[83636]_ , \new_[83639]_ ,
    \new_[83640]_ , \new_[83641]_ , \new_[83644]_ , \new_[83647]_ ,
    \new_[83648]_ , \new_[83651]_ , \new_[83654]_ , \new_[83655]_ ,
    \new_[83656]_ , \new_[83660]_ , \new_[83661]_ , \new_[83664]_ ,
    \new_[83667]_ , \new_[83668]_ , \new_[83669]_ , \new_[83672]_ ,
    \new_[83675]_ , \new_[83676]_ , \new_[83679]_ , \new_[83682]_ ,
    \new_[83683]_ , \new_[83684]_ , \new_[83688]_ , \new_[83689]_ ,
    \new_[83692]_ , \new_[83695]_ , \new_[83696]_ , \new_[83697]_ ,
    \new_[83700]_ , \new_[83703]_ , \new_[83704]_ , \new_[83707]_ ,
    \new_[83710]_ , \new_[83711]_ , \new_[83712]_ , \new_[83716]_ ,
    \new_[83717]_ , \new_[83720]_ , \new_[83723]_ , \new_[83724]_ ,
    \new_[83725]_ , \new_[83728]_ , \new_[83731]_ , \new_[83732]_ ,
    \new_[83735]_ , \new_[83738]_ , \new_[83739]_ , \new_[83740]_ ,
    \new_[83744]_ , \new_[83745]_ , \new_[83748]_ , \new_[83751]_ ,
    \new_[83752]_ , \new_[83753]_ , \new_[83756]_ , \new_[83759]_ ,
    \new_[83760]_ , \new_[83763]_ , \new_[83766]_ , \new_[83767]_ ,
    \new_[83768]_ , \new_[83772]_ , \new_[83773]_ , \new_[83776]_ ,
    \new_[83779]_ , \new_[83780]_ , \new_[83781]_ , \new_[83784]_ ,
    \new_[83787]_ , \new_[83788]_ , \new_[83791]_ , \new_[83794]_ ,
    \new_[83795]_ , \new_[83796]_ , \new_[83800]_ , \new_[83801]_ ,
    \new_[83804]_ , \new_[83807]_ , \new_[83808]_ , \new_[83809]_ ,
    \new_[83812]_ , \new_[83815]_ , \new_[83816]_ , \new_[83819]_ ,
    \new_[83822]_ , \new_[83823]_ , \new_[83824]_ , \new_[83828]_ ,
    \new_[83829]_ , \new_[83832]_ , \new_[83835]_ , \new_[83836]_ ,
    \new_[83837]_ , \new_[83840]_ , \new_[83843]_ , \new_[83844]_ ,
    \new_[83847]_ , \new_[83850]_ , \new_[83851]_ , \new_[83852]_ ,
    \new_[83856]_ , \new_[83857]_ , \new_[83860]_ , \new_[83863]_ ,
    \new_[83864]_ , \new_[83865]_ , \new_[83868]_ , \new_[83871]_ ,
    \new_[83872]_ , \new_[83875]_ , \new_[83878]_ , \new_[83879]_ ,
    \new_[83880]_ , \new_[83884]_ , \new_[83885]_ , \new_[83888]_ ,
    \new_[83891]_ , \new_[83892]_ , \new_[83893]_ , \new_[83896]_ ,
    \new_[83899]_ , \new_[83900]_ , \new_[83903]_ , \new_[83906]_ ,
    \new_[83907]_ , \new_[83908]_ , \new_[83912]_ , \new_[83913]_ ,
    \new_[83916]_ , \new_[83919]_ , \new_[83920]_ , \new_[83921]_ ,
    \new_[83924]_ , \new_[83927]_ , \new_[83928]_ , \new_[83931]_ ,
    \new_[83934]_ , \new_[83935]_ , \new_[83936]_ , \new_[83940]_ ,
    \new_[83941]_ , \new_[83944]_ , \new_[83947]_ , \new_[83948]_ ,
    \new_[83949]_ , \new_[83952]_ , \new_[83955]_ , \new_[83956]_ ,
    \new_[83959]_ , \new_[83962]_ , \new_[83963]_ , \new_[83964]_ ,
    \new_[83968]_ , \new_[83969]_ , \new_[83972]_ , \new_[83975]_ ,
    \new_[83976]_ , \new_[83977]_ , \new_[83980]_ , \new_[83983]_ ,
    \new_[83984]_ , \new_[83987]_ , \new_[83990]_ , \new_[83991]_ ,
    \new_[83992]_ , \new_[83996]_ , \new_[83997]_ , \new_[84000]_ ,
    \new_[84003]_ , \new_[84004]_ , \new_[84005]_ , \new_[84008]_ ,
    \new_[84011]_ , \new_[84012]_ , \new_[84015]_ , \new_[84018]_ ,
    \new_[84019]_ , \new_[84020]_ , \new_[84024]_ , \new_[84025]_ ,
    \new_[84028]_ , \new_[84031]_ , \new_[84032]_ , \new_[84033]_ ,
    \new_[84036]_ , \new_[84039]_ , \new_[84040]_ , \new_[84043]_ ,
    \new_[84046]_ , \new_[84047]_ , \new_[84048]_ , \new_[84052]_ ,
    \new_[84053]_ , \new_[84056]_ , \new_[84059]_ , \new_[84060]_ ,
    \new_[84061]_ , \new_[84064]_ , \new_[84067]_ , \new_[84068]_ ,
    \new_[84071]_ , \new_[84074]_ , \new_[84075]_ , \new_[84076]_ ,
    \new_[84080]_ , \new_[84081]_ , \new_[84084]_ , \new_[84087]_ ,
    \new_[84088]_ , \new_[84089]_ , \new_[84092]_ , \new_[84095]_ ,
    \new_[84096]_ , \new_[84099]_ , \new_[84102]_ , \new_[84103]_ ,
    \new_[84104]_ , \new_[84108]_ , \new_[84109]_ , \new_[84112]_ ,
    \new_[84115]_ , \new_[84116]_ , \new_[84117]_ , \new_[84120]_ ,
    \new_[84123]_ , \new_[84124]_ , \new_[84127]_ , \new_[84130]_ ,
    \new_[84131]_ , \new_[84132]_ , \new_[84136]_ , \new_[84137]_ ,
    \new_[84140]_ , \new_[84143]_ , \new_[84144]_ , \new_[84145]_ ,
    \new_[84148]_ , \new_[84151]_ , \new_[84152]_ , \new_[84155]_ ,
    \new_[84158]_ , \new_[84159]_ , \new_[84160]_ , \new_[84164]_ ,
    \new_[84165]_ , \new_[84168]_ , \new_[84171]_ , \new_[84172]_ ,
    \new_[84173]_ , \new_[84176]_ , \new_[84179]_ , \new_[84180]_ ,
    \new_[84183]_ , \new_[84186]_ , \new_[84187]_ , \new_[84188]_ ,
    \new_[84192]_ , \new_[84193]_ , \new_[84196]_ , \new_[84199]_ ,
    \new_[84200]_ , \new_[84201]_ , \new_[84204]_ , \new_[84207]_ ,
    \new_[84208]_ , \new_[84211]_ , \new_[84214]_ , \new_[84215]_ ,
    \new_[84216]_ , \new_[84220]_ , \new_[84221]_ , \new_[84224]_ ,
    \new_[84227]_ , \new_[84228]_ , \new_[84229]_ , \new_[84232]_ ,
    \new_[84235]_ , \new_[84236]_ , \new_[84239]_ , \new_[84242]_ ,
    \new_[84243]_ , \new_[84244]_ , \new_[84248]_ , \new_[84249]_ ,
    \new_[84252]_ , \new_[84255]_ , \new_[84256]_ , \new_[84257]_ ,
    \new_[84260]_ , \new_[84263]_ , \new_[84264]_ , \new_[84267]_ ,
    \new_[84270]_ , \new_[84271]_ , \new_[84272]_ , \new_[84276]_ ,
    \new_[84277]_ , \new_[84280]_ , \new_[84283]_ , \new_[84284]_ ,
    \new_[84285]_ , \new_[84288]_ , \new_[84291]_ , \new_[84292]_ ,
    \new_[84295]_ , \new_[84298]_ , \new_[84299]_ , \new_[84300]_ ,
    \new_[84304]_ , \new_[84305]_ , \new_[84308]_ , \new_[84311]_ ,
    \new_[84312]_ , \new_[84313]_ , \new_[84316]_ , \new_[84319]_ ,
    \new_[84320]_ , \new_[84323]_ , \new_[84326]_ , \new_[84327]_ ,
    \new_[84328]_ , \new_[84332]_ , \new_[84333]_ , \new_[84336]_ ,
    \new_[84339]_ , \new_[84340]_ , \new_[84341]_ , \new_[84344]_ ,
    \new_[84347]_ , \new_[84348]_ , \new_[84351]_ , \new_[84354]_ ,
    \new_[84355]_ , \new_[84356]_ , \new_[84360]_ , \new_[84361]_ ,
    \new_[84364]_ , \new_[84367]_ , \new_[84368]_ , \new_[84369]_ ,
    \new_[84372]_ , \new_[84375]_ , \new_[84376]_ , \new_[84379]_ ,
    \new_[84382]_ , \new_[84383]_ , \new_[84384]_ , \new_[84388]_ ,
    \new_[84389]_ , \new_[84392]_ , \new_[84395]_ , \new_[84396]_ ,
    \new_[84397]_ , \new_[84400]_ , \new_[84403]_ , \new_[84404]_ ,
    \new_[84407]_ , \new_[84410]_ , \new_[84411]_ , \new_[84412]_ ,
    \new_[84416]_ , \new_[84417]_ , \new_[84420]_ , \new_[84423]_ ,
    \new_[84424]_ , \new_[84425]_ , \new_[84428]_ , \new_[84431]_ ,
    \new_[84432]_ , \new_[84435]_ , \new_[84438]_ , \new_[84439]_ ,
    \new_[84440]_ , \new_[84444]_ , \new_[84445]_ , \new_[84448]_ ,
    \new_[84451]_ , \new_[84452]_ , \new_[84453]_ , \new_[84456]_ ,
    \new_[84459]_ , \new_[84460]_ , \new_[84463]_ , \new_[84466]_ ,
    \new_[84467]_ , \new_[84468]_ , \new_[84472]_ , \new_[84473]_ ,
    \new_[84476]_ , \new_[84479]_ , \new_[84480]_ , \new_[84481]_ ,
    \new_[84484]_ , \new_[84487]_ , \new_[84488]_ , \new_[84491]_ ,
    \new_[84494]_ , \new_[84495]_ , \new_[84496]_ , \new_[84500]_ ,
    \new_[84501]_ , \new_[84504]_ , \new_[84507]_ , \new_[84508]_ ,
    \new_[84509]_ , \new_[84512]_ , \new_[84515]_ , \new_[84516]_ ,
    \new_[84519]_ , \new_[84522]_ , \new_[84523]_ , \new_[84524]_ ,
    \new_[84528]_ , \new_[84529]_ , \new_[84532]_ , \new_[84535]_ ,
    \new_[84536]_ , \new_[84537]_ , \new_[84540]_ , \new_[84543]_ ,
    \new_[84544]_ , \new_[84547]_ , \new_[84550]_ , \new_[84551]_ ,
    \new_[84552]_ , \new_[84556]_ , \new_[84557]_ , \new_[84560]_ ,
    \new_[84563]_ , \new_[84564]_ , \new_[84565]_ , \new_[84568]_ ,
    \new_[84571]_ , \new_[84572]_ , \new_[84575]_ , \new_[84578]_ ,
    \new_[84579]_ , \new_[84580]_ , \new_[84584]_ , \new_[84585]_ ,
    \new_[84588]_ , \new_[84591]_ , \new_[84592]_ , \new_[84593]_ ,
    \new_[84596]_ , \new_[84599]_ , \new_[84600]_ , \new_[84603]_ ,
    \new_[84606]_ , \new_[84607]_ , \new_[84608]_ , \new_[84612]_ ,
    \new_[84613]_ , \new_[84616]_ , \new_[84619]_ , \new_[84620]_ ,
    \new_[84621]_ , \new_[84624]_ , \new_[84627]_ , \new_[84628]_ ,
    \new_[84631]_ , \new_[84634]_ , \new_[84635]_ , \new_[84636]_ ,
    \new_[84640]_ , \new_[84641]_ , \new_[84644]_ , \new_[84647]_ ,
    \new_[84648]_ , \new_[84649]_ , \new_[84652]_ , \new_[84655]_ ,
    \new_[84656]_ , \new_[84659]_ , \new_[84662]_ , \new_[84663]_ ,
    \new_[84664]_ , \new_[84668]_ , \new_[84669]_ , \new_[84672]_ ,
    \new_[84675]_ , \new_[84676]_ , \new_[84677]_ , \new_[84680]_ ,
    \new_[84683]_ , \new_[84684]_ , \new_[84687]_ , \new_[84690]_ ,
    \new_[84691]_ , \new_[84692]_ , \new_[84696]_ , \new_[84697]_ ,
    \new_[84700]_ , \new_[84703]_ , \new_[84704]_ , \new_[84705]_ ,
    \new_[84708]_ , \new_[84711]_ , \new_[84712]_ , \new_[84715]_ ,
    \new_[84718]_ , \new_[84719]_ , \new_[84720]_ , \new_[84724]_ ,
    \new_[84725]_ , \new_[84728]_ , \new_[84731]_ , \new_[84732]_ ,
    \new_[84733]_ , \new_[84736]_ , \new_[84739]_ , \new_[84740]_ ,
    \new_[84743]_ , \new_[84746]_ , \new_[84747]_ , \new_[84748]_ ,
    \new_[84752]_ , \new_[84753]_ , \new_[84756]_ , \new_[84759]_ ,
    \new_[84760]_ , \new_[84761]_ , \new_[84764]_ , \new_[84767]_ ,
    \new_[84768]_ , \new_[84771]_ , \new_[84774]_ , \new_[84775]_ ,
    \new_[84776]_ , \new_[84780]_ , \new_[84781]_ , \new_[84784]_ ,
    \new_[84787]_ , \new_[84788]_ , \new_[84789]_ , \new_[84792]_ ,
    \new_[84795]_ , \new_[84796]_ , \new_[84799]_ , \new_[84802]_ ,
    \new_[84803]_ , \new_[84804]_ , \new_[84808]_ , \new_[84809]_ ,
    \new_[84812]_ , \new_[84815]_ , \new_[84816]_ , \new_[84817]_ ,
    \new_[84820]_ , \new_[84823]_ , \new_[84824]_ , \new_[84827]_ ,
    \new_[84830]_ , \new_[84831]_ , \new_[84832]_ , \new_[84836]_ ,
    \new_[84837]_ , \new_[84840]_ , \new_[84843]_ , \new_[84844]_ ,
    \new_[84845]_ , \new_[84848]_ , \new_[84851]_ , \new_[84852]_ ,
    \new_[84855]_ , \new_[84858]_ , \new_[84859]_ , \new_[84860]_ ,
    \new_[84864]_ , \new_[84865]_ , \new_[84868]_ , \new_[84871]_ ,
    \new_[84872]_ , \new_[84873]_ , \new_[84876]_ , \new_[84879]_ ,
    \new_[84880]_ , \new_[84883]_ , \new_[84886]_ , \new_[84887]_ ,
    \new_[84888]_ , \new_[84892]_ , \new_[84893]_ , \new_[84896]_ ,
    \new_[84899]_ , \new_[84900]_ , \new_[84901]_ , \new_[84904]_ ,
    \new_[84907]_ , \new_[84908]_ , \new_[84911]_ , \new_[84914]_ ,
    \new_[84915]_ , \new_[84916]_ , \new_[84920]_ , \new_[84921]_ ,
    \new_[84924]_ , \new_[84927]_ , \new_[84928]_ , \new_[84929]_ ,
    \new_[84932]_ , \new_[84935]_ , \new_[84936]_ , \new_[84939]_ ,
    \new_[84942]_ , \new_[84943]_ , \new_[84944]_ , \new_[84948]_ ,
    \new_[84949]_ , \new_[84952]_ , \new_[84955]_ , \new_[84956]_ ,
    \new_[84957]_ , \new_[84960]_ , \new_[84963]_ , \new_[84964]_ ,
    \new_[84967]_ , \new_[84970]_ , \new_[84971]_ , \new_[84972]_ ,
    \new_[84976]_ , \new_[84977]_ , \new_[84980]_ , \new_[84983]_ ,
    \new_[84984]_ , \new_[84985]_ , \new_[84988]_ , \new_[84991]_ ,
    \new_[84992]_ , \new_[84995]_ , \new_[84998]_ , \new_[84999]_ ,
    \new_[85000]_ , \new_[85004]_ , \new_[85005]_ , \new_[85008]_ ,
    \new_[85011]_ , \new_[85012]_ , \new_[85013]_ , \new_[85016]_ ,
    \new_[85019]_ , \new_[85020]_ , \new_[85023]_ , \new_[85026]_ ,
    \new_[85027]_ , \new_[85028]_ , \new_[85032]_ , \new_[85033]_ ,
    \new_[85036]_ , \new_[85039]_ , \new_[85040]_ , \new_[85041]_ ,
    \new_[85044]_ , \new_[85047]_ , \new_[85048]_ , \new_[85051]_ ,
    \new_[85054]_ , \new_[85055]_ , \new_[85056]_ , \new_[85060]_ ,
    \new_[85061]_ , \new_[85064]_ , \new_[85067]_ , \new_[85068]_ ,
    \new_[85069]_ , \new_[85072]_ , \new_[85075]_ , \new_[85076]_ ,
    \new_[85079]_ , \new_[85082]_ , \new_[85083]_ , \new_[85084]_ ,
    \new_[85088]_ , \new_[85089]_ , \new_[85092]_ , \new_[85095]_ ,
    \new_[85096]_ , \new_[85097]_ , \new_[85100]_ , \new_[85103]_ ,
    \new_[85104]_ , \new_[85107]_ , \new_[85110]_ , \new_[85111]_ ,
    \new_[85112]_ , \new_[85116]_ , \new_[85117]_ , \new_[85120]_ ,
    \new_[85123]_ , \new_[85124]_ , \new_[85125]_ , \new_[85128]_ ,
    \new_[85131]_ , \new_[85132]_ , \new_[85135]_ , \new_[85138]_ ,
    \new_[85139]_ , \new_[85140]_ , \new_[85144]_ , \new_[85145]_ ,
    \new_[85148]_ , \new_[85151]_ , \new_[85152]_ , \new_[85153]_ ,
    \new_[85156]_ , \new_[85159]_ , \new_[85160]_ , \new_[85163]_ ,
    \new_[85166]_ , \new_[85167]_ , \new_[85168]_ , \new_[85172]_ ,
    \new_[85173]_ , \new_[85176]_ , \new_[85179]_ , \new_[85180]_ ,
    \new_[85181]_ , \new_[85184]_ , \new_[85187]_ , \new_[85188]_ ,
    \new_[85191]_ , \new_[85194]_ , \new_[85195]_ , \new_[85196]_ ,
    \new_[85200]_ , \new_[85201]_ , \new_[85204]_ , \new_[85207]_ ,
    \new_[85208]_ , \new_[85209]_ , \new_[85212]_ , \new_[85215]_ ,
    \new_[85216]_ , \new_[85219]_ , \new_[85222]_ , \new_[85223]_ ,
    \new_[85224]_ , \new_[85228]_ , \new_[85229]_ , \new_[85232]_ ,
    \new_[85235]_ , \new_[85236]_ , \new_[85237]_ , \new_[85240]_ ,
    \new_[85243]_ , \new_[85244]_ , \new_[85247]_ , \new_[85250]_ ,
    \new_[85251]_ , \new_[85252]_ , \new_[85256]_ , \new_[85257]_ ,
    \new_[85260]_ , \new_[85263]_ , \new_[85264]_ , \new_[85265]_ ,
    \new_[85268]_ , \new_[85271]_ , \new_[85272]_ , \new_[85275]_ ,
    \new_[85278]_ , \new_[85279]_ , \new_[85280]_ , \new_[85284]_ ,
    \new_[85285]_ , \new_[85288]_ , \new_[85291]_ , \new_[85292]_ ,
    \new_[85293]_ , \new_[85296]_ , \new_[85299]_ , \new_[85300]_ ,
    \new_[85303]_ , \new_[85306]_ , \new_[85307]_ , \new_[85308]_ ,
    \new_[85312]_ , \new_[85313]_ , \new_[85316]_ , \new_[85319]_ ,
    \new_[85320]_ , \new_[85321]_ , \new_[85324]_ , \new_[85327]_ ,
    \new_[85328]_ , \new_[85331]_ , \new_[85334]_ , \new_[85335]_ ,
    \new_[85336]_ , \new_[85340]_ , \new_[85341]_ , \new_[85344]_ ,
    \new_[85347]_ , \new_[85348]_ , \new_[85349]_ , \new_[85352]_ ,
    \new_[85355]_ , \new_[85356]_ , \new_[85359]_ , \new_[85362]_ ,
    \new_[85363]_ , \new_[85364]_ , \new_[85368]_ , \new_[85369]_ ,
    \new_[85372]_ , \new_[85375]_ , \new_[85376]_ , \new_[85377]_ ,
    \new_[85380]_ , \new_[85383]_ , \new_[85384]_ , \new_[85387]_ ,
    \new_[85390]_ , \new_[85391]_ , \new_[85392]_ , \new_[85396]_ ,
    \new_[85397]_ , \new_[85400]_ , \new_[85403]_ , \new_[85404]_ ,
    \new_[85405]_ , \new_[85408]_ , \new_[85411]_ , \new_[85412]_ ,
    \new_[85415]_ , \new_[85418]_ , \new_[85419]_ , \new_[85420]_ ,
    \new_[85424]_ , \new_[85425]_ , \new_[85428]_ , \new_[85431]_ ,
    \new_[85432]_ , \new_[85433]_ , \new_[85436]_ , \new_[85439]_ ,
    \new_[85440]_ , \new_[85443]_ , \new_[85446]_ , \new_[85447]_ ,
    \new_[85448]_ , \new_[85452]_ , \new_[85453]_ , \new_[85456]_ ,
    \new_[85459]_ , \new_[85460]_ , \new_[85461]_ , \new_[85464]_ ,
    \new_[85467]_ , \new_[85468]_ , \new_[85471]_ , \new_[85474]_ ,
    \new_[85475]_ , \new_[85476]_ , \new_[85480]_ , \new_[85481]_ ,
    \new_[85484]_ , \new_[85487]_ , \new_[85488]_ , \new_[85489]_ ,
    \new_[85492]_ , \new_[85495]_ , \new_[85496]_ , \new_[85499]_ ,
    \new_[85502]_ , \new_[85503]_ , \new_[85504]_ , \new_[85508]_ ,
    \new_[85509]_ , \new_[85512]_ , \new_[85515]_ , \new_[85516]_ ,
    \new_[85517]_ , \new_[85520]_ , \new_[85523]_ , \new_[85524]_ ,
    \new_[85527]_ , \new_[85530]_ , \new_[85531]_ , \new_[85532]_ ,
    \new_[85536]_ , \new_[85537]_ , \new_[85540]_ , \new_[85543]_ ,
    \new_[85544]_ , \new_[85545]_ , \new_[85548]_ , \new_[85551]_ ,
    \new_[85552]_ , \new_[85555]_ , \new_[85558]_ , \new_[85559]_ ,
    \new_[85560]_ , \new_[85564]_ , \new_[85565]_ , \new_[85568]_ ,
    \new_[85571]_ , \new_[85572]_ , \new_[85573]_ , \new_[85576]_ ,
    \new_[85579]_ , \new_[85580]_ , \new_[85583]_ , \new_[85586]_ ,
    \new_[85587]_ , \new_[85588]_ , \new_[85592]_ , \new_[85593]_ ,
    \new_[85596]_ , \new_[85599]_ , \new_[85600]_ , \new_[85601]_ ,
    \new_[85604]_ , \new_[85607]_ , \new_[85608]_ , \new_[85611]_ ,
    \new_[85614]_ , \new_[85615]_ , \new_[85616]_ , \new_[85620]_ ,
    \new_[85621]_ , \new_[85624]_ , \new_[85627]_ , \new_[85628]_ ,
    \new_[85629]_ , \new_[85632]_ , \new_[85635]_ , \new_[85636]_ ,
    \new_[85639]_ , \new_[85642]_ , \new_[85643]_ , \new_[85644]_ ,
    \new_[85648]_ , \new_[85649]_ , \new_[85652]_ , \new_[85655]_ ,
    \new_[85656]_ , \new_[85657]_ , \new_[85660]_ , \new_[85663]_ ,
    \new_[85664]_ , \new_[85667]_ , \new_[85670]_ , \new_[85671]_ ,
    \new_[85672]_ , \new_[85676]_ , \new_[85677]_ , \new_[85680]_ ,
    \new_[85683]_ , \new_[85684]_ , \new_[85685]_ , \new_[85688]_ ,
    \new_[85691]_ , \new_[85692]_ , \new_[85695]_ , \new_[85698]_ ,
    \new_[85699]_ , \new_[85700]_ , \new_[85704]_ , \new_[85705]_ ,
    \new_[85708]_ , \new_[85711]_ , \new_[85712]_ , \new_[85713]_ ,
    \new_[85716]_ , \new_[85719]_ , \new_[85720]_ , \new_[85723]_ ,
    \new_[85726]_ , \new_[85727]_ , \new_[85728]_ , \new_[85732]_ ,
    \new_[85733]_ , \new_[85736]_ , \new_[85739]_ , \new_[85740]_ ,
    \new_[85741]_ , \new_[85744]_ , \new_[85747]_ , \new_[85748]_ ,
    \new_[85751]_ , \new_[85754]_ , \new_[85755]_ , \new_[85756]_ ,
    \new_[85760]_ , \new_[85761]_ , \new_[85764]_ , \new_[85767]_ ,
    \new_[85768]_ , \new_[85769]_ , \new_[85772]_ , \new_[85775]_ ,
    \new_[85776]_ , \new_[85779]_ , \new_[85782]_ , \new_[85783]_ ,
    \new_[85784]_ , \new_[85788]_ , \new_[85789]_ , \new_[85792]_ ,
    \new_[85795]_ , \new_[85796]_ , \new_[85797]_ , \new_[85800]_ ,
    \new_[85803]_ , \new_[85804]_ , \new_[85807]_ , \new_[85810]_ ,
    \new_[85811]_ , \new_[85812]_ , \new_[85816]_ , \new_[85817]_ ,
    \new_[85820]_ , \new_[85823]_ , \new_[85824]_ , \new_[85825]_ ,
    \new_[85828]_ , \new_[85831]_ , \new_[85832]_ , \new_[85835]_ ,
    \new_[85838]_ , \new_[85839]_ , \new_[85840]_ , \new_[85844]_ ,
    \new_[85845]_ , \new_[85848]_ , \new_[85851]_ , \new_[85852]_ ,
    \new_[85853]_ , \new_[85856]_ , \new_[85859]_ , \new_[85860]_ ,
    \new_[85863]_ , \new_[85866]_ , \new_[85867]_ , \new_[85868]_ ,
    \new_[85872]_ , \new_[85873]_ , \new_[85876]_ , \new_[85879]_ ,
    \new_[85880]_ , \new_[85881]_ , \new_[85884]_ , \new_[85887]_ ,
    \new_[85888]_ , \new_[85891]_ , \new_[85894]_ , \new_[85895]_ ,
    \new_[85896]_ , \new_[85900]_ , \new_[85901]_ , \new_[85904]_ ,
    \new_[85907]_ , \new_[85908]_ , \new_[85909]_ , \new_[85912]_ ,
    \new_[85915]_ , \new_[85916]_ , \new_[85919]_ , \new_[85922]_ ,
    \new_[85923]_ , \new_[85924]_ , \new_[85928]_ , \new_[85929]_ ,
    \new_[85932]_ , \new_[85935]_ , \new_[85936]_ , \new_[85937]_ ,
    \new_[85940]_ , \new_[85943]_ , \new_[85944]_ , \new_[85947]_ ,
    \new_[85950]_ , \new_[85951]_ , \new_[85952]_ , \new_[85956]_ ,
    \new_[85957]_ , \new_[85960]_ , \new_[85963]_ , \new_[85964]_ ,
    \new_[85965]_ , \new_[85968]_ , \new_[85971]_ , \new_[85972]_ ,
    \new_[85975]_ , \new_[85978]_ , \new_[85979]_ , \new_[85980]_ ,
    \new_[85984]_ , \new_[85985]_ , \new_[85988]_ , \new_[85991]_ ,
    \new_[85992]_ , \new_[85993]_ , \new_[85996]_ , \new_[85999]_ ,
    \new_[86000]_ , \new_[86003]_ , \new_[86006]_ , \new_[86007]_ ,
    \new_[86008]_ , \new_[86012]_ , \new_[86013]_ , \new_[86016]_ ,
    \new_[86019]_ , \new_[86020]_ , \new_[86021]_ , \new_[86024]_ ,
    \new_[86027]_ , \new_[86028]_ , \new_[86031]_ , \new_[86034]_ ,
    \new_[86035]_ , \new_[86036]_ , \new_[86040]_ , \new_[86041]_ ,
    \new_[86044]_ , \new_[86047]_ , \new_[86048]_ , \new_[86049]_ ,
    \new_[86052]_ , \new_[86055]_ , \new_[86056]_ , \new_[86059]_ ,
    \new_[86062]_ , \new_[86063]_ , \new_[86064]_ , \new_[86068]_ ,
    \new_[86069]_ , \new_[86072]_ , \new_[86075]_ , \new_[86076]_ ,
    \new_[86077]_ , \new_[86080]_ , \new_[86083]_ , \new_[86084]_ ,
    \new_[86087]_ , \new_[86090]_ , \new_[86091]_ , \new_[86092]_ ,
    \new_[86096]_ , \new_[86097]_ , \new_[86100]_ , \new_[86103]_ ,
    \new_[86104]_ , \new_[86105]_ , \new_[86108]_ , \new_[86111]_ ,
    \new_[86112]_ , \new_[86115]_ , \new_[86118]_ , \new_[86119]_ ,
    \new_[86120]_ , \new_[86124]_ , \new_[86125]_ , \new_[86128]_ ,
    \new_[86131]_ , \new_[86132]_ , \new_[86133]_ , \new_[86136]_ ,
    \new_[86139]_ , \new_[86140]_ , \new_[86143]_ , \new_[86146]_ ,
    \new_[86147]_ , \new_[86148]_ , \new_[86152]_ , \new_[86153]_ ,
    \new_[86156]_ , \new_[86159]_ , \new_[86160]_ , \new_[86161]_ ,
    \new_[86164]_ , \new_[86167]_ , \new_[86168]_ , \new_[86171]_ ,
    \new_[86174]_ , \new_[86175]_ , \new_[86176]_ , \new_[86180]_ ,
    \new_[86181]_ , \new_[86184]_ , \new_[86187]_ , \new_[86188]_ ,
    \new_[86189]_ , \new_[86192]_ , \new_[86195]_ , \new_[86196]_ ,
    \new_[86199]_ , \new_[86202]_ , \new_[86203]_ , \new_[86204]_ ,
    \new_[86208]_ , \new_[86209]_ , \new_[86212]_ , \new_[86215]_ ,
    \new_[86216]_ , \new_[86217]_ , \new_[86220]_ , \new_[86223]_ ,
    \new_[86224]_ , \new_[86227]_ , \new_[86230]_ , \new_[86231]_ ,
    \new_[86232]_ , \new_[86236]_ , \new_[86237]_ , \new_[86240]_ ,
    \new_[86243]_ , \new_[86244]_ , \new_[86245]_ , \new_[86248]_ ,
    \new_[86251]_ , \new_[86252]_ , \new_[86255]_ , \new_[86258]_ ,
    \new_[86259]_ , \new_[86260]_ , \new_[86264]_ , \new_[86265]_ ,
    \new_[86268]_ , \new_[86271]_ , \new_[86272]_ , \new_[86273]_ ,
    \new_[86276]_ , \new_[86279]_ , \new_[86280]_ , \new_[86283]_ ,
    \new_[86286]_ , \new_[86287]_ , \new_[86288]_ , \new_[86292]_ ,
    \new_[86293]_ , \new_[86296]_ , \new_[86299]_ , \new_[86300]_ ,
    \new_[86301]_ , \new_[86304]_ , \new_[86307]_ , \new_[86308]_ ,
    \new_[86311]_ , \new_[86314]_ , \new_[86315]_ , \new_[86316]_ ,
    \new_[86320]_ , \new_[86321]_ , \new_[86324]_ , \new_[86327]_ ,
    \new_[86328]_ , \new_[86329]_ , \new_[86332]_ , \new_[86335]_ ,
    \new_[86336]_ , \new_[86339]_ , \new_[86342]_ , \new_[86343]_ ,
    \new_[86344]_ , \new_[86348]_ , \new_[86349]_ , \new_[86352]_ ,
    \new_[86355]_ , \new_[86356]_ , \new_[86357]_ , \new_[86360]_ ,
    \new_[86363]_ , \new_[86364]_ , \new_[86367]_ , \new_[86370]_ ,
    \new_[86371]_ , \new_[86372]_ , \new_[86376]_ , \new_[86377]_ ,
    \new_[86380]_ , \new_[86383]_ , \new_[86384]_ , \new_[86385]_ ,
    \new_[86388]_ , \new_[86391]_ , \new_[86392]_ , \new_[86395]_ ,
    \new_[86398]_ , \new_[86399]_ , \new_[86400]_ , \new_[86404]_ ,
    \new_[86405]_ , \new_[86408]_ , \new_[86411]_ , \new_[86412]_ ,
    \new_[86413]_ , \new_[86416]_ , \new_[86419]_ , \new_[86420]_ ,
    \new_[86423]_ , \new_[86426]_ , \new_[86427]_ , \new_[86428]_ ,
    \new_[86432]_ , \new_[86433]_ , \new_[86436]_ , \new_[86439]_ ,
    \new_[86440]_ , \new_[86441]_ , \new_[86444]_ , \new_[86447]_ ,
    \new_[86448]_ , \new_[86451]_ , \new_[86454]_ , \new_[86455]_ ,
    \new_[86456]_ , \new_[86460]_ , \new_[86461]_ , \new_[86464]_ ,
    \new_[86467]_ , \new_[86468]_ , \new_[86469]_ , \new_[86472]_ ,
    \new_[86475]_ , \new_[86476]_ , \new_[86479]_ , \new_[86482]_ ,
    \new_[86483]_ , \new_[86484]_ , \new_[86488]_ , \new_[86489]_ ,
    \new_[86492]_ , \new_[86495]_ , \new_[86496]_ , \new_[86497]_ ,
    \new_[86500]_ , \new_[86503]_ , \new_[86504]_ , \new_[86507]_ ,
    \new_[86510]_ , \new_[86511]_ , \new_[86512]_ , \new_[86516]_ ,
    \new_[86517]_ , \new_[86520]_ , \new_[86523]_ , \new_[86524]_ ,
    \new_[86525]_ , \new_[86528]_ , \new_[86531]_ , \new_[86532]_ ,
    \new_[86535]_ , \new_[86538]_ , \new_[86539]_ , \new_[86540]_ ,
    \new_[86544]_ , \new_[86545]_ , \new_[86548]_ , \new_[86551]_ ,
    \new_[86552]_ , \new_[86553]_ , \new_[86556]_ , \new_[86559]_ ,
    \new_[86560]_ , \new_[86563]_ , \new_[86566]_ , \new_[86567]_ ,
    \new_[86568]_ , \new_[86572]_ , \new_[86573]_ , \new_[86576]_ ,
    \new_[86579]_ , \new_[86580]_ , \new_[86581]_ , \new_[86584]_ ,
    \new_[86587]_ , \new_[86588]_ , \new_[86591]_ , \new_[86594]_ ,
    \new_[86595]_ , \new_[86596]_ , \new_[86600]_ , \new_[86601]_ ,
    \new_[86604]_ , \new_[86607]_ , \new_[86608]_ , \new_[86609]_ ,
    \new_[86612]_ , \new_[86615]_ , \new_[86616]_ , \new_[86619]_ ,
    \new_[86622]_ , \new_[86623]_ , \new_[86624]_ , \new_[86628]_ ,
    \new_[86629]_ , \new_[86632]_ , \new_[86635]_ , \new_[86636]_ ,
    \new_[86637]_ , \new_[86640]_ , \new_[86643]_ , \new_[86644]_ ,
    \new_[86647]_ , \new_[86650]_ , \new_[86651]_ , \new_[86652]_ ,
    \new_[86656]_ , \new_[86657]_ , \new_[86660]_ , \new_[86663]_ ,
    \new_[86664]_ , \new_[86665]_ , \new_[86668]_ , \new_[86671]_ ,
    \new_[86672]_ , \new_[86675]_ , \new_[86678]_ , \new_[86679]_ ,
    \new_[86680]_ , \new_[86684]_ , \new_[86685]_ , \new_[86688]_ ,
    \new_[86691]_ , \new_[86692]_ , \new_[86693]_ , \new_[86696]_ ,
    \new_[86699]_ , \new_[86700]_ , \new_[86703]_ , \new_[86706]_ ,
    \new_[86707]_ , \new_[86708]_ , \new_[86712]_ , \new_[86713]_ ,
    \new_[86716]_ , \new_[86719]_ , \new_[86720]_ , \new_[86721]_ ,
    \new_[86724]_ , \new_[86727]_ , \new_[86728]_ , \new_[86731]_ ,
    \new_[86734]_ , \new_[86735]_ , \new_[86736]_ , \new_[86740]_ ,
    \new_[86741]_ , \new_[86744]_ , \new_[86747]_ , \new_[86748]_ ,
    \new_[86749]_ , \new_[86752]_ , \new_[86755]_ , \new_[86756]_ ,
    \new_[86759]_ , \new_[86762]_ , \new_[86763]_ , \new_[86764]_ ,
    \new_[86768]_ , \new_[86769]_ , \new_[86772]_ , \new_[86775]_ ,
    \new_[86776]_ , \new_[86777]_ , \new_[86780]_ , \new_[86783]_ ,
    \new_[86784]_ , \new_[86787]_ , \new_[86790]_ , \new_[86791]_ ,
    \new_[86792]_ , \new_[86796]_ , \new_[86797]_ , \new_[86800]_ ,
    \new_[86803]_ , \new_[86804]_ , \new_[86805]_ , \new_[86808]_ ,
    \new_[86811]_ , \new_[86812]_ , \new_[86815]_ , \new_[86818]_ ,
    \new_[86819]_ , \new_[86820]_ , \new_[86824]_ , \new_[86825]_ ,
    \new_[86828]_ , \new_[86831]_ , \new_[86832]_ , \new_[86833]_ ,
    \new_[86836]_ , \new_[86839]_ , \new_[86840]_ , \new_[86843]_ ,
    \new_[86846]_ , \new_[86847]_ , \new_[86848]_ , \new_[86852]_ ,
    \new_[86853]_ , \new_[86856]_ , \new_[86859]_ , \new_[86860]_ ,
    \new_[86861]_ , \new_[86864]_ , \new_[86867]_ , \new_[86868]_ ,
    \new_[86871]_ , \new_[86874]_ , \new_[86875]_ , \new_[86876]_ ,
    \new_[86880]_ , \new_[86881]_ , \new_[86884]_ , \new_[86887]_ ,
    \new_[86888]_ , \new_[86889]_ , \new_[86892]_ , \new_[86895]_ ,
    \new_[86896]_ , \new_[86899]_ , \new_[86902]_ , \new_[86903]_ ,
    \new_[86904]_ , \new_[86908]_ , \new_[86909]_ , \new_[86912]_ ,
    \new_[86915]_ , \new_[86916]_ , \new_[86917]_ , \new_[86920]_ ,
    \new_[86923]_ , \new_[86924]_ , \new_[86927]_ , \new_[86930]_ ,
    \new_[86931]_ , \new_[86932]_ , \new_[86936]_ , \new_[86937]_ ,
    \new_[86940]_ , \new_[86943]_ , \new_[86944]_ , \new_[86945]_ ,
    \new_[86948]_ , \new_[86951]_ , \new_[86952]_ , \new_[86955]_ ,
    \new_[86958]_ , \new_[86959]_ , \new_[86960]_ , \new_[86964]_ ,
    \new_[86965]_ , \new_[86968]_ , \new_[86971]_ , \new_[86972]_ ,
    \new_[86973]_ , \new_[86976]_ , \new_[86979]_ , \new_[86980]_ ,
    \new_[86983]_ , \new_[86986]_ , \new_[86987]_ , \new_[86988]_ ,
    \new_[86992]_ , \new_[86993]_ , \new_[86996]_ , \new_[86999]_ ,
    \new_[87000]_ , \new_[87001]_ , \new_[87004]_ , \new_[87007]_ ,
    \new_[87008]_ , \new_[87011]_ , \new_[87014]_ , \new_[87015]_ ,
    \new_[87016]_ , \new_[87020]_ , \new_[87021]_ , \new_[87024]_ ,
    \new_[87027]_ , \new_[87028]_ , \new_[87029]_ , \new_[87032]_ ,
    \new_[87035]_ , \new_[87036]_ , \new_[87039]_ , \new_[87042]_ ,
    \new_[87043]_ , \new_[87044]_ , \new_[87048]_ , \new_[87049]_ ,
    \new_[87052]_ , \new_[87055]_ , \new_[87056]_ , \new_[87057]_ ,
    \new_[87060]_ , \new_[87063]_ , \new_[87064]_ , \new_[87067]_ ,
    \new_[87070]_ , \new_[87071]_ , \new_[87072]_ , \new_[87076]_ ,
    \new_[87077]_ , \new_[87080]_ , \new_[87083]_ , \new_[87084]_ ,
    \new_[87085]_ , \new_[87088]_ , \new_[87091]_ , \new_[87092]_ ,
    \new_[87095]_ , \new_[87098]_ , \new_[87099]_ , \new_[87100]_ ,
    \new_[87104]_ , \new_[87105]_ , \new_[87108]_ , \new_[87111]_ ,
    \new_[87112]_ , \new_[87113]_ , \new_[87116]_ , \new_[87119]_ ,
    \new_[87120]_ , \new_[87123]_ , \new_[87126]_ , \new_[87127]_ ,
    \new_[87128]_ , \new_[87132]_ , \new_[87133]_ , \new_[87136]_ ,
    \new_[87139]_ , \new_[87140]_ , \new_[87141]_ , \new_[87144]_ ,
    \new_[87147]_ , \new_[87148]_ , \new_[87151]_ , \new_[87154]_ ,
    \new_[87155]_ , \new_[87156]_ , \new_[87160]_ , \new_[87161]_ ,
    \new_[87164]_ , \new_[87167]_ , \new_[87168]_ , \new_[87169]_ ,
    \new_[87172]_ , \new_[87175]_ , \new_[87176]_ , \new_[87179]_ ,
    \new_[87182]_ , \new_[87183]_ , \new_[87184]_ , \new_[87188]_ ,
    \new_[87189]_ , \new_[87192]_ , \new_[87195]_ , \new_[87196]_ ,
    \new_[87197]_ , \new_[87200]_ , \new_[87203]_ , \new_[87204]_ ,
    \new_[87207]_ , \new_[87210]_ , \new_[87211]_ , \new_[87212]_ ,
    \new_[87216]_ , \new_[87217]_ , \new_[87220]_ , \new_[87223]_ ,
    \new_[87224]_ , \new_[87225]_ , \new_[87228]_ , \new_[87231]_ ,
    \new_[87232]_ , \new_[87235]_ , \new_[87238]_ , \new_[87239]_ ,
    \new_[87240]_ , \new_[87244]_ , \new_[87245]_ , \new_[87248]_ ,
    \new_[87251]_ , \new_[87252]_ , \new_[87253]_ , \new_[87256]_ ,
    \new_[87259]_ , \new_[87260]_ , \new_[87263]_ , \new_[87266]_ ,
    \new_[87267]_ , \new_[87268]_ , \new_[87272]_ , \new_[87273]_ ,
    \new_[87276]_ , \new_[87279]_ , \new_[87280]_ , \new_[87281]_ ,
    \new_[87284]_ , \new_[87287]_ , \new_[87288]_ , \new_[87291]_ ,
    \new_[87294]_ , \new_[87295]_ , \new_[87296]_ , \new_[87300]_ ,
    \new_[87301]_ , \new_[87304]_ , \new_[87307]_ , \new_[87308]_ ,
    \new_[87309]_ , \new_[87312]_ , \new_[87315]_ , \new_[87316]_ ,
    \new_[87319]_ , \new_[87322]_ , \new_[87323]_ , \new_[87324]_ ,
    \new_[87328]_ , \new_[87329]_ , \new_[87332]_ , \new_[87335]_ ,
    \new_[87336]_ , \new_[87337]_ , \new_[87340]_ , \new_[87343]_ ,
    \new_[87344]_ , \new_[87347]_ , \new_[87350]_ , \new_[87351]_ ,
    \new_[87352]_ , \new_[87356]_ , \new_[87357]_ , \new_[87360]_ ,
    \new_[87363]_ , \new_[87364]_ , \new_[87365]_ , \new_[87368]_ ,
    \new_[87371]_ , \new_[87372]_ , \new_[87375]_ , \new_[87378]_ ,
    \new_[87379]_ , \new_[87380]_ , \new_[87384]_ , \new_[87385]_ ,
    \new_[87388]_ , \new_[87391]_ , \new_[87392]_ , \new_[87393]_ ,
    \new_[87396]_ , \new_[87399]_ , \new_[87400]_ , \new_[87403]_ ,
    \new_[87406]_ , \new_[87407]_ , \new_[87408]_ , \new_[87412]_ ,
    \new_[87413]_ , \new_[87416]_ , \new_[87419]_ , \new_[87420]_ ,
    \new_[87421]_ , \new_[87424]_ , \new_[87427]_ , \new_[87428]_ ,
    \new_[87431]_ , \new_[87434]_ , \new_[87435]_ , \new_[87436]_ ,
    \new_[87440]_ , \new_[87441]_ , \new_[87444]_ , \new_[87447]_ ,
    \new_[87448]_ , \new_[87449]_ , \new_[87452]_ , \new_[87455]_ ,
    \new_[87456]_ , \new_[87459]_ , \new_[87462]_ , \new_[87463]_ ,
    \new_[87464]_ , \new_[87468]_ , \new_[87469]_ , \new_[87472]_ ,
    \new_[87475]_ , \new_[87476]_ , \new_[87477]_ , \new_[87480]_ ,
    \new_[87483]_ , \new_[87484]_ , \new_[87487]_ , \new_[87490]_ ,
    \new_[87491]_ , \new_[87492]_ , \new_[87496]_ , \new_[87497]_ ,
    \new_[87500]_ , \new_[87503]_ , \new_[87504]_ , \new_[87505]_ ,
    \new_[87508]_ , \new_[87511]_ , \new_[87512]_ , \new_[87515]_ ,
    \new_[87518]_ , \new_[87519]_ , \new_[87520]_ , \new_[87524]_ ,
    \new_[87525]_ , \new_[87528]_ , \new_[87531]_ , \new_[87532]_ ,
    \new_[87533]_ , \new_[87536]_ , \new_[87539]_ , \new_[87540]_ ,
    \new_[87543]_ , \new_[87546]_ , \new_[87547]_ , \new_[87548]_ ,
    \new_[87552]_ , \new_[87553]_ , \new_[87556]_ , \new_[87559]_ ,
    \new_[87560]_ , \new_[87561]_ , \new_[87564]_ , \new_[87567]_ ,
    \new_[87568]_ , \new_[87571]_ , \new_[87574]_ , \new_[87575]_ ,
    \new_[87576]_ , \new_[87580]_ , \new_[87581]_ , \new_[87584]_ ,
    \new_[87587]_ , \new_[87588]_ , \new_[87589]_ , \new_[87592]_ ,
    \new_[87595]_ , \new_[87596]_ , \new_[87599]_ , \new_[87602]_ ,
    \new_[87603]_ , \new_[87604]_ , \new_[87608]_ , \new_[87609]_ ,
    \new_[87612]_ , \new_[87615]_ , \new_[87616]_ , \new_[87617]_ ,
    \new_[87620]_ , \new_[87623]_ , \new_[87624]_ , \new_[87627]_ ,
    \new_[87630]_ , \new_[87631]_ , \new_[87632]_ , \new_[87636]_ ,
    \new_[87637]_ , \new_[87640]_ , \new_[87643]_ , \new_[87644]_ ,
    \new_[87645]_ , \new_[87648]_ , \new_[87651]_ , \new_[87652]_ ,
    \new_[87655]_ , \new_[87658]_ , \new_[87659]_ , \new_[87660]_ ,
    \new_[87664]_ , \new_[87665]_ , \new_[87668]_ , \new_[87671]_ ,
    \new_[87672]_ , \new_[87673]_ , \new_[87676]_ , \new_[87679]_ ,
    \new_[87680]_ , \new_[87683]_ , \new_[87686]_ , \new_[87687]_ ,
    \new_[87688]_ , \new_[87692]_ , \new_[87693]_ , \new_[87696]_ ,
    \new_[87699]_ , \new_[87700]_ , \new_[87701]_ , \new_[87704]_ ,
    \new_[87707]_ , \new_[87708]_ , \new_[87711]_ , \new_[87714]_ ,
    \new_[87715]_ , \new_[87716]_ , \new_[87720]_ , \new_[87721]_ ,
    \new_[87724]_ , \new_[87727]_ , \new_[87728]_ , \new_[87729]_ ,
    \new_[87732]_ , \new_[87735]_ , \new_[87736]_ , \new_[87739]_ ,
    \new_[87742]_ , \new_[87743]_ , \new_[87744]_ , \new_[87748]_ ,
    \new_[87749]_ , \new_[87752]_ , \new_[87755]_ , \new_[87756]_ ,
    \new_[87757]_ , \new_[87760]_ , \new_[87763]_ , \new_[87764]_ ,
    \new_[87767]_ , \new_[87770]_ , \new_[87771]_ , \new_[87772]_ ,
    \new_[87776]_ , \new_[87777]_ , \new_[87780]_ , \new_[87783]_ ,
    \new_[87784]_ , \new_[87785]_ , \new_[87788]_ , \new_[87791]_ ,
    \new_[87792]_ , \new_[87795]_ , \new_[87798]_ , \new_[87799]_ ,
    \new_[87800]_ , \new_[87804]_ , \new_[87805]_ , \new_[87808]_ ,
    \new_[87811]_ , \new_[87812]_ , \new_[87813]_ , \new_[87816]_ ,
    \new_[87819]_ , \new_[87820]_ , \new_[87823]_ , \new_[87826]_ ,
    \new_[87827]_ , \new_[87828]_ , \new_[87832]_ , \new_[87833]_ ,
    \new_[87836]_ , \new_[87839]_ , \new_[87840]_ , \new_[87841]_ ,
    \new_[87844]_ , \new_[87847]_ , \new_[87848]_ , \new_[87851]_ ,
    \new_[87854]_ , \new_[87855]_ , \new_[87856]_ , \new_[87860]_ ,
    \new_[87861]_ , \new_[87864]_ , \new_[87867]_ , \new_[87868]_ ,
    \new_[87869]_ , \new_[87872]_ , \new_[87875]_ , \new_[87876]_ ,
    \new_[87879]_ , \new_[87882]_ , \new_[87883]_ , \new_[87884]_ ,
    \new_[87888]_ , \new_[87889]_ , \new_[87892]_ , \new_[87895]_ ,
    \new_[87896]_ , \new_[87897]_ , \new_[87900]_ , \new_[87903]_ ,
    \new_[87904]_ , \new_[87907]_ , \new_[87910]_ , \new_[87911]_ ,
    \new_[87912]_ , \new_[87916]_ , \new_[87917]_ , \new_[87920]_ ,
    \new_[87923]_ , \new_[87924]_ , \new_[87925]_ , \new_[87928]_ ,
    \new_[87931]_ , \new_[87932]_ , \new_[87935]_ , \new_[87938]_ ,
    \new_[87939]_ , \new_[87940]_ , \new_[87944]_ , \new_[87945]_ ,
    \new_[87948]_ , \new_[87951]_ , \new_[87952]_ , \new_[87953]_ ,
    \new_[87956]_ , \new_[87959]_ , \new_[87960]_ , \new_[87963]_ ,
    \new_[87966]_ , \new_[87967]_ , \new_[87968]_ , \new_[87972]_ ,
    \new_[87973]_ , \new_[87976]_ , \new_[87979]_ , \new_[87980]_ ,
    \new_[87981]_ , \new_[87984]_ , \new_[87987]_ , \new_[87988]_ ,
    \new_[87991]_ , \new_[87994]_ , \new_[87995]_ , \new_[87996]_ ,
    \new_[88000]_ , \new_[88001]_ , \new_[88004]_ , \new_[88007]_ ,
    \new_[88008]_ , \new_[88009]_ , \new_[88012]_ , \new_[88015]_ ,
    \new_[88016]_ , \new_[88019]_ , \new_[88022]_ , \new_[88023]_ ,
    \new_[88024]_ , \new_[88028]_ , \new_[88029]_ , \new_[88032]_ ,
    \new_[88035]_ , \new_[88036]_ , \new_[88037]_ , \new_[88040]_ ,
    \new_[88043]_ , \new_[88044]_ , \new_[88047]_ , \new_[88050]_ ,
    \new_[88051]_ , \new_[88052]_ , \new_[88056]_ , \new_[88057]_ ,
    \new_[88060]_ , \new_[88063]_ , \new_[88064]_ , \new_[88065]_ ,
    \new_[88068]_ , \new_[88071]_ , \new_[88072]_ , \new_[88075]_ ,
    \new_[88078]_ , \new_[88079]_ , \new_[88080]_ , \new_[88084]_ ,
    \new_[88085]_ , \new_[88088]_ , \new_[88091]_ , \new_[88092]_ ,
    \new_[88093]_ , \new_[88096]_ , \new_[88099]_ , \new_[88100]_ ,
    \new_[88103]_ , \new_[88106]_ , \new_[88107]_ , \new_[88108]_ ,
    \new_[88112]_ , \new_[88113]_ , \new_[88116]_ , \new_[88119]_ ,
    \new_[88120]_ , \new_[88121]_ , \new_[88124]_ , \new_[88127]_ ,
    \new_[88128]_ , \new_[88131]_ , \new_[88134]_ , \new_[88135]_ ,
    \new_[88136]_ , \new_[88140]_ , \new_[88141]_ , \new_[88144]_ ,
    \new_[88147]_ , \new_[88148]_ , \new_[88149]_ , \new_[88152]_ ,
    \new_[88155]_ , \new_[88156]_ , \new_[88159]_ , \new_[88162]_ ,
    \new_[88163]_ , \new_[88164]_ , \new_[88168]_ , \new_[88169]_ ,
    \new_[88172]_ , \new_[88175]_ , \new_[88176]_ , \new_[88177]_ ,
    \new_[88180]_ , \new_[88183]_ , \new_[88184]_ , \new_[88187]_ ,
    \new_[88190]_ , \new_[88191]_ , \new_[88192]_ , \new_[88196]_ ,
    \new_[88197]_ , \new_[88200]_ , \new_[88203]_ , \new_[88204]_ ,
    \new_[88205]_ , \new_[88208]_ , \new_[88211]_ , \new_[88212]_ ,
    \new_[88215]_ , \new_[88218]_ , \new_[88219]_ , \new_[88220]_ ,
    \new_[88224]_ , \new_[88225]_ , \new_[88228]_ , \new_[88231]_ ,
    \new_[88232]_ , \new_[88233]_ , \new_[88236]_ , \new_[88239]_ ,
    \new_[88240]_ , \new_[88243]_ , \new_[88246]_ , \new_[88247]_ ,
    \new_[88248]_ , \new_[88252]_ , \new_[88253]_ , \new_[88256]_ ,
    \new_[88259]_ , \new_[88260]_ , \new_[88261]_ , \new_[88264]_ ,
    \new_[88267]_ , \new_[88268]_ , \new_[88271]_ , \new_[88274]_ ,
    \new_[88275]_ , \new_[88276]_ , \new_[88280]_ , \new_[88281]_ ,
    \new_[88284]_ , \new_[88287]_ , \new_[88288]_ , \new_[88289]_ ,
    \new_[88292]_ , \new_[88295]_ , \new_[88296]_ , \new_[88299]_ ,
    \new_[88302]_ , \new_[88303]_ , \new_[88304]_ , \new_[88308]_ ,
    \new_[88309]_ , \new_[88312]_ , \new_[88315]_ , \new_[88316]_ ,
    \new_[88317]_ , \new_[88320]_ , \new_[88323]_ , \new_[88324]_ ,
    \new_[88327]_ , \new_[88330]_ , \new_[88331]_ , \new_[88332]_ ,
    \new_[88336]_ , \new_[88337]_ , \new_[88340]_ , \new_[88343]_ ,
    \new_[88344]_ , \new_[88345]_ , \new_[88348]_ , \new_[88351]_ ,
    \new_[88352]_ , \new_[88355]_ , \new_[88358]_ , \new_[88359]_ ,
    \new_[88360]_ , \new_[88364]_ , \new_[88365]_ , \new_[88368]_ ,
    \new_[88371]_ , \new_[88372]_ , \new_[88373]_ , \new_[88376]_ ,
    \new_[88379]_ , \new_[88380]_ , \new_[88383]_ , \new_[88386]_ ,
    \new_[88387]_ , \new_[88388]_ , \new_[88392]_ , \new_[88393]_ ,
    \new_[88396]_ , \new_[88399]_ , \new_[88400]_ , \new_[88401]_ ,
    \new_[88404]_ , \new_[88407]_ , \new_[88408]_ , \new_[88411]_ ,
    \new_[88414]_ , \new_[88415]_ , \new_[88416]_ , \new_[88420]_ ,
    \new_[88421]_ , \new_[88424]_ , \new_[88427]_ , \new_[88428]_ ,
    \new_[88429]_ , \new_[88432]_ , \new_[88435]_ , \new_[88436]_ ,
    \new_[88439]_ , \new_[88442]_ , \new_[88443]_ , \new_[88444]_ ,
    \new_[88448]_ , \new_[88449]_ , \new_[88452]_ , \new_[88455]_ ,
    \new_[88456]_ , \new_[88457]_ , \new_[88460]_ , \new_[88463]_ ,
    \new_[88464]_ , \new_[88467]_ , \new_[88470]_ , \new_[88471]_ ,
    \new_[88472]_ , \new_[88476]_ , \new_[88477]_ , \new_[88480]_ ,
    \new_[88483]_ , \new_[88484]_ , \new_[88485]_ , \new_[88488]_ ,
    \new_[88491]_ , \new_[88492]_ , \new_[88495]_ , \new_[88498]_ ,
    \new_[88499]_ , \new_[88500]_ , \new_[88504]_ , \new_[88505]_ ,
    \new_[88508]_ , \new_[88511]_ , \new_[88512]_ , \new_[88513]_ ,
    \new_[88516]_ , \new_[88519]_ , \new_[88520]_ , \new_[88523]_ ,
    \new_[88526]_ , \new_[88527]_ , \new_[88528]_ , \new_[88532]_ ,
    \new_[88533]_ , \new_[88536]_ , \new_[88539]_ , \new_[88540]_ ,
    \new_[88541]_ , \new_[88544]_ , \new_[88547]_ , \new_[88548]_ ,
    \new_[88551]_ , \new_[88554]_ , \new_[88555]_ , \new_[88556]_ ,
    \new_[88560]_ , \new_[88561]_ , \new_[88564]_ , \new_[88567]_ ,
    \new_[88568]_ , \new_[88569]_ , \new_[88572]_ , \new_[88575]_ ,
    \new_[88576]_ , \new_[88579]_ , \new_[88582]_ , \new_[88583]_ ,
    \new_[88584]_ , \new_[88588]_ , \new_[88589]_ , \new_[88592]_ ,
    \new_[88595]_ , \new_[88596]_ , \new_[88597]_ , \new_[88600]_ ,
    \new_[88603]_ , \new_[88604]_ , \new_[88607]_ , \new_[88610]_ ,
    \new_[88611]_ , \new_[88612]_ , \new_[88616]_ , \new_[88617]_ ,
    \new_[88620]_ , \new_[88623]_ , \new_[88624]_ , \new_[88625]_ ,
    \new_[88628]_ , \new_[88631]_ , \new_[88632]_ , \new_[88635]_ ,
    \new_[88638]_ , \new_[88639]_ , \new_[88640]_ , \new_[88644]_ ,
    \new_[88645]_ , \new_[88648]_ , \new_[88651]_ , \new_[88652]_ ,
    \new_[88653]_ , \new_[88656]_ , \new_[88659]_ , \new_[88660]_ ,
    \new_[88663]_ , \new_[88666]_ , \new_[88667]_ , \new_[88668]_ ,
    \new_[88672]_ , \new_[88673]_ , \new_[88676]_ , \new_[88679]_ ,
    \new_[88680]_ , \new_[88681]_ , \new_[88684]_ , \new_[88687]_ ,
    \new_[88688]_ , \new_[88691]_ , \new_[88694]_ , \new_[88695]_ ,
    \new_[88696]_ , \new_[88700]_ , \new_[88701]_ , \new_[88704]_ ,
    \new_[88707]_ , \new_[88708]_ , \new_[88709]_ , \new_[88712]_ ,
    \new_[88715]_ , \new_[88716]_ , \new_[88719]_ , \new_[88722]_ ,
    \new_[88723]_ , \new_[88724]_ , \new_[88728]_ , \new_[88729]_ ,
    \new_[88732]_ , \new_[88735]_ , \new_[88736]_ , \new_[88737]_ ,
    \new_[88740]_ , \new_[88743]_ , \new_[88744]_ , \new_[88747]_ ,
    \new_[88750]_ , \new_[88751]_ , \new_[88752]_ , \new_[88756]_ ,
    \new_[88757]_ , \new_[88760]_ , \new_[88763]_ , \new_[88764]_ ,
    \new_[88765]_ , \new_[88768]_ , \new_[88771]_ , \new_[88772]_ ,
    \new_[88775]_ , \new_[88778]_ , \new_[88779]_ , \new_[88780]_ ,
    \new_[88784]_ , \new_[88785]_ , \new_[88788]_ , \new_[88791]_ ,
    \new_[88792]_ , \new_[88793]_ , \new_[88796]_ , \new_[88799]_ ,
    \new_[88800]_ , \new_[88803]_ , \new_[88806]_ , \new_[88807]_ ,
    \new_[88808]_ , \new_[88812]_ , \new_[88813]_ , \new_[88816]_ ,
    \new_[88819]_ , \new_[88820]_ , \new_[88821]_ , \new_[88824]_ ,
    \new_[88827]_ , \new_[88828]_ , \new_[88831]_ , \new_[88834]_ ,
    \new_[88835]_ , \new_[88836]_ , \new_[88840]_ , \new_[88841]_ ,
    \new_[88844]_ , \new_[88847]_ , \new_[88848]_ , \new_[88849]_ ,
    \new_[88852]_ , \new_[88855]_ , \new_[88856]_ , \new_[88859]_ ,
    \new_[88862]_ , \new_[88863]_ , \new_[88864]_ , \new_[88868]_ ,
    \new_[88869]_ , \new_[88872]_ , \new_[88875]_ , \new_[88876]_ ,
    \new_[88877]_ , \new_[88880]_ , \new_[88883]_ , \new_[88884]_ ,
    \new_[88887]_ , \new_[88890]_ , \new_[88891]_ , \new_[88892]_ ,
    \new_[88896]_ , \new_[88897]_ , \new_[88900]_ , \new_[88903]_ ,
    \new_[88904]_ , \new_[88905]_ , \new_[88908]_ , \new_[88911]_ ,
    \new_[88912]_ , \new_[88915]_ , \new_[88918]_ , \new_[88919]_ ,
    \new_[88920]_ , \new_[88924]_ , \new_[88925]_ , \new_[88928]_ ,
    \new_[88931]_ , \new_[88932]_ , \new_[88933]_ , \new_[88936]_ ,
    \new_[88939]_ , \new_[88940]_ , \new_[88943]_ , \new_[88946]_ ,
    \new_[88947]_ , \new_[88948]_ , \new_[88952]_ , \new_[88953]_ ,
    \new_[88956]_ , \new_[88959]_ , \new_[88960]_ , \new_[88961]_ ,
    \new_[88964]_ , \new_[88967]_ , \new_[88968]_ , \new_[88971]_ ,
    \new_[88974]_ , \new_[88975]_ , \new_[88976]_ , \new_[88980]_ ,
    \new_[88981]_ , \new_[88984]_ , \new_[88987]_ , \new_[88988]_ ,
    \new_[88989]_ , \new_[88992]_ , \new_[88995]_ , \new_[88996]_ ,
    \new_[88999]_ , \new_[89002]_ , \new_[89003]_ , \new_[89004]_ ,
    \new_[89008]_ , \new_[89009]_ , \new_[89012]_ , \new_[89015]_ ,
    \new_[89016]_ , \new_[89017]_ , \new_[89020]_ , \new_[89023]_ ,
    \new_[89024]_ , \new_[89027]_ , \new_[89030]_ , \new_[89031]_ ,
    \new_[89032]_ , \new_[89036]_ , \new_[89037]_ , \new_[89040]_ ,
    \new_[89043]_ , \new_[89044]_ , \new_[89045]_ , \new_[89048]_ ,
    \new_[89051]_ , \new_[89052]_ , \new_[89055]_ , \new_[89058]_ ,
    \new_[89059]_ , \new_[89060]_ , \new_[89064]_ , \new_[89065]_ ,
    \new_[89068]_ , \new_[89071]_ , \new_[89072]_ , \new_[89073]_ ,
    \new_[89076]_ , \new_[89079]_ , \new_[89080]_ , \new_[89083]_ ,
    \new_[89086]_ , \new_[89087]_ , \new_[89088]_ , \new_[89092]_ ,
    \new_[89093]_ , \new_[89096]_ , \new_[89099]_ , \new_[89100]_ ,
    \new_[89101]_ , \new_[89104]_ , \new_[89107]_ , \new_[89108]_ ,
    \new_[89111]_ , \new_[89114]_ , \new_[89115]_ , \new_[89116]_ ,
    \new_[89120]_ , \new_[89121]_ , \new_[89124]_ , \new_[89127]_ ,
    \new_[89128]_ , \new_[89129]_ , \new_[89132]_ , \new_[89135]_ ,
    \new_[89136]_ , \new_[89139]_ , \new_[89142]_ , \new_[89143]_ ,
    \new_[89144]_ , \new_[89148]_ , \new_[89149]_ , \new_[89152]_ ,
    \new_[89155]_ , \new_[89156]_ , \new_[89157]_ , \new_[89160]_ ,
    \new_[89163]_ , \new_[89164]_ , \new_[89167]_ , \new_[89170]_ ,
    \new_[89171]_ , \new_[89172]_ , \new_[89176]_ , \new_[89177]_ ,
    \new_[89180]_ , \new_[89183]_ , \new_[89184]_ , \new_[89185]_ ,
    \new_[89188]_ , \new_[89191]_ , \new_[89192]_ , \new_[89195]_ ,
    \new_[89198]_ , \new_[89199]_ , \new_[89200]_ , \new_[89204]_ ,
    \new_[89205]_ , \new_[89208]_ , \new_[89211]_ , \new_[89212]_ ,
    \new_[89213]_ , \new_[89216]_ , \new_[89219]_ , \new_[89220]_ ,
    \new_[89223]_ , \new_[89226]_ , \new_[89227]_ , \new_[89228]_ ,
    \new_[89232]_ , \new_[89233]_ , \new_[89236]_ , \new_[89239]_ ,
    \new_[89240]_ , \new_[89241]_ , \new_[89244]_ , \new_[89247]_ ,
    \new_[89248]_ , \new_[89251]_ , \new_[89254]_ , \new_[89255]_ ,
    \new_[89256]_ , \new_[89260]_ , \new_[89261]_ , \new_[89264]_ ,
    \new_[89267]_ , \new_[89268]_ , \new_[89269]_ , \new_[89272]_ ,
    \new_[89275]_ , \new_[89276]_ , \new_[89279]_ , \new_[89282]_ ,
    \new_[89283]_ , \new_[89284]_ , \new_[89288]_ , \new_[89289]_ ,
    \new_[89292]_ , \new_[89295]_ , \new_[89296]_ , \new_[89297]_ ,
    \new_[89300]_ , \new_[89303]_ , \new_[89304]_ , \new_[89307]_ ,
    \new_[89310]_ , \new_[89311]_ , \new_[89312]_ , \new_[89316]_ ,
    \new_[89317]_ , \new_[89320]_ , \new_[89323]_ , \new_[89324]_ ,
    \new_[89325]_ , \new_[89328]_ , \new_[89331]_ , \new_[89332]_ ,
    \new_[89335]_ , \new_[89338]_ , \new_[89339]_ , \new_[89340]_ ,
    \new_[89344]_ , \new_[89345]_ , \new_[89348]_ , \new_[89351]_ ,
    \new_[89352]_ , \new_[89353]_ , \new_[89356]_ , \new_[89359]_ ,
    \new_[89360]_ , \new_[89363]_ , \new_[89366]_ , \new_[89367]_ ,
    \new_[89368]_ , \new_[89372]_ , \new_[89373]_ , \new_[89376]_ ,
    \new_[89379]_ , \new_[89380]_ , \new_[89381]_ , \new_[89384]_ ,
    \new_[89387]_ , \new_[89388]_ , \new_[89391]_ , \new_[89394]_ ,
    \new_[89395]_ , \new_[89396]_ , \new_[89400]_ , \new_[89401]_ ,
    \new_[89404]_ , \new_[89407]_ , \new_[89408]_ , \new_[89409]_ ,
    \new_[89412]_ , \new_[89415]_ , \new_[89416]_ , \new_[89419]_ ,
    \new_[89422]_ , \new_[89423]_ , \new_[89424]_ , \new_[89428]_ ,
    \new_[89429]_ , \new_[89432]_ , \new_[89435]_ , \new_[89436]_ ,
    \new_[89437]_ , \new_[89440]_ , \new_[89443]_ , \new_[89444]_ ,
    \new_[89447]_ , \new_[89450]_ , \new_[89451]_ , \new_[89452]_ ,
    \new_[89456]_ , \new_[89457]_ , \new_[89460]_ , \new_[89463]_ ,
    \new_[89464]_ , \new_[89465]_ , \new_[89468]_ , \new_[89471]_ ,
    \new_[89472]_ , \new_[89475]_ , \new_[89478]_ , \new_[89479]_ ,
    \new_[89480]_ , \new_[89484]_ , \new_[89485]_ , \new_[89488]_ ,
    \new_[89491]_ , \new_[89492]_ , \new_[89493]_ , \new_[89496]_ ,
    \new_[89499]_ , \new_[89500]_ , \new_[89503]_ , \new_[89506]_ ,
    \new_[89507]_ , \new_[89508]_ , \new_[89511]_ , \new_[89514]_ ,
    \new_[89515]_ , \new_[89518]_ , \new_[89521]_ , \new_[89522]_ ,
    \new_[89523]_ , \new_[89526]_ , \new_[89529]_ , \new_[89530]_ ,
    \new_[89533]_ , \new_[89536]_ , \new_[89537]_ , \new_[89538]_ ,
    \new_[89541]_ , \new_[89544]_ , \new_[89545]_ , \new_[89548]_ ,
    \new_[89551]_ , \new_[89552]_ , \new_[89553]_ , \new_[89556]_ ,
    \new_[89559]_ , \new_[89560]_ , \new_[89563]_ , \new_[89566]_ ,
    \new_[89567]_ , \new_[89568]_ , \new_[89571]_ , \new_[89574]_ ,
    \new_[89575]_ , \new_[89578]_ , \new_[89581]_ , \new_[89582]_ ,
    \new_[89583]_ , \new_[89586]_ , \new_[89589]_ , \new_[89590]_ ,
    \new_[89593]_ , \new_[89596]_ , \new_[89597]_ , \new_[89598]_ ,
    \new_[89601]_ , \new_[89604]_ , \new_[89605]_ , \new_[89608]_ ,
    \new_[89611]_ , \new_[89612]_ , \new_[89613]_ , \new_[89616]_ ,
    \new_[89619]_ , \new_[89620]_ , \new_[89623]_ , \new_[89626]_ ,
    \new_[89627]_ , \new_[89628]_ , \new_[89631]_ , \new_[89634]_ ,
    \new_[89635]_ , \new_[89638]_ , \new_[89641]_ , \new_[89642]_ ,
    \new_[89643]_ , \new_[89646]_ , \new_[89649]_ , \new_[89650]_ ,
    \new_[89653]_ , \new_[89656]_ , \new_[89657]_ , \new_[89658]_ ,
    \new_[89661]_ , \new_[89664]_ , \new_[89665]_ , \new_[89668]_ ,
    \new_[89671]_ , \new_[89672]_ , \new_[89673]_ , \new_[89676]_ ,
    \new_[89679]_ , \new_[89680]_ , \new_[89683]_ , \new_[89686]_ ,
    \new_[89687]_ , \new_[89688]_ , \new_[89691]_ , \new_[89694]_ ,
    \new_[89695]_ , \new_[89698]_ , \new_[89701]_ , \new_[89702]_ ,
    \new_[89703]_ , \new_[89706]_ , \new_[89709]_ , \new_[89710]_ ,
    \new_[89713]_ , \new_[89716]_ , \new_[89717]_ , \new_[89718]_ ,
    \new_[89721]_ , \new_[89724]_ , \new_[89725]_ , \new_[89728]_ ,
    \new_[89731]_ , \new_[89732]_ , \new_[89733]_ , \new_[89736]_ ,
    \new_[89739]_ , \new_[89740]_ , \new_[89743]_ , \new_[89746]_ ,
    \new_[89747]_ , \new_[89748]_ , \new_[89751]_ , \new_[89754]_ ,
    \new_[89755]_ , \new_[89758]_ , \new_[89761]_ , \new_[89762]_ ,
    \new_[89763]_ , \new_[89766]_ , \new_[89769]_ , \new_[89770]_ ,
    \new_[89773]_ , \new_[89776]_ , \new_[89777]_ , \new_[89778]_ ,
    \new_[89781]_ , \new_[89784]_ , \new_[89785]_ , \new_[89788]_ ,
    \new_[89791]_ , \new_[89792]_ , \new_[89793]_ , \new_[89796]_ ,
    \new_[89799]_ , \new_[89800]_ , \new_[89803]_ , \new_[89806]_ ,
    \new_[89807]_ , \new_[89808]_ , \new_[89811]_ , \new_[89814]_ ,
    \new_[89815]_ , \new_[89818]_ , \new_[89821]_ , \new_[89822]_ ,
    \new_[89823]_ , \new_[89826]_ , \new_[89829]_ , \new_[89830]_ ,
    \new_[89833]_ , \new_[89836]_ , \new_[89837]_ , \new_[89838]_ ,
    \new_[89841]_ , \new_[89844]_ , \new_[89845]_ , \new_[89848]_ ,
    \new_[89851]_ , \new_[89852]_ , \new_[89853]_ , \new_[89856]_ ,
    \new_[89859]_ , \new_[89860]_ , \new_[89863]_ , \new_[89866]_ ,
    \new_[89867]_ , \new_[89868]_ , \new_[89871]_ , \new_[89874]_ ,
    \new_[89875]_ , \new_[89878]_ , \new_[89881]_ , \new_[89882]_ ,
    \new_[89883]_ , \new_[89886]_ , \new_[89889]_ , \new_[89890]_ ,
    \new_[89893]_ , \new_[89896]_ , \new_[89897]_ , \new_[89898]_ ,
    \new_[89901]_ , \new_[89904]_ , \new_[89905]_ , \new_[89908]_ ,
    \new_[89911]_ , \new_[89912]_ , \new_[89913]_ , \new_[89916]_ ,
    \new_[89919]_ , \new_[89920]_ , \new_[89923]_ , \new_[89926]_ ,
    \new_[89927]_ , \new_[89928]_ , \new_[89931]_ , \new_[89934]_ ,
    \new_[89935]_ , \new_[89938]_ , \new_[89941]_ , \new_[89942]_ ,
    \new_[89943]_ , \new_[89946]_ , \new_[89949]_ , \new_[89950]_ ,
    \new_[89953]_ , \new_[89956]_ , \new_[89957]_ , \new_[89958]_ ,
    \new_[89961]_ , \new_[89964]_ , \new_[89965]_ , \new_[89968]_ ,
    \new_[89971]_ , \new_[89972]_ , \new_[89973]_ , \new_[89976]_ ,
    \new_[89979]_ , \new_[89980]_ , \new_[89983]_ , \new_[89986]_ ,
    \new_[89987]_ , \new_[89988]_ , \new_[89991]_ , \new_[89994]_ ,
    \new_[89995]_ , \new_[89998]_ , \new_[90001]_ , \new_[90002]_ ,
    \new_[90003]_ , \new_[90006]_ , \new_[90009]_ , \new_[90010]_ ,
    \new_[90013]_ , \new_[90016]_ , \new_[90017]_ , \new_[90018]_ ,
    \new_[90021]_ , \new_[90024]_ , \new_[90025]_ , \new_[90028]_ ,
    \new_[90031]_ , \new_[90032]_ , \new_[90033]_ , \new_[90036]_ ,
    \new_[90039]_ , \new_[90040]_ , \new_[90043]_ , \new_[90046]_ ,
    \new_[90047]_ , \new_[90048]_ , \new_[90051]_ , \new_[90054]_ ,
    \new_[90055]_ , \new_[90058]_ , \new_[90061]_ , \new_[90062]_ ,
    \new_[90063]_ , \new_[90066]_ , \new_[90069]_ , \new_[90070]_ ,
    \new_[90073]_ , \new_[90076]_ , \new_[90077]_ , \new_[90078]_ ,
    \new_[90081]_ , \new_[90084]_ , \new_[90085]_ , \new_[90088]_ ,
    \new_[90091]_ , \new_[90092]_ , \new_[90093]_ , \new_[90096]_ ,
    \new_[90099]_ , \new_[90100]_ , \new_[90103]_ , \new_[90106]_ ,
    \new_[90107]_ , \new_[90108]_ , \new_[90111]_ , \new_[90114]_ ,
    \new_[90115]_ , \new_[90118]_ , \new_[90121]_ , \new_[90122]_ ,
    \new_[90123]_ , \new_[90126]_ , \new_[90129]_ , \new_[90130]_ ,
    \new_[90133]_ , \new_[90136]_ , \new_[90137]_ , \new_[90138]_ ,
    \new_[90141]_ , \new_[90144]_ , \new_[90145]_ , \new_[90148]_ ,
    \new_[90151]_ , \new_[90152]_ , \new_[90153]_ , \new_[90156]_ ,
    \new_[90159]_ , \new_[90160]_ , \new_[90163]_ , \new_[90166]_ ,
    \new_[90167]_ , \new_[90168]_ , \new_[90171]_ , \new_[90174]_ ,
    \new_[90175]_ , \new_[90178]_ , \new_[90181]_ , \new_[90182]_ ,
    \new_[90183]_ , \new_[90186]_ , \new_[90189]_ , \new_[90190]_ ,
    \new_[90193]_ , \new_[90196]_ , \new_[90197]_ , \new_[90198]_ ,
    \new_[90201]_ , \new_[90204]_ , \new_[90205]_ , \new_[90208]_ ,
    \new_[90211]_ , \new_[90212]_ , \new_[90213]_ , \new_[90216]_ ,
    \new_[90219]_ , \new_[90220]_ , \new_[90223]_ , \new_[90226]_ ,
    \new_[90227]_ , \new_[90228]_ , \new_[90231]_ , \new_[90234]_ ,
    \new_[90235]_ , \new_[90238]_ , \new_[90241]_ , \new_[90242]_ ,
    \new_[90243]_ , \new_[90246]_ , \new_[90249]_ , \new_[90250]_ ,
    \new_[90253]_ , \new_[90256]_ , \new_[90257]_ , \new_[90258]_ ,
    \new_[90261]_ , \new_[90264]_ , \new_[90265]_ , \new_[90268]_ ,
    \new_[90271]_ , \new_[90272]_ , \new_[90273]_ , \new_[90276]_ ,
    \new_[90279]_ , \new_[90280]_ , \new_[90283]_ , \new_[90286]_ ,
    \new_[90287]_ , \new_[90288]_ , \new_[90291]_ , \new_[90294]_ ,
    \new_[90295]_ , \new_[90298]_ , \new_[90301]_ , \new_[90302]_ ,
    \new_[90303]_ , \new_[90306]_ , \new_[90309]_ , \new_[90310]_ ,
    \new_[90313]_ , \new_[90316]_ , \new_[90317]_ , \new_[90318]_ ,
    \new_[90321]_ , \new_[90324]_ , \new_[90325]_ , \new_[90328]_ ,
    \new_[90331]_ , \new_[90332]_ , \new_[90333]_ , \new_[90336]_ ,
    \new_[90339]_ , \new_[90340]_ , \new_[90343]_ , \new_[90346]_ ,
    \new_[90347]_ , \new_[90348]_ , \new_[90351]_ , \new_[90354]_ ,
    \new_[90355]_ , \new_[90358]_ , \new_[90361]_ , \new_[90362]_ ,
    \new_[90363]_ , \new_[90366]_ , \new_[90369]_ , \new_[90370]_ ,
    \new_[90373]_ , \new_[90376]_ , \new_[90377]_ , \new_[90378]_ ,
    \new_[90381]_ , \new_[90384]_ , \new_[90385]_ , \new_[90388]_ ,
    \new_[90391]_ , \new_[90392]_ , \new_[90393]_ , \new_[90396]_ ,
    \new_[90399]_ , \new_[90400]_ , \new_[90403]_ , \new_[90406]_ ,
    \new_[90407]_ , \new_[90408]_ , \new_[90411]_ , \new_[90414]_ ,
    \new_[90415]_ , \new_[90418]_ , \new_[90421]_ , \new_[90422]_ ,
    \new_[90423]_ , \new_[90426]_ , \new_[90429]_ , \new_[90430]_ ,
    \new_[90433]_ , \new_[90436]_ , \new_[90437]_ , \new_[90438]_ ,
    \new_[90441]_ , \new_[90444]_ , \new_[90445]_ , \new_[90448]_ ,
    \new_[90451]_ , \new_[90452]_ , \new_[90453]_ , \new_[90456]_ ,
    \new_[90459]_ , \new_[90460]_ , \new_[90463]_ , \new_[90466]_ ,
    \new_[90467]_ , \new_[90468]_ , \new_[90471]_ , \new_[90474]_ ,
    \new_[90475]_ , \new_[90478]_ , \new_[90481]_ , \new_[90482]_ ,
    \new_[90483]_ , \new_[90486]_ , \new_[90489]_ , \new_[90490]_ ,
    \new_[90493]_ , \new_[90496]_ , \new_[90497]_ , \new_[90498]_ ,
    \new_[90501]_ , \new_[90504]_ , \new_[90505]_ , \new_[90508]_ ,
    \new_[90511]_ , \new_[90512]_ , \new_[90513]_ , \new_[90516]_ ,
    \new_[90519]_ , \new_[90520]_ , \new_[90523]_ , \new_[90526]_ ,
    \new_[90527]_ , \new_[90528]_ , \new_[90531]_ , \new_[90534]_ ,
    \new_[90535]_ , \new_[90538]_ , \new_[90541]_ , \new_[90542]_ ,
    \new_[90543]_ , \new_[90546]_ , \new_[90549]_ , \new_[90550]_ ,
    \new_[90553]_ , \new_[90556]_ , \new_[90557]_ , \new_[90558]_ ,
    \new_[90561]_ , \new_[90564]_ , \new_[90565]_ , \new_[90568]_ ,
    \new_[90571]_ , \new_[90572]_ , \new_[90573]_ , \new_[90576]_ ,
    \new_[90579]_ , \new_[90580]_ , \new_[90583]_ , \new_[90586]_ ,
    \new_[90587]_ , \new_[90588]_ , \new_[90591]_ , \new_[90594]_ ,
    \new_[90595]_ , \new_[90598]_ , \new_[90601]_ , \new_[90602]_ ,
    \new_[90603]_ , \new_[90606]_ , \new_[90609]_ , \new_[90610]_ ,
    \new_[90613]_ , \new_[90616]_ , \new_[90617]_ , \new_[90618]_ ,
    \new_[90621]_ , \new_[90624]_ , \new_[90625]_ , \new_[90628]_ ,
    \new_[90631]_ , \new_[90632]_ , \new_[90633]_ , \new_[90636]_ ,
    \new_[90639]_ , \new_[90640]_ , \new_[90643]_ , \new_[90646]_ ,
    \new_[90647]_ , \new_[90648]_ , \new_[90651]_ , \new_[90654]_ ,
    \new_[90655]_ , \new_[90658]_ , \new_[90661]_ , \new_[90662]_ ,
    \new_[90663]_ , \new_[90666]_ , \new_[90669]_ , \new_[90670]_ ,
    \new_[90673]_ , \new_[90676]_ , \new_[90677]_ , \new_[90678]_ ,
    \new_[90681]_ , \new_[90684]_ , \new_[90685]_ , \new_[90688]_ ,
    \new_[90691]_ , \new_[90692]_ , \new_[90693]_ , \new_[90696]_ ,
    \new_[90699]_ , \new_[90700]_ , \new_[90703]_ , \new_[90706]_ ,
    \new_[90707]_ , \new_[90708]_ , \new_[90711]_ , \new_[90714]_ ,
    \new_[90715]_ , \new_[90718]_ , \new_[90721]_ , \new_[90722]_ ,
    \new_[90723]_ , \new_[90726]_ , \new_[90729]_ , \new_[90730]_ ,
    \new_[90733]_ , \new_[90736]_ , \new_[90737]_ , \new_[90738]_ ,
    \new_[90741]_ , \new_[90744]_ , \new_[90745]_ , \new_[90748]_ ,
    \new_[90751]_ , \new_[90752]_ , \new_[90753]_ , \new_[90756]_ ,
    \new_[90759]_ , \new_[90760]_ , \new_[90763]_ , \new_[90766]_ ,
    \new_[90767]_ , \new_[90768]_ , \new_[90771]_ , \new_[90774]_ ,
    \new_[90775]_ , \new_[90778]_ , \new_[90781]_ , \new_[90782]_ ,
    \new_[90783]_ , \new_[90786]_ , \new_[90789]_ , \new_[90790]_ ,
    \new_[90793]_ , \new_[90796]_ , \new_[90797]_ , \new_[90798]_ ,
    \new_[90801]_ , \new_[90804]_ , \new_[90805]_ , \new_[90808]_ ,
    \new_[90811]_ , \new_[90812]_ , \new_[90813]_ , \new_[90816]_ ,
    \new_[90819]_ , \new_[90820]_ , \new_[90823]_ , \new_[90826]_ ,
    \new_[90827]_ , \new_[90828]_ , \new_[90831]_ , \new_[90834]_ ,
    \new_[90835]_ , \new_[90838]_ , \new_[90841]_ , \new_[90842]_ ,
    \new_[90843]_ , \new_[90846]_ , \new_[90849]_ , \new_[90850]_ ,
    \new_[90853]_ , \new_[90856]_ , \new_[90857]_ , \new_[90858]_ ,
    \new_[90861]_ , \new_[90864]_ , \new_[90865]_ , \new_[90868]_ ,
    \new_[90871]_ , \new_[90872]_ , \new_[90873]_ , \new_[90876]_ ,
    \new_[90879]_ , \new_[90880]_ , \new_[90883]_ , \new_[90886]_ ,
    \new_[90887]_ , \new_[90888]_ , \new_[90891]_ , \new_[90894]_ ,
    \new_[90895]_ , \new_[90898]_ , \new_[90901]_ , \new_[90902]_ ,
    \new_[90903]_ , \new_[90906]_ , \new_[90909]_ , \new_[90910]_ ,
    \new_[90913]_ , \new_[90916]_ , \new_[90917]_ , \new_[90918]_ ,
    \new_[90921]_ , \new_[90924]_ , \new_[90925]_ , \new_[90928]_ ,
    \new_[90931]_ , \new_[90932]_ , \new_[90933]_ , \new_[90936]_ ,
    \new_[90939]_ , \new_[90940]_ , \new_[90943]_ , \new_[90946]_ ,
    \new_[90947]_ , \new_[90948]_ , \new_[90951]_ , \new_[90954]_ ,
    \new_[90955]_ , \new_[90958]_ , \new_[90961]_ , \new_[90962]_ ,
    \new_[90963]_ , \new_[90966]_ , \new_[90969]_ , \new_[90970]_ ,
    \new_[90973]_ , \new_[90976]_ , \new_[90977]_ , \new_[90978]_ ,
    \new_[90981]_ , \new_[90984]_ , \new_[90985]_ , \new_[90988]_ ,
    \new_[90991]_ , \new_[90992]_ , \new_[90993]_ , \new_[90996]_ ,
    \new_[90999]_ , \new_[91000]_ , \new_[91003]_ , \new_[91006]_ ,
    \new_[91007]_ , \new_[91008]_ , \new_[91011]_ , \new_[91014]_ ,
    \new_[91015]_ , \new_[91018]_ , \new_[91021]_ , \new_[91022]_ ,
    \new_[91023]_ , \new_[91026]_ , \new_[91029]_ , \new_[91030]_ ,
    \new_[91033]_ , \new_[91036]_ , \new_[91037]_ , \new_[91038]_ ,
    \new_[91041]_ , \new_[91044]_ , \new_[91045]_ , \new_[91048]_ ,
    \new_[91051]_ , \new_[91052]_ , \new_[91053]_ , \new_[91056]_ ,
    \new_[91059]_ , \new_[91060]_ , \new_[91063]_ , \new_[91066]_ ,
    \new_[91067]_ , \new_[91068]_ , \new_[91071]_ , \new_[91074]_ ,
    \new_[91075]_ , \new_[91078]_ , \new_[91081]_ , \new_[91082]_ ,
    \new_[91083]_ , \new_[91086]_ , \new_[91089]_ , \new_[91090]_ ,
    \new_[91093]_ , \new_[91096]_ , \new_[91097]_ , \new_[91098]_ ,
    \new_[91101]_ , \new_[91104]_ , \new_[91105]_ , \new_[91108]_ ,
    \new_[91111]_ , \new_[91112]_ , \new_[91113]_ , \new_[91116]_ ,
    \new_[91119]_ , \new_[91120]_ , \new_[91123]_ , \new_[91126]_ ,
    \new_[91127]_ , \new_[91128]_ , \new_[91131]_ , \new_[91134]_ ,
    \new_[91135]_ , \new_[91138]_ , \new_[91141]_ , \new_[91142]_ ,
    \new_[91143]_ , \new_[91146]_ , \new_[91149]_ , \new_[91150]_ ,
    \new_[91153]_ , \new_[91156]_ , \new_[91157]_ , \new_[91158]_ ,
    \new_[91161]_ , \new_[91164]_ , \new_[91165]_ , \new_[91168]_ ,
    \new_[91171]_ , \new_[91172]_ , \new_[91173]_ , \new_[91176]_ ,
    \new_[91179]_ , \new_[91180]_ , \new_[91183]_ , \new_[91186]_ ,
    \new_[91187]_ , \new_[91188]_ , \new_[91191]_ , \new_[91194]_ ,
    \new_[91195]_ , \new_[91198]_ , \new_[91201]_ , \new_[91202]_ ,
    \new_[91203]_ , \new_[91206]_ , \new_[91209]_ , \new_[91210]_ ,
    \new_[91213]_ , \new_[91216]_ , \new_[91217]_ , \new_[91218]_ ,
    \new_[91221]_ , \new_[91224]_ , \new_[91225]_ , \new_[91228]_ ,
    \new_[91231]_ , \new_[91232]_ , \new_[91233]_ , \new_[91236]_ ,
    \new_[91239]_ , \new_[91240]_ , \new_[91243]_ , \new_[91246]_ ,
    \new_[91247]_ , \new_[91248]_ , \new_[91251]_ , \new_[91254]_ ,
    \new_[91255]_ , \new_[91258]_ , \new_[91261]_ , \new_[91262]_ ,
    \new_[91263]_ , \new_[91266]_ , \new_[91269]_ , \new_[91270]_ ,
    \new_[91273]_ , \new_[91276]_ , \new_[91277]_ , \new_[91278]_ ,
    \new_[91281]_ , \new_[91284]_ , \new_[91285]_ , \new_[91288]_ ,
    \new_[91291]_ , \new_[91292]_ , \new_[91293]_ , \new_[91296]_ ,
    \new_[91299]_ , \new_[91300]_ , \new_[91303]_ , \new_[91306]_ ,
    \new_[91307]_ , \new_[91308]_ , \new_[91311]_ , \new_[91314]_ ,
    \new_[91315]_ , \new_[91318]_ , \new_[91321]_ , \new_[91322]_ ,
    \new_[91323]_ , \new_[91326]_ , \new_[91329]_ , \new_[91330]_ ,
    \new_[91333]_ , \new_[91336]_ , \new_[91337]_ , \new_[91338]_ ,
    \new_[91341]_ , \new_[91344]_ , \new_[91345]_ , \new_[91348]_ ,
    \new_[91351]_ , \new_[91352]_ , \new_[91353]_ , \new_[91356]_ ,
    \new_[91359]_ , \new_[91360]_ , \new_[91363]_ , \new_[91366]_ ,
    \new_[91367]_ , \new_[91368]_ , \new_[91371]_ , \new_[91374]_ ,
    \new_[91375]_ , \new_[91378]_ , \new_[91381]_ , \new_[91382]_ ,
    \new_[91383]_ , \new_[91386]_ , \new_[91389]_ , \new_[91390]_ ,
    \new_[91393]_ , \new_[91396]_ , \new_[91397]_ , \new_[91398]_ ,
    \new_[91401]_ , \new_[91404]_ , \new_[91405]_ , \new_[91408]_ ,
    \new_[91411]_ , \new_[91412]_ , \new_[91413]_ , \new_[91416]_ ,
    \new_[91419]_ , \new_[91420]_ , \new_[91423]_ , \new_[91426]_ ,
    \new_[91427]_ , \new_[91428]_ , \new_[91431]_ , \new_[91434]_ ,
    \new_[91435]_ , \new_[91438]_ , \new_[91441]_ , \new_[91442]_ ,
    \new_[91443]_ , \new_[91446]_ , \new_[91449]_ , \new_[91450]_ ,
    \new_[91453]_ , \new_[91456]_ , \new_[91457]_ , \new_[91458]_ ,
    \new_[91461]_ , \new_[91464]_ , \new_[91465]_ , \new_[91468]_ ,
    \new_[91471]_ , \new_[91472]_ , \new_[91473]_ , \new_[91476]_ ,
    \new_[91479]_ , \new_[91480]_ , \new_[91483]_ , \new_[91486]_ ,
    \new_[91487]_ , \new_[91488]_ , \new_[91491]_ , \new_[91494]_ ,
    \new_[91495]_ , \new_[91498]_ , \new_[91501]_ , \new_[91502]_ ,
    \new_[91503]_ , \new_[91506]_ , \new_[91509]_ , \new_[91510]_ ,
    \new_[91513]_ , \new_[91516]_ , \new_[91517]_ , \new_[91518]_ ,
    \new_[91521]_ , \new_[91524]_ , \new_[91525]_ , \new_[91528]_ ,
    \new_[91531]_ , \new_[91532]_ , \new_[91533]_ , \new_[91536]_ ,
    \new_[91539]_ , \new_[91540]_ , \new_[91543]_ , \new_[91546]_ ,
    \new_[91547]_ , \new_[91548]_ , \new_[91551]_ , \new_[91554]_ ,
    \new_[91555]_ , \new_[91558]_ , \new_[91561]_ , \new_[91562]_ ,
    \new_[91563]_ , \new_[91566]_ , \new_[91569]_ , \new_[91570]_ ,
    \new_[91573]_ , \new_[91576]_ , \new_[91577]_ , \new_[91578]_ ,
    \new_[91581]_ , \new_[91584]_ , \new_[91585]_ , \new_[91588]_ ,
    \new_[91591]_ , \new_[91592]_ , \new_[91593]_ , \new_[91596]_ ,
    \new_[91599]_ , \new_[91600]_ , \new_[91603]_ , \new_[91606]_ ,
    \new_[91607]_ , \new_[91608]_ , \new_[91611]_ , \new_[91614]_ ,
    \new_[91615]_ , \new_[91618]_ , \new_[91621]_ , \new_[91622]_ ,
    \new_[91623]_ , \new_[91626]_ , \new_[91629]_ , \new_[91630]_ ,
    \new_[91633]_ , \new_[91636]_ , \new_[91637]_ , \new_[91638]_ ,
    \new_[91641]_ , \new_[91644]_ , \new_[91645]_ , \new_[91648]_ ,
    \new_[91651]_ , \new_[91652]_ , \new_[91653]_ , \new_[91656]_ ,
    \new_[91659]_ , \new_[91660]_ , \new_[91663]_ , \new_[91666]_ ,
    \new_[91667]_ , \new_[91668]_ , \new_[91671]_ , \new_[91674]_ ,
    \new_[91675]_ , \new_[91678]_ , \new_[91681]_ , \new_[91682]_ ,
    \new_[91683]_ , \new_[91686]_ , \new_[91689]_ , \new_[91690]_ ,
    \new_[91693]_ , \new_[91696]_ , \new_[91697]_ , \new_[91698]_ ,
    \new_[91701]_ , \new_[91704]_ , \new_[91705]_ , \new_[91708]_ ,
    \new_[91711]_ , \new_[91712]_ , \new_[91713]_ , \new_[91716]_ ,
    \new_[91719]_ , \new_[91720]_ , \new_[91723]_ , \new_[91726]_ ,
    \new_[91727]_ , \new_[91728]_ , \new_[91731]_ , \new_[91734]_ ,
    \new_[91735]_ , \new_[91738]_ , \new_[91741]_ , \new_[91742]_ ,
    \new_[91743]_ , \new_[91746]_ , \new_[91749]_ , \new_[91750]_ ,
    \new_[91753]_ , \new_[91756]_ , \new_[91757]_ , \new_[91758]_ ,
    \new_[91761]_ , \new_[91764]_ , \new_[91765]_ , \new_[91768]_ ,
    \new_[91771]_ , \new_[91772]_ , \new_[91773]_ , \new_[91776]_ ,
    \new_[91779]_ , \new_[91780]_ , \new_[91783]_ , \new_[91786]_ ,
    \new_[91787]_ , \new_[91788]_ , \new_[91791]_ , \new_[91794]_ ,
    \new_[91795]_ , \new_[91798]_ , \new_[91801]_ , \new_[91802]_ ,
    \new_[91803]_ , \new_[91806]_ , \new_[91809]_ , \new_[91810]_ ,
    \new_[91813]_ , \new_[91816]_ , \new_[91817]_ , \new_[91818]_ ,
    \new_[91821]_ , \new_[91824]_ , \new_[91825]_ , \new_[91828]_ ,
    \new_[91831]_ , \new_[91832]_ , \new_[91833]_ , \new_[91836]_ ,
    \new_[91839]_ , \new_[91840]_ , \new_[91843]_ , \new_[91846]_ ,
    \new_[91847]_ , \new_[91848]_ , \new_[91851]_ , \new_[91854]_ ,
    \new_[91855]_ , \new_[91858]_ , \new_[91861]_ , \new_[91862]_ ,
    \new_[91863]_ , \new_[91866]_ , \new_[91869]_ , \new_[91870]_ ,
    \new_[91873]_ , \new_[91876]_ , \new_[91877]_ , \new_[91878]_ ,
    \new_[91881]_ , \new_[91884]_ , \new_[91885]_ , \new_[91888]_ ,
    \new_[91891]_ , \new_[91892]_ , \new_[91893]_ , \new_[91896]_ ,
    \new_[91899]_ , \new_[91900]_ , \new_[91903]_ , \new_[91906]_ ,
    \new_[91907]_ , \new_[91908]_ , \new_[91911]_ , \new_[91914]_ ,
    \new_[91915]_ , \new_[91918]_ , \new_[91921]_ , \new_[91922]_ ,
    \new_[91923]_ , \new_[91926]_ , \new_[91929]_ , \new_[91930]_ ,
    \new_[91933]_ , \new_[91936]_ , \new_[91937]_ , \new_[91938]_ ,
    \new_[91941]_ , \new_[91944]_ , \new_[91945]_ , \new_[91948]_ ,
    \new_[91951]_ , \new_[91952]_ , \new_[91953]_ , \new_[91956]_ ,
    \new_[91959]_ , \new_[91960]_ , \new_[91963]_ , \new_[91966]_ ,
    \new_[91967]_ , \new_[91968]_ , \new_[91971]_ , \new_[91974]_ ,
    \new_[91975]_ , \new_[91978]_ , \new_[91981]_ , \new_[91982]_ ,
    \new_[91983]_ , \new_[91986]_ , \new_[91989]_ , \new_[91990]_ ,
    \new_[91993]_ , \new_[91996]_ , \new_[91997]_ , \new_[91998]_ ,
    \new_[92001]_ , \new_[92004]_ , \new_[92005]_ , \new_[92008]_ ,
    \new_[92011]_ , \new_[92012]_ , \new_[92013]_ , \new_[92016]_ ,
    \new_[92019]_ , \new_[92020]_ , \new_[92023]_ , \new_[92026]_ ,
    \new_[92027]_ , \new_[92028]_ , \new_[92031]_ , \new_[92034]_ ,
    \new_[92035]_ , \new_[92038]_ , \new_[92041]_ , \new_[92042]_ ,
    \new_[92043]_ , \new_[92046]_ , \new_[92049]_ , \new_[92050]_ ,
    \new_[92053]_ , \new_[92056]_ , \new_[92057]_ , \new_[92058]_ ,
    \new_[92061]_ , \new_[92064]_ , \new_[92065]_ , \new_[92068]_ ,
    \new_[92071]_ , \new_[92072]_ , \new_[92073]_ , \new_[92076]_ ,
    \new_[92079]_ , \new_[92080]_ , \new_[92083]_ , \new_[92086]_ ,
    \new_[92087]_ , \new_[92088]_ , \new_[92091]_ , \new_[92094]_ ,
    \new_[92095]_ , \new_[92098]_ , \new_[92101]_ , \new_[92102]_ ,
    \new_[92103]_ , \new_[92106]_ , \new_[92109]_ , \new_[92110]_ ,
    \new_[92113]_ , \new_[92116]_ , \new_[92117]_ , \new_[92118]_ ,
    \new_[92121]_ , \new_[92124]_ , \new_[92125]_ , \new_[92128]_ ,
    \new_[92131]_ , \new_[92132]_ , \new_[92133]_ , \new_[92136]_ ,
    \new_[92139]_ , \new_[92140]_ , \new_[92143]_ , \new_[92146]_ ,
    \new_[92147]_ , \new_[92148]_ , \new_[92151]_ , \new_[92154]_ ,
    \new_[92155]_ , \new_[92158]_ , \new_[92161]_ , \new_[92162]_ ,
    \new_[92163]_ , \new_[92166]_ , \new_[92169]_ , \new_[92170]_ ,
    \new_[92173]_ , \new_[92176]_ , \new_[92177]_ , \new_[92178]_ ,
    \new_[92181]_ , \new_[92184]_ , \new_[92185]_ , \new_[92188]_ ,
    \new_[92191]_ , \new_[92192]_ , \new_[92193]_ , \new_[92196]_ ,
    \new_[92199]_ , \new_[92200]_ , \new_[92203]_ , \new_[92206]_ ,
    \new_[92207]_ , \new_[92208]_ , \new_[92211]_ , \new_[92214]_ ,
    \new_[92215]_ , \new_[92218]_ , \new_[92221]_ , \new_[92222]_ ,
    \new_[92223]_ , \new_[92226]_ , \new_[92229]_ , \new_[92230]_ ,
    \new_[92233]_ , \new_[92236]_ , \new_[92237]_ , \new_[92238]_ ,
    \new_[92241]_ , \new_[92244]_ , \new_[92245]_ , \new_[92248]_ ,
    \new_[92251]_ , \new_[92252]_ , \new_[92253]_ , \new_[92256]_ ,
    \new_[92259]_ , \new_[92260]_ , \new_[92263]_ , \new_[92266]_ ,
    \new_[92267]_ , \new_[92268]_ , \new_[92271]_ , \new_[92274]_ ,
    \new_[92275]_ , \new_[92278]_ , \new_[92281]_ , \new_[92282]_ ,
    \new_[92283]_ , \new_[92286]_ , \new_[92289]_ , \new_[92290]_ ,
    \new_[92293]_ , \new_[92296]_ , \new_[92297]_ , \new_[92298]_ ,
    \new_[92301]_ , \new_[92304]_ , \new_[92305]_ , \new_[92308]_ ,
    \new_[92311]_ , \new_[92312]_ , \new_[92313]_ , \new_[92316]_ ,
    \new_[92319]_ , \new_[92320]_ , \new_[92323]_ , \new_[92326]_ ,
    \new_[92327]_ , \new_[92328]_ , \new_[92331]_ , \new_[92334]_ ,
    \new_[92335]_ , \new_[92338]_ , \new_[92341]_ , \new_[92342]_ ,
    \new_[92343]_ , \new_[92346]_ , \new_[92349]_ , \new_[92350]_ ,
    \new_[92353]_ , \new_[92356]_ , \new_[92357]_ , \new_[92358]_ ,
    \new_[92361]_ , \new_[92364]_ , \new_[92365]_ , \new_[92368]_ ,
    \new_[92371]_ , \new_[92372]_ , \new_[92373]_ , \new_[92376]_ ,
    \new_[92379]_ , \new_[92380]_ , \new_[92383]_ , \new_[92386]_ ,
    \new_[92387]_ , \new_[92388]_ , \new_[92391]_ , \new_[92394]_ ,
    \new_[92395]_ , \new_[92398]_ , \new_[92401]_ , \new_[92402]_ ,
    \new_[92403]_ , \new_[92406]_ , \new_[92409]_ , \new_[92410]_ ,
    \new_[92413]_ , \new_[92416]_ , \new_[92417]_ , \new_[92418]_ ,
    \new_[92421]_ , \new_[92424]_ , \new_[92425]_ , \new_[92428]_ ,
    \new_[92431]_ , \new_[92432]_ , \new_[92433]_ , \new_[92436]_ ,
    \new_[92439]_ , \new_[92440]_ , \new_[92443]_ , \new_[92446]_ ,
    \new_[92447]_ , \new_[92448]_ , \new_[92451]_ , \new_[92454]_ ,
    \new_[92455]_ , \new_[92458]_ , \new_[92461]_ , \new_[92462]_ ,
    \new_[92463]_ , \new_[92466]_ , \new_[92469]_ , \new_[92470]_ ,
    \new_[92473]_ , \new_[92476]_ , \new_[92477]_ , \new_[92478]_ ,
    \new_[92481]_ , \new_[92484]_ , \new_[92485]_ , \new_[92488]_ ,
    \new_[92491]_ , \new_[92492]_ , \new_[92493]_ , \new_[92496]_ ,
    \new_[92499]_ , \new_[92500]_ , \new_[92503]_ , \new_[92506]_ ,
    \new_[92507]_ , \new_[92508]_ , \new_[92511]_ , \new_[92514]_ ,
    \new_[92515]_ , \new_[92518]_ , \new_[92521]_ , \new_[92522]_ ,
    \new_[92523]_ , \new_[92526]_ , \new_[92529]_ , \new_[92530]_ ,
    \new_[92533]_ , \new_[92536]_ , \new_[92537]_ , \new_[92538]_ ,
    \new_[92541]_ , \new_[92544]_ , \new_[92545]_ , \new_[92548]_ ,
    \new_[92551]_ , \new_[92552]_ , \new_[92553]_ , \new_[92556]_ ,
    \new_[92559]_ , \new_[92560]_ , \new_[92563]_ , \new_[92566]_ ,
    \new_[92567]_ , \new_[92568]_ , \new_[92571]_ , \new_[92574]_ ,
    \new_[92575]_ , \new_[92578]_ , \new_[92581]_ , \new_[92582]_ ,
    \new_[92583]_ , \new_[92586]_ , \new_[92589]_ , \new_[92590]_ ,
    \new_[92593]_ , \new_[92596]_ , \new_[92597]_ , \new_[92598]_ ,
    \new_[92601]_ , \new_[92604]_ , \new_[92605]_ , \new_[92608]_ ,
    \new_[92611]_ , \new_[92612]_ , \new_[92613]_ , \new_[92616]_ ,
    \new_[92619]_ , \new_[92620]_ , \new_[92623]_ , \new_[92626]_ ,
    \new_[92627]_ , \new_[92628]_ , \new_[92631]_ , \new_[92634]_ ,
    \new_[92635]_ , \new_[92638]_ , \new_[92641]_ , \new_[92642]_ ,
    \new_[92643]_ , \new_[92646]_ , \new_[92649]_ , \new_[92650]_ ,
    \new_[92653]_ , \new_[92656]_ , \new_[92657]_ , \new_[92658]_ ,
    \new_[92661]_ , \new_[92664]_ , \new_[92665]_ , \new_[92668]_ ,
    \new_[92671]_ , \new_[92672]_ , \new_[92673]_ , \new_[92676]_ ,
    \new_[92679]_ , \new_[92680]_ , \new_[92683]_ , \new_[92686]_ ,
    \new_[92687]_ , \new_[92688]_ , \new_[92691]_ , \new_[92694]_ ,
    \new_[92695]_ , \new_[92698]_ , \new_[92701]_ , \new_[92702]_ ,
    \new_[92703]_ , \new_[92706]_ , \new_[92709]_ , \new_[92710]_ ,
    \new_[92713]_ , \new_[92716]_ , \new_[92717]_ , \new_[92718]_ ,
    \new_[92721]_ , \new_[92724]_ , \new_[92725]_ , \new_[92728]_ ,
    \new_[92731]_ , \new_[92732]_ , \new_[92733]_ , \new_[92736]_ ,
    \new_[92739]_ , \new_[92740]_ , \new_[92743]_ , \new_[92746]_ ,
    \new_[92747]_ , \new_[92748]_ , \new_[92751]_ , \new_[92754]_ ,
    \new_[92755]_ , \new_[92758]_ , \new_[92761]_ , \new_[92762]_ ,
    \new_[92763]_ , \new_[92766]_ , \new_[92769]_ , \new_[92770]_ ,
    \new_[92773]_ , \new_[92776]_ , \new_[92777]_ , \new_[92778]_ ,
    \new_[92781]_ , \new_[92784]_ , \new_[92785]_ , \new_[92788]_ ,
    \new_[92791]_ , \new_[92792]_ , \new_[92793]_ , \new_[92796]_ ,
    \new_[92799]_ , \new_[92800]_ , \new_[92803]_ , \new_[92806]_ ,
    \new_[92807]_ , \new_[92808]_ , \new_[92811]_ , \new_[92814]_ ,
    \new_[92815]_ , \new_[92818]_ , \new_[92821]_ , \new_[92822]_ ,
    \new_[92823]_ , \new_[92826]_ , \new_[92829]_ , \new_[92830]_ ,
    \new_[92833]_ , \new_[92836]_ , \new_[92837]_ , \new_[92838]_ ,
    \new_[92841]_ , \new_[92844]_ , \new_[92845]_ , \new_[92848]_ ,
    \new_[92851]_ , \new_[92852]_ , \new_[92853]_ , \new_[92856]_ ,
    \new_[92859]_ , \new_[92860]_ , \new_[92863]_ , \new_[92866]_ ,
    \new_[92867]_ , \new_[92868]_ , \new_[92871]_ , \new_[92874]_ ,
    \new_[92875]_ , \new_[92878]_ , \new_[92881]_ , \new_[92882]_ ,
    \new_[92883]_ , \new_[92886]_ , \new_[92889]_ , \new_[92890]_ ,
    \new_[92893]_ , \new_[92896]_ , \new_[92897]_ , \new_[92898]_ ,
    \new_[92901]_ , \new_[92904]_ , \new_[92905]_ , \new_[92908]_ ,
    \new_[92911]_ , \new_[92912]_ , \new_[92913]_ , \new_[92916]_ ,
    \new_[92919]_ , \new_[92920]_ , \new_[92923]_ , \new_[92926]_ ,
    \new_[92927]_ , \new_[92928]_ , \new_[92931]_ , \new_[92934]_ ,
    \new_[92935]_ , \new_[92938]_ , \new_[92941]_ , \new_[92942]_ ,
    \new_[92943]_ , \new_[92946]_ , \new_[92949]_ , \new_[92950]_ ,
    \new_[92953]_ , \new_[92956]_ , \new_[92957]_ , \new_[92958]_ ,
    \new_[92961]_ , \new_[92964]_ , \new_[92965]_ , \new_[92968]_ ,
    \new_[92971]_ , \new_[92972]_ , \new_[92973]_ , \new_[92976]_ ,
    \new_[92979]_ , \new_[92980]_ , \new_[92983]_ , \new_[92986]_ ,
    \new_[92987]_ , \new_[92988]_ , \new_[92991]_ , \new_[92994]_ ,
    \new_[92995]_ , \new_[92998]_ , \new_[93001]_ , \new_[93002]_ ,
    \new_[93003]_ , \new_[93006]_ , \new_[93009]_ , \new_[93010]_ ,
    \new_[93013]_ , \new_[93016]_ , \new_[93017]_ , \new_[93018]_ ,
    \new_[93021]_ , \new_[93024]_ , \new_[93025]_ , \new_[93028]_ ,
    \new_[93031]_ , \new_[93032]_ , \new_[93033]_ , \new_[93036]_ ,
    \new_[93039]_ , \new_[93040]_ , \new_[93043]_ , \new_[93046]_ ,
    \new_[93047]_ , \new_[93048]_ , \new_[93051]_ , \new_[93054]_ ,
    \new_[93055]_ , \new_[93058]_ , \new_[93061]_ , \new_[93062]_ ,
    \new_[93063]_ , \new_[93066]_ , \new_[93069]_ , \new_[93070]_ ,
    \new_[93073]_ , \new_[93076]_ , \new_[93077]_ , \new_[93078]_ ,
    \new_[93081]_ , \new_[93084]_ , \new_[93085]_ , \new_[93088]_ ,
    \new_[93091]_ , \new_[93092]_ , \new_[93093]_ , \new_[93096]_ ,
    \new_[93099]_ , \new_[93100]_ , \new_[93103]_ , \new_[93106]_ ,
    \new_[93107]_ , \new_[93108]_ , \new_[93111]_ , \new_[93114]_ ,
    \new_[93115]_ , \new_[93118]_ , \new_[93121]_ , \new_[93122]_ ,
    \new_[93123]_ , \new_[93126]_ , \new_[93129]_ , \new_[93130]_ ,
    \new_[93133]_ , \new_[93136]_ , \new_[93137]_ , \new_[93138]_ ,
    \new_[93141]_ , \new_[93144]_ , \new_[93145]_ , \new_[93148]_ ,
    \new_[93151]_ , \new_[93152]_ , \new_[93153]_ , \new_[93156]_ ,
    \new_[93159]_ , \new_[93160]_ , \new_[93163]_ , \new_[93166]_ ,
    \new_[93167]_ , \new_[93168]_ , \new_[93171]_ , \new_[93174]_ ,
    \new_[93175]_ , \new_[93178]_ , \new_[93181]_ , \new_[93182]_ ,
    \new_[93183]_ , \new_[93186]_ , \new_[93189]_ , \new_[93190]_ ,
    \new_[93193]_ , \new_[93196]_ , \new_[93197]_ , \new_[93198]_ ,
    \new_[93201]_ , \new_[93204]_ , \new_[93205]_ , \new_[93208]_ ,
    \new_[93211]_ , \new_[93212]_ , \new_[93213]_ , \new_[93216]_ ,
    \new_[93219]_ , \new_[93220]_ , \new_[93223]_ , \new_[93226]_ ,
    \new_[93227]_ , \new_[93228]_ , \new_[93231]_ , \new_[93234]_ ,
    \new_[93235]_ , \new_[93238]_ , \new_[93241]_ , \new_[93242]_ ,
    \new_[93243]_ , \new_[93246]_ , \new_[93249]_ , \new_[93250]_ ,
    \new_[93253]_ , \new_[93256]_ , \new_[93257]_ , \new_[93258]_ ,
    \new_[93261]_ , \new_[93264]_ , \new_[93265]_ , \new_[93268]_ ,
    \new_[93271]_ , \new_[93272]_ , \new_[93273]_ , \new_[93276]_ ,
    \new_[93279]_ , \new_[93280]_ , \new_[93283]_ , \new_[93286]_ ,
    \new_[93287]_ , \new_[93288]_ , \new_[93291]_ , \new_[93294]_ ,
    \new_[93295]_ , \new_[93298]_ , \new_[93301]_ , \new_[93302]_ ,
    \new_[93303]_ , \new_[93306]_ , \new_[93309]_ , \new_[93310]_ ,
    \new_[93313]_ , \new_[93316]_ , \new_[93317]_ , \new_[93318]_ ,
    \new_[93321]_ , \new_[93324]_ , \new_[93325]_ , \new_[93328]_ ,
    \new_[93331]_ , \new_[93332]_ , \new_[93333]_ , \new_[93336]_ ,
    \new_[93339]_ , \new_[93340]_ , \new_[93343]_ , \new_[93346]_ ,
    \new_[93347]_ , \new_[93348]_ , \new_[93351]_ , \new_[93354]_ ,
    \new_[93355]_ , \new_[93358]_ , \new_[93361]_ , \new_[93362]_ ,
    \new_[93363]_ , \new_[93366]_ , \new_[93369]_ , \new_[93370]_ ,
    \new_[93373]_ , \new_[93376]_ , \new_[93377]_ , \new_[93378]_ ,
    \new_[93381]_ , \new_[93384]_ , \new_[93385]_ , \new_[93388]_ ,
    \new_[93391]_ , \new_[93392]_ , \new_[93393]_ , \new_[93396]_ ,
    \new_[93399]_ , \new_[93400]_ , \new_[93403]_ , \new_[93406]_ ,
    \new_[93407]_ , \new_[93408]_ , \new_[93411]_ , \new_[93414]_ ,
    \new_[93415]_ , \new_[93418]_ , \new_[93421]_ , \new_[93422]_ ,
    \new_[93423]_ , \new_[93426]_ , \new_[93429]_ , \new_[93430]_ ,
    \new_[93433]_ , \new_[93436]_ , \new_[93437]_ , \new_[93438]_ ,
    \new_[93441]_ , \new_[93444]_ , \new_[93445]_ , \new_[93448]_ ,
    \new_[93451]_ , \new_[93452]_ , \new_[93453]_ , \new_[93456]_ ,
    \new_[93459]_ , \new_[93460]_ , \new_[93463]_ , \new_[93466]_ ,
    \new_[93467]_ , \new_[93468]_ , \new_[93471]_ , \new_[93474]_ ,
    \new_[93475]_ , \new_[93478]_ , \new_[93481]_ , \new_[93482]_ ,
    \new_[93483]_ , \new_[93486]_ , \new_[93489]_ , \new_[93490]_ ,
    \new_[93493]_ , \new_[93496]_ , \new_[93497]_ , \new_[93498]_ ,
    \new_[93501]_ , \new_[93504]_ , \new_[93505]_ , \new_[93508]_ ,
    \new_[93511]_ , \new_[93512]_ , \new_[93513]_ , \new_[93516]_ ,
    \new_[93519]_ , \new_[93520]_ , \new_[93523]_ , \new_[93526]_ ,
    \new_[93527]_ , \new_[93528]_ , \new_[93531]_ , \new_[93534]_ ,
    \new_[93535]_ , \new_[93538]_ , \new_[93541]_ , \new_[93542]_ ,
    \new_[93543]_ , \new_[93546]_ , \new_[93549]_ , \new_[93550]_ ,
    \new_[93553]_ , \new_[93556]_ , \new_[93557]_ , \new_[93558]_ ,
    \new_[93561]_ , \new_[93564]_ , \new_[93565]_ , \new_[93568]_ ,
    \new_[93571]_ , \new_[93572]_ , \new_[93573]_ , \new_[93576]_ ,
    \new_[93579]_ , \new_[93580]_ , \new_[93583]_ , \new_[93586]_ ,
    \new_[93587]_ , \new_[93588]_ , \new_[93591]_ , \new_[93594]_ ,
    \new_[93595]_ , \new_[93598]_ , \new_[93601]_ , \new_[93602]_ ,
    \new_[93603]_ , \new_[93606]_ , \new_[93609]_ , \new_[93610]_ ,
    \new_[93613]_ , \new_[93616]_ , \new_[93617]_ , \new_[93618]_ ,
    \new_[93621]_ , \new_[93624]_ , \new_[93625]_ , \new_[93628]_ ,
    \new_[93631]_ , \new_[93632]_ , \new_[93633]_ , \new_[93636]_ ,
    \new_[93639]_ , \new_[93640]_ , \new_[93643]_ , \new_[93646]_ ,
    \new_[93647]_ , \new_[93648]_ , \new_[93651]_ , \new_[93654]_ ,
    \new_[93655]_ , \new_[93658]_ , \new_[93661]_ , \new_[93662]_ ,
    \new_[93663]_ , \new_[93666]_ , \new_[93669]_ , \new_[93670]_ ,
    \new_[93673]_ , \new_[93676]_ , \new_[93677]_ , \new_[93678]_ ,
    \new_[93681]_ , \new_[93684]_ , \new_[93685]_ , \new_[93688]_ ,
    \new_[93691]_ , \new_[93692]_ , \new_[93693]_ , \new_[93696]_ ,
    \new_[93699]_ , \new_[93700]_ , \new_[93703]_ , \new_[93706]_ ,
    \new_[93707]_ , \new_[93708]_ , \new_[93711]_ , \new_[93714]_ ,
    \new_[93715]_ , \new_[93718]_ , \new_[93721]_ , \new_[93722]_ ,
    \new_[93723]_ , \new_[93726]_ , \new_[93729]_ , \new_[93730]_ ,
    \new_[93733]_ , \new_[93736]_ , \new_[93737]_ , \new_[93738]_ ,
    \new_[93741]_ , \new_[93744]_ , \new_[93745]_ , \new_[93748]_ ,
    \new_[93751]_ , \new_[93752]_ , \new_[93753]_ , \new_[93756]_ ,
    \new_[93759]_ , \new_[93760]_ , \new_[93763]_ , \new_[93766]_ ,
    \new_[93767]_ , \new_[93768]_ , \new_[93771]_ , \new_[93774]_ ,
    \new_[93775]_ , \new_[93778]_ , \new_[93781]_ , \new_[93782]_ ,
    \new_[93783]_ , \new_[93786]_ , \new_[93789]_ , \new_[93790]_ ,
    \new_[93793]_ , \new_[93796]_ , \new_[93797]_ , \new_[93798]_ ,
    \new_[93801]_ , \new_[93804]_ , \new_[93805]_ , \new_[93808]_ ,
    \new_[93811]_ , \new_[93812]_ , \new_[93813]_ , \new_[93816]_ ,
    \new_[93819]_ , \new_[93820]_ , \new_[93823]_ , \new_[93826]_ ,
    \new_[93827]_ , \new_[93828]_ , \new_[93831]_ , \new_[93834]_ ,
    \new_[93835]_ , \new_[93838]_ , \new_[93841]_ , \new_[93842]_ ,
    \new_[93843]_ , \new_[93846]_ , \new_[93849]_ , \new_[93850]_ ,
    \new_[93853]_ , \new_[93856]_ , \new_[93857]_ , \new_[93858]_ ,
    \new_[93861]_ , \new_[93864]_ , \new_[93865]_ , \new_[93868]_ ,
    \new_[93871]_ , \new_[93872]_ , \new_[93873]_ , \new_[93876]_ ,
    \new_[93879]_ , \new_[93880]_ , \new_[93883]_ , \new_[93886]_ ,
    \new_[93887]_ , \new_[93888]_ , \new_[93891]_ , \new_[93894]_ ,
    \new_[93895]_ , \new_[93898]_ , \new_[93901]_ , \new_[93902]_ ,
    \new_[93903]_ , \new_[93906]_ , \new_[93909]_ , \new_[93910]_ ,
    \new_[93913]_ , \new_[93916]_ , \new_[93917]_ , \new_[93918]_ ,
    \new_[93921]_ , \new_[93924]_ , \new_[93925]_ , \new_[93928]_ ,
    \new_[93931]_ , \new_[93932]_ , \new_[93933]_ , \new_[93936]_ ,
    \new_[93939]_ , \new_[93940]_ , \new_[93943]_ , \new_[93946]_ ,
    \new_[93947]_ , \new_[93948]_ , \new_[93951]_ , \new_[93954]_ ,
    \new_[93955]_ , \new_[93958]_ , \new_[93961]_ , \new_[93962]_ ,
    \new_[93963]_ , \new_[93966]_ , \new_[93969]_ , \new_[93970]_ ,
    \new_[93973]_ , \new_[93976]_ , \new_[93977]_ , \new_[93978]_ ,
    \new_[93981]_ , \new_[93984]_ , \new_[93985]_ , \new_[93988]_ ,
    \new_[93991]_ , \new_[93992]_ , \new_[93993]_ , \new_[93996]_ ,
    \new_[93999]_ , \new_[94000]_ , \new_[94003]_ , \new_[94006]_ ,
    \new_[94007]_ , \new_[94008]_ , \new_[94011]_ , \new_[94014]_ ,
    \new_[94015]_ , \new_[94018]_ , \new_[94021]_ , \new_[94022]_ ,
    \new_[94023]_ , \new_[94026]_ , \new_[94029]_ , \new_[94030]_ ,
    \new_[94033]_ , \new_[94036]_ , \new_[94037]_ , \new_[94038]_ ,
    \new_[94041]_ , \new_[94044]_ , \new_[94045]_ , \new_[94048]_ ,
    \new_[94051]_ , \new_[94052]_ , \new_[94053]_ , \new_[94056]_ ,
    \new_[94059]_ , \new_[94060]_ , \new_[94063]_ , \new_[94066]_ ,
    \new_[94067]_ , \new_[94068]_ , \new_[94071]_ , \new_[94074]_ ,
    \new_[94075]_ , \new_[94078]_ , \new_[94081]_ , \new_[94082]_ ,
    \new_[94083]_ , \new_[94086]_ , \new_[94089]_ , \new_[94090]_ ,
    \new_[94093]_ , \new_[94096]_ , \new_[94097]_ , \new_[94098]_ ,
    \new_[94101]_ , \new_[94104]_ , \new_[94105]_ , \new_[94108]_ ,
    \new_[94111]_ , \new_[94112]_ , \new_[94113]_ , \new_[94116]_ ,
    \new_[94119]_ , \new_[94120]_ , \new_[94123]_ , \new_[94126]_ ,
    \new_[94127]_ , \new_[94128]_ , \new_[94131]_ , \new_[94134]_ ,
    \new_[94135]_ , \new_[94138]_ , \new_[94141]_ , \new_[94142]_ ,
    \new_[94143]_ , \new_[94146]_ , \new_[94149]_ , \new_[94150]_ ,
    \new_[94153]_ , \new_[94156]_ , \new_[94157]_ , \new_[94158]_ ,
    \new_[94161]_ , \new_[94164]_ , \new_[94165]_ , \new_[94168]_ ,
    \new_[94171]_ , \new_[94172]_ , \new_[94173]_ , \new_[94176]_ ,
    \new_[94179]_ , \new_[94180]_ , \new_[94183]_ , \new_[94186]_ ,
    \new_[94187]_ , \new_[94188]_ , \new_[94191]_ , \new_[94194]_ ,
    \new_[94195]_ , \new_[94198]_ , \new_[94201]_ , \new_[94202]_ ,
    \new_[94203]_ , \new_[94206]_ , \new_[94209]_ , \new_[94210]_ ,
    \new_[94213]_ , \new_[94216]_ , \new_[94217]_ , \new_[94218]_ ,
    \new_[94221]_ , \new_[94224]_ , \new_[94225]_ , \new_[94228]_ ,
    \new_[94231]_ , \new_[94232]_ , \new_[94233]_ , \new_[94236]_ ,
    \new_[94239]_ , \new_[94240]_ , \new_[94243]_ , \new_[94246]_ ,
    \new_[94247]_ , \new_[94248]_ , \new_[94251]_ , \new_[94254]_ ,
    \new_[94255]_ , \new_[94258]_ , \new_[94261]_ , \new_[94262]_ ,
    \new_[94263]_ , \new_[94266]_ , \new_[94269]_ , \new_[94270]_ ,
    \new_[94273]_ , \new_[94276]_ , \new_[94277]_ , \new_[94278]_ ,
    \new_[94281]_ , \new_[94284]_ , \new_[94285]_ , \new_[94288]_ ,
    \new_[94291]_ , \new_[94292]_ , \new_[94293]_ , \new_[94296]_ ,
    \new_[94299]_ , \new_[94300]_ , \new_[94303]_ , \new_[94306]_ ,
    \new_[94307]_ , \new_[94308]_ , \new_[94311]_ , \new_[94314]_ ,
    \new_[94315]_ , \new_[94318]_ , \new_[94321]_ , \new_[94322]_ ,
    \new_[94323]_ , \new_[94326]_ , \new_[94329]_ , \new_[94330]_ ,
    \new_[94333]_ , \new_[94336]_ , \new_[94337]_ , \new_[94338]_ ,
    \new_[94341]_ , \new_[94344]_ , \new_[94345]_ , \new_[94348]_ ,
    \new_[94351]_ , \new_[94352]_ , \new_[94353]_ , \new_[94356]_ ,
    \new_[94359]_ , \new_[94360]_ , \new_[94363]_ , \new_[94366]_ ,
    \new_[94367]_ , \new_[94368]_ , \new_[94371]_ , \new_[94374]_ ,
    \new_[94375]_ , \new_[94378]_ , \new_[94381]_ , \new_[94382]_ ,
    \new_[94383]_ , \new_[94386]_ , \new_[94389]_ , \new_[94390]_ ,
    \new_[94393]_ , \new_[94396]_ , \new_[94397]_ , \new_[94398]_ ,
    \new_[94401]_ , \new_[94404]_ , \new_[94405]_ , \new_[94408]_ ,
    \new_[94411]_ , \new_[94412]_ , \new_[94413]_ , \new_[94416]_ ,
    \new_[94419]_ , \new_[94420]_ , \new_[94423]_ , \new_[94426]_ ,
    \new_[94427]_ , \new_[94428]_ , \new_[94431]_ , \new_[94434]_ ,
    \new_[94435]_ , \new_[94438]_ , \new_[94441]_ , \new_[94442]_ ,
    \new_[94443]_ , \new_[94446]_ , \new_[94449]_ , \new_[94450]_ ,
    \new_[94453]_ , \new_[94456]_ , \new_[94457]_ , \new_[94458]_ ,
    \new_[94461]_ , \new_[94464]_ , \new_[94465]_ , \new_[94468]_ ,
    \new_[94471]_ , \new_[94472]_ , \new_[94473]_ , \new_[94476]_ ,
    \new_[94479]_ , \new_[94480]_ , \new_[94483]_ , \new_[94486]_ ,
    \new_[94487]_ , \new_[94488]_ , \new_[94491]_ , \new_[94494]_ ,
    \new_[94495]_ , \new_[94498]_ , \new_[94501]_ , \new_[94502]_ ,
    \new_[94503]_ , \new_[94506]_ , \new_[94509]_ , \new_[94510]_ ,
    \new_[94513]_ , \new_[94516]_ , \new_[94517]_ , \new_[94518]_ ,
    \new_[94521]_ , \new_[94524]_ , \new_[94525]_ , \new_[94528]_ ,
    \new_[94531]_ , \new_[94532]_ , \new_[94533]_ , \new_[94536]_ ,
    \new_[94539]_ , \new_[94540]_ , \new_[94543]_ , \new_[94546]_ ,
    \new_[94547]_ , \new_[94548]_ , \new_[94551]_ , \new_[94554]_ ,
    \new_[94555]_ , \new_[94558]_ , \new_[94561]_ , \new_[94562]_ ,
    \new_[94563]_ , \new_[94566]_ , \new_[94569]_ , \new_[94570]_ ,
    \new_[94573]_ , \new_[94576]_ , \new_[94577]_ , \new_[94578]_ ,
    \new_[94581]_ , \new_[94584]_ , \new_[94585]_ , \new_[94588]_ ,
    \new_[94591]_ , \new_[94592]_ , \new_[94593]_ , \new_[94596]_ ,
    \new_[94599]_ , \new_[94600]_ , \new_[94603]_ , \new_[94606]_ ,
    \new_[94607]_ , \new_[94608]_ , \new_[94611]_ , \new_[94614]_ ,
    \new_[94615]_ , \new_[94618]_ , \new_[94621]_ , \new_[94622]_ ,
    \new_[94623]_ , \new_[94626]_ , \new_[94629]_ , \new_[94630]_ ,
    \new_[94633]_ , \new_[94636]_ , \new_[94637]_ , \new_[94638]_ ,
    \new_[94641]_ , \new_[94644]_ , \new_[94645]_ , \new_[94648]_ ,
    \new_[94651]_ , \new_[94652]_ , \new_[94653]_ , \new_[94656]_ ,
    \new_[94659]_ , \new_[94660]_ , \new_[94663]_ , \new_[94666]_ ,
    \new_[94667]_ , \new_[94668]_ , \new_[94671]_ , \new_[94674]_ ,
    \new_[94675]_ , \new_[94678]_ , \new_[94681]_ , \new_[94682]_ ,
    \new_[94683]_ , \new_[94686]_ , \new_[94689]_ , \new_[94690]_ ,
    \new_[94693]_ , \new_[94696]_ , \new_[94697]_ , \new_[94698]_ ,
    \new_[94701]_ , \new_[94704]_ , \new_[94705]_ , \new_[94708]_ ,
    \new_[94711]_ , \new_[94712]_ , \new_[94713]_ , \new_[94716]_ ,
    \new_[94719]_ , \new_[94720]_ , \new_[94723]_ , \new_[94726]_ ,
    \new_[94727]_ , \new_[94728]_ , \new_[94731]_ , \new_[94734]_ ,
    \new_[94735]_ , \new_[94738]_ , \new_[94741]_ , \new_[94742]_ ,
    \new_[94743]_ , \new_[94746]_ , \new_[94749]_ , \new_[94750]_ ,
    \new_[94753]_ , \new_[94756]_ , \new_[94757]_ , \new_[94758]_ ,
    \new_[94761]_ , \new_[94764]_ , \new_[94765]_ , \new_[94768]_ ,
    \new_[94771]_ , \new_[94772]_ , \new_[94773]_ , \new_[94776]_ ,
    \new_[94779]_ , \new_[94780]_ , \new_[94783]_ , \new_[94786]_ ,
    \new_[94787]_ , \new_[94788]_ , \new_[94791]_ , \new_[94794]_ ,
    \new_[94795]_ , \new_[94798]_ , \new_[94801]_ , \new_[94802]_ ,
    \new_[94803]_ , \new_[94806]_ , \new_[94809]_ , \new_[94810]_ ,
    \new_[94813]_ , \new_[94816]_ , \new_[94817]_ , \new_[94818]_ ,
    \new_[94821]_ , \new_[94824]_ , \new_[94825]_ , \new_[94828]_ ,
    \new_[94831]_ , \new_[94832]_ , \new_[94833]_ , \new_[94836]_ ,
    \new_[94839]_ , \new_[94840]_ , \new_[94843]_ , \new_[94846]_ ,
    \new_[94847]_ , \new_[94848]_ , \new_[94851]_ , \new_[94854]_ ,
    \new_[94855]_ , \new_[94858]_ , \new_[94861]_ , \new_[94862]_ ,
    \new_[94863]_ , \new_[94866]_ , \new_[94869]_ , \new_[94870]_ ,
    \new_[94873]_ , \new_[94876]_ , \new_[94877]_ , \new_[94878]_ ,
    \new_[94881]_ , \new_[94884]_ , \new_[94885]_ , \new_[94888]_ ,
    \new_[94891]_ , \new_[94892]_ , \new_[94893]_ , \new_[94896]_ ,
    \new_[94899]_ , \new_[94900]_ , \new_[94903]_ , \new_[94906]_ ,
    \new_[94907]_ , \new_[94908]_ , \new_[94911]_ , \new_[94914]_ ,
    \new_[94915]_ , \new_[94918]_ , \new_[94921]_ , \new_[94922]_ ,
    \new_[94923]_ , \new_[94926]_ , \new_[94929]_ , \new_[94930]_ ,
    \new_[94933]_ , \new_[94936]_ , \new_[94937]_ , \new_[94938]_ ,
    \new_[94941]_ , \new_[94944]_ , \new_[94945]_ , \new_[94948]_ ,
    \new_[94951]_ , \new_[94952]_ , \new_[94953]_ , \new_[94956]_ ,
    \new_[94959]_ , \new_[94960]_ , \new_[94963]_ , \new_[94966]_ ,
    \new_[94967]_ , \new_[94968]_ , \new_[94971]_ , \new_[94974]_ ,
    \new_[94975]_ , \new_[94978]_ , \new_[94981]_ , \new_[94982]_ ,
    \new_[94983]_ , \new_[94986]_ , \new_[94989]_ , \new_[94990]_ ,
    \new_[94993]_ , \new_[94996]_ , \new_[94997]_ , \new_[94998]_ ,
    \new_[95001]_ , \new_[95004]_ , \new_[95005]_ , \new_[95008]_ ,
    \new_[95011]_ , \new_[95012]_ , \new_[95013]_ , \new_[95016]_ ,
    \new_[95019]_ , \new_[95020]_ , \new_[95023]_ , \new_[95026]_ ,
    \new_[95027]_ , \new_[95028]_ , \new_[95031]_ , \new_[95034]_ ,
    \new_[95035]_ , \new_[95038]_ , \new_[95041]_ , \new_[95042]_ ,
    \new_[95043]_ , \new_[95046]_ , \new_[95049]_ , \new_[95050]_ ,
    \new_[95053]_ , \new_[95056]_ , \new_[95057]_ , \new_[95058]_ ,
    \new_[95061]_ , \new_[95064]_ , \new_[95065]_ , \new_[95068]_ ,
    \new_[95071]_ , \new_[95072]_ , \new_[95073]_ , \new_[95076]_ ,
    \new_[95079]_ , \new_[95080]_ , \new_[95083]_ , \new_[95086]_ ,
    \new_[95087]_ , \new_[95088]_ , \new_[95091]_ , \new_[95094]_ ,
    \new_[95095]_ , \new_[95098]_ , \new_[95101]_ , \new_[95102]_ ,
    \new_[95103]_ , \new_[95106]_ , \new_[95109]_ , \new_[95110]_ ,
    \new_[95113]_ , \new_[95116]_ , \new_[95117]_ , \new_[95118]_ ,
    \new_[95121]_ , \new_[95124]_ , \new_[95125]_ , \new_[95128]_ ,
    \new_[95131]_ , \new_[95132]_ , \new_[95133]_ , \new_[95136]_ ,
    \new_[95139]_ , \new_[95140]_ , \new_[95143]_ , \new_[95146]_ ,
    \new_[95147]_ , \new_[95148]_ , \new_[95151]_ , \new_[95154]_ ,
    \new_[95155]_ , \new_[95158]_ , \new_[95161]_ , \new_[95162]_ ,
    \new_[95163]_ , \new_[95166]_ , \new_[95169]_ , \new_[95170]_ ,
    \new_[95173]_ , \new_[95176]_ , \new_[95177]_ , \new_[95178]_ ,
    \new_[95181]_ , \new_[95184]_ , \new_[95185]_ , \new_[95188]_ ,
    \new_[95191]_ , \new_[95192]_ , \new_[95193]_ , \new_[95196]_ ,
    \new_[95199]_ , \new_[95200]_ , \new_[95203]_ , \new_[95206]_ ,
    \new_[95207]_ , \new_[95208]_ , \new_[95211]_ , \new_[95214]_ ,
    \new_[95215]_ , \new_[95218]_ , \new_[95221]_ , \new_[95222]_ ,
    \new_[95223]_ , \new_[95226]_ , \new_[95229]_ , \new_[95230]_ ,
    \new_[95233]_ , \new_[95236]_ , \new_[95237]_ , \new_[95238]_ ,
    \new_[95241]_ , \new_[95244]_ , \new_[95245]_ , \new_[95248]_ ,
    \new_[95251]_ , \new_[95252]_ , \new_[95253]_ , \new_[95256]_ ,
    \new_[95259]_ , \new_[95260]_ , \new_[95263]_ , \new_[95266]_ ,
    \new_[95267]_ , \new_[95268]_ , \new_[95271]_ , \new_[95274]_ ,
    \new_[95275]_ , \new_[95278]_ , \new_[95281]_ , \new_[95282]_ ,
    \new_[95283]_ , \new_[95286]_ , \new_[95289]_ , \new_[95290]_ ,
    \new_[95293]_ , \new_[95296]_ , \new_[95297]_ , \new_[95298]_ ,
    \new_[95301]_ , \new_[95304]_ , \new_[95305]_ , \new_[95308]_ ,
    \new_[95311]_ , \new_[95312]_ , \new_[95313]_ , \new_[95316]_ ,
    \new_[95319]_ , \new_[95320]_ , \new_[95323]_ , \new_[95326]_ ,
    \new_[95327]_ , \new_[95328]_ , \new_[95331]_ , \new_[95334]_ ,
    \new_[95335]_ , \new_[95338]_ , \new_[95341]_ , \new_[95342]_ ,
    \new_[95343]_ , \new_[95346]_ , \new_[95349]_ , \new_[95350]_ ,
    \new_[95353]_ , \new_[95356]_ , \new_[95357]_ , \new_[95358]_ ,
    \new_[95361]_ , \new_[95364]_ , \new_[95365]_ , \new_[95368]_ ,
    \new_[95371]_ , \new_[95372]_ , \new_[95373]_ , \new_[95376]_ ,
    \new_[95379]_ , \new_[95380]_ , \new_[95383]_ , \new_[95386]_ ,
    \new_[95387]_ , \new_[95388]_ , \new_[95391]_ , \new_[95394]_ ,
    \new_[95395]_ , \new_[95398]_ , \new_[95401]_ , \new_[95402]_ ,
    \new_[95403]_ , \new_[95406]_ , \new_[95409]_ , \new_[95410]_ ,
    \new_[95413]_ , \new_[95416]_ , \new_[95417]_ , \new_[95418]_ ,
    \new_[95421]_ , \new_[95424]_ , \new_[95425]_ , \new_[95428]_ ,
    \new_[95431]_ , \new_[95432]_ , \new_[95433]_ , \new_[95436]_ ,
    \new_[95439]_ , \new_[95440]_ , \new_[95443]_ , \new_[95446]_ ,
    \new_[95447]_ , \new_[95448]_ , \new_[95451]_ , \new_[95454]_ ,
    \new_[95455]_ , \new_[95458]_ , \new_[95461]_ , \new_[95462]_ ,
    \new_[95463]_ , \new_[95466]_ , \new_[95469]_ , \new_[95470]_ ,
    \new_[95473]_ , \new_[95476]_ , \new_[95477]_ , \new_[95478]_ ,
    \new_[95481]_ , \new_[95484]_ , \new_[95485]_ , \new_[95488]_ ,
    \new_[95491]_ , \new_[95492]_ , \new_[95493]_ , \new_[95496]_ ,
    \new_[95499]_ , \new_[95500]_ , \new_[95503]_ , \new_[95506]_ ,
    \new_[95507]_ , \new_[95508]_ , \new_[95511]_ , \new_[95514]_ ,
    \new_[95515]_ , \new_[95518]_ , \new_[95521]_ , \new_[95522]_ ,
    \new_[95523]_ , \new_[95526]_ , \new_[95529]_ , \new_[95530]_ ,
    \new_[95533]_ , \new_[95536]_ , \new_[95537]_ , \new_[95538]_ ,
    \new_[95541]_ , \new_[95544]_ , \new_[95545]_ , \new_[95548]_ ,
    \new_[95551]_ , \new_[95552]_ , \new_[95553]_ , \new_[95556]_ ,
    \new_[95559]_ , \new_[95560]_ , \new_[95563]_ , \new_[95566]_ ,
    \new_[95567]_ , \new_[95568]_ , \new_[95571]_ , \new_[95574]_ ,
    \new_[95575]_ , \new_[95578]_ , \new_[95581]_ , \new_[95582]_ ,
    \new_[95583]_ , \new_[95586]_ , \new_[95589]_ , \new_[95590]_ ,
    \new_[95593]_ , \new_[95596]_ , \new_[95597]_ , \new_[95598]_ ,
    \new_[95601]_ , \new_[95604]_ , \new_[95605]_ , \new_[95608]_ ,
    \new_[95611]_ , \new_[95612]_ , \new_[95613]_ , \new_[95616]_ ,
    \new_[95619]_ , \new_[95620]_ , \new_[95623]_ , \new_[95626]_ ,
    \new_[95627]_ , \new_[95628]_ , \new_[95631]_ , \new_[95634]_ ,
    \new_[95635]_ , \new_[95638]_ , \new_[95641]_ , \new_[95642]_ ,
    \new_[95643]_ , \new_[95646]_ , \new_[95649]_ , \new_[95650]_ ,
    \new_[95653]_ , \new_[95656]_ , \new_[95657]_ , \new_[95658]_ ,
    \new_[95661]_ , \new_[95664]_ , \new_[95665]_ , \new_[95668]_ ,
    \new_[95671]_ , \new_[95672]_ , \new_[95673]_ , \new_[95676]_ ,
    \new_[95679]_ , \new_[95680]_ , \new_[95683]_ , \new_[95686]_ ,
    \new_[95687]_ , \new_[95688]_ , \new_[95691]_ , \new_[95694]_ ,
    \new_[95695]_ , \new_[95698]_ , \new_[95701]_ , \new_[95702]_ ,
    \new_[95703]_ , \new_[95706]_ , \new_[95709]_ , \new_[95710]_ ,
    \new_[95713]_ , \new_[95716]_ , \new_[95717]_ , \new_[95718]_ ,
    \new_[95721]_ , \new_[95724]_ , \new_[95725]_ , \new_[95728]_ ,
    \new_[95731]_ , \new_[95732]_ , \new_[95733]_ , \new_[95736]_ ,
    \new_[95739]_ , \new_[95740]_ , \new_[95743]_ , \new_[95746]_ ,
    \new_[95747]_ , \new_[95748]_ , \new_[95751]_ , \new_[95754]_ ,
    \new_[95755]_ , \new_[95758]_ , \new_[95761]_ , \new_[95762]_ ,
    \new_[95763]_ , \new_[95766]_ , \new_[95769]_ , \new_[95770]_ ,
    \new_[95773]_ , \new_[95776]_ , \new_[95777]_ , \new_[95778]_ ,
    \new_[95781]_ , \new_[95784]_ , \new_[95785]_ , \new_[95788]_ ,
    \new_[95791]_ , \new_[95792]_ , \new_[95793]_ , \new_[95796]_ ,
    \new_[95799]_ , \new_[95800]_ , \new_[95803]_ , \new_[95806]_ ,
    \new_[95807]_ , \new_[95808]_ , \new_[95811]_ , \new_[95814]_ ,
    \new_[95815]_ , \new_[95818]_ , \new_[95821]_ , \new_[95822]_ ,
    \new_[95823]_ , \new_[95826]_ , \new_[95829]_ , \new_[95830]_ ,
    \new_[95833]_ , \new_[95836]_ , \new_[95837]_ , \new_[95838]_ ,
    \new_[95841]_ , \new_[95844]_ , \new_[95845]_ , \new_[95848]_ ,
    \new_[95851]_ , \new_[95852]_ , \new_[95853]_ , \new_[95856]_ ,
    \new_[95859]_ , \new_[95860]_ , \new_[95863]_ , \new_[95866]_ ,
    \new_[95867]_ , \new_[95868]_ , \new_[95871]_ , \new_[95874]_ ,
    \new_[95875]_ , \new_[95878]_ , \new_[95881]_ , \new_[95882]_ ,
    \new_[95883]_ , \new_[95886]_ , \new_[95889]_ , \new_[95890]_ ,
    \new_[95893]_ , \new_[95896]_ , \new_[95897]_ , \new_[95898]_ ,
    \new_[95901]_ , \new_[95904]_ , \new_[95905]_ , \new_[95908]_ ,
    \new_[95911]_ , \new_[95912]_ , \new_[95913]_ , \new_[95916]_ ,
    \new_[95919]_ , \new_[95920]_ , \new_[95923]_ , \new_[95926]_ ,
    \new_[95927]_ , \new_[95928]_ , \new_[95931]_ , \new_[95934]_ ,
    \new_[95935]_ , \new_[95938]_ , \new_[95941]_ , \new_[95942]_ ,
    \new_[95943]_ , \new_[95946]_ , \new_[95949]_ , \new_[95950]_ ,
    \new_[95953]_ , \new_[95956]_ , \new_[95957]_ , \new_[95958]_ ,
    \new_[95961]_ , \new_[95964]_ , \new_[95965]_ , \new_[95968]_ ,
    \new_[95971]_ , \new_[95972]_ , \new_[95973]_ , \new_[95976]_ ,
    \new_[95979]_ , \new_[95980]_ , \new_[95983]_ , \new_[95986]_ ,
    \new_[95987]_ , \new_[95988]_ , \new_[95991]_ , \new_[95994]_ ,
    \new_[95995]_ , \new_[95998]_ , \new_[96001]_ , \new_[96002]_ ,
    \new_[96003]_ , \new_[96006]_ , \new_[96009]_ , \new_[96010]_ ,
    \new_[96013]_ , \new_[96016]_ , \new_[96017]_ , \new_[96018]_ ,
    \new_[96021]_ , \new_[96024]_ , \new_[96025]_ , \new_[96028]_ ,
    \new_[96031]_ , \new_[96032]_ , \new_[96033]_ , \new_[96036]_ ,
    \new_[96039]_ , \new_[96040]_ , \new_[96043]_ , \new_[96046]_ ,
    \new_[96047]_ , \new_[96048]_ , \new_[96051]_ , \new_[96054]_ ,
    \new_[96055]_ , \new_[96058]_ , \new_[96061]_ , \new_[96062]_ ,
    \new_[96063]_ , \new_[96066]_ , \new_[96069]_ , \new_[96070]_ ,
    \new_[96073]_ , \new_[96076]_ , \new_[96077]_ , \new_[96078]_ ,
    \new_[96081]_ , \new_[96084]_ , \new_[96085]_ , \new_[96088]_ ,
    \new_[96091]_ , \new_[96092]_ , \new_[96093]_ , \new_[96096]_ ,
    \new_[96099]_ , \new_[96100]_ , \new_[96103]_ , \new_[96106]_ ,
    \new_[96107]_ , \new_[96108]_ , \new_[96111]_ , \new_[96114]_ ,
    \new_[96115]_ , \new_[96118]_ , \new_[96121]_ , \new_[96122]_ ,
    \new_[96123]_ , \new_[96126]_ , \new_[96129]_ , \new_[96130]_ ,
    \new_[96133]_ , \new_[96136]_ , \new_[96137]_ , \new_[96138]_ ,
    \new_[96141]_ , \new_[96144]_ , \new_[96145]_ , \new_[96148]_ ,
    \new_[96151]_ , \new_[96152]_ , \new_[96153]_ , \new_[96156]_ ,
    \new_[96159]_ , \new_[96160]_ , \new_[96163]_ , \new_[96166]_ ,
    \new_[96167]_ , \new_[96168]_ , \new_[96171]_ , \new_[96174]_ ,
    \new_[96175]_ , \new_[96178]_ , \new_[96181]_ , \new_[96182]_ ,
    \new_[96183]_ , \new_[96186]_ , \new_[96189]_ , \new_[96190]_ ,
    \new_[96193]_ , \new_[96196]_ , \new_[96197]_ , \new_[96198]_ ,
    \new_[96201]_ , \new_[96204]_ , \new_[96205]_ , \new_[96208]_ ,
    \new_[96211]_ , \new_[96212]_ , \new_[96213]_ , \new_[96216]_ ,
    \new_[96219]_ , \new_[96220]_ , \new_[96223]_ , \new_[96226]_ ,
    \new_[96227]_ , \new_[96228]_ , \new_[96231]_ , \new_[96234]_ ,
    \new_[96235]_ , \new_[96238]_ , \new_[96241]_ , \new_[96242]_ ,
    \new_[96243]_ , \new_[96246]_ , \new_[96249]_ , \new_[96250]_ ,
    \new_[96253]_ , \new_[96256]_ , \new_[96257]_ , \new_[96258]_ ,
    \new_[96261]_ , \new_[96264]_ , \new_[96265]_ , \new_[96268]_ ,
    \new_[96271]_ , \new_[96272]_ , \new_[96273]_ , \new_[96276]_ ,
    \new_[96279]_ , \new_[96280]_ , \new_[96283]_ , \new_[96286]_ ,
    \new_[96287]_ , \new_[96288]_ , \new_[96291]_ , \new_[96294]_ ,
    \new_[96295]_ , \new_[96298]_ , \new_[96301]_ , \new_[96302]_ ,
    \new_[96303]_ , \new_[96306]_ , \new_[96309]_ , \new_[96310]_ ,
    \new_[96313]_ , \new_[96316]_ , \new_[96317]_ , \new_[96318]_ ,
    \new_[96321]_ , \new_[96324]_ , \new_[96325]_ , \new_[96328]_ ,
    \new_[96331]_ , \new_[96332]_ , \new_[96333]_ , \new_[96336]_ ,
    \new_[96339]_ , \new_[96340]_ , \new_[96343]_ , \new_[96346]_ ,
    \new_[96347]_ , \new_[96348]_ , \new_[96351]_ , \new_[96354]_ ,
    \new_[96355]_ , \new_[96358]_ , \new_[96361]_ , \new_[96362]_ ,
    \new_[96363]_ , \new_[96366]_ , \new_[96369]_ , \new_[96370]_ ,
    \new_[96373]_ , \new_[96376]_ , \new_[96377]_ , \new_[96378]_ ,
    \new_[96381]_ , \new_[96384]_ , \new_[96385]_ , \new_[96388]_ ,
    \new_[96391]_ , \new_[96392]_ , \new_[96393]_ , \new_[96396]_ ,
    \new_[96399]_ , \new_[96400]_ , \new_[96403]_ , \new_[96406]_ ,
    \new_[96407]_ , \new_[96408]_ , \new_[96411]_ , \new_[96414]_ ,
    \new_[96415]_ , \new_[96418]_ , \new_[96421]_ , \new_[96422]_ ,
    \new_[96423]_ , \new_[96426]_ , \new_[96429]_ , \new_[96430]_ ,
    \new_[96433]_ , \new_[96436]_ , \new_[96437]_ , \new_[96438]_ ,
    \new_[96441]_ , \new_[96444]_ , \new_[96445]_ , \new_[96448]_ ,
    \new_[96451]_ , \new_[96452]_ , \new_[96453]_ , \new_[96456]_ ,
    \new_[96459]_ , \new_[96460]_ , \new_[96463]_ , \new_[96466]_ ,
    \new_[96467]_ , \new_[96468]_ , \new_[96471]_ , \new_[96474]_ ,
    \new_[96475]_ , \new_[96478]_ , \new_[96481]_ , \new_[96482]_ ,
    \new_[96483]_ , \new_[96486]_ , \new_[96489]_ , \new_[96490]_ ,
    \new_[96493]_ , \new_[96496]_ , \new_[96497]_ , \new_[96498]_ ,
    \new_[96501]_ , \new_[96504]_ , \new_[96505]_ , \new_[96508]_ ,
    \new_[96511]_ , \new_[96512]_ , \new_[96513]_ , \new_[96516]_ ,
    \new_[96519]_ , \new_[96520]_ , \new_[96523]_ , \new_[96526]_ ,
    \new_[96527]_ , \new_[96528]_ , \new_[96531]_ , \new_[96534]_ ,
    \new_[96535]_ , \new_[96538]_ , \new_[96541]_ , \new_[96542]_ ,
    \new_[96543]_ , \new_[96546]_ , \new_[96549]_ , \new_[96550]_ ,
    \new_[96553]_ , \new_[96556]_ , \new_[96557]_ , \new_[96558]_ ,
    \new_[96561]_ , \new_[96564]_ , \new_[96565]_ , \new_[96568]_ ,
    \new_[96571]_ , \new_[96572]_ , \new_[96573]_ , \new_[96576]_ ,
    \new_[96579]_ , \new_[96580]_ , \new_[96583]_ , \new_[96586]_ ,
    \new_[96587]_ , \new_[96588]_ , \new_[96591]_ , \new_[96594]_ ,
    \new_[96595]_ , \new_[96598]_ , \new_[96601]_ , \new_[96602]_ ,
    \new_[96603]_ , \new_[96606]_ , \new_[96609]_ , \new_[96610]_ ,
    \new_[96613]_ , \new_[96616]_ , \new_[96617]_ , \new_[96618]_ ,
    \new_[96621]_ , \new_[96624]_ , \new_[96625]_ , \new_[96628]_ ,
    \new_[96631]_ , \new_[96632]_ , \new_[96633]_ , \new_[96636]_ ,
    \new_[96639]_ , \new_[96640]_ , \new_[96643]_ , \new_[96646]_ ,
    \new_[96647]_ , \new_[96648]_ , \new_[96651]_ , \new_[96654]_ ,
    \new_[96655]_ , \new_[96658]_ , \new_[96661]_ , \new_[96662]_ ,
    \new_[96663]_ , \new_[96666]_ , \new_[96669]_ , \new_[96670]_ ,
    \new_[96673]_ , \new_[96676]_ , \new_[96677]_ , \new_[96678]_ ,
    \new_[96681]_ , \new_[96684]_ , \new_[96685]_ , \new_[96688]_ ,
    \new_[96691]_ , \new_[96692]_ , \new_[96693]_ , \new_[96696]_ ,
    \new_[96699]_ , \new_[96700]_ , \new_[96703]_ , \new_[96706]_ ,
    \new_[96707]_ , \new_[96708]_ , \new_[96711]_ , \new_[96714]_ ,
    \new_[96715]_ , \new_[96718]_ , \new_[96721]_ , \new_[96722]_ ,
    \new_[96723]_ , \new_[96726]_ , \new_[96729]_ , \new_[96730]_ ,
    \new_[96733]_ , \new_[96736]_ , \new_[96737]_ , \new_[96738]_ ,
    \new_[96741]_ , \new_[96744]_ , \new_[96745]_ , \new_[96748]_ ,
    \new_[96751]_ , \new_[96752]_ , \new_[96753]_ , \new_[96756]_ ,
    \new_[96759]_ , \new_[96760]_ , \new_[96763]_ , \new_[96766]_ ,
    \new_[96767]_ , \new_[96768]_ , \new_[96771]_ , \new_[96774]_ ,
    \new_[96775]_ , \new_[96778]_ , \new_[96781]_ , \new_[96782]_ ,
    \new_[96783]_ , \new_[96786]_ , \new_[96789]_ , \new_[96790]_ ,
    \new_[96793]_ , \new_[96796]_ , \new_[96797]_ , \new_[96798]_ ,
    \new_[96801]_ , \new_[96804]_ , \new_[96805]_ , \new_[96808]_ ,
    \new_[96811]_ , \new_[96812]_ , \new_[96813]_ , \new_[96816]_ ,
    \new_[96819]_ , \new_[96820]_ , \new_[96823]_ , \new_[96826]_ ,
    \new_[96827]_ , \new_[96828]_ , \new_[96831]_ , \new_[96834]_ ,
    \new_[96835]_ , \new_[96838]_ , \new_[96841]_ , \new_[96842]_ ,
    \new_[96843]_ , \new_[96846]_ , \new_[96849]_ , \new_[96850]_ ,
    \new_[96853]_ , \new_[96856]_ , \new_[96857]_ , \new_[96858]_ ,
    \new_[96861]_ , \new_[96864]_ , \new_[96865]_ , \new_[96868]_ ,
    \new_[96871]_ , \new_[96872]_ , \new_[96873]_ , \new_[96876]_ ,
    \new_[96879]_ , \new_[96880]_ , \new_[96883]_ , \new_[96886]_ ,
    \new_[96887]_ , \new_[96888]_ , \new_[96891]_ , \new_[96894]_ ,
    \new_[96895]_ , \new_[96898]_ , \new_[96901]_ , \new_[96902]_ ,
    \new_[96903]_ , \new_[96906]_ , \new_[96909]_ , \new_[96910]_ ,
    \new_[96913]_ , \new_[96916]_ , \new_[96917]_ , \new_[96918]_ ,
    \new_[96921]_ , \new_[96924]_ , \new_[96925]_ , \new_[96928]_ ,
    \new_[96931]_ , \new_[96932]_ , \new_[96933]_ , \new_[96936]_ ,
    \new_[96939]_ , \new_[96940]_ , \new_[96943]_ , \new_[96946]_ ,
    \new_[96947]_ , \new_[96948]_ , \new_[96951]_ , \new_[96954]_ ,
    \new_[96955]_ , \new_[96958]_ , \new_[96961]_ , \new_[96962]_ ,
    \new_[96963]_ , \new_[96966]_ , \new_[96969]_ , \new_[96970]_ ,
    \new_[96973]_ , \new_[96976]_ , \new_[96977]_ , \new_[96978]_ ,
    \new_[96981]_ , \new_[96984]_ , \new_[96985]_ , \new_[96988]_ ,
    \new_[96991]_ , \new_[96992]_ , \new_[96993]_ , \new_[96996]_ ,
    \new_[96999]_ , \new_[97000]_ , \new_[97003]_ , \new_[97006]_ ,
    \new_[97007]_ , \new_[97008]_ , \new_[97011]_ , \new_[97014]_ ,
    \new_[97015]_ , \new_[97018]_ , \new_[97021]_ , \new_[97022]_ ,
    \new_[97023]_ , \new_[97026]_ , \new_[97029]_ , \new_[97030]_ ,
    \new_[97033]_ , \new_[97036]_ , \new_[97037]_ , \new_[97038]_ ,
    \new_[97041]_ , \new_[97044]_ , \new_[97045]_ , \new_[97048]_ ,
    \new_[97051]_ , \new_[97052]_ , \new_[97053]_ , \new_[97056]_ ,
    \new_[97059]_ , \new_[97060]_ , \new_[97063]_ , \new_[97066]_ ,
    \new_[97067]_ , \new_[97068]_ , \new_[97071]_ , \new_[97074]_ ,
    \new_[97075]_ , \new_[97078]_ , \new_[97081]_ , \new_[97082]_ ,
    \new_[97083]_ , \new_[97086]_ , \new_[97089]_ , \new_[97090]_ ,
    \new_[97093]_ , \new_[97096]_ , \new_[97097]_ , \new_[97098]_ ,
    \new_[97101]_ , \new_[97104]_ , \new_[97105]_ , \new_[97108]_ ,
    \new_[97111]_ , \new_[97112]_ , \new_[97113]_ , \new_[97116]_ ,
    \new_[97119]_ , \new_[97120]_ , \new_[97123]_ , \new_[97126]_ ,
    \new_[97127]_ , \new_[97128]_ , \new_[97131]_ , \new_[97134]_ ,
    \new_[97135]_ , \new_[97138]_ , \new_[97141]_ , \new_[97142]_ ,
    \new_[97143]_ , \new_[97146]_ , \new_[97149]_ , \new_[97150]_ ,
    \new_[97153]_ , \new_[97156]_ , \new_[97157]_ , \new_[97158]_ ,
    \new_[97161]_ , \new_[97164]_ , \new_[97165]_ , \new_[97168]_ ,
    \new_[97171]_ , \new_[97172]_ , \new_[97173]_ , \new_[97176]_ ,
    \new_[97179]_ , \new_[97180]_ , \new_[97183]_ , \new_[97186]_ ,
    \new_[97187]_ , \new_[97188]_ , \new_[97191]_ , \new_[97194]_ ,
    \new_[97195]_ , \new_[97198]_ , \new_[97201]_ , \new_[97202]_ ,
    \new_[97203]_ , \new_[97206]_ , \new_[97209]_ , \new_[97210]_ ,
    \new_[97213]_ , \new_[97216]_ , \new_[97217]_ , \new_[97218]_ ,
    \new_[97221]_ , \new_[97224]_ , \new_[97225]_ , \new_[97228]_ ,
    \new_[97231]_ , \new_[97232]_ , \new_[97233]_ , \new_[97236]_ ,
    \new_[97239]_ , \new_[97240]_ , \new_[97243]_ , \new_[97246]_ ,
    \new_[97247]_ , \new_[97248]_ , \new_[97251]_ , \new_[97254]_ ,
    \new_[97255]_ , \new_[97258]_ , \new_[97261]_ , \new_[97262]_ ,
    \new_[97263]_ , \new_[97266]_ , \new_[97269]_ , \new_[97270]_ ,
    \new_[97273]_ , \new_[97276]_ , \new_[97277]_ , \new_[97278]_ ,
    \new_[97281]_ , \new_[97284]_ , \new_[97285]_ , \new_[97288]_ ,
    \new_[97291]_ , \new_[97292]_ , \new_[97293]_ , \new_[97296]_ ,
    \new_[97299]_ , \new_[97300]_ , \new_[97303]_ , \new_[97306]_ ,
    \new_[97307]_ , \new_[97308]_ , \new_[97311]_ , \new_[97314]_ ,
    \new_[97315]_ , \new_[97318]_ , \new_[97321]_ , \new_[97322]_ ,
    \new_[97323]_ , \new_[97326]_ , \new_[97329]_ , \new_[97330]_ ,
    \new_[97333]_ , \new_[97336]_ , \new_[97337]_ , \new_[97338]_ ,
    \new_[97341]_ , \new_[97344]_ , \new_[97345]_ , \new_[97348]_ ,
    \new_[97351]_ , \new_[97352]_ , \new_[97353]_ , \new_[97356]_ ,
    \new_[97359]_ , \new_[97360]_ , \new_[97363]_ , \new_[97366]_ ,
    \new_[97367]_ , \new_[97368]_ , \new_[97371]_ , \new_[97374]_ ,
    \new_[97375]_ , \new_[97378]_ , \new_[97381]_ , \new_[97382]_ ,
    \new_[97383]_ , \new_[97386]_ , \new_[97389]_ , \new_[97390]_ ,
    \new_[97393]_ , \new_[97396]_ , \new_[97397]_ , \new_[97398]_ ,
    \new_[97401]_ , \new_[97404]_ , \new_[97405]_ , \new_[97408]_ ,
    \new_[97411]_ , \new_[97412]_ , \new_[97413]_ , \new_[97416]_ ,
    \new_[97419]_ , \new_[97420]_ , \new_[97423]_ , \new_[97426]_ ,
    \new_[97427]_ , \new_[97428]_ , \new_[97431]_ , \new_[97434]_ ,
    \new_[97435]_ , \new_[97438]_ , \new_[97441]_ , \new_[97442]_ ,
    \new_[97443]_ , \new_[97446]_ , \new_[97449]_ , \new_[97450]_ ,
    \new_[97453]_ , \new_[97456]_ , \new_[97457]_ , \new_[97458]_ ,
    \new_[97461]_ , \new_[97464]_ , \new_[97465]_ , \new_[97468]_ ,
    \new_[97471]_ , \new_[97472]_ , \new_[97473]_ , \new_[97476]_ ,
    \new_[97479]_ , \new_[97480]_ , \new_[97483]_ , \new_[97486]_ ,
    \new_[97487]_ , \new_[97488]_ , \new_[97491]_ , \new_[97494]_ ,
    \new_[97495]_ , \new_[97498]_ , \new_[97501]_ , \new_[97502]_ ,
    \new_[97503]_ , \new_[97506]_ , \new_[97509]_ , \new_[97510]_ ,
    \new_[97513]_ , \new_[97516]_ , \new_[97517]_ , \new_[97518]_ ,
    \new_[97521]_ , \new_[97524]_ , \new_[97525]_ , \new_[97528]_ ,
    \new_[97531]_ , \new_[97532]_ , \new_[97533]_ , \new_[97536]_ ,
    \new_[97539]_ , \new_[97540]_ , \new_[97543]_ , \new_[97546]_ ,
    \new_[97547]_ , \new_[97548]_ , \new_[97551]_ , \new_[97554]_ ,
    \new_[97555]_ , \new_[97558]_ , \new_[97561]_ , \new_[97562]_ ,
    \new_[97563]_ , \new_[97566]_ , \new_[97569]_ , \new_[97570]_ ,
    \new_[97573]_ , \new_[97576]_ , \new_[97577]_ , \new_[97578]_ ,
    \new_[97581]_ , \new_[97584]_ , \new_[97585]_ , \new_[97588]_ ,
    \new_[97591]_ , \new_[97592]_ , \new_[97593]_ , \new_[97596]_ ,
    \new_[97599]_ , \new_[97600]_ , \new_[97603]_ , \new_[97606]_ ,
    \new_[97607]_ , \new_[97608]_ , \new_[97611]_ , \new_[97614]_ ,
    \new_[97615]_ , \new_[97618]_ , \new_[97621]_ , \new_[97622]_ ,
    \new_[97623]_ , \new_[97626]_ , \new_[97629]_ , \new_[97630]_ ,
    \new_[97633]_ , \new_[97636]_ , \new_[97637]_ , \new_[97638]_ ,
    \new_[97641]_ , \new_[97644]_ , \new_[97645]_ , \new_[97648]_ ,
    \new_[97651]_ , \new_[97652]_ , \new_[97653]_ , \new_[97656]_ ,
    \new_[97659]_ , \new_[97660]_ , \new_[97663]_ , \new_[97666]_ ,
    \new_[97667]_ , \new_[97668]_ , \new_[97671]_ , \new_[97674]_ ,
    \new_[97675]_ , \new_[97678]_ , \new_[97681]_ , \new_[97682]_ ,
    \new_[97683]_ , \new_[97686]_ , \new_[97689]_ , \new_[97690]_ ,
    \new_[97693]_ , \new_[97696]_ , \new_[97697]_ , \new_[97698]_ ,
    \new_[97701]_ , \new_[97704]_ , \new_[97705]_ , \new_[97708]_ ,
    \new_[97711]_ , \new_[97712]_ , \new_[97713]_ , \new_[97716]_ ,
    \new_[97719]_ , \new_[97720]_ , \new_[97723]_ , \new_[97726]_ ,
    \new_[97727]_ , \new_[97728]_ , \new_[97731]_ , \new_[97734]_ ,
    \new_[97735]_ , \new_[97738]_ , \new_[97741]_ , \new_[97742]_ ,
    \new_[97743]_ , \new_[97746]_ , \new_[97749]_ , \new_[97750]_ ,
    \new_[97753]_ , \new_[97756]_ , \new_[97757]_ , \new_[97758]_ ,
    \new_[97761]_ , \new_[97764]_ , \new_[97765]_ , \new_[97768]_ ,
    \new_[97771]_ , \new_[97772]_ , \new_[97773]_ , \new_[97776]_ ,
    \new_[97779]_ , \new_[97780]_ , \new_[97783]_ , \new_[97786]_ ,
    \new_[97787]_ , \new_[97788]_ , \new_[97791]_ , \new_[97794]_ ,
    \new_[97795]_ , \new_[97798]_ , \new_[97801]_ , \new_[97802]_ ,
    \new_[97803]_ , \new_[97806]_ , \new_[97809]_ , \new_[97810]_ ,
    \new_[97813]_ , \new_[97816]_ , \new_[97817]_ , \new_[97818]_ ,
    \new_[97821]_ , \new_[97824]_ , \new_[97825]_ , \new_[97828]_ ,
    \new_[97831]_ , \new_[97832]_ , \new_[97833]_ , \new_[97836]_ ,
    \new_[97839]_ , \new_[97840]_ , \new_[97843]_ , \new_[97846]_ ,
    \new_[97847]_ , \new_[97848]_ , \new_[97851]_ , \new_[97854]_ ,
    \new_[97855]_ , \new_[97858]_ , \new_[97861]_ , \new_[97862]_ ,
    \new_[97863]_ , \new_[97866]_ , \new_[97869]_ , \new_[97870]_ ,
    \new_[97873]_ , \new_[97876]_ , \new_[97877]_ , \new_[97878]_ ,
    \new_[97881]_ , \new_[97884]_ , \new_[97885]_ , \new_[97888]_ ,
    \new_[97891]_ , \new_[97892]_ , \new_[97893]_ , \new_[97896]_ ,
    \new_[97899]_ , \new_[97900]_ , \new_[97903]_ , \new_[97906]_ ,
    \new_[97907]_ , \new_[97908]_ , \new_[97911]_ , \new_[97914]_ ,
    \new_[97915]_ , \new_[97918]_ , \new_[97921]_ , \new_[97922]_ ,
    \new_[97923]_ , \new_[97926]_ , \new_[97929]_ , \new_[97930]_ ,
    \new_[97933]_ , \new_[97936]_ , \new_[97937]_ , \new_[97938]_ ,
    \new_[97941]_ , \new_[97944]_ , \new_[97945]_ , \new_[97948]_ ,
    \new_[97951]_ , \new_[97952]_ , \new_[97953]_ , \new_[97956]_ ,
    \new_[97959]_ , \new_[97960]_ , \new_[97963]_ , \new_[97966]_ ,
    \new_[97967]_ , \new_[97968]_ , \new_[97971]_ , \new_[97974]_ ,
    \new_[97975]_ , \new_[97978]_ , \new_[97981]_ , \new_[97982]_ ,
    \new_[97983]_ , \new_[97986]_ , \new_[97989]_ , \new_[97990]_ ,
    \new_[97993]_ , \new_[97996]_ , \new_[97997]_ , \new_[97998]_ ,
    \new_[98001]_ , \new_[98004]_ , \new_[98005]_ , \new_[98008]_ ,
    \new_[98011]_ , \new_[98012]_ , \new_[98013]_ , \new_[98016]_ ,
    \new_[98019]_ , \new_[98020]_ , \new_[98023]_ , \new_[98026]_ ,
    \new_[98027]_ , \new_[98028]_ , \new_[98031]_ , \new_[98034]_ ,
    \new_[98035]_ , \new_[98038]_ , \new_[98041]_ , \new_[98042]_ ,
    \new_[98043]_ , \new_[98046]_ , \new_[98049]_ , \new_[98050]_ ,
    \new_[98053]_ , \new_[98056]_ , \new_[98057]_ , \new_[98058]_ ,
    \new_[98061]_ , \new_[98064]_ , \new_[98065]_ , \new_[98068]_ ,
    \new_[98071]_ , \new_[98072]_ , \new_[98073]_ , \new_[98076]_ ,
    \new_[98079]_ , \new_[98080]_ , \new_[98083]_ , \new_[98086]_ ,
    \new_[98087]_ , \new_[98088]_ , \new_[98091]_ , \new_[98094]_ ,
    \new_[98095]_ , \new_[98098]_ , \new_[98101]_ , \new_[98102]_ ,
    \new_[98103]_ , \new_[98106]_ , \new_[98109]_ , \new_[98110]_ ,
    \new_[98113]_ , \new_[98116]_ , \new_[98117]_ , \new_[98118]_ ,
    \new_[98121]_ , \new_[98124]_ , \new_[98125]_ , \new_[98128]_ ,
    \new_[98131]_ , \new_[98132]_ , \new_[98133]_ , \new_[98136]_ ,
    \new_[98139]_ , \new_[98140]_ , \new_[98143]_ , \new_[98146]_ ,
    \new_[98147]_ , \new_[98148]_ , \new_[98151]_ , \new_[98154]_ ,
    \new_[98155]_ , \new_[98158]_ , \new_[98161]_ , \new_[98162]_ ,
    \new_[98163]_ , \new_[98166]_ , \new_[98169]_ , \new_[98170]_ ,
    \new_[98173]_ , \new_[98176]_ , \new_[98177]_ , \new_[98178]_ ,
    \new_[98181]_ , \new_[98184]_ , \new_[98185]_ , \new_[98188]_ ,
    \new_[98191]_ , \new_[98192]_ , \new_[98193]_ , \new_[98196]_ ,
    \new_[98199]_ , \new_[98200]_ , \new_[98203]_ , \new_[98206]_ ,
    \new_[98207]_ , \new_[98208]_ , \new_[98211]_ , \new_[98214]_ ,
    \new_[98215]_ , \new_[98218]_ , \new_[98221]_ , \new_[98222]_ ,
    \new_[98223]_ , \new_[98226]_ , \new_[98229]_ , \new_[98230]_ ,
    \new_[98233]_ , \new_[98236]_ , \new_[98237]_ , \new_[98238]_ ,
    \new_[98241]_ , \new_[98244]_ , \new_[98245]_ , \new_[98248]_ ,
    \new_[98251]_ , \new_[98252]_ , \new_[98253]_ , \new_[98256]_ ,
    \new_[98259]_ , \new_[98260]_ , \new_[98263]_ , \new_[98266]_ ,
    \new_[98267]_ , \new_[98268]_ , \new_[98271]_ , \new_[98274]_ ,
    \new_[98275]_ , \new_[98278]_ , \new_[98281]_ , \new_[98282]_ ,
    \new_[98283]_ , \new_[98286]_ , \new_[98289]_ , \new_[98290]_ ,
    \new_[98293]_ , \new_[98296]_ , \new_[98297]_ , \new_[98298]_ ,
    \new_[98301]_ , \new_[98304]_ , \new_[98305]_ , \new_[98308]_ ,
    \new_[98311]_ , \new_[98312]_ , \new_[98313]_ , \new_[98316]_ ,
    \new_[98319]_ , \new_[98320]_ , \new_[98323]_ , \new_[98326]_ ,
    \new_[98327]_ , \new_[98328]_ , \new_[98331]_ , \new_[98334]_ ,
    \new_[98335]_ , \new_[98338]_ , \new_[98341]_ , \new_[98342]_ ,
    \new_[98343]_ , \new_[98346]_ , \new_[98349]_ , \new_[98350]_ ,
    \new_[98353]_ , \new_[98356]_ , \new_[98357]_ , \new_[98358]_ ,
    \new_[98361]_ , \new_[98364]_ , \new_[98365]_ , \new_[98368]_ ,
    \new_[98371]_ , \new_[98372]_ , \new_[98373]_ , \new_[98376]_ ,
    \new_[98379]_ , \new_[98380]_ , \new_[98383]_ , \new_[98386]_ ,
    \new_[98387]_ , \new_[98388]_ , \new_[98391]_ , \new_[98394]_ ,
    \new_[98395]_ , \new_[98398]_ , \new_[98401]_ , \new_[98402]_ ,
    \new_[98403]_ , \new_[98406]_ , \new_[98409]_ , \new_[98410]_ ,
    \new_[98413]_ , \new_[98417]_ , \new_[98418]_ , \new_[98419]_ ,
    \new_[98420]_ , \new_[98423]_ , \new_[98426]_ , \new_[98427]_ ,
    \new_[98430]_ , \new_[98433]_ , \new_[98434]_ , \new_[98435]_ ,
    \new_[98438]_ , \new_[98441]_ , \new_[98442]_ , \new_[98445]_ ,
    \new_[98449]_ , \new_[98450]_ , \new_[98451]_ , \new_[98452]_ ,
    \new_[98455]_ , \new_[98458]_ , \new_[98459]_ , \new_[98462]_ ,
    \new_[98465]_ , \new_[98466]_ , \new_[98467]_ , \new_[98470]_ ,
    \new_[98473]_ , \new_[98474]_ , \new_[98477]_ , \new_[98481]_ ,
    \new_[98482]_ , \new_[98483]_ , \new_[98484]_ , \new_[98487]_ ,
    \new_[98490]_ , \new_[98491]_ , \new_[98494]_ , \new_[98497]_ ,
    \new_[98498]_ , \new_[98499]_ , \new_[98502]_ , \new_[98505]_ ,
    \new_[98506]_ , \new_[98509]_ , \new_[98513]_ , \new_[98514]_ ,
    \new_[98515]_ , \new_[98516]_ , \new_[98519]_ , \new_[98522]_ ,
    \new_[98523]_ , \new_[98526]_ , \new_[98529]_ , \new_[98530]_ ,
    \new_[98531]_ , \new_[98534]_ , \new_[98537]_ , \new_[98538]_ ,
    \new_[98541]_ , \new_[98545]_ , \new_[98546]_ , \new_[98547]_ ,
    \new_[98548]_ , \new_[98551]_ , \new_[98554]_ , \new_[98555]_ ,
    \new_[98558]_ , \new_[98561]_ , \new_[98562]_ , \new_[98563]_ ,
    \new_[98566]_ , \new_[98569]_ , \new_[98570]_ , \new_[98573]_ ,
    \new_[98577]_ , \new_[98578]_ , \new_[98579]_ , \new_[98580]_ ,
    \new_[98583]_ , \new_[98586]_ , \new_[98587]_ , \new_[98590]_ ,
    \new_[98593]_ , \new_[98594]_ , \new_[98595]_ , \new_[98598]_ ,
    \new_[98601]_ , \new_[98602]_ , \new_[98605]_ , \new_[98609]_ ,
    \new_[98610]_ , \new_[98611]_ , \new_[98612]_ , \new_[98615]_ ,
    \new_[98618]_ , \new_[98619]_ , \new_[98622]_ , \new_[98625]_ ,
    \new_[98626]_ , \new_[98627]_ , \new_[98630]_ , \new_[98633]_ ,
    \new_[98634]_ , \new_[98637]_ , \new_[98641]_ , \new_[98642]_ ,
    \new_[98643]_ , \new_[98644]_ , \new_[98647]_ , \new_[98650]_ ,
    \new_[98651]_ , \new_[98654]_ , \new_[98657]_ , \new_[98658]_ ,
    \new_[98659]_ , \new_[98662]_ , \new_[98665]_ , \new_[98666]_ ,
    \new_[98669]_ , \new_[98673]_ , \new_[98674]_ , \new_[98675]_ ,
    \new_[98676]_ , \new_[98679]_ , \new_[98682]_ , \new_[98683]_ ,
    \new_[98686]_ , \new_[98689]_ , \new_[98690]_ , \new_[98691]_ ,
    \new_[98694]_ , \new_[98697]_ , \new_[98698]_ , \new_[98701]_ ,
    \new_[98705]_ , \new_[98706]_ , \new_[98707]_ , \new_[98708]_ ,
    \new_[98711]_ , \new_[98714]_ , \new_[98715]_ , \new_[98718]_ ,
    \new_[98721]_ , \new_[98722]_ , \new_[98723]_ , \new_[98726]_ ,
    \new_[98729]_ , \new_[98730]_ , \new_[98733]_ , \new_[98737]_ ,
    \new_[98738]_ , \new_[98739]_ , \new_[98740]_ , \new_[98743]_ ,
    \new_[98746]_ , \new_[98747]_ , \new_[98750]_ , \new_[98753]_ ,
    \new_[98754]_ , \new_[98755]_ , \new_[98758]_ , \new_[98761]_ ,
    \new_[98762]_ , \new_[98765]_ , \new_[98769]_ , \new_[98770]_ ,
    \new_[98771]_ , \new_[98772]_ , \new_[98775]_ , \new_[98778]_ ,
    \new_[98779]_ , \new_[98782]_ , \new_[98785]_ , \new_[98786]_ ,
    \new_[98787]_ , \new_[98790]_ , \new_[98793]_ , \new_[98794]_ ,
    \new_[98797]_ , \new_[98801]_ , \new_[98802]_ , \new_[98803]_ ,
    \new_[98804]_ , \new_[98807]_ , \new_[98810]_ , \new_[98811]_ ,
    \new_[98814]_ , \new_[98817]_ , \new_[98818]_ , \new_[98819]_ ,
    \new_[98822]_ , \new_[98825]_ , \new_[98826]_ , \new_[98829]_ ,
    \new_[98833]_ , \new_[98834]_ , \new_[98835]_ , \new_[98836]_ ,
    \new_[98839]_ , \new_[98842]_ , \new_[98843]_ , \new_[98846]_ ,
    \new_[98849]_ , \new_[98850]_ , \new_[98851]_ , \new_[98854]_ ,
    \new_[98857]_ , \new_[98858]_ , \new_[98861]_ , \new_[98865]_ ,
    \new_[98866]_ , \new_[98867]_ , \new_[98868]_ , \new_[98871]_ ,
    \new_[98874]_ , \new_[98875]_ , \new_[98878]_ , \new_[98881]_ ,
    \new_[98882]_ , \new_[98883]_ , \new_[98886]_ , \new_[98889]_ ,
    \new_[98890]_ , \new_[98893]_ , \new_[98897]_ , \new_[98898]_ ,
    \new_[98899]_ , \new_[98900]_ , \new_[98903]_ , \new_[98906]_ ,
    \new_[98907]_ , \new_[98910]_ , \new_[98913]_ , \new_[98914]_ ,
    \new_[98915]_ , \new_[98918]_ , \new_[98921]_ , \new_[98922]_ ,
    \new_[98925]_ , \new_[98929]_ , \new_[98930]_ , \new_[98931]_ ,
    \new_[98932]_ , \new_[98935]_ , \new_[98938]_ , \new_[98939]_ ,
    \new_[98942]_ , \new_[98945]_ , \new_[98946]_ , \new_[98947]_ ,
    \new_[98950]_ , \new_[98953]_ , \new_[98954]_ , \new_[98957]_ ,
    \new_[98961]_ , \new_[98962]_ , \new_[98963]_ , \new_[98964]_ ,
    \new_[98967]_ , \new_[98970]_ , \new_[98971]_ , \new_[98974]_ ,
    \new_[98977]_ , \new_[98978]_ , \new_[98979]_ , \new_[98982]_ ,
    \new_[98985]_ , \new_[98986]_ , \new_[98989]_ , \new_[98993]_ ,
    \new_[98994]_ , \new_[98995]_ , \new_[98996]_ , \new_[98999]_ ,
    \new_[99002]_ , \new_[99003]_ , \new_[99006]_ , \new_[99009]_ ,
    \new_[99010]_ , \new_[99011]_ , \new_[99014]_ , \new_[99017]_ ,
    \new_[99018]_ , \new_[99021]_ , \new_[99025]_ , \new_[99026]_ ,
    \new_[99027]_ , \new_[99028]_ , \new_[99031]_ , \new_[99034]_ ,
    \new_[99035]_ , \new_[99038]_ , \new_[99041]_ , \new_[99042]_ ,
    \new_[99043]_ , \new_[99046]_ , \new_[99049]_ , \new_[99050]_ ,
    \new_[99053]_ , \new_[99057]_ , \new_[99058]_ , \new_[99059]_ ,
    \new_[99060]_ , \new_[99063]_ , \new_[99066]_ , \new_[99067]_ ,
    \new_[99070]_ , \new_[99073]_ , \new_[99074]_ , \new_[99075]_ ,
    \new_[99078]_ , \new_[99081]_ , \new_[99082]_ , \new_[99085]_ ,
    \new_[99089]_ , \new_[99090]_ , \new_[99091]_ , \new_[99092]_ ,
    \new_[99095]_ , \new_[99098]_ , \new_[99099]_ , \new_[99102]_ ,
    \new_[99105]_ , \new_[99106]_ , \new_[99107]_ , \new_[99110]_ ,
    \new_[99113]_ , \new_[99114]_ , \new_[99117]_ , \new_[99121]_ ,
    \new_[99122]_ , \new_[99123]_ , \new_[99124]_ , \new_[99127]_ ,
    \new_[99130]_ , \new_[99131]_ , \new_[99134]_ , \new_[99137]_ ,
    \new_[99138]_ , \new_[99139]_ , \new_[99142]_ , \new_[99145]_ ,
    \new_[99146]_ , \new_[99149]_ , \new_[99153]_ , \new_[99154]_ ,
    \new_[99155]_ , \new_[99156]_ , \new_[99159]_ , \new_[99162]_ ,
    \new_[99163]_ , \new_[99166]_ , \new_[99169]_ , \new_[99170]_ ,
    \new_[99171]_ , \new_[99174]_ , \new_[99177]_ , \new_[99178]_ ,
    \new_[99181]_ , \new_[99185]_ , \new_[99186]_ , \new_[99187]_ ,
    \new_[99188]_ , \new_[99191]_ , \new_[99194]_ , \new_[99195]_ ,
    \new_[99198]_ , \new_[99201]_ , \new_[99202]_ , \new_[99203]_ ,
    \new_[99206]_ , \new_[99209]_ , \new_[99210]_ , \new_[99213]_ ,
    \new_[99217]_ , \new_[99218]_ , \new_[99219]_ , \new_[99220]_ ,
    \new_[99223]_ , \new_[99226]_ , \new_[99227]_ , \new_[99230]_ ,
    \new_[99233]_ , \new_[99234]_ , \new_[99235]_ , \new_[99238]_ ,
    \new_[99241]_ , \new_[99242]_ , \new_[99245]_ , \new_[99249]_ ,
    \new_[99250]_ , \new_[99251]_ , \new_[99252]_ , \new_[99255]_ ,
    \new_[99258]_ , \new_[99259]_ , \new_[99262]_ , \new_[99265]_ ,
    \new_[99266]_ , \new_[99267]_ , \new_[99270]_ , \new_[99273]_ ,
    \new_[99274]_ , \new_[99277]_ , \new_[99281]_ , \new_[99282]_ ,
    \new_[99283]_ , \new_[99284]_ , \new_[99287]_ , \new_[99290]_ ,
    \new_[99291]_ , \new_[99294]_ , \new_[99297]_ , \new_[99298]_ ,
    \new_[99299]_ , \new_[99302]_ , \new_[99305]_ , \new_[99306]_ ,
    \new_[99309]_ , \new_[99313]_ , \new_[99314]_ , \new_[99315]_ ,
    \new_[99316]_ , \new_[99319]_ , \new_[99322]_ , \new_[99323]_ ,
    \new_[99326]_ , \new_[99329]_ , \new_[99330]_ , \new_[99331]_ ,
    \new_[99334]_ , \new_[99337]_ , \new_[99338]_ , \new_[99341]_ ,
    \new_[99345]_ , \new_[99346]_ , \new_[99347]_ , \new_[99348]_ ,
    \new_[99351]_ , \new_[99354]_ , \new_[99355]_ , \new_[99358]_ ,
    \new_[99361]_ , \new_[99362]_ , \new_[99363]_ , \new_[99366]_ ,
    \new_[99369]_ , \new_[99370]_ , \new_[99373]_ , \new_[99377]_ ,
    \new_[99378]_ , \new_[99379]_ , \new_[99380]_ , \new_[99383]_ ,
    \new_[99386]_ , \new_[99387]_ , \new_[99390]_ , \new_[99393]_ ,
    \new_[99394]_ , \new_[99395]_ , \new_[99398]_ , \new_[99401]_ ,
    \new_[99402]_ , \new_[99405]_ , \new_[99409]_ , \new_[99410]_ ,
    \new_[99411]_ , \new_[99412]_ , \new_[99415]_ , \new_[99418]_ ,
    \new_[99419]_ , \new_[99422]_ , \new_[99425]_ , \new_[99426]_ ,
    \new_[99427]_ , \new_[99430]_ , \new_[99433]_ , \new_[99434]_ ,
    \new_[99437]_ , \new_[99441]_ , \new_[99442]_ , \new_[99443]_ ,
    \new_[99444]_ , \new_[99447]_ , \new_[99450]_ , \new_[99451]_ ,
    \new_[99454]_ , \new_[99457]_ , \new_[99458]_ , \new_[99459]_ ,
    \new_[99462]_ , \new_[99465]_ , \new_[99466]_ , \new_[99469]_ ,
    \new_[99473]_ , \new_[99474]_ , \new_[99475]_ , \new_[99476]_ ,
    \new_[99479]_ , \new_[99482]_ , \new_[99483]_ , \new_[99486]_ ,
    \new_[99489]_ , \new_[99490]_ , \new_[99491]_ , \new_[99494]_ ,
    \new_[99497]_ , \new_[99498]_ , \new_[99501]_ , \new_[99505]_ ,
    \new_[99506]_ , \new_[99507]_ , \new_[99508]_ , \new_[99511]_ ,
    \new_[99514]_ , \new_[99515]_ , \new_[99518]_ , \new_[99521]_ ,
    \new_[99522]_ , \new_[99523]_ , \new_[99526]_ , \new_[99529]_ ,
    \new_[99530]_ , \new_[99533]_ , \new_[99537]_ , \new_[99538]_ ,
    \new_[99539]_ , \new_[99540]_ , \new_[99543]_ , \new_[99546]_ ,
    \new_[99547]_ , \new_[99550]_ , \new_[99553]_ , \new_[99554]_ ,
    \new_[99555]_ , \new_[99558]_ , \new_[99561]_ , \new_[99562]_ ,
    \new_[99565]_ , \new_[99569]_ , \new_[99570]_ , \new_[99571]_ ,
    \new_[99572]_ , \new_[99575]_ , \new_[99578]_ , \new_[99579]_ ,
    \new_[99582]_ , \new_[99585]_ , \new_[99586]_ , \new_[99587]_ ,
    \new_[99590]_ , \new_[99593]_ , \new_[99594]_ , \new_[99597]_ ,
    \new_[99601]_ , \new_[99602]_ , \new_[99603]_ , \new_[99604]_ ,
    \new_[99607]_ , \new_[99610]_ , \new_[99611]_ , \new_[99614]_ ,
    \new_[99617]_ , \new_[99618]_ , \new_[99619]_ , \new_[99622]_ ,
    \new_[99625]_ , \new_[99626]_ , \new_[99629]_ , \new_[99633]_ ,
    \new_[99634]_ , \new_[99635]_ , \new_[99636]_ , \new_[99639]_ ,
    \new_[99642]_ , \new_[99643]_ , \new_[99646]_ , \new_[99649]_ ,
    \new_[99650]_ , \new_[99651]_ , \new_[99654]_ , \new_[99657]_ ,
    \new_[99658]_ , \new_[99661]_ , \new_[99665]_ , \new_[99666]_ ,
    \new_[99667]_ , \new_[99668]_ , \new_[99671]_ , \new_[99674]_ ,
    \new_[99675]_ , \new_[99678]_ , \new_[99681]_ , \new_[99682]_ ,
    \new_[99683]_ , \new_[99686]_ , \new_[99689]_ , \new_[99690]_ ,
    \new_[99693]_ , \new_[99697]_ , \new_[99698]_ , \new_[99699]_ ,
    \new_[99700]_ , \new_[99703]_ , \new_[99706]_ , \new_[99707]_ ,
    \new_[99710]_ , \new_[99713]_ , \new_[99714]_ , \new_[99715]_ ,
    \new_[99718]_ , \new_[99721]_ , \new_[99722]_ , \new_[99725]_ ,
    \new_[99729]_ , \new_[99730]_ , \new_[99731]_ , \new_[99732]_ ,
    \new_[99735]_ , \new_[99738]_ , \new_[99739]_ , \new_[99742]_ ,
    \new_[99745]_ , \new_[99746]_ , \new_[99747]_ , \new_[99750]_ ,
    \new_[99753]_ , \new_[99754]_ , \new_[99757]_ , \new_[99761]_ ,
    \new_[99762]_ , \new_[99763]_ , \new_[99764]_ , \new_[99767]_ ,
    \new_[99770]_ , \new_[99771]_ , \new_[99774]_ , \new_[99777]_ ,
    \new_[99778]_ , \new_[99779]_ , \new_[99782]_ , \new_[99785]_ ,
    \new_[99786]_ , \new_[99789]_ , \new_[99793]_ , \new_[99794]_ ,
    \new_[99795]_ , \new_[99796]_ , \new_[99799]_ , \new_[99802]_ ,
    \new_[99803]_ , \new_[99806]_ , \new_[99809]_ , \new_[99810]_ ,
    \new_[99811]_ , \new_[99814]_ , \new_[99817]_ , \new_[99818]_ ,
    \new_[99821]_ , \new_[99825]_ , \new_[99826]_ , \new_[99827]_ ,
    \new_[99828]_ , \new_[99831]_ , \new_[99834]_ , \new_[99835]_ ,
    \new_[99838]_ , \new_[99841]_ , \new_[99842]_ , \new_[99843]_ ,
    \new_[99846]_ , \new_[99849]_ , \new_[99850]_ , \new_[99853]_ ,
    \new_[99857]_ , \new_[99858]_ , \new_[99859]_ , \new_[99860]_ ,
    \new_[99863]_ , \new_[99866]_ , \new_[99867]_ , \new_[99870]_ ,
    \new_[99873]_ , \new_[99874]_ , \new_[99875]_ , \new_[99878]_ ,
    \new_[99881]_ , \new_[99882]_ , \new_[99885]_ , \new_[99889]_ ,
    \new_[99890]_ , \new_[99891]_ , \new_[99892]_ , \new_[99895]_ ,
    \new_[99898]_ , \new_[99899]_ , \new_[99902]_ , \new_[99905]_ ,
    \new_[99906]_ , \new_[99907]_ , \new_[99910]_ , \new_[99913]_ ,
    \new_[99914]_ , \new_[99917]_ , \new_[99921]_ , \new_[99922]_ ,
    \new_[99923]_ , \new_[99924]_ , \new_[99927]_ , \new_[99930]_ ,
    \new_[99931]_ , \new_[99934]_ , \new_[99937]_ , \new_[99938]_ ,
    \new_[99939]_ , \new_[99942]_ , \new_[99945]_ , \new_[99946]_ ,
    \new_[99949]_ , \new_[99953]_ , \new_[99954]_ , \new_[99955]_ ,
    \new_[99956]_ , \new_[99959]_ , \new_[99962]_ , \new_[99963]_ ,
    \new_[99966]_ , \new_[99969]_ , \new_[99970]_ , \new_[99971]_ ,
    \new_[99974]_ , \new_[99977]_ , \new_[99978]_ , \new_[99981]_ ,
    \new_[99985]_ , \new_[99986]_ , \new_[99987]_ , \new_[99988]_ ,
    \new_[99991]_ , \new_[99994]_ , \new_[99995]_ , \new_[99998]_ ,
    \new_[100001]_ , \new_[100002]_ , \new_[100003]_ , \new_[100006]_ ,
    \new_[100009]_ , \new_[100010]_ , \new_[100013]_ , \new_[100017]_ ,
    \new_[100018]_ , \new_[100019]_ , \new_[100020]_ , \new_[100023]_ ,
    \new_[100026]_ , \new_[100027]_ , \new_[100030]_ , \new_[100033]_ ,
    \new_[100034]_ , \new_[100035]_ , \new_[100038]_ , \new_[100041]_ ,
    \new_[100042]_ , \new_[100045]_ , \new_[100049]_ , \new_[100050]_ ,
    \new_[100051]_ , \new_[100052]_ , \new_[100055]_ , \new_[100058]_ ,
    \new_[100059]_ , \new_[100062]_ , \new_[100065]_ , \new_[100066]_ ,
    \new_[100067]_ , \new_[100070]_ , \new_[100073]_ , \new_[100074]_ ,
    \new_[100077]_ , \new_[100081]_ , \new_[100082]_ , \new_[100083]_ ,
    \new_[100084]_ , \new_[100087]_ , \new_[100090]_ , \new_[100091]_ ,
    \new_[100094]_ , \new_[100097]_ , \new_[100098]_ , \new_[100099]_ ,
    \new_[100102]_ , \new_[100105]_ , \new_[100106]_ , \new_[100109]_ ,
    \new_[100113]_ , \new_[100114]_ , \new_[100115]_ , \new_[100116]_ ,
    \new_[100119]_ , \new_[100122]_ , \new_[100123]_ , \new_[100126]_ ,
    \new_[100129]_ , \new_[100130]_ , \new_[100131]_ , \new_[100134]_ ,
    \new_[100137]_ , \new_[100138]_ , \new_[100141]_ , \new_[100145]_ ,
    \new_[100146]_ , \new_[100147]_ , \new_[100148]_ , \new_[100151]_ ,
    \new_[100154]_ , \new_[100155]_ , \new_[100158]_ , \new_[100161]_ ,
    \new_[100162]_ , \new_[100163]_ , \new_[100166]_ , \new_[100169]_ ,
    \new_[100170]_ , \new_[100173]_ , \new_[100177]_ , \new_[100178]_ ,
    \new_[100179]_ , \new_[100180]_ , \new_[100183]_ , \new_[100186]_ ,
    \new_[100187]_ , \new_[100190]_ , \new_[100193]_ , \new_[100194]_ ,
    \new_[100195]_ , \new_[100198]_ , \new_[100201]_ , \new_[100202]_ ,
    \new_[100205]_ , \new_[100209]_ , \new_[100210]_ , \new_[100211]_ ,
    \new_[100212]_ , \new_[100215]_ , \new_[100218]_ , \new_[100219]_ ,
    \new_[100222]_ , \new_[100225]_ , \new_[100226]_ , \new_[100227]_ ,
    \new_[100230]_ , \new_[100233]_ , \new_[100234]_ , \new_[100237]_ ,
    \new_[100241]_ , \new_[100242]_ , \new_[100243]_ , \new_[100244]_ ,
    \new_[100247]_ , \new_[100250]_ , \new_[100251]_ , \new_[100254]_ ,
    \new_[100257]_ , \new_[100258]_ , \new_[100259]_ , \new_[100262]_ ,
    \new_[100265]_ , \new_[100266]_ , \new_[100269]_ , \new_[100273]_ ,
    \new_[100274]_ , \new_[100275]_ , \new_[100276]_ , \new_[100279]_ ,
    \new_[100282]_ , \new_[100283]_ , \new_[100286]_ , \new_[100289]_ ,
    \new_[100290]_ , \new_[100291]_ , \new_[100294]_ , \new_[100297]_ ,
    \new_[100298]_ , \new_[100301]_ , \new_[100305]_ , \new_[100306]_ ,
    \new_[100307]_ , \new_[100308]_ , \new_[100311]_ , \new_[100314]_ ,
    \new_[100315]_ , \new_[100318]_ , \new_[100321]_ , \new_[100322]_ ,
    \new_[100323]_ , \new_[100326]_ , \new_[100329]_ , \new_[100330]_ ,
    \new_[100333]_ , \new_[100337]_ , \new_[100338]_ , \new_[100339]_ ,
    \new_[100340]_ , \new_[100343]_ , \new_[100346]_ , \new_[100347]_ ,
    \new_[100350]_ , \new_[100353]_ , \new_[100354]_ , \new_[100355]_ ,
    \new_[100358]_ , \new_[100361]_ , \new_[100362]_ , \new_[100365]_ ,
    \new_[100369]_ , \new_[100370]_ , \new_[100371]_ , \new_[100372]_ ,
    \new_[100375]_ , \new_[100378]_ , \new_[100379]_ , \new_[100382]_ ,
    \new_[100385]_ , \new_[100386]_ , \new_[100387]_ , \new_[100390]_ ,
    \new_[100393]_ , \new_[100394]_ , \new_[100397]_ , \new_[100401]_ ,
    \new_[100402]_ , \new_[100403]_ , \new_[100404]_ , \new_[100407]_ ,
    \new_[100410]_ , \new_[100411]_ , \new_[100414]_ , \new_[100417]_ ,
    \new_[100418]_ , \new_[100419]_ , \new_[100422]_ , \new_[100425]_ ,
    \new_[100426]_ , \new_[100429]_ , \new_[100433]_ , \new_[100434]_ ,
    \new_[100435]_ , \new_[100436]_ , \new_[100439]_ , \new_[100442]_ ,
    \new_[100443]_ , \new_[100446]_ , \new_[100449]_ , \new_[100450]_ ,
    \new_[100451]_ , \new_[100454]_ , \new_[100457]_ , \new_[100458]_ ,
    \new_[100461]_ , \new_[100465]_ , \new_[100466]_ , \new_[100467]_ ,
    \new_[100468]_ , \new_[100471]_ , \new_[100474]_ , \new_[100475]_ ,
    \new_[100478]_ , \new_[100481]_ , \new_[100482]_ , \new_[100483]_ ,
    \new_[100486]_ , \new_[100489]_ , \new_[100490]_ , \new_[100493]_ ,
    \new_[100497]_ , \new_[100498]_ , \new_[100499]_ , \new_[100500]_ ,
    \new_[100503]_ , \new_[100506]_ , \new_[100507]_ , \new_[100510]_ ,
    \new_[100513]_ , \new_[100514]_ , \new_[100515]_ , \new_[100518]_ ,
    \new_[100521]_ , \new_[100522]_ , \new_[100525]_ , \new_[100529]_ ,
    \new_[100530]_ , \new_[100531]_ , \new_[100532]_ , \new_[100535]_ ,
    \new_[100538]_ , \new_[100539]_ , \new_[100542]_ , \new_[100545]_ ,
    \new_[100546]_ , \new_[100547]_ , \new_[100550]_ , \new_[100553]_ ,
    \new_[100554]_ , \new_[100557]_ , \new_[100561]_ , \new_[100562]_ ,
    \new_[100563]_ , \new_[100564]_ , \new_[100567]_ , \new_[100570]_ ,
    \new_[100571]_ , \new_[100574]_ , \new_[100577]_ , \new_[100578]_ ,
    \new_[100579]_ , \new_[100582]_ , \new_[100585]_ , \new_[100586]_ ,
    \new_[100589]_ , \new_[100593]_ , \new_[100594]_ , \new_[100595]_ ,
    \new_[100596]_ , \new_[100599]_ , \new_[100602]_ , \new_[100603]_ ,
    \new_[100606]_ , \new_[100609]_ , \new_[100610]_ , \new_[100611]_ ,
    \new_[100614]_ , \new_[100617]_ , \new_[100618]_ , \new_[100621]_ ,
    \new_[100625]_ , \new_[100626]_ , \new_[100627]_ , \new_[100628]_ ,
    \new_[100631]_ , \new_[100634]_ , \new_[100635]_ , \new_[100638]_ ,
    \new_[100641]_ , \new_[100642]_ , \new_[100643]_ , \new_[100646]_ ,
    \new_[100649]_ , \new_[100650]_ , \new_[100653]_ , \new_[100657]_ ,
    \new_[100658]_ , \new_[100659]_ , \new_[100660]_ , \new_[100663]_ ,
    \new_[100666]_ , \new_[100667]_ , \new_[100670]_ , \new_[100673]_ ,
    \new_[100674]_ , \new_[100675]_ , \new_[100678]_ , \new_[100681]_ ,
    \new_[100682]_ , \new_[100685]_ , \new_[100689]_ , \new_[100690]_ ,
    \new_[100691]_ , \new_[100692]_ , \new_[100695]_ , \new_[100698]_ ,
    \new_[100699]_ , \new_[100702]_ , \new_[100705]_ , \new_[100706]_ ,
    \new_[100707]_ , \new_[100710]_ , \new_[100713]_ , \new_[100714]_ ,
    \new_[100717]_ , \new_[100721]_ , \new_[100722]_ , \new_[100723]_ ,
    \new_[100724]_ , \new_[100727]_ , \new_[100730]_ , \new_[100731]_ ,
    \new_[100734]_ , \new_[100737]_ , \new_[100738]_ , \new_[100739]_ ,
    \new_[100742]_ , \new_[100745]_ , \new_[100746]_ , \new_[100749]_ ,
    \new_[100753]_ , \new_[100754]_ , \new_[100755]_ , \new_[100756]_ ,
    \new_[100759]_ , \new_[100762]_ , \new_[100763]_ , \new_[100766]_ ,
    \new_[100769]_ , \new_[100770]_ , \new_[100771]_ , \new_[100774]_ ,
    \new_[100777]_ , \new_[100778]_ , \new_[100781]_ , \new_[100785]_ ,
    \new_[100786]_ , \new_[100787]_ , \new_[100788]_ , \new_[100791]_ ,
    \new_[100794]_ , \new_[100795]_ , \new_[100798]_ , \new_[100801]_ ,
    \new_[100802]_ , \new_[100803]_ , \new_[100806]_ , \new_[100809]_ ,
    \new_[100810]_ , \new_[100813]_ , \new_[100817]_ , \new_[100818]_ ,
    \new_[100819]_ , \new_[100820]_ , \new_[100823]_ , \new_[100826]_ ,
    \new_[100827]_ , \new_[100830]_ , \new_[100833]_ , \new_[100834]_ ,
    \new_[100835]_ , \new_[100838]_ , \new_[100841]_ , \new_[100842]_ ,
    \new_[100845]_ , \new_[100849]_ , \new_[100850]_ , \new_[100851]_ ,
    \new_[100852]_ , \new_[100855]_ , \new_[100858]_ , \new_[100859]_ ,
    \new_[100862]_ , \new_[100865]_ , \new_[100866]_ , \new_[100867]_ ,
    \new_[100870]_ , \new_[100873]_ , \new_[100874]_ , \new_[100877]_ ,
    \new_[100881]_ , \new_[100882]_ , \new_[100883]_ , \new_[100884]_ ,
    \new_[100887]_ , \new_[100890]_ , \new_[100891]_ , \new_[100894]_ ,
    \new_[100897]_ , \new_[100898]_ , \new_[100899]_ , \new_[100902]_ ,
    \new_[100905]_ , \new_[100906]_ , \new_[100909]_ , \new_[100913]_ ,
    \new_[100914]_ , \new_[100915]_ , \new_[100916]_ , \new_[100919]_ ,
    \new_[100922]_ , \new_[100923]_ , \new_[100926]_ , \new_[100929]_ ,
    \new_[100930]_ , \new_[100931]_ , \new_[100934]_ , \new_[100937]_ ,
    \new_[100938]_ , \new_[100941]_ , \new_[100945]_ , \new_[100946]_ ,
    \new_[100947]_ , \new_[100948]_ , \new_[100951]_ , \new_[100954]_ ,
    \new_[100955]_ , \new_[100958]_ , \new_[100962]_ , \new_[100963]_ ,
    \new_[100964]_ , \new_[100965]_ , \new_[100968]_ , \new_[100971]_ ,
    \new_[100972]_ , \new_[100975]_ , \new_[100979]_ , \new_[100980]_ ,
    \new_[100981]_ , \new_[100982]_ , \new_[100985]_ , \new_[100988]_ ,
    \new_[100989]_ , \new_[100992]_ , \new_[100996]_ , \new_[100997]_ ,
    \new_[100998]_ , \new_[100999]_ , \new_[101002]_ , \new_[101005]_ ,
    \new_[101006]_ , \new_[101009]_ , \new_[101013]_ , \new_[101014]_ ,
    \new_[101015]_ , \new_[101016]_ , \new_[101019]_ , \new_[101022]_ ,
    \new_[101023]_ , \new_[101026]_ , \new_[101030]_ , \new_[101031]_ ,
    \new_[101032]_ , \new_[101033]_ , \new_[101036]_ , \new_[101039]_ ,
    \new_[101040]_ , \new_[101043]_ , \new_[101047]_ , \new_[101048]_ ,
    \new_[101049]_ , \new_[101050]_ , \new_[101053]_ , \new_[101056]_ ,
    \new_[101057]_ , \new_[101060]_ , \new_[101064]_ , \new_[101065]_ ,
    \new_[101066]_ , \new_[101067]_ , \new_[101070]_ , \new_[101073]_ ,
    \new_[101074]_ , \new_[101077]_ , \new_[101081]_ , \new_[101082]_ ,
    \new_[101083]_ , \new_[101084]_ , \new_[101087]_ , \new_[101090]_ ,
    \new_[101091]_ , \new_[101094]_ , \new_[101098]_ , \new_[101099]_ ,
    \new_[101100]_ , \new_[101101]_ , \new_[101104]_ , \new_[101107]_ ,
    \new_[101108]_ , \new_[101111]_ , \new_[101115]_ , \new_[101116]_ ,
    \new_[101117]_ , \new_[101118]_ , \new_[101121]_ , \new_[101124]_ ,
    \new_[101125]_ , \new_[101128]_ , \new_[101132]_ , \new_[101133]_ ,
    \new_[101134]_ , \new_[101135]_ , \new_[101138]_ , \new_[101141]_ ,
    \new_[101142]_ , \new_[101145]_ , \new_[101149]_ , \new_[101150]_ ,
    \new_[101151]_ , \new_[101152]_ , \new_[101155]_ , \new_[101158]_ ,
    \new_[101159]_ , \new_[101162]_ , \new_[101166]_ , \new_[101167]_ ,
    \new_[101168]_ , \new_[101169]_ , \new_[101172]_ , \new_[101175]_ ,
    \new_[101176]_ , \new_[101179]_ , \new_[101183]_ , \new_[101184]_ ,
    \new_[101185]_ , \new_[101186]_ , \new_[101189]_ , \new_[101192]_ ,
    \new_[101193]_ , \new_[101196]_ , \new_[101200]_ , \new_[101201]_ ,
    \new_[101202]_ , \new_[101203]_ , \new_[101206]_ , \new_[101209]_ ,
    \new_[101210]_ , \new_[101213]_ , \new_[101217]_ , \new_[101218]_ ,
    \new_[101219]_ , \new_[101220]_ ;
  assign A139 = \new_[11104]_  | \new_[7403]_ ;
  assign \new_[1]_  = \new_[101220]_  & \new_[101203]_ ;
  assign \new_[2]_  = \new_[101186]_  & \new_[101169]_ ;
  assign \new_[3]_  = \new_[101152]_  & \new_[101135]_ ;
  assign \new_[4]_  = \new_[101118]_  & \new_[101101]_ ;
  assign \new_[5]_  = \new_[101084]_  & \new_[101067]_ ;
  assign \new_[6]_  = \new_[101050]_  & \new_[101033]_ ;
  assign \new_[7]_  = \new_[101016]_  & \new_[100999]_ ;
  assign \new_[8]_  = \new_[100982]_  & \new_[100965]_ ;
  assign \new_[9]_  = \new_[100948]_  & \new_[100931]_ ;
  assign \new_[10]_  = \new_[100916]_  & \new_[100899]_ ;
  assign \new_[11]_  = \new_[100884]_  & \new_[100867]_ ;
  assign \new_[12]_  = \new_[100852]_  & \new_[100835]_ ;
  assign \new_[13]_  = \new_[100820]_  & \new_[100803]_ ;
  assign \new_[14]_  = \new_[100788]_  & \new_[100771]_ ;
  assign \new_[15]_  = \new_[100756]_  & \new_[100739]_ ;
  assign \new_[16]_  = \new_[100724]_  & \new_[100707]_ ;
  assign \new_[17]_  = \new_[100692]_  & \new_[100675]_ ;
  assign \new_[18]_  = \new_[100660]_  & \new_[100643]_ ;
  assign \new_[19]_  = \new_[100628]_  & \new_[100611]_ ;
  assign \new_[20]_  = \new_[100596]_  & \new_[100579]_ ;
  assign \new_[21]_  = \new_[100564]_  & \new_[100547]_ ;
  assign \new_[22]_  = \new_[100532]_  & \new_[100515]_ ;
  assign \new_[23]_  = \new_[100500]_  & \new_[100483]_ ;
  assign \new_[24]_  = \new_[100468]_  & \new_[100451]_ ;
  assign \new_[25]_  = \new_[100436]_  & \new_[100419]_ ;
  assign \new_[26]_  = \new_[100404]_  & \new_[100387]_ ;
  assign \new_[27]_  = \new_[100372]_  & \new_[100355]_ ;
  assign \new_[28]_  = \new_[100340]_  & \new_[100323]_ ;
  assign \new_[29]_  = \new_[100308]_  & \new_[100291]_ ;
  assign \new_[30]_  = \new_[100276]_  & \new_[100259]_ ;
  assign \new_[31]_  = \new_[100244]_  & \new_[100227]_ ;
  assign \new_[32]_  = \new_[100212]_  & \new_[100195]_ ;
  assign \new_[33]_  = \new_[100180]_  & \new_[100163]_ ;
  assign \new_[34]_  = \new_[100148]_  & \new_[100131]_ ;
  assign \new_[35]_  = \new_[100116]_  & \new_[100099]_ ;
  assign \new_[36]_  = \new_[100084]_  & \new_[100067]_ ;
  assign \new_[37]_  = \new_[100052]_  & \new_[100035]_ ;
  assign \new_[38]_  = \new_[100020]_  & \new_[100003]_ ;
  assign \new_[39]_  = \new_[99988]_  & \new_[99971]_ ;
  assign \new_[40]_  = \new_[99956]_  & \new_[99939]_ ;
  assign \new_[41]_  = \new_[99924]_  & \new_[99907]_ ;
  assign \new_[42]_  = \new_[99892]_  & \new_[99875]_ ;
  assign \new_[43]_  = \new_[99860]_  & \new_[99843]_ ;
  assign \new_[44]_  = \new_[99828]_  & \new_[99811]_ ;
  assign \new_[45]_  = \new_[99796]_  & \new_[99779]_ ;
  assign \new_[46]_  = \new_[99764]_  & \new_[99747]_ ;
  assign \new_[47]_  = \new_[99732]_  & \new_[99715]_ ;
  assign \new_[48]_  = \new_[99700]_  & \new_[99683]_ ;
  assign \new_[49]_  = \new_[99668]_  & \new_[99651]_ ;
  assign \new_[50]_  = \new_[99636]_  & \new_[99619]_ ;
  assign \new_[51]_  = \new_[99604]_  & \new_[99587]_ ;
  assign \new_[52]_  = \new_[99572]_  & \new_[99555]_ ;
  assign \new_[53]_  = \new_[99540]_  & \new_[99523]_ ;
  assign \new_[54]_  = \new_[99508]_  & \new_[99491]_ ;
  assign \new_[55]_  = \new_[99476]_  & \new_[99459]_ ;
  assign \new_[56]_  = \new_[99444]_  & \new_[99427]_ ;
  assign \new_[57]_  = \new_[99412]_  & \new_[99395]_ ;
  assign \new_[58]_  = \new_[99380]_  & \new_[99363]_ ;
  assign \new_[59]_  = \new_[99348]_  & \new_[99331]_ ;
  assign \new_[60]_  = \new_[99316]_  & \new_[99299]_ ;
  assign \new_[61]_  = \new_[99284]_  & \new_[99267]_ ;
  assign \new_[62]_  = \new_[99252]_  & \new_[99235]_ ;
  assign \new_[63]_  = \new_[99220]_  & \new_[99203]_ ;
  assign \new_[64]_  = \new_[99188]_  & \new_[99171]_ ;
  assign \new_[65]_  = \new_[99156]_  & \new_[99139]_ ;
  assign \new_[66]_  = \new_[99124]_  & \new_[99107]_ ;
  assign \new_[67]_  = \new_[99092]_  & \new_[99075]_ ;
  assign \new_[68]_  = \new_[99060]_  & \new_[99043]_ ;
  assign \new_[69]_  = \new_[99028]_  & \new_[99011]_ ;
  assign \new_[70]_  = \new_[98996]_  & \new_[98979]_ ;
  assign \new_[71]_  = \new_[98964]_  & \new_[98947]_ ;
  assign \new_[72]_  = \new_[98932]_  & \new_[98915]_ ;
  assign \new_[73]_  = \new_[98900]_  & \new_[98883]_ ;
  assign \new_[74]_  = \new_[98868]_  & \new_[98851]_ ;
  assign \new_[75]_  = \new_[98836]_  & \new_[98819]_ ;
  assign \new_[76]_  = \new_[98804]_  & \new_[98787]_ ;
  assign \new_[77]_  = \new_[98772]_  & \new_[98755]_ ;
  assign \new_[78]_  = \new_[98740]_  & \new_[98723]_ ;
  assign \new_[79]_  = \new_[98708]_  & \new_[98691]_ ;
  assign \new_[80]_  = \new_[98676]_  & \new_[98659]_ ;
  assign \new_[81]_  = \new_[98644]_  & \new_[98627]_ ;
  assign \new_[82]_  = \new_[98612]_  & \new_[98595]_ ;
  assign \new_[83]_  = \new_[98580]_  & \new_[98563]_ ;
  assign \new_[84]_  = \new_[98548]_  & \new_[98531]_ ;
  assign \new_[85]_  = \new_[98516]_  & \new_[98499]_ ;
  assign \new_[86]_  = \new_[98484]_  & \new_[98467]_ ;
  assign \new_[87]_  = \new_[98452]_  & \new_[98435]_ ;
  assign \new_[88]_  = \new_[98420]_  & \new_[98403]_ ;
  assign \new_[89]_  = \new_[98388]_  & \new_[98373]_ ;
  assign \new_[90]_  = \new_[98358]_  & \new_[98343]_ ;
  assign \new_[91]_  = \new_[98328]_  & \new_[98313]_ ;
  assign \new_[92]_  = \new_[98298]_  & \new_[98283]_ ;
  assign \new_[93]_  = \new_[98268]_  & \new_[98253]_ ;
  assign \new_[94]_  = \new_[98238]_  & \new_[98223]_ ;
  assign \new_[95]_  = \new_[98208]_  & \new_[98193]_ ;
  assign \new_[96]_  = \new_[98178]_  & \new_[98163]_ ;
  assign \new_[97]_  = \new_[98148]_  & \new_[98133]_ ;
  assign \new_[98]_  = \new_[98118]_  & \new_[98103]_ ;
  assign \new_[99]_  = \new_[98088]_  & \new_[98073]_ ;
  assign \new_[100]_  = \new_[98058]_  & \new_[98043]_ ;
  assign \new_[101]_  = \new_[98028]_  & \new_[98013]_ ;
  assign \new_[102]_  = \new_[97998]_  & \new_[97983]_ ;
  assign \new_[103]_  = \new_[97968]_  & \new_[97953]_ ;
  assign \new_[104]_  = \new_[97938]_  & \new_[97923]_ ;
  assign \new_[105]_  = \new_[97908]_  & \new_[97893]_ ;
  assign \new_[106]_  = \new_[97878]_  & \new_[97863]_ ;
  assign \new_[107]_  = \new_[97848]_  & \new_[97833]_ ;
  assign \new_[108]_  = \new_[97818]_  & \new_[97803]_ ;
  assign \new_[109]_  = \new_[97788]_  & \new_[97773]_ ;
  assign \new_[110]_  = \new_[97758]_  & \new_[97743]_ ;
  assign \new_[111]_  = \new_[97728]_  & \new_[97713]_ ;
  assign \new_[112]_  = \new_[97698]_  & \new_[97683]_ ;
  assign \new_[113]_  = \new_[97668]_  & \new_[97653]_ ;
  assign \new_[114]_  = \new_[97638]_  & \new_[97623]_ ;
  assign \new_[115]_  = \new_[97608]_  & \new_[97593]_ ;
  assign \new_[116]_  = \new_[97578]_  & \new_[97563]_ ;
  assign \new_[117]_  = \new_[97548]_  & \new_[97533]_ ;
  assign \new_[118]_  = \new_[97518]_  & \new_[97503]_ ;
  assign \new_[119]_  = \new_[97488]_  & \new_[97473]_ ;
  assign \new_[120]_  = \new_[97458]_  & \new_[97443]_ ;
  assign \new_[121]_  = \new_[97428]_  & \new_[97413]_ ;
  assign \new_[122]_  = \new_[97398]_  & \new_[97383]_ ;
  assign \new_[123]_  = \new_[97368]_  & \new_[97353]_ ;
  assign \new_[124]_  = \new_[97338]_  & \new_[97323]_ ;
  assign \new_[125]_  = \new_[97308]_  & \new_[97293]_ ;
  assign \new_[126]_  = \new_[97278]_  & \new_[97263]_ ;
  assign \new_[127]_  = \new_[97248]_  & \new_[97233]_ ;
  assign \new_[128]_  = \new_[97218]_  & \new_[97203]_ ;
  assign \new_[129]_  = \new_[97188]_  & \new_[97173]_ ;
  assign \new_[130]_  = \new_[97158]_  & \new_[97143]_ ;
  assign \new_[131]_  = \new_[97128]_  & \new_[97113]_ ;
  assign \new_[132]_  = \new_[97098]_  & \new_[97083]_ ;
  assign \new_[133]_  = \new_[97068]_  & \new_[97053]_ ;
  assign \new_[134]_  = \new_[97038]_  & \new_[97023]_ ;
  assign \new_[135]_  = \new_[97008]_  & \new_[96993]_ ;
  assign \new_[136]_  = \new_[96978]_  & \new_[96963]_ ;
  assign \new_[137]_  = \new_[96948]_  & \new_[96933]_ ;
  assign \new_[138]_  = \new_[96918]_  & \new_[96903]_ ;
  assign \new_[139]_  = \new_[96888]_  & \new_[96873]_ ;
  assign \new_[140]_  = \new_[96858]_  & \new_[96843]_ ;
  assign \new_[141]_  = \new_[96828]_  & \new_[96813]_ ;
  assign \new_[142]_  = \new_[96798]_  & \new_[96783]_ ;
  assign \new_[143]_  = \new_[96768]_  & \new_[96753]_ ;
  assign \new_[144]_  = \new_[96738]_  & \new_[96723]_ ;
  assign \new_[145]_  = \new_[96708]_  & \new_[96693]_ ;
  assign \new_[146]_  = \new_[96678]_  & \new_[96663]_ ;
  assign \new_[147]_  = \new_[96648]_  & \new_[96633]_ ;
  assign \new_[148]_  = \new_[96618]_  & \new_[96603]_ ;
  assign \new_[149]_  = \new_[96588]_  & \new_[96573]_ ;
  assign \new_[150]_  = \new_[96558]_  & \new_[96543]_ ;
  assign \new_[151]_  = \new_[96528]_  & \new_[96513]_ ;
  assign \new_[152]_  = \new_[96498]_  & \new_[96483]_ ;
  assign \new_[153]_  = \new_[96468]_  & \new_[96453]_ ;
  assign \new_[154]_  = \new_[96438]_  & \new_[96423]_ ;
  assign \new_[155]_  = \new_[96408]_  & \new_[96393]_ ;
  assign \new_[156]_  = \new_[96378]_  & \new_[96363]_ ;
  assign \new_[157]_  = \new_[96348]_  & \new_[96333]_ ;
  assign \new_[158]_  = \new_[96318]_  & \new_[96303]_ ;
  assign \new_[159]_  = \new_[96288]_  & \new_[96273]_ ;
  assign \new_[160]_  = \new_[96258]_  & \new_[96243]_ ;
  assign \new_[161]_  = \new_[96228]_  & \new_[96213]_ ;
  assign \new_[162]_  = \new_[96198]_  & \new_[96183]_ ;
  assign \new_[163]_  = \new_[96168]_  & \new_[96153]_ ;
  assign \new_[164]_  = \new_[96138]_  & \new_[96123]_ ;
  assign \new_[165]_  = \new_[96108]_  & \new_[96093]_ ;
  assign \new_[166]_  = \new_[96078]_  & \new_[96063]_ ;
  assign \new_[167]_  = \new_[96048]_  & \new_[96033]_ ;
  assign \new_[168]_  = \new_[96018]_  & \new_[96003]_ ;
  assign \new_[169]_  = \new_[95988]_  & \new_[95973]_ ;
  assign \new_[170]_  = \new_[95958]_  & \new_[95943]_ ;
  assign \new_[171]_  = \new_[95928]_  & \new_[95913]_ ;
  assign \new_[172]_  = \new_[95898]_  & \new_[95883]_ ;
  assign \new_[173]_  = \new_[95868]_  & \new_[95853]_ ;
  assign \new_[174]_  = \new_[95838]_  & \new_[95823]_ ;
  assign \new_[175]_  = \new_[95808]_  & \new_[95793]_ ;
  assign \new_[176]_  = \new_[95778]_  & \new_[95763]_ ;
  assign \new_[177]_  = \new_[95748]_  & \new_[95733]_ ;
  assign \new_[178]_  = \new_[95718]_  & \new_[95703]_ ;
  assign \new_[179]_  = \new_[95688]_  & \new_[95673]_ ;
  assign \new_[180]_  = \new_[95658]_  & \new_[95643]_ ;
  assign \new_[181]_  = \new_[95628]_  & \new_[95613]_ ;
  assign \new_[182]_  = \new_[95598]_  & \new_[95583]_ ;
  assign \new_[183]_  = \new_[95568]_  & \new_[95553]_ ;
  assign \new_[184]_  = \new_[95538]_  & \new_[95523]_ ;
  assign \new_[185]_  = \new_[95508]_  & \new_[95493]_ ;
  assign \new_[186]_  = \new_[95478]_  & \new_[95463]_ ;
  assign \new_[187]_  = \new_[95448]_  & \new_[95433]_ ;
  assign \new_[188]_  = \new_[95418]_  & \new_[95403]_ ;
  assign \new_[189]_  = \new_[95388]_  & \new_[95373]_ ;
  assign \new_[190]_  = \new_[95358]_  & \new_[95343]_ ;
  assign \new_[191]_  = \new_[95328]_  & \new_[95313]_ ;
  assign \new_[192]_  = \new_[95298]_  & \new_[95283]_ ;
  assign \new_[193]_  = \new_[95268]_  & \new_[95253]_ ;
  assign \new_[194]_  = \new_[95238]_  & \new_[95223]_ ;
  assign \new_[195]_  = \new_[95208]_  & \new_[95193]_ ;
  assign \new_[196]_  = \new_[95178]_  & \new_[95163]_ ;
  assign \new_[197]_  = \new_[95148]_  & \new_[95133]_ ;
  assign \new_[198]_  = \new_[95118]_  & \new_[95103]_ ;
  assign \new_[199]_  = \new_[95088]_  & \new_[95073]_ ;
  assign \new_[200]_  = \new_[95058]_  & \new_[95043]_ ;
  assign \new_[201]_  = \new_[95028]_  & \new_[95013]_ ;
  assign \new_[202]_  = \new_[94998]_  & \new_[94983]_ ;
  assign \new_[203]_  = \new_[94968]_  & \new_[94953]_ ;
  assign \new_[204]_  = \new_[94938]_  & \new_[94923]_ ;
  assign \new_[205]_  = \new_[94908]_  & \new_[94893]_ ;
  assign \new_[206]_  = \new_[94878]_  & \new_[94863]_ ;
  assign \new_[207]_  = \new_[94848]_  & \new_[94833]_ ;
  assign \new_[208]_  = \new_[94818]_  & \new_[94803]_ ;
  assign \new_[209]_  = \new_[94788]_  & \new_[94773]_ ;
  assign \new_[210]_  = \new_[94758]_  & \new_[94743]_ ;
  assign \new_[211]_  = \new_[94728]_  & \new_[94713]_ ;
  assign \new_[212]_  = \new_[94698]_  & \new_[94683]_ ;
  assign \new_[213]_  = \new_[94668]_  & \new_[94653]_ ;
  assign \new_[214]_  = \new_[94638]_  & \new_[94623]_ ;
  assign \new_[215]_  = \new_[94608]_  & \new_[94593]_ ;
  assign \new_[216]_  = \new_[94578]_  & \new_[94563]_ ;
  assign \new_[217]_  = \new_[94548]_  & \new_[94533]_ ;
  assign \new_[218]_  = \new_[94518]_  & \new_[94503]_ ;
  assign \new_[219]_  = \new_[94488]_  & \new_[94473]_ ;
  assign \new_[220]_  = \new_[94458]_  & \new_[94443]_ ;
  assign \new_[221]_  = \new_[94428]_  & \new_[94413]_ ;
  assign \new_[222]_  = \new_[94398]_  & \new_[94383]_ ;
  assign \new_[223]_  = \new_[94368]_  & \new_[94353]_ ;
  assign \new_[224]_  = \new_[94338]_  & \new_[94323]_ ;
  assign \new_[225]_  = \new_[94308]_  & \new_[94293]_ ;
  assign \new_[226]_  = \new_[94278]_  & \new_[94263]_ ;
  assign \new_[227]_  = \new_[94248]_  & \new_[94233]_ ;
  assign \new_[228]_  = \new_[94218]_  & \new_[94203]_ ;
  assign \new_[229]_  = \new_[94188]_  & \new_[94173]_ ;
  assign \new_[230]_  = \new_[94158]_  & \new_[94143]_ ;
  assign \new_[231]_  = \new_[94128]_  & \new_[94113]_ ;
  assign \new_[232]_  = \new_[94098]_  & \new_[94083]_ ;
  assign \new_[233]_  = \new_[94068]_  & \new_[94053]_ ;
  assign \new_[234]_  = \new_[94038]_  & \new_[94023]_ ;
  assign \new_[235]_  = \new_[94008]_  & \new_[93993]_ ;
  assign \new_[236]_  = \new_[93978]_  & \new_[93963]_ ;
  assign \new_[237]_  = \new_[93948]_  & \new_[93933]_ ;
  assign \new_[238]_  = \new_[93918]_  & \new_[93903]_ ;
  assign \new_[239]_  = \new_[93888]_  & \new_[93873]_ ;
  assign \new_[240]_  = \new_[93858]_  & \new_[93843]_ ;
  assign \new_[241]_  = \new_[93828]_  & \new_[93813]_ ;
  assign \new_[242]_  = \new_[93798]_  & \new_[93783]_ ;
  assign \new_[243]_  = \new_[93768]_  & \new_[93753]_ ;
  assign \new_[244]_  = \new_[93738]_  & \new_[93723]_ ;
  assign \new_[245]_  = \new_[93708]_  & \new_[93693]_ ;
  assign \new_[246]_  = \new_[93678]_  & \new_[93663]_ ;
  assign \new_[247]_  = \new_[93648]_  & \new_[93633]_ ;
  assign \new_[248]_  = \new_[93618]_  & \new_[93603]_ ;
  assign \new_[249]_  = \new_[93588]_  & \new_[93573]_ ;
  assign \new_[250]_  = \new_[93558]_  & \new_[93543]_ ;
  assign \new_[251]_  = \new_[93528]_  & \new_[93513]_ ;
  assign \new_[252]_  = \new_[93498]_  & \new_[93483]_ ;
  assign \new_[253]_  = \new_[93468]_  & \new_[93453]_ ;
  assign \new_[254]_  = \new_[93438]_  & \new_[93423]_ ;
  assign \new_[255]_  = \new_[93408]_  & \new_[93393]_ ;
  assign \new_[256]_  = \new_[93378]_  & \new_[93363]_ ;
  assign \new_[257]_  = \new_[93348]_  & \new_[93333]_ ;
  assign \new_[258]_  = \new_[93318]_  & \new_[93303]_ ;
  assign \new_[259]_  = \new_[93288]_  & \new_[93273]_ ;
  assign \new_[260]_  = \new_[93258]_  & \new_[93243]_ ;
  assign \new_[261]_  = \new_[93228]_  & \new_[93213]_ ;
  assign \new_[262]_  = \new_[93198]_  & \new_[93183]_ ;
  assign \new_[263]_  = \new_[93168]_  & \new_[93153]_ ;
  assign \new_[264]_  = \new_[93138]_  & \new_[93123]_ ;
  assign \new_[265]_  = \new_[93108]_  & \new_[93093]_ ;
  assign \new_[266]_  = \new_[93078]_  & \new_[93063]_ ;
  assign \new_[267]_  = \new_[93048]_  & \new_[93033]_ ;
  assign \new_[268]_  = \new_[93018]_  & \new_[93003]_ ;
  assign \new_[269]_  = \new_[92988]_  & \new_[92973]_ ;
  assign \new_[270]_  = \new_[92958]_  & \new_[92943]_ ;
  assign \new_[271]_  = \new_[92928]_  & \new_[92913]_ ;
  assign \new_[272]_  = \new_[92898]_  & \new_[92883]_ ;
  assign \new_[273]_  = \new_[92868]_  & \new_[92853]_ ;
  assign \new_[274]_  = \new_[92838]_  & \new_[92823]_ ;
  assign \new_[275]_  = \new_[92808]_  & \new_[92793]_ ;
  assign \new_[276]_  = \new_[92778]_  & \new_[92763]_ ;
  assign \new_[277]_  = \new_[92748]_  & \new_[92733]_ ;
  assign \new_[278]_  = \new_[92718]_  & \new_[92703]_ ;
  assign \new_[279]_  = \new_[92688]_  & \new_[92673]_ ;
  assign \new_[280]_  = \new_[92658]_  & \new_[92643]_ ;
  assign \new_[281]_  = \new_[92628]_  & \new_[92613]_ ;
  assign \new_[282]_  = \new_[92598]_  & \new_[92583]_ ;
  assign \new_[283]_  = \new_[92568]_  & \new_[92553]_ ;
  assign \new_[284]_  = \new_[92538]_  & \new_[92523]_ ;
  assign \new_[285]_  = \new_[92508]_  & \new_[92493]_ ;
  assign \new_[286]_  = \new_[92478]_  & \new_[92463]_ ;
  assign \new_[287]_  = \new_[92448]_  & \new_[92433]_ ;
  assign \new_[288]_  = \new_[92418]_  & \new_[92403]_ ;
  assign \new_[289]_  = \new_[92388]_  & \new_[92373]_ ;
  assign \new_[290]_  = \new_[92358]_  & \new_[92343]_ ;
  assign \new_[291]_  = \new_[92328]_  & \new_[92313]_ ;
  assign \new_[292]_  = \new_[92298]_  & \new_[92283]_ ;
  assign \new_[293]_  = \new_[92268]_  & \new_[92253]_ ;
  assign \new_[294]_  = \new_[92238]_  & \new_[92223]_ ;
  assign \new_[295]_  = \new_[92208]_  & \new_[92193]_ ;
  assign \new_[296]_  = \new_[92178]_  & \new_[92163]_ ;
  assign \new_[297]_  = \new_[92148]_  & \new_[92133]_ ;
  assign \new_[298]_  = \new_[92118]_  & \new_[92103]_ ;
  assign \new_[299]_  = \new_[92088]_  & \new_[92073]_ ;
  assign \new_[300]_  = \new_[92058]_  & \new_[92043]_ ;
  assign \new_[301]_  = \new_[92028]_  & \new_[92013]_ ;
  assign \new_[302]_  = \new_[91998]_  & \new_[91983]_ ;
  assign \new_[303]_  = \new_[91968]_  & \new_[91953]_ ;
  assign \new_[304]_  = \new_[91938]_  & \new_[91923]_ ;
  assign \new_[305]_  = \new_[91908]_  & \new_[91893]_ ;
  assign \new_[306]_  = \new_[91878]_  & \new_[91863]_ ;
  assign \new_[307]_  = \new_[91848]_  & \new_[91833]_ ;
  assign \new_[308]_  = \new_[91818]_  & \new_[91803]_ ;
  assign \new_[309]_  = \new_[91788]_  & \new_[91773]_ ;
  assign \new_[310]_  = \new_[91758]_  & \new_[91743]_ ;
  assign \new_[311]_  = \new_[91728]_  & \new_[91713]_ ;
  assign \new_[312]_  = \new_[91698]_  & \new_[91683]_ ;
  assign \new_[313]_  = \new_[91668]_  & \new_[91653]_ ;
  assign \new_[314]_  = \new_[91638]_  & \new_[91623]_ ;
  assign \new_[315]_  = \new_[91608]_  & \new_[91593]_ ;
  assign \new_[316]_  = \new_[91578]_  & \new_[91563]_ ;
  assign \new_[317]_  = \new_[91548]_  & \new_[91533]_ ;
  assign \new_[318]_  = \new_[91518]_  & \new_[91503]_ ;
  assign \new_[319]_  = \new_[91488]_  & \new_[91473]_ ;
  assign \new_[320]_  = \new_[91458]_  & \new_[91443]_ ;
  assign \new_[321]_  = \new_[91428]_  & \new_[91413]_ ;
  assign \new_[322]_  = \new_[91398]_  & \new_[91383]_ ;
  assign \new_[323]_  = \new_[91368]_  & \new_[91353]_ ;
  assign \new_[324]_  = \new_[91338]_  & \new_[91323]_ ;
  assign \new_[325]_  = \new_[91308]_  & \new_[91293]_ ;
  assign \new_[326]_  = \new_[91278]_  & \new_[91263]_ ;
  assign \new_[327]_  = \new_[91248]_  & \new_[91233]_ ;
  assign \new_[328]_  = \new_[91218]_  & \new_[91203]_ ;
  assign \new_[329]_  = \new_[91188]_  & \new_[91173]_ ;
  assign \new_[330]_  = \new_[91158]_  & \new_[91143]_ ;
  assign \new_[331]_  = \new_[91128]_  & \new_[91113]_ ;
  assign \new_[332]_  = \new_[91098]_  & \new_[91083]_ ;
  assign \new_[333]_  = \new_[91068]_  & \new_[91053]_ ;
  assign \new_[334]_  = \new_[91038]_  & \new_[91023]_ ;
  assign \new_[335]_  = \new_[91008]_  & \new_[90993]_ ;
  assign \new_[336]_  = \new_[90978]_  & \new_[90963]_ ;
  assign \new_[337]_  = \new_[90948]_  & \new_[90933]_ ;
  assign \new_[338]_  = \new_[90918]_  & \new_[90903]_ ;
  assign \new_[339]_  = \new_[90888]_  & \new_[90873]_ ;
  assign \new_[340]_  = \new_[90858]_  & \new_[90843]_ ;
  assign \new_[341]_  = \new_[90828]_  & \new_[90813]_ ;
  assign \new_[342]_  = \new_[90798]_  & \new_[90783]_ ;
  assign \new_[343]_  = \new_[90768]_  & \new_[90753]_ ;
  assign \new_[344]_  = \new_[90738]_  & \new_[90723]_ ;
  assign \new_[345]_  = \new_[90708]_  & \new_[90693]_ ;
  assign \new_[346]_  = \new_[90678]_  & \new_[90663]_ ;
  assign \new_[347]_  = \new_[90648]_  & \new_[90633]_ ;
  assign \new_[348]_  = \new_[90618]_  & \new_[90603]_ ;
  assign \new_[349]_  = \new_[90588]_  & \new_[90573]_ ;
  assign \new_[350]_  = \new_[90558]_  & \new_[90543]_ ;
  assign \new_[351]_  = \new_[90528]_  & \new_[90513]_ ;
  assign \new_[352]_  = \new_[90498]_  & \new_[90483]_ ;
  assign \new_[353]_  = \new_[90468]_  & \new_[90453]_ ;
  assign \new_[354]_  = \new_[90438]_  & \new_[90423]_ ;
  assign \new_[355]_  = \new_[90408]_  & \new_[90393]_ ;
  assign \new_[356]_  = \new_[90378]_  & \new_[90363]_ ;
  assign \new_[357]_  = \new_[90348]_  & \new_[90333]_ ;
  assign \new_[358]_  = \new_[90318]_  & \new_[90303]_ ;
  assign \new_[359]_  = \new_[90288]_  & \new_[90273]_ ;
  assign \new_[360]_  = \new_[90258]_  & \new_[90243]_ ;
  assign \new_[361]_  = \new_[90228]_  & \new_[90213]_ ;
  assign \new_[362]_  = \new_[90198]_  & \new_[90183]_ ;
  assign \new_[363]_  = \new_[90168]_  & \new_[90153]_ ;
  assign \new_[364]_  = \new_[90138]_  & \new_[90123]_ ;
  assign \new_[365]_  = \new_[90108]_  & \new_[90093]_ ;
  assign \new_[366]_  = \new_[90078]_  & \new_[90063]_ ;
  assign \new_[367]_  = \new_[90048]_  & \new_[90033]_ ;
  assign \new_[368]_  = \new_[90018]_  & \new_[90003]_ ;
  assign \new_[369]_  = \new_[89988]_  & \new_[89973]_ ;
  assign \new_[370]_  = \new_[89958]_  & \new_[89943]_ ;
  assign \new_[371]_  = \new_[89928]_  & \new_[89913]_ ;
  assign \new_[372]_  = \new_[89898]_  & \new_[89883]_ ;
  assign \new_[373]_  = \new_[89868]_  & \new_[89853]_ ;
  assign \new_[374]_  = \new_[89838]_  & \new_[89823]_ ;
  assign \new_[375]_  = \new_[89808]_  & \new_[89793]_ ;
  assign \new_[376]_  = \new_[89778]_  & \new_[89763]_ ;
  assign \new_[377]_  = \new_[89748]_  & \new_[89733]_ ;
  assign \new_[378]_  = \new_[89718]_  & \new_[89703]_ ;
  assign \new_[379]_  = \new_[89688]_  & \new_[89673]_ ;
  assign \new_[380]_  = \new_[89658]_  & \new_[89643]_ ;
  assign \new_[381]_  = \new_[89628]_  & \new_[89613]_ ;
  assign \new_[382]_  = \new_[89598]_  & \new_[89583]_ ;
  assign \new_[383]_  = \new_[89568]_  & \new_[89553]_ ;
  assign \new_[384]_  = \new_[89538]_  & \new_[89523]_ ;
  assign \new_[385]_  = \new_[89508]_  & \new_[89493]_ ;
  assign \new_[386]_  = \new_[89480]_  & \new_[89465]_ ;
  assign \new_[387]_  = \new_[89452]_  & \new_[89437]_ ;
  assign \new_[388]_  = \new_[89424]_  & \new_[89409]_ ;
  assign \new_[389]_  = \new_[89396]_  & \new_[89381]_ ;
  assign \new_[390]_  = \new_[89368]_  & \new_[89353]_ ;
  assign \new_[391]_  = \new_[89340]_  & \new_[89325]_ ;
  assign \new_[392]_  = \new_[89312]_  & \new_[89297]_ ;
  assign \new_[393]_  = \new_[89284]_  & \new_[89269]_ ;
  assign \new_[394]_  = \new_[89256]_  & \new_[89241]_ ;
  assign \new_[395]_  = \new_[89228]_  & \new_[89213]_ ;
  assign \new_[396]_  = \new_[89200]_  & \new_[89185]_ ;
  assign \new_[397]_  = \new_[89172]_  & \new_[89157]_ ;
  assign \new_[398]_  = \new_[89144]_  & \new_[89129]_ ;
  assign \new_[399]_  = \new_[89116]_  & \new_[89101]_ ;
  assign \new_[400]_  = \new_[89088]_  & \new_[89073]_ ;
  assign \new_[401]_  = \new_[89060]_  & \new_[89045]_ ;
  assign \new_[402]_  = \new_[89032]_  & \new_[89017]_ ;
  assign \new_[403]_  = \new_[89004]_  & \new_[88989]_ ;
  assign \new_[404]_  = \new_[88976]_  & \new_[88961]_ ;
  assign \new_[405]_  = \new_[88948]_  & \new_[88933]_ ;
  assign \new_[406]_  = \new_[88920]_  & \new_[88905]_ ;
  assign \new_[407]_  = \new_[88892]_  & \new_[88877]_ ;
  assign \new_[408]_  = \new_[88864]_  & \new_[88849]_ ;
  assign \new_[409]_  = \new_[88836]_  & \new_[88821]_ ;
  assign \new_[410]_  = \new_[88808]_  & \new_[88793]_ ;
  assign \new_[411]_  = \new_[88780]_  & \new_[88765]_ ;
  assign \new_[412]_  = \new_[88752]_  & \new_[88737]_ ;
  assign \new_[413]_  = \new_[88724]_  & \new_[88709]_ ;
  assign \new_[414]_  = \new_[88696]_  & \new_[88681]_ ;
  assign \new_[415]_  = \new_[88668]_  & \new_[88653]_ ;
  assign \new_[416]_  = \new_[88640]_  & \new_[88625]_ ;
  assign \new_[417]_  = \new_[88612]_  & \new_[88597]_ ;
  assign \new_[418]_  = \new_[88584]_  & \new_[88569]_ ;
  assign \new_[419]_  = \new_[88556]_  & \new_[88541]_ ;
  assign \new_[420]_  = \new_[88528]_  & \new_[88513]_ ;
  assign \new_[421]_  = \new_[88500]_  & \new_[88485]_ ;
  assign \new_[422]_  = \new_[88472]_  & \new_[88457]_ ;
  assign \new_[423]_  = \new_[88444]_  & \new_[88429]_ ;
  assign \new_[424]_  = \new_[88416]_  & \new_[88401]_ ;
  assign \new_[425]_  = \new_[88388]_  & \new_[88373]_ ;
  assign \new_[426]_  = \new_[88360]_  & \new_[88345]_ ;
  assign \new_[427]_  = \new_[88332]_  & \new_[88317]_ ;
  assign \new_[428]_  = \new_[88304]_  & \new_[88289]_ ;
  assign \new_[429]_  = \new_[88276]_  & \new_[88261]_ ;
  assign \new_[430]_  = \new_[88248]_  & \new_[88233]_ ;
  assign \new_[431]_  = \new_[88220]_  & \new_[88205]_ ;
  assign \new_[432]_  = \new_[88192]_  & \new_[88177]_ ;
  assign \new_[433]_  = \new_[88164]_  & \new_[88149]_ ;
  assign \new_[434]_  = \new_[88136]_  & \new_[88121]_ ;
  assign \new_[435]_  = \new_[88108]_  & \new_[88093]_ ;
  assign \new_[436]_  = \new_[88080]_  & \new_[88065]_ ;
  assign \new_[437]_  = \new_[88052]_  & \new_[88037]_ ;
  assign \new_[438]_  = \new_[88024]_  & \new_[88009]_ ;
  assign \new_[439]_  = \new_[87996]_  & \new_[87981]_ ;
  assign \new_[440]_  = \new_[87968]_  & \new_[87953]_ ;
  assign \new_[441]_  = \new_[87940]_  & \new_[87925]_ ;
  assign \new_[442]_  = \new_[87912]_  & \new_[87897]_ ;
  assign \new_[443]_  = \new_[87884]_  & \new_[87869]_ ;
  assign \new_[444]_  = \new_[87856]_  & \new_[87841]_ ;
  assign \new_[445]_  = \new_[87828]_  & \new_[87813]_ ;
  assign \new_[446]_  = \new_[87800]_  & \new_[87785]_ ;
  assign \new_[447]_  = \new_[87772]_  & \new_[87757]_ ;
  assign \new_[448]_  = \new_[87744]_  & \new_[87729]_ ;
  assign \new_[449]_  = \new_[87716]_  & \new_[87701]_ ;
  assign \new_[450]_  = \new_[87688]_  & \new_[87673]_ ;
  assign \new_[451]_  = \new_[87660]_  & \new_[87645]_ ;
  assign \new_[452]_  = \new_[87632]_  & \new_[87617]_ ;
  assign \new_[453]_  = \new_[87604]_  & \new_[87589]_ ;
  assign \new_[454]_  = \new_[87576]_  & \new_[87561]_ ;
  assign \new_[455]_  = \new_[87548]_  & \new_[87533]_ ;
  assign \new_[456]_  = \new_[87520]_  & \new_[87505]_ ;
  assign \new_[457]_  = \new_[87492]_  & \new_[87477]_ ;
  assign \new_[458]_  = \new_[87464]_  & \new_[87449]_ ;
  assign \new_[459]_  = \new_[87436]_  & \new_[87421]_ ;
  assign \new_[460]_  = \new_[87408]_  & \new_[87393]_ ;
  assign \new_[461]_  = \new_[87380]_  & \new_[87365]_ ;
  assign \new_[462]_  = \new_[87352]_  & \new_[87337]_ ;
  assign \new_[463]_  = \new_[87324]_  & \new_[87309]_ ;
  assign \new_[464]_  = \new_[87296]_  & \new_[87281]_ ;
  assign \new_[465]_  = \new_[87268]_  & \new_[87253]_ ;
  assign \new_[466]_  = \new_[87240]_  & \new_[87225]_ ;
  assign \new_[467]_  = \new_[87212]_  & \new_[87197]_ ;
  assign \new_[468]_  = \new_[87184]_  & \new_[87169]_ ;
  assign \new_[469]_  = \new_[87156]_  & \new_[87141]_ ;
  assign \new_[470]_  = \new_[87128]_  & \new_[87113]_ ;
  assign \new_[471]_  = \new_[87100]_  & \new_[87085]_ ;
  assign \new_[472]_  = \new_[87072]_  & \new_[87057]_ ;
  assign \new_[473]_  = \new_[87044]_  & \new_[87029]_ ;
  assign \new_[474]_  = \new_[87016]_  & \new_[87001]_ ;
  assign \new_[475]_  = \new_[86988]_  & \new_[86973]_ ;
  assign \new_[476]_  = \new_[86960]_  & \new_[86945]_ ;
  assign \new_[477]_  = \new_[86932]_  & \new_[86917]_ ;
  assign \new_[478]_  = \new_[86904]_  & \new_[86889]_ ;
  assign \new_[479]_  = \new_[86876]_  & \new_[86861]_ ;
  assign \new_[480]_  = \new_[86848]_  & \new_[86833]_ ;
  assign \new_[481]_  = \new_[86820]_  & \new_[86805]_ ;
  assign \new_[482]_  = \new_[86792]_  & \new_[86777]_ ;
  assign \new_[483]_  = \new_[86764]_  & \new_[86749]_ ;
  assign \new_[484]_  = \new_[86736]_  & \new_[86721]_ ;
  assign \new_[485]_  = \new_[86708]_  & \new_[86693]_ ;
  assign \new_[486]_  = \new_[86680]_  & \new_[86665]_ ;
  assign \new_[487]_  = \new_[86652]_  & \new_[86637]_ ;
  assign \new_[488]_  = \new_[86624]_  & \new_[86609]_ ;
  assign \new_[489]_  = \new_[86596]_  & \new_[86581]_ ;
  assign \new_[490]_  = \new_[86568]_  & \new_[86553]_ ;
  assign \new_[491]_  = \new_[86540]_  & \new_[86525]_ ;
  assign \new_[492]_  = \new_[86512]_  & \new_[86497]_ ;
  assign \new_[493]_  = \new_[86484]_  & \new_[86469]_ ;
  assign \new_[494]_  = \new_[86456]_  & \new_[86441]_ ;
  assign \new_[495]_  = \new_[86428]_  & \new_[86413]_ ;
  assign \new_[496]_  = \new_[86400]_  & \new_[86385]_ ;
  assign \new_[497]_  = \new_[86372]_  & \new_[86357]_ ;
  assign \new_[498]_  = \new_[86344]_  & \new_[86329]_ ;
  assign \new_[499]_  = \new_[86316]_  & \new_[86301]_ ;
  assign \new_[500]_  = \new_[86288]_  & \new_[86273]_ ;
  assign \new_[501]_  = \new_[86260]_  & \new_[86245]_ ;
  assign \new_[502]_  = \new_[86232]_  & \new_[86217]_ ;
  assign \new_[503]_  = \new_[86204]_  & \new_[86189]_ ;
  assign \new_[504]_  = \new_[86176]_  & \new_[86161]_ ;
  assign \new_[505]_  = \new_[86148]_  & \new_[86133]_ ;
  assign \new_[506]_  = \new_[86120]_  & \new_[86105]_ ;
  assign \new_[507]_  = \new_[86092]_  & \new_[86077]_ ;
  assign \new_[508]_  = \new_[86064]_  & \new_[86049]_ ;
  assign \new_[509]_  = \new_[86036]_  & \new_[86021]_ ;
  assign \new_[510]_  = \new_[86008]_  & \new_[85993]_ ;
  assign \new_[511]_  = \new_[85980]_  & \new_[85965]_ ;
  assign \new_[512]_  = \new_[85952]_  & \new_[85937]_ ;
  assign \new_[513]_  = \new_[85924]_  & \new_[85909]_ ;
  assign \new_[514]_  = \new_[85896]_  & \new_[85881]_ ;
  assign \new_[515]_  = \new_[85868]_  & \new_[85853]_ ;
  assign \new_[516]_  = \new_[85840]_  & \new_[85825]_ ;
  assign \new_[517]_  = \new_[85812]_  & \new_[85797]_ ;
  assign \new_[518]_  = \new_[85784]_  & \new_[85769]_ ;
  assign \new_[519]_  = \new_[85756]_  & \new_[85741]_ ;
  assign \new_[520]_  = \new_[85728]_  & \new_[85713]_ ;
  assign \new_[521]_  = \new_[85700]_  & \new_[85685]_ ;
  assign \new_[522]_  = \new_[85672]_  & \new_[85657]_ ;
  assign \new_[523]_  = \new_[85644]_  & \new_[85629]_ ;
  assign \new_[524]_  = \new_[85616]_  & \new_[85601]_ ;
  assign \new_[525]_  = \new_[85588]_  & \new_[85573]_ ;
  assign \new_[526]_  = \new_[85560]_  & \new_[85545]_ ;
  assign \new_[527]_  = \new_[85532]_  & \new_[85517]_ ;
  assign \new_[528]_  = \new_[85504]_  & \new_[85489]_ ;
  assign \new_[529]_  = \new_[85476]_  & \new_[85461]_ ;
  assign \new_[530]_  = \new_[85448]_  & \new_[85433]_ ;
  assign \new_[531]_  = \new_[85420]_  & \new_[85405]_ ;
  assign \new_[532]_  = \new_[85392]_  & \new_[85377]_ ;
  assign \new_[533]_  = \new_[85364]_  & \new_[85349]_ ;
  assign \new_[534]_  = \new_[85336]_  & \new_[85321]_ ;
  assign \new_[535]_  = \new_[85308]_  & \new_[85293]_ ;
  assign \new_[536]_  = \new_[85280]_  & \new_[85265]_ ;
  assign \new_[537]_  = \new_[85252]_  & \new_[85237]_ ;
  assign \new_[538]_  = \new_[85224]_  & \new_[85209]_ ;
  assign \new_[539]_  = \new_[85196]_  & \new_[85181]_ ;
  assign \new_[540]_  = \new_[85168]_  & \new_[85153]_ ;
  assign \new_[541]_  = \new_[85140]_  & \new_[85125]_ ;
  assign \new_[542]_  = \new_[85112]_  & \new_[85097]_ ;
  assign \new_[543]_  = \new_[85084]_  & \new_[85069]_ ;
  assign \new_[544]_  = \new_[85056]_  & \new_[85041]_ ;
  assign \new_[545]_  = \new_[85028]_  & \new_[85013]_ ;
  assign \new_[546]_  = \new_[85000]_  & \new_[84985]_ ;
  assign \new_[547]_  = \new_[84972]_  & \new_[84957]_ ;
  assign \new_[548]_  = \new_[84944]_  & \new_[84929]_ ;
  assign \new_[549]_  = \new_[84916]_  & \new_[84901]_ ;
  assign \new_[550]_  = \new_[84888]_  & \new_[84873]_ ;
  assign \new_[551]_  = \new_[84860]_  & \new_[84845]_ ;
  assign \new_[552]_  = \new_[84832]_  & \new_[84817]_ ;
  assign \new_[553]_  = \new_[84804]_  & \new_[84789]_ ;
  assign \new_[554]_  = \new_[84776]_  & \new_[84761]_ ;
  assign \new_[555]_  = \new_[84748]_  & \new_[84733]_ ;
  assign \new_[556]_  = \new_[84720]_  & \new_[84705]_ ;
  assign \new_[557]_  = \new_[84692]_  & \new_[84677]_ ;
  assign \new_[558]_  = \new_[84664]_  & \new_[84649]_ ;
  assign \new_[559]_  = \new_[84636]_  & \new_[84621]_ ;
  assign \new_[560]_  = \new_[84608]_  & \new_[84593]_ ;
  assign \new_[561]_  = \new_[84580]_  & \new_[84565]_ ;
  assign \new_[562]_  = \new_[84552]_  & \new_[84537]_ ;
  assign \new_[563]_  = \new_[84524]_  & \new_[84509]_ ;
  assign \new_[564]_  = \new_[84496]_  & \new_[84481]_ ;
  assign \new_[565]_  = \new_[84468]_  & \new_[84453]_ ;
  assign \new_[566]_  = \new_[84440]_  & \new_[84425]_ ;
  assign \new_[567]_  = \new_[84412]_  & \new_[84397]_ ;
  assign \new_[568]_  = \new_[84384]_  & \new_[84369]_ ;
  assign \new_[569]_  = \new_[84356]_  & \new_[84341]_ ;
  assign \new_[570]_  = \new_[84328]_  & \new_[84313]_ ;
  assign \new_[571]_  = \new_[84300]_  & \new_[84285]_ ;
  assign \new_[572]_  = \new_[84272]_  & \new_[84257]_ ;
  assign \new_[573]_  = \new_[84244]_  & \new_[84229]_ ;
  assign \new_[574]_  = \new_[84216]_  & \new_[84201]_ ;
  assign \new_[575]_  = \new_[84188]_  & \new_[84173]_ ;
  assign \new_[576]_  = \new_[84160]_  & \new_[84145]_ ;
  assign \new_[577]_  = \new_[84132]_  & \new_[84117]_ ;
  assign \new_[578]_  = \new_[84104]_  & \new_[84089]_ ;
  assign \new_[579]_  = \new_[84076]_  & \new_[84061]_ ;
  assign \new_[580]_  = \new_[84048]_  & \new_[84033]_ ;
  assign \new_[581]_  = \new_[84020]_  & \new_[84005]_ ;
  assign \new_[582]_  = \new_[83992]_  & \new_[83977]_ ;
  assign \new_[583]_  = \new_[83964]_  & \new_[83949]_ ;
  assign \new_[584]_  = \new_[83936]_  & \new_[83921]_ ;
  assign \new_[585]_  = \new_[83908]_  & \new_[83893]_ ;
  assign \new_[586]_  = \new_[83880]_  & \new_[83865]_ ;
  assign \new_[587]_  = \new_[83852]_  & \new_[83837]_ ;
  assign \new_[588]_  = \new_[83824]_  & \new_[83809]_ ;
  assign \new_[589]_  = \new_[83796]_  & \new_[83781]_ ;
  assign \new_[590]_  = \new_[83768]_  & \new_[83753]_ ;
  assign \new_[591]_  = \new_[83740]_  & \new_[83725]_ ;
  assign \new_[592]_  = \new_[83712]_  & \new_[83697]_ ;
  assign \new_[593]_  = \new_[83684]_  & \new_[83669]_ ;
  assign \new_[594]_  = \new_[83656]_  & \new_[83641]_ ;
  assign \new_[595]_  = \new_[83628]_  & \new_[83613]_ ;
  assign \new_[596]_  = \new_[83600]_  & \new_[83585]_ ;
  assign \new_[597]_  = \new_[83572]_  & \new_[83557]_ ;
  assign \new_[598]_  = \new_[83544]_  & \new_[83529]_ ;
  assign \new_[599]_  = \new_[83516]_  & \new_[83501]_ ;
  assign \new_[600]_  = \new_[83488]_  & \new_[83473]_ ;
  assign \new_[601]_  = \new_[83460]_  & \new_[83445]_ ;
  assign \new_[602]_  = \new_[83432]_  & \new_[83417]_ ;
  assign \new_[603]_  = \new_[83404]_  & \new_[83389]_ ;
  assign \new_[604]_  = \new_[83376]_  & \new_[83361]_ ;
  assign \new_[605]_  = \new_[83348]_  & \new_[83333]_ ;
  assign \new_[606]_  = \new_[83320]_  & \new_[83305]_ ;
  assign \new_[607]_  = \new_[83292]_  & \new_[83277]_ ;
  assign \new_[608]_  = \new_[83264]_  & \new_[83249]_ ;
  assign \new_[609]_  = \new_[83236]_  & \new_[83221]_ ;
  assign \new_[610]_  = \new_[83208]_  & \new_[83193]_ ;
  assign \new_[611]_  = \new_[83180]_  & \new_[83165]_ ;
  assign \new_[612]_  = \new_[83152]_  & \new_[83137]_ ;
  assign \new_[613]_  = \new_[83124]_  & \new_[83109]_ ;
  assign \new_[614]_  = \new_[83096]_  & \new_[83081]_ ;
  assign \new_[615]_  = \new_[83068]_  & \new_[83053]_ ;
  assign \new_[616]_  = \new_[83040]_  & \new_[83025]_ ;
  assign \new_[617]_  = \new_[83012]_  & \new_[82997]_ ;
  assign \new_[618]_  = \new_[82984]_  & \new_[82969]_ ;
  assign \new_[619]_  = \new_[82956]_  & \new_[82941]_ ;
  assign \new_[620]_  = \new_[82928]_  & \new_[82913]_ ;
  assign \new_[621]_  = \new_[82900]_  & \new_[82885]_ ;
  assign \new_[622]_  = \new_[82872]_  & \new_[82857]_ ;
  assign \new_[623]_  = \new_[82844]_  & \new_[82829]_ ;
  assign \new_[624]_  = \new_[82816]_  & \new_[82801]_ ;
  assign \new_[625]_  = \new_[82788]_  & \new_[82773]_ ;
  assign \new_[626]_  = \new_[82760]_  & \new_[82745]_ ;
  assign \new_[627]_  = \new_[82732]_  & \new_[82717]_ ;
  assign \new_[628]_  = \new_[82704]_  & \new_[82689]_ ;
  assign \new_[629]_  = \new_[82676]_  & \new_[82661]_ ;
  assign \new_[630]_  = \new_[82648]_  & \new_[82633]_ ;
  assign \new_[631]_  = \new_[82620]_  & \new_[82605]_ ;
  assign \new_[632]_  = \new_[82592]_  & \new_[82577]_ ;
  assign \new_[633]_  = \new_[82564]_  & \new_[82549]_ ;
  assign \new_[634]_  = \new_[82536]_  & \new_[82521]_ ;
  assign \new_[635]_  = \new_[82508]_  & \new_[82493]_ ;
  assign \new_[636]_  = \new_[82480]_  & \new_[82465]_ ;
  assign \new_[637]_  = \new_[82452]_  & \new_[82437]_ ;
  assign \new_[638]_  = \new_[82424]_  & \new_[82409]_ ;
  assign \new_[639]_  = \new_[82396]_  & \new_[82381]_ ;
  assign \new_[640]_  = \new_[82368]_  & \new_[82353]_ ;
  assign \new_[641]_  = \new_[82340]_  & \new_[82325]_ ;
  assign \new_[642]_  = \new_[82312]_  & \new_[82297]_ ;
  assign \new_[643]_  = \new_[82284]_  & \new_[82269]_ ;
  assign \new_[644]_  = \new_[82256]_  & \new_[82241]_ ;
  assign \new_[645]_  = \new_[82228]_  & \new_[82213]_ ;
  assign \new_[646]_  = \new_[82200]_  & \new_[82185]_ ;
  assign \new_[647]_  = \new_[82172]_  & \new_[82157]_ ;
  assign \new_[648]_  = \new_[82144]_  & \new_[82129]_ ;
  assign \new_[649]_  = \new_[82116]_  & \new_[82101]_ ;
  assign \new_[650]_  = \new_[82088]_  & \new_[82073]_ ;
  assign \new_[651]_  = \new_[82060]_  & \new_[82045]_ ;
  assign \new_[652]_  = \new_[82032]_  & \new_[82017]_ ;
  assign \new_[653]_  = \new_[82004]_  & \new_[81989]_ ;
  assign \new_[654]_  = \new_[81976]_  & \new_[81961]_ ;
  assign \new_[655]_  = \new_[81948]_  & \new_[81933]_ ;
  assign \new_[656]_  = \new_[81920]_  & \new_[81905]_ ;
  assign \new_[657]_  = \new_[81892]_  & \new_[81877]_ ;
  assign \new_[658]_  = \new_[81864]_  & \new_[81849]_ ;
  assign \new_[659]_  = \new_[81836]_  & \new_[81821]_ ;
  assign \new_[660]_  = \new_[81808]_  & \new_[81793]_ ;
  assign \new_[661]_  = \new_[81780]_  & \new_[81765]_ ;
  assign \new_[662]_  = \new_[81752]_  & \new_[81737]_ ;
  assign \new_[663]_  = \new_[81724]_  & \new_[81709]_ ;
  assign \new_[664]_  = \new_[81696]_  & \new_[81681]_ ;
  assign \new_[665]_  = \new_[81668]_  & \new_[81653]_ ;
  assign \new_[666]_  = \new_[81640]_  & \new_[81625]_ ;
  assign \new_[667]_  = \new_[81612]_  & \new_[81597]_ ;
  assign \new_[668]_  = \new_[81584]_  & \new_[81569]_ ;
  assign \new_[669]_  = \new_[81556]_  & \new_[81541]_ ;
  assign \new_[670]_  = \new_[81528]_  & \new_[81513]_ ;
  assign \new_[671]_  = \new_[81500]_  & \new_[81485]_ ;
  assign \new_[672]_  = \new_[81472]_  & \new_[81457]_ ;
  assign \new_[673]_  = \new_[81444]_  & \new_[81429]_ ;
  assign \new_[674]_  = \new_[81416]_  & \new_[81401]_ ;
  assign \new_[675]_  = \new_[81388]_  & \new_[81373]_ ;
  assign \new_[676]_  = \new_[81360]_  & \new_[81345]_ ;
  assign \new_[677]_  = \new_[81332]_  & \new_[81317]_ ;
  assign \new_[678]_  = \new_[81304]_  & \new_[81289]_ ;
  assign \new_[679]_  = \new_[81276]_  & \new_[81261]_ ;
  assign \new_[680]_  = \new_[81248]_  & \new_[81233]_ ;
  assign \new_[681]_  = \new_[81220]_  & \new_[81205]_ ;
  assign \new_[682]_  = \new_[81192]_  & \new_[81177]_ ;
  assign \new_[683]_  = \new_[81164]_  & \new_[81149]_ ;
  assign \new_[684]_  = \new_[81136]_  & \new_[81121]_ ;
  assign \new_[685]_  = \new_[81108]_  & \new_[81093]_ ;
  assign \new_[686]_  = \new_[81080]_  & \new_[81065]_ ;
  assign \new_[687]_  = \new_[81052]_  & \new_[81037]_ ;
  assign \new_[688]_  = \new_[81024]_  & \new_[81009]_ ;
  assign \new_[689]_  = \new_[80996]_  & \new_[80981]_ ;
  assign \new_[690]_  = \new_[80968]_  & \new_[80953]_ ;
  assign \new_[691]_  = \new_[80940]_  & \new_[80925]_ ;
  assign \new_[692]_  = \new_[80912]_  & \new_[80897]_ ;
  assign \new_[693]_  = \new_[80884]_  & \new_[80869]_ ;
  assign \new_[694]_  = \new_[80856]_  & \new_[80841]_ ;
  assign \new_[695]_  = \new_[80828]_  & \new_[80813]_ ;
  assign \new_[696]_  = \new_[80800]_  & \new_[80785]_ ;
  assign \new_[697]_  = \new_[80772]_  & \new_[80757]_ ;
  assign \new_[698]_  = \new_[80744]_  & \new_[80729]_ ;
  assign \new_[699]_  = \new_[80716]_  & \new_[80701]_ ;
  assign \new_[700]_  = \new_[80688]_  & \new_[80673]_ ;
  assign \new_[701]_  = \new_[80660]_  & \new_[80645]_ ;
  assign \new_[702]_  = \new_[80632]_  & \new_[80617]_ ;
  assign \new_[703]_  = \new_[80604]_  & \new_[80589]_ ;
  assign \new_[704]_  = \new_[80576]_  & \new_[80561]_ ;
  assign \new_[705]_  = \new_[80548]_  & \new_[80533]_ ;
  assign \new_[706]_  = \new_[80520]_  & \new_[80505]_ ;
  assign \new_[707]_  = \new_[80492]_  & \new_[80477]_ ;
  assign \new_[708]_  = \new_[80464]_  & \new_[80449]_ ;
  assign \new_[709]_  = \new_[80436]_  & \new_[80421]_ ;
  assign \new_[710]_  = \new_[80408]_  & \new_[80393]_ ;
  assign \new_[711]_  = \new_[80380]_  & \new_[80365]_ ;
  assign \new_[712]_  = \new_[80352]_  & \new_[80337]_ ;
  assign \new_[713]_  = \new_[80324]_  & \new_[80309]_ ;
  assign \new_[714]_  = \new_[80296]_  & \new_[80281]_ ;
  assign \new_[715]_  = \new_[80268]_  & \new_[80253]_ ;
  assign \new_[716]_  = \new_[80240]_  & \new_[80225]_ ;
  assign \new_[717]_  = \new_[80212]_  & \new_[80197]_ ;
  assign \new_[718]_  = \new_[80184]_  & \new_[80169]_ ;
  assign \new_[719]_  = \new_[80156]_  & \new_[80141]_ ;
  assign \new_[720]_  = \new_[80128]_  & \new_[80113]_ ;
  assign \new_[721]_  = \new_[80100]_  & \new_[80085]_ ;
  assign \new_[722]_  = \new_[80072]_  & \new_[80057]_ ;
  assign \new_[723]_  = \new_[80044]_  & \new_[80029]_ ;
  assign \new_[724]_  = \new_[80016]_  & \new_[80001]_ ;
  assign \new_[725]_  = \new_[79988]_  & \new_[79973]_ ;
  assign \new_[726]_  = \new_[79960]_  & \new_[79945]_ ;
  assign \new_[727]_  = \new_[79932]_  & \new_[79917]_ ;
  assign \new_[728]_  = \new_[79904]_  & \new_[79889]_ ;
  assign \new_[729]_  = \new_[79876]_  & \new_[79861]_ ;
  assign \new_[730]_  = \new_[79848]_  & \new_[79833]_ ;
  assign \new_[731]_  = \new_[79820]_  & \new_[79805]_ ;
  assign \new_[732]_  = \new_[79792]_  & \new_[79777]_ ;
  assign \new_[733]_  = \new_[79764]_  & \new_[79749]_ ;
  assign \new_[734]_  = \new_[79736]_  & \new_[79721]_ ;
  assign \new_[735]_  = \new_[79708]_  & \new_[79693]_ ;
  assign \new_[736]_  = \new_[79680]_  & \new_[79665]_ ;
  assign \new_[737]_  = \new_[79652]_  & \new_[79637]_ ;
  assign \new_[738]_  = \new_[79624]_  & \new_[79609]_ ;
  assign \new_[739]_  = \new_[79596]_  & \new_[79581]_ ;
  assign \new_[740]_  = \new_[79568]_  & \new_[79553]_ ;
  assign \new_[741]_  = \new_[79540]_  & \new_[79525]_ ;
  assign \new_[742]_  = \new_[79512]_  & \new_[79497]_ ;
  assign \new_[743]_  = \new_[79484]_  & \new_[79469]_ ;
  assign \new_[744]_  = \new_[79456]_  & \new_[79441]_ ;
  assign \new_[745]_  = \new_[79428]_  & \new_[79413]_ ;
  assign \new_[746]_  = \new_[79400]_  & \new_[79385]_ ;
  assign \new_[747]_  = \new_[79372]_  & \new_[79357]_ ;
  assign \new_[748]_  = \new_[79344]_  & \new_[79329]_ ;
  assign \new_[749]_  = \new_[79316]_  & \new_[79301]_ ;
  assign \new_[750]_  = \new_[79288]_  & \new_[79273]_ ;
  assign \new_[751]_  = \new_[79260]_  & \new_[79245]_ ;
  assign \new_[752]_  = \new_[79232]_  & \new_[79217]_ ;
  assign \new_[753]_  = \new_[79204]_  & \new_[79189]_ ;
  assign \new_[754]_  = \new_[79176]_  & \new_[79161]_ ;
  assign \new_[755]_  = \new_[79148]_  & \new_[79133]_ ;
  assign \new_[756]_  = \new_[79120]_  & \new_[79105]_ ;
  assign \new_[757]_  = \new_[79092]_  & \new_[79077]_ ;
  assign \new_[758]_  = \new_[79064]_  & \new_[79049]_ ;
  assign \new_[759]_  = \new_[79036]_  & \new_[79021]_ ;
  assign \new_[760]_  = \new_[79008]_  & \new_[78993]_ ;
  assign \new_[761]_  = \new_[78980]_  & \new_[78965]_ ;
  assign \new_[762]_  = \new_[78952]_  & \new_[78937]_ ;
  assign \new_[763]_  = \new_[78924]_  & \new_[78909]_ ;
  assign \new_[764]_  = \new_[78896]_  & \new_[78881]_ ;
  assign \new_[765]_  = \new_[78868]_  & \new_[78853]_ ;
  assign \new_[766]_  = \new_[78840]_  & \new_[78825]_ ;
  assign \new_[767]_  = \new_[78812]_  & \new_[78797]_ ;
  assign \new_[768]_  = \new_[78784]_  & \new_[78769]_ ;
  assign \new_[769]_  = \new_[78756]_  & \new_[78741]_ ;
  assign \new_[770]_  = \new_[78728]_  & \new_[78713]_ ;
  assign \new_[771]_  = \new_[78700]_  & \new_[78685]_ ;
  assign \new_[772]_  = \new_[78672]_  & \new_[78657]_ ;
  assign \new_[773]_  = \new_[78644]_  & \new_[78629]_ ;
  assign \new_[774]_  = \new_[78616]_  & \new_[78601]_ ;
  assign \new_[775]_  = \new_[78588]_  & \new_[78573]_ ;
  assign \new_[776]_  = \new_[78560]_  & \new_[78545]_ ;
  assign \new_[777]_  = \new_[78532]_  & \new_[78517]_ ;
  assign \new_[778]_  = \new_[78504]_  & \new_[78489]_ ;
  assign \new_[779]_  = \new_[78476]_  & \new_[78461]_ ;
  assign \new_[780]_  = \new_[78448]_  & \new_[78433]_ ;
  assign \new_[781]_  = \new_[78420]_  & \new_[78405]_ ;
  assign \new_[782]_  = \new_[78392]_  & \new_[78377]_ ;
  assign \new_[783]_  = \new_[78364]_  & \new_[78349]_ ;
  assign \new_[784]_  = \new_[78336]_  & \new_[78321]_ ;
  assign \new_[785]_  = \new_[78308]_  & \new_[78293]_ ;
  assign \new_[786]_  = \new_[78280]_  & \new_[78265]_ ;
  assign \new_[787]_  = \new_[78252]_  & \new_[78237]_ ;
  assign \new_[788]_  = \new_[78224]_  & \new_[78209]_ ;
  assign \new_[789]_  = \new_[78196]_  & \new_[78181]_ ;
  assign \new_[790]_  = \new_[78168]_  & \new_[78153]_ ;
  assign \new_[791]_  = \new_[78140]_  & \new_[78125]_ ;
  assign \new_[792]_  = \new_[78112]_  & \new_[78097]_ ;
  assign \new_[793]_  = \new_[78084]_  & \new_[78069]_ ;
  assign \new_[794]_  = \new_[78056]_  & \new_[78041]_ ;
  assign \new_[795]_  = \new_[78028]_  & \new_[78013]_ ;
  assign \new_[796]_  = \new_[78000]_  & \new_[77985]_ ;
  assign \new_[797]_  = \new_[77972]_  & \new_[77957]_ ;
  assign \new_[798]_  = \new_[77944]_  & \new_[77929]_ ;
  assign \new_[799]_  = \new_[77916]_  & \new_[77901]_ ;
  assign \new_[800]_  = \new_[77888]_  & \new_[77873]_ ;
  assign \new_[801]_  = \new_[77860]_  & \new_[77845]_ ;
  assign \new_[802]_  = \new_[77832]_  & \new_[77817]_ ;
  assign \new_[803]_  = \new_[77804]_  & \new_[77789]_ ;
  assign \new_[804]_  = \new_[77776]_  & \new_[77761]_ ;
  assign \new_[805]_  = \new_[77748]_  & \new_[77733]_ ;
  assign \new_[806]_  = \new_[77720]_  & \new_[77705]_ ;
  assign \new_[807]_  = \new_[77692]_  & \new_[77677]_ ;
  assign \new_[808]_  = \new_[77664]_  & \new_[77649]_ ;
  assign \new_[809]_  = \new_[77636]_  & \new_[77621]_ ;
  assign \new_[810]_  = \new_[77608]_  & \new_[77593]_ ;
  assign \new_[811]_  = \new_[77580]_  & \new_[77565]_ ;
  assign \new_[812]_  = \new_[77552]_  & \new_[77537]_ ;
  assign \new_[813]_  = \new_[77524]_  & \new_[77509]_ ;
  assign \new_[814]_  = \new_[77496]_  & \new_[77481]_ ;
  assign \new_[815]_  = \new_[77468]_  & \new_[77453]_ ;
  assign \new_[816]_  = \new_[77440]_  & \new_[77425]_ ;
  assign \new_[817]_  = \new_[77412]_  & \new_[77397]_ ;
  assign \new_[818]_  = \new_[77384]_  & \new_[77369]_ ;
  assign \new_[819]_  = \new_[77356]_  & \new_[77341]_ ;
  assign \new_[820]_  = \new_[77328]_  & \new_[77313]_ ;
  assign \new_[821]_  = \new_[77300]_  & \new_[77285]_ ;
  assign \new_[822]_  = \new_[77272]_  & \new_[77257]_ ;
  assign \new_[823]_  = \new_[77244]_  & \new_[77229]_ ;
  assign \new_[824]_  = \new_[77216]_  & \new_[77201]_ ;
  assign \new_[825]_  = \new_[77188]_  & \new_[77173]_ ;
  assign \new_[826]_  = \new_[77160]_  & \new_[77145]_ ;
  assign \new_[827]_  = \new_[77132]_  & \new_[77117]_ ;
  assign \new_[828]_  = \new_[77104]_  & \new_[77089]_ ;
  assign \new_[829]_  = \new_[77076]_  & \new_[77061]_ ;
  assign \new_[830]_  = \new_[77048]_  & \new_[77033]_ ;
  assign \new_[831]_  = \new_[77020]_  & \new_[77005]_ ;
  assign \new_[832]_  = \new_[76992]_  & \new_[76977]_ ;
  assign \new_[833]_  = \new_[76964]_  & \new_[76949]_ ;
  assign \new_[834]_  = \new_[76936]_  & \new_[76921]_ ;
  assign \new_[835]_  = \new_[76908]_  & \new_[76893]_ ;
  assign \new_[836]_  = \new_[76880]_  & \new_[76865]_ ;
  assign \new_[837]_  = \new_[76852]_  & \new_[76837]_ ;
  assign \new_[838]_  = \new_[76824]_  & \new_[76809]_ ;
  assign \new_[839]_  = \new_[76796]_  & \new_[76781]_ ;
  assign \new_[840]_  = \new_[76768]_  & \new_[76753]_ ;
  assign \new_[841]_  = \new_[76740]_  & \new_[76725]_ ;
  assign \new_[842]_  = \new_[76712]_  & \new_[76697]_ ;
  assign \new_[843]_  = \new_[76684]_  & \new_[76669]_ ;
  assign \new_[844]_  = \new_[76656]_  & \new_[76641]_ ;
  assign \new_[845]_  = \new_[76628]_  & \new_[76613]_ ;
  assign \new_[846]_  = \new_[76600]_  & \new_[76585]_ ;
  assign \new_[847]_  = \new_[76572]_  & \new_[76557]_ ;
  assign \new_[848]_  = \new_[76544]_  & \new_[76529]_ ;
  assign \new_[849]_  = \new_[76516]_  & \new_[76501]_ ;
  assign \new_[850]_  = \new_[76488]_  & \new_[76473]_ ;
  assign \new_[851]_  = \new_[76460]_  & \new_[76445]_ ;
  assign \new_[852]_  = \new_[76432]_  & \new_[76417]_ ;
  assign \new_[853]_  = \new_[76404]_  & \new_[76389]_ ;
  assign \new_[854]_  = \new_[76376]_  & \new_[76361]_ ;
  assign \new_[855]_  = \new_[76348]_  & \new_[76333]_ ;
  assign \new_[856]_  = \new_[76320]_  & \new_[76305]_ ;
  assign \new_[857]_  = \new_[76292]_  & \new_[76277]_ ;
  assign \new_[858]_  = \new_[76264]_  & \new_[76249]_ ;
  assign \new_[859]_  = \new_[76236]_  & \new_[76221]_ ;
  assign \new_[860]_  = \new_[76208]_  & \new_[76193]_ ;
  assign \new_[861]_  = \new_[76180]_  & \new_[76165]_ ;
  assign \new_[862]_  = \new_[76152]_  & \new_[76137]_ ;
  assign \new_[863]_  = \new_[76124]_  & \new_[76109]_ ;
  assign \new_[864]_  = \new_[76096]_  & \new_[76081]_ ;
  assign \new_[865]_  = \new_[76068]_  & \new_[76053]_ ;
  assign \new_[866]_  = \new_[76040]_  & \new_[76025]_ ;
  assign \new_[867]_  = \new_[76012]_  & \new_[75997]_ ;
  assign \new_[868]_  = \new_[75984]_  & \new_[75969]_ ;
  assign \new_[869]_  = \new_[75956]_  & \new_[75941]_ ;
  assign \new_[870]_  = \new_[75928]_  & \new_[75913]_ ;
  assign \new_[871]_  = \new_[75900]_  & \new_[75885]_ ;
  assign \new_[872]_  = \new_[75872]_  & \new_[75857]_ ;
  assign \new_[873]_  = \new_[75844]_  & \new_[75829]_ ;
  assign \new_[874]_  = \new_[75816]_  & \new_[75801]_ ;
  assign \new_[875]_  = \new_[75788]_  & \new_[75773]_ ;
  assign \new_[876]_  = \new_[75760]_  & \new_[75745]_ ;
  assign \new_[877]_  = \new_[75732]_  & \new_[75717]_ ;
  assign \new_[878]_  = \new_[75704]_  & \new_[75689]_ ;
  assign \new_[879]_  = \new_[75676]_  & \new_[75661]_ ;
  assign \new_[880]_  = \new_[75648]_  & \new_[75633]_ ;
  assign \new_[881]_  = \new_[75620]_  & \new_[75605]_ ;
  assign \new_[882]_  = \new_[75592]_  & \new_[75577]_ ;
  assign \new_[883]_  = \new_[75564]_  & \new_[75549]_ ;
  assign \new_[884]_  = \new_[75536]_  & \new_[75521]_ ;
  assign \new_[885]_  = \new_[75508]_  & \new_[75493]_ ;
  assign \new_[886]_  = \new_[75480]_  & \new_[75465]_ ;
  assign \new_[887]_  = \new_[75452]_  & \new_[75437]_ ;
  assign \new_[888]_  = \new_[75424]_  & \new_[75409]_ ;
  assign \new_[889]_  = \new_[75396]_  & \new_[75381]_ ;
  assign \new_[890]_  = \new_[75368]_  & \new_[75353]_ ;
  assign \new_[891]_  = \new_[75340]_  & \new_[75325]_ ;
  assign \new_[892]_  = \new_[75312]_  & \new_[75297]_ ;
  assign \new_[893]_  = \new_[75284]_  & \new_[75269]_ ;
  assign \new_[894]_  = \new_[75256]_  & \new_[75241]_ ;
  assign \new_[895]_  = \new_[75228]_  & \new_[75213]_ ;
  assign \new_[896]_  = \new_[75200]_  & \new_[75185]_ ;
  assign \new_[897]_  = \new_[75172]_  & \new_[75157]_ ;
  assign \new_[898]_  = \new_[75144]_  & \new_[75129]_ ;
  assign \new_[899]_  = \new_[75116]_  & \new_[75101]_ ;
  assign \new_[900]_  = \new_[75088]_  & \new_[75073]_ ;
  assign \new_[901]_  = \new_[75060]_  & \new_[75045]_ ;
  assign \new_[902]_  = \new_[75032]_  & \new_[75017]_ ;
  assign \new_[903]_  = \new_[75004]_  & \new_[74989]_ ;
  assign \new_[904]_  = \new_[74976]_  & \new_[74961]_ ;
  assign \new_[905]_  = \new_[74948]_  & \new_[74933]_ ;
  assign \new_[906]_  = \new_[74920]_  & \new_[74905]_ ;
  assign \new_[907]_  = \new_[74892]_  & \new_[74877]_ ;
  assign \new_[908]_  = \new_[74864]_  & \new_[74849]_ ;
  assign \new_[909]_  = \new_[74836]_  & \new_[74821]_ ;
  assign \new_[910]_  = \new_[74808]_  & \new_[74793]_ ;
  assign \new_[911]_  = \new_[74780]_  & \new_[74765]_ ;
  assign \new_[912]_  = \new_[74752]_  & \new_[74737]_ ;
  assign \new_[913]_  = \new_[74724]_  & \new_[74709]_ ;
  assign \new_[914]_  = \new_[74696]_  & \new_[74681]_ ;
  assign \new_[915]_  = \new_[74668]_  & \new_[74653]_ ;
  assign \new_[916]_  = \new_[74640]_  & \new_[74625]_ ;
  assign \new_[917]_  = \new_[74612]_  & \new_[74597]_ ;
  assign \new_[918]_  = \new_[74584]_  & \new_[74569]_ ;
  assign \new_[919]_  = \new_[74556]_  & \new_[74541]_ ;
  assign \new_[920]_  = \new_[74528]_  & \new_[74513]_ ;
  assign \new_[921]_  = \new_[74500]_  & \new_[74485]_ ;
  assign \new_[922]_  = \new_[74472]_  & \new_[74457]_ ;
  assign \new_[923]_  = \new_[74444]_  & \new_[74429]_ ;
  assign \new_[924]_  = \new_[74416]_  & \new_[74401]_ ;
  assign \new_[925]_  = \new_[74388]_  & \new_[74373]_ ;
  assign \new_[926]_  = \new_[74360]_  & \new_[74345]_ ;
  assign \new_[927]_  = \new_[74332]_  & \new_[74317]_ ;
  assign \new_[928]_  = \new_[74304]_  & \new_[74289]_ ;
  assign \new_[929]_  = \new_[74276]_  & \new_[74263]_ ;
  assign \new_[930]_  = \new_[74250]_  & \new_[74237]_ ;
  assign \new_[931]_  = \new_[74224]_  & \new_[74211]_ ;
  assign \new_[932]_  = \new_[74198]_  & \new_[74185]_ ;
  assign \new_[933]_  = \new_[74172]_  & \new_[74159]_ ;
  assign \new_[934]_  = \new_[74146]_  & \new_[74133]_ ;
  assign \new_[935]_  = \new_[74120]_  & \new_[74107]_ ;
  assign \new_[936]_  = \new_[74094]_  & \new_[74081]_ ;
  assign \new_[937]_  = \new_[74068]_  & \new_[74055]_ ;
  assign \new_[938]_  = \new_[74042]_  & \new_[74029]_ ;
  assign \new_[939]_  = \new_[74016]_  & \new_[74003]_ ;
  assign \new_[940]_  = \new_[73990]_  & \new_[73977]_ ;
  assign \new_[941]_  = \new_[73964]_  & \new_[73951]_ ;
  assign \new_[942]_  = \new_[73938]_  & \new_[73925]_ ;
  assign \new_[943]_  = \new_[73912]_  & \new_[73899]_ ;
  assign \new_[944]_  = \new_[73886]_  & \new_[73873]_ ;
  assign \new_[945]_  = \new_[73860]_  & \new_[73847]_ ;
  assign \new_[946]_  = \new_[73834]_  & \new_[73821]_ ;
  assign \new_[947]_  = \new_[73808]_  & \new_[73795]_ ;
  assign \new_[948]_  = \new_[73782]_  & \new_[73769]_ ;
  assign \new_[949]_  = \new_[73756]_  & \new_[73743]_ ;
  assign \new_[950]_  = \new_[73730]_  & \new_[73717]_ ;
  assign \new_[951]_  = \new_[73704]_  & \new_[73691]_ ;
  assign \new_[952]_  = \new_[73678]_  & \new_[73665]_ ;
  assign \new_[953]_  = \new_[73652]_  & \new_[73639]_ ;
  assign \new_[954]_  = \new_[73626]_  & \new_[73613]_ ;
  assign \new_[955]_  = \new_[73600]_  & \new_[73587]_ ;
  assign \new_[956]_  = \new_[73574]_  & \new_[73561]_ ;
  assign \new_[957]_  = \new_[73548]_  & \new_[73535]_ ;
  assign \new_[958]_  = \new_[73522]_  & \new_[73509]_ ;
  assign \new_[959]_  = \new_[73496]_  & \new_[73483]_ ;
  assign \new_[960]_  = \new_[73470]_  & \new_[73457]_ ;
  assign \new_[961]_  = \new_[73444]_  & \new_[73431]_ ;
  assign \new_[962]_  = \new_[73418]_  & \new_[73405]_ ;
  assign \new_[963]_  = \new_[73392]_  & \new_[73379]_ ;
  assign \new_[964]_  = \new_[73366]_  & \new_[73353]_ ;
  assign \new_[965]_  = \new_[73340]_  & \new_[73327]_ ;
  assign \new_[966]_  = \new_[73314]_  & \new_[73301]_ ;
  assign \new_[967]_  = \new_[73288]_  & \new_[73275]_ ;
  assign \new_[968]_  = \new_[73262]_  & \new_[73249]_ ;
  assign \new_[969]_  = \new_[73236]_  & \new_[73223]_ ;
  assign \new_[970]_  = \new_[73210]_  & \new_[73197]_ ;
  assign \new_[971]_  = \new_[73184]_  & \new_[73171]_ ;
  assign \new_[972]_  = \new_[73158]_  & \new_[73145]_ ;
  assign \new_[973]_  = \new_[73132]_  & \new_[73119]_ ;
  assign \new_[974]_  = \new_[73106]_  & \new_[73093]_ ;
  assign \new_[975]_  = \new_[73080]_  & \new_[73067]_ ;
  assign \new_[976]_  = \new_[73054]_  & \new_[73041]_ ;
  assign \new_[977]_  = \new_[73028]_  & \new_[73015]_ ;
  assign \new_[978]_  = \new_[73002]_  & \new_[72989]_ ;
  assign \new_[979]_  = \new_[72976]_  & \new_[72963]_ ;
  assign \new_[980]_  = \new_[72950]_  & \new_[72937]_ ;
  assign \new_[981]_  = \new_[72924]_  & \new_[72911]_ ;
  assign \new_[982]_  = \new_[72898]_  & \new_[72885]_ ;
  assign \new_[983]_  = \new_[72872]_  & \new_[72859]_ ;
  assign \new_[984]_  = \new_[72846]_  & \new_[72833]_ ;
  assign \new_[985]_  = \new_[72820]_  & \new_[72807]_ ;
  assign \new_[986]_  = \new_[72794]_  & \new_[72781]_ ;
  assign \new_[987]_  = \new_[72768]_  & \new_[72755]_ ;
  assign \new_[988]_  = \new_[72742]_  & \new_[72729]_ ;
  assign \new_[989]_  = \new_[72716]_  & \new_[72703]_ ;
  assign \new_[990]_  = \new_[72690]_  & \new_[72677]_ ;
  assign \new_[991]_  = \new_[72664]_  & \new_[72651]_ ;
  assign \new_[992]_  = \new_[72638]_  & \new_[72625]_ ;
  assign \new_[993]_  = \new_[72612]_  & \new_[72599]_ ;
  assign \new_[994]_  = \new_[72586]_  & \new_[72573]_ ;
  assign \new_[995]_  = \new_[72560]_  & \new_[72547]_ ;
  assign \new_[996]_  = \new_[72534]_  & \new_[72521]_ ;
  assign \new_[997]_  = \new_[72508]_  & \new_[72495]_ ;
  assign \new_[998]_  = \new_[72482]_  & \new_[72469]_ ;
  assign \new_[999]_  = \new_[72456]_  & \new_[72443]_ ;
  assign \new_[1000]_  = \new_[72430]_  & \new_[72417]_ ;
  assign \new_[1001]_  = \new_[72404]_  & \new_[72391]_ ;
  assign \new_[1002]_  = \new_[72378]_  & \new_[72365]_ ;
  assign \new_[1003]_  = \new_[72352]_  & \new_[72339]_ ;
  assign \new_[1004]_  = \new_[72326]_  & \new_[72313]_ ;
  assign \new_[1005]_  = \new_[72300]_  & \new_[72287]_ ;
  assign \new_[1006]_  = \new_[72274]_  & \new_[72261]_ ;
  assign \new_[1007]_  = \new_[72248]_  & \new_[72235]_ ;
  assign \new_[1008]_  = \new_[72222]_  & \new_[72209]_ ;
  assign \new_[1009]_  = \new_[72196]_  & \new_[72183]_ ;
  assign \new_[1010]_  = \new_[72170]_  & \new_[72157]_ ;
  assign \new_[1011]_  = \new_[72144]_  & \new_[72131]_ ;
  assign \new_[1012]_  = \new_[72118]_  & \new_[72105]_ ;
  assign \new_[1013]_  = \new_[72092]_  & \new_[72079]_ ;
  assign \new_[1014]_  = \new_[72066]_  & \new_[72053]_ ;
  assign \new_[1015]_  = \new_[72040]_  & \new_[72027]_ ;
  assign \new_[1016]_  = \new_[72014]_  & \new_[72001]_ ;
  assign \new_[1017]_  = \new_[71988]_  & \new_[71975]_ ;
  assign \new_[1018]_  = \new_[71962]_  & \new_[71949]_ ;
  assign \new_[1019]_  = \new_[71936]_  & \new_[71923]_ ;
  assign \new_[1020]_  = \new_[71910]_  & \new_[71897]_ ;
  assign \new_[1021]_  = \new_[71884]_  & \new_[71871]_ ;
  assign \new_[1022]_  = \new_[71858]_  & \new_[71845]_ ;
  assign \new_[1023]_  = \new_[71832]_  & \new_[71819]_ ;
  assign \new_[1024]_  = \new_[71806]_  & \new_[71793]_ ;
  assign \new_[1025]_  = \new_[71780]_  & \new_[71767]_ ;
  assign \new_[1026]_  = \new_[71754]_  & \new_[71741]_ ;
  assign \new_[1027]_  = \new_[71728]_  & \new_[71715]_ ;
  assign \new_[1028]_  = \new_[71702]_  & \new_[71689]_ ;
  assign \new_[1029]_  = \new_[71676]_  & \new_[71663]_ ;
  assign \new_[1030]_  = \new_[71650]_  & \new_[71637]_ ;
  assign \new_[1031]_  = \new_[71624]_  & \new_[71611]_ ;
  assign \new_[1032]_  = \new_[71598]_  & \new_[71585]_ ;
  assign \new_[1033]_  = \new_[71572]_  & \new_[71559]_ ;
  assign \new_[1034]_  = \new_[71546]_  & \new_[71533]_ ;
  assign \new_[1035]_  = \new_[71520]_  & \new_[71507]_ ;
  assign \new_[1036]_  = \new_[71494]_  & \new_[71481]_ ;
  assign \new_[1037]_  = \new_[71468]_  & \new_[71455]_ ;
  assign \new_[1038]_  = \new_[71442]_  & \new_[71429]_ ;
  assign \new_[1039]_  = \new_[71416]_  & \new_[71403]_ ;
  assign \new_[1040]_  = \new_[71390]_  & \new_[71377]_ ;
  assign \new_[1041]_  = \new_[71364]_  & \new_[71351]_ ;
  assign \new_[1042]_  = \new_[71338]_  & \new_[71325]_ ;
  assign \new_[1043]_  = \new_[71312]_  & \new_[71299]_ ;
  assign \new_[1044]_  = \new_[71286]_  & \new_[71273]_ ;
  assign \new_[1045]_  = \new_[71260]_  & \new_[71247]_ ;
  assign \new_[1046]_  = \new_[71234]_  & \new_[71221]_ ;
  assign \new_[1047]_  = \new_[71208]_  & \new_[71195]_ ;
  assign \new_[1048]_  = \new_[71182]_  & \new_[71169]_ ;
  assign \new_[1049]_  = \new_[71156]_  & \new_[71143]_ ;
  assign \new_[1050]_  = \new_[71130]_  & \new_[71117]_ ;
  assign \new_[1051]_  = \new_[71104]_  & \new_[71091]_ ;
  assign \new_[1052]_  = \new_[71078]_  & \new_[71065]_ ;
  assign \new_[1053]_  = \new_[71052]_  & \new_[71039]_ ;
  assign \new_[1054]_  = \new_[71026]_  & \new_[71013]_ ;
  assign \new_[1055]_  = \new_[71000]_  & \new_[70987]_ ;
  assign \new_[1056]_  = \new_[70974]_  & \new_[70961]_ ;
  assign \new_[1057]_  = \new_[70948]_  & \new_[70935]_ ;
  assign \new_[1058]_  = \new_[70922]_  & \new_[70909]_ ;
  assign \new_[1059]_  = \new_[70896]_  & \new_[70883]_ ;
  assign \new_[1060]_  = \new_[70870]_  & \new_[70857]_ ;
  assign \new_[1061]_  = \new_[70844]_  & \new_[70831]_ ;
  assign \new_[1062]_  = \new_[70818]_  & \new_[70805]_ ;
  assign \new_[1063]_  = \new_[70792]_  & \new_[70779]_ ;
  assign \new_[1064]_  = \new_[70766]_  & \new_[70753]_ ;
  assign \new_[1065]_  = \new_[70740]_  & \new_[70727]_ ;
  assign \new_[1066]_  = \new_[70714]_  & \new_[70701]_ ;
  assign \new_[1067]_  = \new_[70688]_  & \new_[70675]_ ;
  assign \new_[1068]_  = \new_[70662]_  & \new_[70649]_ ;
  assign \new_[1069]_  = \new_[70636]_  & \new_[70623]_ ;
  assign \new_[1070]_  = \new_[70610]_  & \new_[70597]_ ;
  assign \new_[1071]_  = \new_[70584]_  & \new_[70571]_ ;
  assign \new_[1072]_  = \new_[70558]_  & \new_[70545]_ ;
  assign \new_[1073]_  = \new_[70532]_  & \new_[70519]_ ;
  assign \new_[1074]_  = \new_[70506]_  & \new_[70493]_ ;
  assign \new_[1075]_  = \new_[70480]_  & \new_[70467]_ ;
  assign \new_[1076]_  = \new_[70454]_  & \new_[70441]_ ;
  assign \new_[1077]_  = \new_[70428]_  & \new_[70415]_ ;
  assign \new_[1078]_  = \new_[70402]_  & \new_[70389]_ ;
  assign \new_[1079]_  = \new_[70376]_  & \new_[70363]_ ;
  assign \new_[1080]_  = \new_[70350]_  & \new_[70337]_ ;
  assign \new_[1081]_  = \new_[70324]_  & \new_[70311]_ ;
  assign \new_[1082]_  = \new_[70298]_  & \new_[70285]_ ;
  assign \new_[1083]_  = \new_[70272]_  & \new_[70259]_ ;
  assign \new_[1084]_  = \new_[70246]_  & \new_[70233]_ ;
  assign \new_[1085]_  = \new_[70220]_  & \new_[70207]_ ;
  assign \new_[1086]_  = \new_[70194]_  & \new_[70181]_ ;
  assign \new_[1087]_  = \new_[70168]_  & \new_[70155]_ ;
  assign \new_[1088]_  = \new_[70142]_  & \new_[70129]_ ;
  assign \new_[1089]_  = \new_[70116]_  & \new_[70103]_ ;
  assign \new_[1090]_  = \new_[70090]_  & \new_[70077]_ ;
  assign \new_[1091]_  = \new_[70064]_  & \new_[70051]_ ;
  assign \new_[1092]_  = \new_[70038]_  & \new_[70025]_ ;
  assign \new_[1093]_  = \new_[70012]_  & \new_[69999]_ ;
  assign \new_[1094]_  = \new_[69986]_  & \new_[69973]_ ;
  assign \new_[1095]_  = \new_[69960]_  & \new_[69947]_ ;
  assign \new_[1096]_  = \new_[69934]_  & \new_[69921]_ ;
  assign \new_[1097]_  = \new_[69908]_  & \new_[69895]_ ;
  assign \new_[1098]_  = \new_[69882]_  & \new_[69869]_ ;
  assign \new_[1099]_  = \new_[69856]_  & \new_[69843]_ ;
  assign \new_[1100]_  = \new_[69830]_  & \new_[69817]_ ;
  assign \new_[1101]_  = \new_[69804]_  & \new_[69791]_ ;
  assign \new_[1102]_  = \new_[69778]_  & \new_[69765]_ ;
  assign \new_[1103]_  = \new_[69752]_  & \new_[69739]_ ;
  assign \new_[1104]_  = \new_[69726]_  & \new_[69713]_ ;
  assign \new_[1105]_  = \new_[69700]_  & \new_[69687]_ ;
  assign \new_[1106]_  = \new_[69674]_  & \new_[69661]_ ;
  assign \new_[1107]_  = \new_[69648]_  & \new_[69635]_ ;
  assign \new_[1108]_  = \new_[69622]_  & \new_[69609]_ ;
  assign \new_[1109]_  = \new_[69596]_  & \new_[69583]_ ;
  assign \new_[1110]_  = \new_[69570]_  & \new_[69557]_ ;
  assign \new_[1111]_  = \new_[69544]_  & \new_[69531]_ ;
  assign \new_[1112]_  = \new_[69518]_  & \new_[69505]_ ;
  assign \new_[1113]_  = \new_[69492]_  & \new_[69479]_ ;
  assign \new_[1114]_  = \new_[69466]_  & \new_[69453]_ ;
  assign \new_[1115]_  = \new_[69440]_  & \new_[69427]_ ;
  assign \new_[1116]_  = \new_[69414]_  & \new_[69401]_ ;
  assign \new_[1117]_  = \new_[69388]_  & \new_[69375]_ ;
  assign \new_[1118]_  = \new_[69362]_  & \new_[69349]_ ;
  assign \new_[1119]_  = \new_[69336]_  & \new_[69323]_ ;
  assign \new_[1120]_  = \new_[69310]_  & \new_[69297]_ ;
  assign \new_[1121]_  = \new_[69284]_  & \new_[69271]_ ;
  assign \new_[1122]_  = \new_[69258]_  & \new_[69245]_ ;
  assign \new_[1123]_  = \new_[69232]_  & \new_[69219]_ ;
  assign \new_[1124]_  = \new_[69206]_  & \new_[69193]_ ;
  assign \new_[1125]_  = \new_[69180]_  & \new_[69167]_ ;
  assign \new_[1126]_  = \new_[69154]_  & \new_[69141]_ ;
  assign \new_[1127]_  = \new_[69128]_  & \new_[69115]_ ;
  assign \new_[1128]_  = \new_[69102]_  & \new_[69089]_ ;
  assign \new_[1129]_  = \new_[69076]_  & \new_[69063]_ ;
  assign \new_[1130]_  = \new_[69050]_  & \new_[69037]_ ;
  assign \new_[1131]_  = \new_[69024]_  & \new_[69011]_ ;
  assign \new_[1132]_  = \new_[68998]_  & \new_[68985]_ ;
  assign \new_[1133]_  = \new_[68972]_  & \new_[68959]_ ;
  assign \new_[1134]_  = \new_[68946]_  & \new_[68933]_ ;
  assign \new_[1135]_  = \new_[68920]_  & \new_[68907]_ ;
  assign \new_[1136]_  = \new_[68894]_  & \new_[68881]_ ;
  assign \new_[1137]_  = \new_[68868]_  & \new_[68855]_ ;
  assign \new_[1138]_  = \new_[68842]_  & \new_[68829]_ ;
  assign \new_[1139]_  = \new_[68816]_  & \new_[68803]_ ;
  assign \new_[1140]_  = \new_[68790]_  & \new_[68777]_ ;
  assign \new_[1141]_  = \new_[68764]_  & \new_[68751]_ ;
  assign \new_[1142]_  = \new_[68738]_  & \new_[68725]_ ;
  assign \new_[1143]_  = \new_[68712]_  & \new_[68699]_ ;
  assign \new_[1144]_  = \new_[68686]_  & \new_[68673]_ ;
  assign \new_[1145]_  = \new_[68660]_  & \new_[68647]_ ;
  assign \new_[1146]_  = \new_[68634]_  & \new_[68621]_ ;
  assign \new_[1147]_  = \new_[68608]_  & \new_[68595]_ ;
  assign \new_[1148]_  = \new_[68582]_  & \new_[68569]_ ;
  assign \new_[1149]_  = \new_[68556]_  & \new_[68543]_ ;
  assign \new_[1150]_  = \new_[68530]_  & \new_[68517]_ ;
  assign \new_[1151]_  = \new_[68504]_  & \new_[68491]_ ;
  assign \new_[1152]_  = \new_[68478]_  & \new_[68465]_ ;
  assign \new_[1153]_  = \new_[68452]_  & \new_[68439]_ ;
  assign \new_[1154]_  = \new_[68426]_  & \new_[68413]_ ;
  assign \new_[1155]_  = \new_[68400]_  & \new_[68387]_ ;
  assign \new_[1156]_  = \new_[68374]_  & \new_[68361]_ ;
  assign \new_[1157]_  = \new_[68348]_  & \new_[68335]_ ;
  assign \new_[1158]_  = \new_[68322]_  & \new_[68309]_ ;
  assign \new_[1159]_  = \new_[68296]_  & \new_[68283]_ ;
  assign \new_[1160]_  = \new_[68270]_  & \new_[68257]_ ;
  assign \new_[1161]_  = \new_[68244]_  & \new_[68231]_ ;
  assign \new_[1162]_  = \new_[68218]_  & \new_[68205]_ ;
  assign \new_[1163]_  = \new_[68192]_  & \new_[68179]_ ;
  assign \new_[1164]_  = \new_[68166]_  & \new_[68153]_ ;
  assign \new_[1165]_  = \new_[68140]_  & \new_[68127]_ ;
  assign \new_[1166]_  = \new_[68114]_  & \new_[68101]_ ;
  assign \new_[1167]_  = \new_[68088]_  & \new_[68075]_ ;
  assign \new_[1168]_  = \new_[68062]_  & \new_[68049]_ ;
  assign \new_[1169]_  = \new_[68036]_  & \new_[68023]_ ;
  assign \new_[1170]_  = \new_[68010]_  & \new_[67997]_ ;
  assign \new_[1171]_  = \new_[67984]_  & \new_[67971]_ ;
  assign \new_[1172]_  = \new_[67958]_  & \new_[67945]_ ;
  assign \new_[1173]_  = \new_[67932]_  & \new_[67919]_ ;
  assign \new_[1174]_  = \new_[67906]_  & \new_[67893]_ ;
  assign \new_[1175]_  = \new_[67880]_  & \new_[67867]_ ;
  assign \new_[1176]_  = \new_[67854]_  & \new_[67841]_ ;
  assign \new_[1177]_  = \new_[67828]_  & \new_[67815]_ ;
  assign \new_[1178]_  = \new_[67802]_  & \new_[67789]_ ;
  assign \new_[1179]_  = \new_[67776]_  & \new_[67763]_ ;
  assign \new_[1180]_  = \new_[67750]_  & \new_[67737]_ ;
  assign \new_[1181]_  = \new_[67724]_  & \new_[67711]_ ;
  assign \new_[1182]_  = \new_[67698]_  & \new_[67685]_ ;
  assign \new_[1183]_  = \new_[67672]_  & \new_[67659]_ ;
  assign \new_[1184]_  = \new_[67646]_  & \new_[67633]_ ;
  assign \new_[1185]_  = \new_[67620]_  & \new_[67607]_ ;
  assign \new_[1186]_  = \new_[67594]_  & \new_[67581]_ ;
  assign \new_[1187]_  = \new_[67568]_  & \new_[67555]_ ;
  assign \new_[1188]_  = \new_[67542]_  & \new_[67529]_ ;
  assign \new_[1189]_  = \new_[67516]_  & \new_[67503]_ ;
  assign \new_[1190]_  = \new_[67490]_  & \new_[67477]_ ;
  assign \new_[1191]_  = \new_[67464]_  & \new_[67451]_ ;
  assign \new_[1192]_  = \new_[67438]_  & \new_[67425]_ ;
  assign \new_[1193]_  = \new_[67412]_  & \new_[67399]_ ;
  assign \new_[1194]_  = \new_[67386]_  & \new_[67373]_ ;
  assign \new_[1195]_  = \new_[67360]_  & \new_[67347]_ ;
  assign \new_[1196]_  = \new_[67334]_  & \new_[67321]_ ;
  assign \new_[1197]_  = \new_[67308]_  & \new_[67295]_ ;
  assign \new_[1198]_  = \new_[67282]_  & \new_[67269]_ ;
  assign \new_[1199]_  = \new_[67256]_  & \new_[67243]_ ;
  assign \new_[1200]_  = \new_[67230]_  & \new_[67217]_ ;
  assign \new_[1201]_  = \new_[67204]_  & \new_[67191]_ ;
  assign \new_[1202]_  = \new_[67178]_  & \new_[67165]_ ;
  assign \new_[1203]_  = \new_[67152]_  & \new_[67139]_ ;
  assign \new_[1204]_  = \new_[67126]_  & \new_[67113]_ ;
  assign \new_[1205]_  = \new_[67100]_  & \new_[67087]_ ;
  assign \new_[1206]_  = \new_[67074]_  & \new_[67061]_ ;
  assign \new_[1207]_  = \new_[67048]_  & \new_[67035]_ ;
  assign \new_[1208]_  = \new_[67022]_  & \new_[67009]_ ;
  assign \new_[1209]_  = \new_[66996]_  & \new_[66983]_ ;
  assign \new_[1210]_  = \new_[66970]_  & \new_[66957]_ ;
  assign \new_[1211]_  = \new_[66944]_  & \new_[66931]_ ;
  assign \new_[1212]_  = \new_[66918]_  & \new_[66905]_ ;
  assign \new_[1213]_  = \new_[66892]_  & \new_[66879]_ ;
  assign \new_[1214]_  = \new_[66866]_  & \new_[66853]_ ;
  assign \new_[1215]_  = \new_[66840]_  & \new_[66827]_ ;
  assign \new_[1216]_  = \new_[66814]_  & \new_[66801]_ ;
  assign \new_[1217]_  = \new_[66788]_  & \new_[66775]_ ;
  assign \new_[1218]_  = \new_[66762]_  & \new_[66749]_ ;
  assign \new_[1219]_  = \new_[66736]_  & \new_[66723]_ ;
  assign \new_[1220]_  = \new_[66710]_  & \new_[66697]_ ;
  assign \new_[1221]_  = \new_[66684]_  & \new_[66671]_ ;
  assign \new_[1222]_  = \new_[66658]_  & \new_[66645]_ ;
  assign \new_[1223]_  = \new_[66632]_  & \new_[66619]_ ;
  assign \new_[1224]_  = \new_[66606]_  & \new_[66593]_ ;
  assign \new_[1225]_  = \new_[66580]_  & \new_[66567]_ ;
  assign \new_[1226]_  = \new_[66554]_  & \new_[66541]_ ;
  assign \new_[1227]_  = \new_[66528]_  & \new_[66515]_ ;
  assign \new_[1228]_  = \new_[66502]_  & \new_[66489]_ ;
  assign \new_[1229]_  = \new_[66476]_  & \new_[66463]_ ;
  assign \new_[1230]_  = \new_[66450]_  & \new_[66437]_ ;
  assign \new_[1231]_  = \new_[66424]_  & \new_[66411]_ ;
  assign \new_[1232]_  = \new_[66398]_  & \new_[66385]_ ;
  assign \new_[1233]_  = \new_[66372]_  & \new_[66359]_ ;
  assign \new_[1234]_  = \new_[66346]_  & \new_[66333]_ ;
  assign \new_[1235]_  = \new_[66320]_  & \new_[66307]_ ;
  assign \new_[1236]_  = \new_[66294]_  & \new_[66281]_ ;
  assign \new_[1237]_  = \new_[66268]_  & \new_[66255]_ ;
  assign \new_[1238]_  = \new_[66242]_  & \new_[66229]_ ;
  assign \new_[1239]_  = \new_[66216]_  & \new_[66203]_ ;
  assign \new_[1240]_  = \new_[66190]_  & \new_[66177]_ ;
  assign \new_[1241]_  = \new_[66164]_  & \new_[66151]_ ;
  assign \new_[1242]_  = \new_[66138]_  & \new_[66125]_ ;
  assign \new_[1243]_  = \new_[66112]_  & \new_[66099]_ ;
  assign \new_[1244]_  = \new_[66086]_  & \new_[66073]_ ;
  assign \new_[1245]_  = \new_[66060]_  & \new_[66047]_ ;
  assign \new_[1246]_  = \new_[66034]_  & \new_[66021]_ ;
  assign \new_[1247]_  = \new_[66008]_  & \new_[65995]_ ;
  assign \new_[1248]_  = \new_[65982]_  & \new_[65969]_ ;
  assign \new_[1249]_  = \new_[65956]_  & \new_[65943]_ ;
  assign \new_[1250]_  = \new_[65930]_  & \new_[65917]_ ;
  assign \new_[1251]_  = \new_[65904]_  & \new_[65891]_ ;
  assign \new_[1252]_  = \new_[65878]_  & \new_[65865]_ ;
  assign \new_[1253]_  = \new_[65852]_  & \new_[65839]_ ;
  assign \new_[1254]_  = \new_[65826]_  & \new_[65813]_ ;
  assign \new_[1255]_  = \new_[65800]_  & \new_[65787]_ ;
  assign \new_[1256]_  = \new_[65774]_  & \new_[65761]_ ;
  assign \new_[1257]_  = \new_[65748]_  & \new_[65735]_ ;
  assign \new_[1258]_  = \new_[65722]_  & \new_[65709]_ ;
  assign \new_[1259]_  = \new_[65696]_  & \new_[65683]_ ;
  assign \new_[1260]_  = \new_[65670]_  & \new_[65657]_ ;
  assign \new_[1261]_  = \new_[65644]_  & \new_[65631]_ ;
  assign \new_[1262]_  = \new_[65618]_  & \new_[65605]_ ;
  assign \new_[1263]_  = \new_[65592]_  & \new_[65579]_ ;
  assign \new_[1264]_  = \new_[65566]_  & \new_[65553]_ ;
  assign \new_[1265]_  = \new_[65540]_  & \new_[65527]_ ;
  assign \new_[1266]_  = \new_[65514]_  & \new_[65501]_ ;
  assign \new_[1267]_  = \new_[65488]_  & \new_[65475]_ ;
  assign \new_[1268]_  = \new_[65462]_  & \new_[65449]_ ;
  assign \new_[1269]_  = \new_[65436]_  & \new_[65423]_ ;
  assign \new_[1270]_  = \new_[65410]_  & \new_[65397]_ ;
  assign \new_[1271]_  = \new_[65384]_  & \new_[65371]_ ;
  assign \new_[1272]_  = \new_[65358]_  & \new_[65345]_ ;
  assign \new_[1273]_  = \new_[65332]_  & \new_[65319]_ ;
  assign \new_[1274]_  = \new_[65306]_  & \new_[65293]_ ;
  assign \new_[1275]_  = \new_[65280]_  & \new_[65267]_ ;
  assign \new_[1276]_  = \new_[65254]_  & \new_[65241]_ ;
  assign \new_[1277]_  = \new_[65228]_  & \new_[65215]_ ;
  assign \new_[1278]_  = \new_[65202]_  & \new_[65189]_ ;
  assign \new_[1279]_  = \new_[65176]_  & \new_[65163]_ ;
  assign \new_[1280]_  = \new_[65150]_  & \new_[65137]_ ;
  assign \new_[1281]_  = \new_[65124]_  & \new_[65111]_ ;
  assign \new_[1282]_  = \new_[65098]_  & \new_[65085]_ ;
  assign \new_[1283]_  = \new_[65072]_  & \new_[65059]_ ;
  assign \new_[1284]_  = \new_[65046]_  & \new_[65033]_ ;
  assign \new_[1285]_  = \new_[65020]_  & \new_[65007]_ ;
  assign \new_[1286]_  = \new_[64994]_  & \new_[64981]_ ;
  assign \new_[1287]_  = \new_[64968]_  & \new_[64955]_ ;
  assign \new_[1288]_  = \new_[64942]_  & \new_[64929]_ ;
  assign \new_[1289]_  = \new_[64916]_  & \new_[64903]_ ;
  assign \new_[1290]_  = \new_[64890]_  & \new_[64877]_ ;
  assign \new_[1291]_  = \new_[64864]_  & \new_[64851]_ ;
  assign \new_[1292]_  = \new_[64838]_  & \new_[64825]_ ;
  assign \new_[1293]_  = \new_[64812]_  & \new_[64799]_ ;
  assign \new_[1294]_  = \new_[64786]_  & \new_[64773]_ ;
  assign \new_[1295]_  = \new_[64760]_  & \new_[64747]_ ;
  assign \new_[1296]_  = \new_[64734]_  & \new_[64721]_ ;
  assign \new_[1297]_  = \new_[64708]_  & \new_[64695]_ ;
  assign \new_[1298]_  = \new_[64682]_  & \new_[64669]_ ;
  assign \new_[1299]_  = \new_[64656]_  & \new_[64643]_ ;
  assign \new_[1300]_  = \new_[64630]_  & \new_[64617]_ ;
  assign \new_[1301]_  = \new_[64604]_  & \new_[64591]_ ;
  assign \new_[1302]_  = \new_[64578]_  & \new_[64565]_ ;
  assign \new_[1303]_  = \new_[64552]_  & \new_[64539]_ ;
  assign \new_[1304]_  = \new_[64526]_  & \new_[64513]_ ;
  assign \new_[1305]_  = \new_[64500]_  & \new_[64487]_ ;
  assign \new_[1306]_  = \new_[64474]_  & \new_[64461]_ ;
  assign \new_[1307]_  = \new_[64448]_  & \new_[64435]_ ;
  assign \new_[1308]_  = \new_[64422]_  & \new_[64409]_ ;
  assign \new_[1309]_  = \new_[64396]_  & \new_[64383]_ ;
  assign \new_[1310]_  = \new_[64370]_  & \new_[64357]_ ;
  assign \new_[1311]_  = \new_[64344]_  & \new_[64331]_ ;
  assign \new_[1312]_  = \new_[64318]_  & \new_[64305]_ ;
  assign \new_[1313]_  = \new_[64292]_  & \new_[64279]_ ;
  assign \new_[1314]_  = \new_[64266]_  & \new_[64253]_ ;
  assign \new_[1315]_  = \new_[64240]_  & \new_[64227]_ ;
  assign \new_[1316]_  = \new_[64214]_  & \new_[64201]_ ;
  assign \new_[1317]_  = \new_[64188]_  & \new_[64175]_ ;
  assign \new_[1318]_  = \new_[64162]_  & \new_[64149]_ ;
  assign \new_[1319]_  = \new_[64136]_  & \new_[64123]_ ;
  assign \new_[1320]_  = \new_[64110]_  & \new_[64097]_ ;
  assign \new_[1321]_  = \new_[64084]_  & \new_[64071]_ ;
  assign \new_[1322]_  = \new_[64058]_  & \new_[64045]_ ;
  assign \new_[1323]_  = \new_[64032]_  & \new_[64019]_ ;
  assign \new_[1324]_  = \new_[64006]_  & \new_[63993]_ ;
  assign \new_[1325]_  = \new_[63980]_  & \new_[63967]_ ;
  assign \new_[1326]_  = \new_[63954]_  & \new_[63941]_ ;
  assign \new_[1327]_  = \new_[63928]_  & \new_[63915]_ ;
  assign \new_[1328]_  = \new_[63902]_  & \new_[63889]_ ;
  assign \new_[1329]_  = \new_[63876]_  & \new_[63863]_ ;
  assign \new_[1330]_  = \new_[63850]_  & \new_[63837]_ ;
  assign \new_[1331]_  = \new_[63824]_  & \new_[63811]_ ;
  assign \new_[1332]_  = \new_[63798]_  & \new_[63785]_ ;
  assign \new_[1333]_  = \new_[63772]_  & \new_[63759]_ ;
  assign \new_[1334]_  = \new_[63746]_  & \new_[63733]_ ;
  assign \new_[1335]_  = \new_[63720]_  & \new_[63707]_ ;
  assign \new_[1336]_  = \new_[63694]_  & \new_[63681]_ ;
  assign \new_[1337]_  = \new_[63668]_  & \new_[63655]_ ;
  assign \new_[1338]_  = \new_[63642]_  & \new_[63629]_ ;
  assign \new_[1339]_  = \new_[63616]_  & \new_[63603]_ ;
  assign \new_[1340]_  = \new_[63590]_  & \new_[63577]_ ;
  assign \new_[1341]_  = \new_[63564]_  & \new_[63551]_ ;
  assign \new_[1342]_  = \new_[63538]_  & \new_[63525]_ ;
  assign \new_[1343]_  = \new_[63512]_  & \new_[63499]_ ;
  assign \new_[1344]_  = \new_[63486]_  & \new_[63473]_ ;
  assign \new_[1345]_  = \new_[63460]_  & \new_[63447]_ ;
  assign \new_[1346]_  = \new_[63434]_  & \new_[63421]_ ;
  assign \new_[1347]_  = \new_[63408]_  & \new_[63395]_ ;
  assign \new_[1348]_  = \new_[63382]_  & \new_[63369]_ ;
  assign \new_[1349]_  = \new_[63356]_  & \new_[63343]_ ;
  assign \new_[1350]_  = \new_[63330]_  & \new_[63317]_ ;
  assign \new_[1351]_  = \new_[63304]_  & \new_[63291]_ ;
  assign \new_[1352]_  = \new_[63278]_  & \new_[63265]_ ;
  assign \new_[1353]_  = \new_[63252]_  & \new_[63239]_ ;
  assign \new_[1354]_  = \new_[63226]_  & \new_[63213]_ ;
  assign \new_[1355]_  = \new_[63200]_  & \new_[63187]_ ;
  assign \new_[1356]_  = \new_[63174]_  & \new_[63161]_ ;
  assign \new_[1357]_  = \new_[63148]_  & \new_[63135]_ ;
  assign \new_[1358]_  = \new_[63122]_  & \new_[63109]_ ;
  assign \new_[1359]_  = \new_[63096]_  & \new_[63083]_ ;
  assign \new_[1360]_  = \new_[63070]_  & \new_[63057]_ ;
  assign \new_[1361]_  = \new_[63044]_  & \new_[63031]_ ;
  assign \new_[1362]_  = \new_[63018]_  & \new_[63005]_ ;
  assign \new_[1363]_  = \new_[62992]_  & \new_[62979]_ ;
  assign \new_[1364]_  = \new_[62966]_  & \new_[62953]_ ;
  assign \new_[1365]_  = \new_[62940]_  & \new_[62927]_ ;
  assign \new_[1366]_  = \new_[62914]_  & \new_[62901]_ ;
  assign \new_[1367]_  = \new_[62888]_  & \new_[62875]_ ;
  assign \new_[1368]_  = \new_[62862]_  & \new_[62849]_ ;
  assign \new_[1369]_  = \new_[62836]_  & \new_[62823]_ ;
  assign \new_[1370]_  = \new_[62810]_  & \new_[62797]_ ;
  assign \new_[1371]_  = \new_[62784]_  & \new_[62771]_ ;
  assign \new_[1372]_  = \new_[62758]_  & \new_[62745]_ ;
  assign \new_[1373]_  = \new_[62732]_  & \new_[62719]_ ;
  assign \new_[1374]_  = \new_[62706]_  & \new_[62693]_ ;
  assign \new_[1375]_  = \new_[62680]_  & \new_[62667]_ ;
  assign \new_[1376]_  = \new_[62654]_  & \new_[62641]_ ;
  assign \new_[1377]_  = \new_[62628]_  & \new_[62615]_ ;
  assign \new_[1378]_  = \new_[62602]_  & \new_[62589]_ ;
  assign \new_[1379]_  = \new_[62576]_  & \new_[62563]_ ;
  assign \new_[1380]_  = \new_[62550]_  & \new_[62537]_ ;
  assign \new_[1381]_  = \new_[62524]_  & \new_[62511]_ ;
  assign \new_[1382]_  = \new_[62498]_  & \new_[62485]_ ;
  assign \new_[1383]_  = \new_[62472]_  & \new_[62459]_ ;
  assign \new_[1384]_  = \new_[62446]_  & \new_[62433]_ ;
  assign \new_[1385]_  = \new_[62420]_  & \new_[62407]_ ;
  assign \new_[1386]_  = \new_[62394]_  & \new_[62381]_ ;
  assign \new_[1387]_  = \new_[62368]_  & \new_[62355]_ ;
  assign \new_[1388]_  = \new_[62342]_  & \new_[62329]_ ;
  assign \new_[1389]_  = \new_[62316]_  & \new_[62303]_ ;
  assign \new_[1390]_  = \new_[62290]_  & \new_[62277]_ ;
  assign \new_[1391]_  = \new_[62264]_  & \new_[62251]_ ;
  assign \new_[1392]_  = \new_[62238]_  & \new_[62225]_ ;
  assign \new_[1393]_  = \new_[62212]_  & \new_[62199]_ ;
  assign \new_[1394]_  = \new_[62186]_  & \new_[62173]_ ;
  assign \new_[1395]_  = \new_[62160]_  & \new_[62147]_ ;
  assign \new_[1396]_  = \new_[62134]_  & \new_[62121]_ ;
  assign \new_[1397]_  = \new_[62108]_  & \new_[62095]_ ;
  assign \new_[1398]_  = \new_[62082]_  & \new_[62069]_ ;
  assign \new_[1399]_  = \new_[62056]_  & \new_[62043]_ ;
  assign \new_[1400]_  = \new_[62030]_  & \new_[62017]_ ;
  assign \new_[1401]_  = \new_[62004]_  & \new_[61991]_ ;
  assign \new_[1402]_  = \new_[61978]_  & \new_[61965]_ ;
  assign \new_[1403]_  = \new_[61952]_  & \new_[61939]_ ;
  assign \new_[1404]_  = \new_[61926]_  & \new_[61913]_ ;
  assign \new_[1405]_  = \new_[61900]_  & \new_[61887]_ ;
  assign \new_[1406]_  = \new_[61874]_  & \new_[61861]_ ;
  assign \new_[1407]_  = \new_[61848]_  & \new_[61835]_ ;
  assign \new_[1408]_  = \new_[61822]_  & \new_[61809]_ ;
  assign \new_[1409]_  = \new_[61796]_  & \new_[61783]_ ;
  assign \new_[1410]_  = \new_[61770]_  & \new_[61757]_ ;
  assign \new_[1411]_  = \new_[61744]_  & \new_[61731]_ ;
  assign \new_[1412]_  = \new_[61718]_  & \new_[61705]_ ;
  assign \new_[1413]_  = \new_[61692]_  & \new_[61679]_ ;
  assign \new_[1414]_  = \new_[61666]_  & \new_[61653]_ ;
  assign \new_[1415]_  = \new_[61640]_  & \new_[61627]_ ;
  assign \new_[1416]_  = \new_[61614]_  & \new_[61601]_ ;
  assign \new_[1417]_  = \new_[61588]_  & \new_[61575]_ ;
  assign \new_[1418]_  = \new_[61562]_  & \new_[61549]_ ;
  assign \new_[1419]_  = \new_[61536]_  & \new_[61523]_ ;
  assign \new_[1420]_  = \new_[61510]_  & \new_[61497]_ ;
  assign \new_[1421]_  = \new_[61484]_  & \new_[61471]_ ;
  assign \new_[1422]_  = \new_[61458]_  & \new_[61445]_ ;
  assign \new_[1423]_  = \new_[61432]_  & \new_[61419]_ ;
  assign \new_[1424]_  = \new_[61406]_  & \new_[61393]_ ;
  assign \new_[1425]_  = \new_[61380]_  & \new_[61367]_ ;
  assign \new_[1426]_  = \new_[61354]_  & \new_[61341]_ ;
  assign \new_[1427]_  = \new_[61328]_  & \new_[61315]_ ;
  assign \new_[1428]_  = \new_[61302]_  & \new_[61289]_ ;
  assign \new_[1429]_  = \new_[61276]_  & \new_[61263]_ ;
  assign \new_[1430]_  = \new_[61250]_  & \new_[61237]_ ;
  assign \new_[1431]_  = \new_[61224]_  & \new_[61211]_ ;
  assign \new_[1432]_  = \new_[61198]_  & \new_[61185]_ ;
  assign \new_[1433]_  = \new_[61172]_  & \new_[61159]_ ;
  assign \new_[1434]_  = \new_[61146]_  & \new_[61133]_ ;
  assign \new_[1435]_  = \new_[61120]_  & \new_[61107]_ ;
  assign \new_[1436]_  = \new_[61094]_  & \new_[61081]_ ;
  assign \new_[1437]_  = \new_[61068]_  & \new_[61055]_ ;
  assign \new_[1438]_  = \new_[61042]_  & \new_[61029]_ ;
  assign \new_[1439]_  = \new_[61016]_  & \new_[61003]_ ;
  assign \new_[1440]_  = \new_[60990]_  & \new_[60977]_ ;
  assign \new_[1441]_  = \new_[60964]_  & \new_[60951]_ ;
  assign \new_[1442]_  = \new_[60938]_  & \new_[60925]_ ;
  assign \new_[1443]_  = \new_[60912]_  & \new_[60899]_ ;
  assign \new_[1444]_  = \new_[60886]_  & \new_[60873]_ ;
  assign \new_[1445]_  = \new_[60860]_  & \new_[60847]_ ;
  assign \new_[1446]_  = \new_[60834]_  & \new_[60821]_ ;
  assign \new_[1447]_  = \new_[60808]_  & \new_[60795]_ ;
  assign \new_[1448]_  = \new_[60782]_  & \new_[60769]_ ;
  assign \new_[1449]_  = \new_[60756]_  & \new_[60743]_ ;
  assign \new_[1450]_  = \new_[60730]_  & \new_[60717]_ ;
  assign \new_[1451]_  = \new_[60704]_  & \new_[60691]_ ;
  assign \new_[1452]_  = \new_[60678]_  & \new_[60665]_ ;
  assign \new_[1453]_  = \new_[60652]_  & \new_[60639]_ ;
  assign \new_[1454]_  = \new_[60626]_  & \new_[60613]_ ;
  assign \new_[1455]_  = \new_[60600]_  & \new_[60587]_ ;
  assign \new_[1456]_  = \new_[60574]_  & \new_[60561]_ ;
  assign \new_[1457]_  = \new_[60548]_  & \new_[60535]_ ;
  assign \new_[1458]_  = \new_[60522]_  & \new_[60509]_ ;
  assign \new_[1459]_  = \new_[60496]_  & \new_[60483]_ ;
  assign \new_[1460]_  = \new_[60470]_  & \new_[60457]_ ;
  assign \new_[1461]_  = \new_[60444]_  & \new_[60431]_ ;
  assign \new_[1462]_  = \new_[60418]_  & \new_[60405]_ ;
  assign \new_[1463]_  = \new_[60392]_  & \new_[60379]_ ;
  assign \new_[1464]_  = \new_[60366]_  & \new_[60353]_ ;
  assign \new_[1465]_  = \new_[60340]_  & \new_[60327]_ ;
  assign \new_[1466]_  = \new_[60314]_  & \new_[60301]_ ;
  assign \new_[1467]_  = \new_[60288]_  & \new_[60275]_ ;
  assign \new_[1468]_  = \new_[60262]_  & \new_[60249]_ ;
  assign \new_[1469]_  = \new_[60236]_  & \new_[60223]_ ;
  assign \new_[1470]_  = \new_[60210]_  & \new_[60197]_ ;
  assign \new_[1471]_  = \new_[60184]_  & \new_[60171]_ ;
  assign \new_[1472]_  = \new_[60158]_  & \new_[60145]_ ;
  assign \new_[1473]_  = \new_[60132]_  & \new_[60119]_ ;
  assign \new_[1474]_  = \new_[60106]_  & \new_[60093]_ ;
  assign \new_[1475]_  = \new_[60080]_  & \new_[60067]_ ;
  assign \new_[1476]_  = \new_[60054]_  & \new_[60041]_ ;
  assign \new_[1477]_  = \new_[60028]_  & \new_[60015]_ ;
  assign \new_[1478]_  = \new_[60002]_  & \new_[59989]_ ;
  assign \new_[1479]_  = \new_[59976]_  & \new_[59963]_ ;
  assign \new_[1480]_  = \new_[59950]_  & \new_[59937]_ ;
  assign \new_[1481]_  = \new_[59924]_  & \new_[59911]_ ;
  assign \new_[1482]_  = \new_[59898]_  & \new_[59885]_ ;
  assign \new_[1483]_  = \new_[59872]_  & \new_[59859]_ ;
  assign \new_[1484]_  = \new_[59846]_  & \new_[59833]_ ;
  assign \new_[1485]_  = \new_[59820]_  & \new_[59807]_ ;
  assign \new_[1486]_  = \new_[59794]_  & \new_[59781]_ ;
  assign \new_[1487]_  = \new_[59768]_  & \new_[59755]_ ;
  assign \new_[1488]_  = \new_[59742]_  & \new_[59729]_ ;
  assign \new_[1489]_  = \new_[59716]_  & \new_[59703]_ ;
  assign \new_[1490]_  = \new_[59690]_  & \new_[59677]_ ;
  assign \new_[1491]_  = \new_[59664]_  & \new_[59651]_ ;
  assign \new_[1492]_  = \new_[59638]_  & \new_[59625]_ ;
  assign \new_[1493]_  = \new_[59612]_  & \new_[59599]_ ;
  assign \new_[1494]_  = \new_[59586]_  & \new_[59573]_ ;
  assign \new_[1495]_  = \new_[59560]_  & \new_[59547]_ ;
  assign \new_[1496]_  = \new_[59534]_  & \new_[59521]_ ;
  assign \new_[1497]_  = \new_[59508]_  & \new_[59495]_ ;
  assign \new_[1498]_  = \new_[59482]_  & \new_[59469]_ ;
  assign \new_[1499]_  = \new_[59456]_  & \new_[59443]_ ;
  assign \new_[1500]_  = \new_[59430]_  & \new_[59417]_ ;
  assign \new_[1501]_  = \new_[59404]_  & \new_[59391]_ ;
  assign \new_[1502]_  = \new_[59378]_  & \new_[59365]_ ;
  assign \new_[1503]_  = \new_[59352]_  & \new_[59339]_ ;
  assign \new_[1504]_  = \new_[59326]_  & \new_[59313]_ ;
  assign \new_[1505]_  = \new_[59300]_  & \new_[59287]_ ;
  assign \new_[1506]_  = \new_[59274]_  & \new_[59261]_ ;
  assign \new_[1507]_  = \new_[59248]_  & \new_[59235]_ ;
  assign \new_[1508]_  = \new_[59222]_  & \new_[59209]_ ;
  assign \new_[1509]_  = \new_[59196]_  & \new_[59183]_ ;
  assign \new_[1510]_  = \new_[59170]_  & \new_[59157]_ ;
  assign \new_[1511]_  = \new_[59144]_  & \new_[59131]_ ;
  assign \new_[1512]_  = \new_[59118]_  & \new_[59105]_ ;
  assign \new_[1513]_  = \new_[59092]_  & \new_[59079]_ ;
  assign \new_[1514]_  = \new_[59066]_  & \new_[59053]_ ;
  assign \new_[1515]_  = \new_[59040]_  & \new_[59027]_ ;
  assign \new_[1516]_  = \new_[59014]_  & \new_[59001]_ ;
  assign \new_[1517]_  = \new_[58988]_  & \new_[58975]_ ;
  assign \new_[1518]_  = \new_[58962]_  & \new_[58949]_ ;
  assign \new_[1519]_  = \new_[58936]_  & \new_[58923]_ ;
  assign \new_[1520]_  = \new_[58910]_  & \new_[58897]_ ;
  assign \new_[1521]_  = \new_[58884]_  & \new_[58871]_ ;
  assign \new_[1522]_  = \new_[58858]_  & \new_[58845]_ ;
  assign \new_[1523]_  = \new_[58832]_  & \new_[58819]_ ;
  assign \new_[1524]_  = \new_[58806]_  & \new_[58793]_ ;
  assign \new_[1525]_  = \new_[58780]_  & \new_[58767]_ ;
  assign \new_[1526]_  = \new_[58754]_  & \new_[58741]_ ;
  assign \new_[1527]_  = \new_[58728]_  & \new_[58715]_ ;
  assign \new_[1528]_  = \new_[58702]_  & \new_[58689]_ ;
  assign \new_[1529]_  = \new_[58676]_  & \new_[58663]_ ;
  assign \new_[1530]_  = \new_[58650]_  & \new_[58637]_ ;
  assign \new_[1531]_  = \new_[58624]_  & \new_[58611]_ ;
  assign \new_[1532]_  = \new_[58598]_  & \new_[58585]_ ;
  assign \new_[1533]_  = \new_[58572]_  & \new_[58559]_ ;
  assign \new_[1534]_  = \new_[58546]_  & \new_[58533]_ ;
  assign \new_[1535]_  = \new_[58520]_  & \new_[58507]_ ;
  assign \new_[1536]_  = \new_[58494]_  & \new_[58481]_ ;
  assign \new_[1537]_  = \new_[58468]_  & \new_[58455]_ ;
  assign \new_[1538]_  = \new_[58442]_  & \new_[58429]_ ;
  assign \new_[1539]_  = \new_[58416]_  & \new_[58403]_ ;
  assign \new_[1540]_  = \new_[58390]_  & \new_[58377]_ ;
  assign \new_[1541]_  = \new_[58364]_  & \new_[58351]_ ;
  assign \new_[1542]_  = \new_[58338]_  & \new_[58325]_ ;
  assign \new_[1543]_  = \new_[58312]_  & \new_[58299]_ ;
  assign \new_[1544]_  = \new_[58286]_  & \new_[58273]_ ;
  assign \new_[1545]_  = \new_[58260]_  & \new_[58247]_ ;
  assign \new_[1546]_  = \new_[58234]_  & \new_[58221]_ ;
  assign \new_[1547]_  = \new_[58208]_  & \new_[58195]_ ;
  assign \new_[1548]_  = \new_[58182]_  & \new_[58169]_ ;
  assign \new_[1549]_  = \new_[58156]_  & \new_[58143]_ ;
  assign \new_[1550]_  = \new_[58130]_  & \new_[58117]_ ;
  assign \new_[1551]_  = \new_[58104]_  & \new_[58091]_ ;
  assign \new_[1552]_  = \new_[58078]_  & \new_[58065]_ ;
  assign \new_[1553]_  = \new_[58052]_  & \new_[58039]_ ;
  assign \new_[1554]_  = \new_[58026]_  & \new_[58013]_ ;
  assign \new_[1555]_  = \new_[58000]_  & \new_[57987]_ ;
  assign \new_[1556]_  = \new_[57974]_  & \new_[57961]_ ;
  assign \new_[1557]_  = \new_[57948]_  & \new_[57935]_ ;
  assign \new_[1558]_  = \new_[57922]_  & \new_[57909]_ ;
  assign \new_[1559]_  = \new_[57896]_  & \new_[57883]_ ;
  assign \new_[1560]_  = \new_[57870]_  & \new_[57857]_ ;
  assign \new_[1561]_  = \new_[57844]_  & \new_[57831]_ ;
  assign \new_[1562]_  = \new_[57818]_  & \new_[57805]_ ;
  assign \new_[1563]_  = \new_[57792]_  & \new_[57779]_ ;
  assign \new_[1564]_  = \new_[57766]_  & \new_[57753]_ ;
  assign \new_[1565]_  = \new_[57740]_  & \new_[57727]_ ;
  assign \new_[1566]_  = \new_[57714]_  & \new_[57701]_ ;
  assign \new_[1567]_  = \new_[57688]_  & \new_[57675]_ ;
  assign \new_[1568]_  = \new_[57662]_  & \new_[57649]_ ;
  assign \new_[1569]_  = \new_[57636]_  & \new_[57623]_ ;
  assign \new_[1570]_  = \new_[57610]_  & \new_[57597]_ ;
  assign \new_[1571]_  = \new_[57584]_  & \new_[57571]_ ;
  assign \new_[1572]_  = \new_[57558]_  & \new_[57545]_ ;
  assign \new_[1573]_  = \new_[57532]_  & \new_[57519]_ ;
  assign \new_[1574]_  = \new_[57506]_  & \new_[57493]_ ;
  assign \new_[1575]_  = \new_[57480]_  & \new_[57467]_ ;
  assign \new_[1576]_  = \new_[57454]_  & \new_[57441]_ ;
  assign \new_[1577]_  = \new_[57428]_  & \new_[57415]_ ;
  assign \new_[1578]_  = \new_[57402]_  & \new_[57389]_ ;
  assign \new_[1579]_  = \new_[57376]_  & \new_[57363]_ ;
  assign \new_[1580]_  = \new_[57350]_  & \new_[57337]_ ;
  assign \new_[1581]_  = \new_[57324]_  & \new_[57311]_ ;
  assign \new_[1582]_  = \new_[57298]_  & \new_[57285]_ ;
  assign \new_[1583]_  = \new_[57272]_  & \new_[57259]_ ;
  assign \new_[1584]_  = \new_[57246]_  & \new_[57233]_ ;
  assign \new_[1585]_  = \new_[57220]_  & \new_[57207]_ ;
  assign \new_[1586]_  = \new_[57194]_  & \new_[57181]_ ;
  assign \new_[1587]_  = \new_[57168]_  & \new_[57155]_ ;
  assign \new_[1588]_  = \new_[57142]_  & \new_[57129]_ ;
  assign \new_[1589]_  = \new_[57116]_  & \new_[57103]_ ;
  assign \new_[1590]_  = \new_[57090]_  & \new_[57077]_ ;
  assign \new_[1591]_  = \new_[57064]_  & \new_[57051]_ ;
  assign \new_[1592]_  = \new_[57038]_  & \new_[57025]_ ;
  assign \new_[1593]_  = \new_[57012]_  & \new_[56999]_ ;
  assign \new_[1594]_  = \new_[56986]_  & \new_[56973]_ ;
  assign \new_[1595]_  = \new_[56960]_  & \new_[56947]_ ;
  assign \new_[1596]_  = \new_[56934]_  & \new_[56921]_ ;
  assign \new_[1597]_  = \new_[56908]_  & \new_[56895]_ ;
  assign \new_[1598]_  = \new_[56882]_  & \new_[56869]_ ;
  assign \new_[1599]_  = \new_[56856]_  & \new_[56843]_ ;
  assign \new_[1600]_  = \new_[56830]_  & \new_[56817]_ ;
  assign \new_[1601]_  = \new_[56804]_  & \new_[56791]_ ;
  assign \new_[1602]_  = \new_[56778]_  & \new_[56765]_ ;
  assign \new_[1603]_  = \new_[56752]_  & \new_[56739]_ ;
  assign \new_[1604]_  = \new_[56728]_  & \new_[56715]_ ;
  assign \new_[1605]_  = \new_[56704]_  & \new_[56691]_ ;
  assign \new_[1606]_  = \new_[56680]_  & \new_[56667]_ ;
  assign \new_[1607]_  = \new_[56656]_  & \new_[56643]_ ;
  assign \new_[1608]_  = \new_[56632]_  & \new_[56619]_ ;
  assign \new_[1609]_  = \new_[56608]_  & \new_[56595]_ ;
  assign \new_[1610]_  = \new_[56584]_  & \new_[56571]_ ;
  assign \new_[1611]_  = \new_[56560]_  & \new_[56547]_ ;
  assign \new_[1612]_  = \new_[56536]_  & \new_[56523]_ ;
  assign \new_[1613]_  = \new_[56512]_  & \new_[56499]_ ;
  assign \new_[1614]_  = \new_[56488]_  & \new_[56475]_ ;
  assign \new_[1615]_  = \new_[56464]_  & \new_[56451]_ ;
  assign \new_[1616]_  = \new_[56440]_  & \new_[56427]_ ;
  assign \new_[1617]_  = \new_[56416]_  & \new_[56403]_ ;
  assign \new_[1618]_  = \new_[56392]_  & \new_[56379]_ ;
  assign \new_[1619]_  = \new_[56368]_  & \new_[56355]_ ;
  assign \new_[1620]_  = \new_[56344]_  & \new_[56331]_ ;
  assign \new_[1621]_  = \new_[56320]_  & \new_[56307]_ ;
  assign \new_[1622]_  = \new_[56296]_  & \new_[56283]_ ;
  assign \new_[1623]_  = \new_[56272]_  & \new_[56259]_ ;
  assign \new_[1624]_  = \new_[56248]_  & \new_[56235]_ ;
  assign \new_[1625]_  = \new_[56224]_  & \new_[56211]_ ;
  assign \new_[1626]_  = \new_[56200]_  & \new_[56187]_ ;
  assign \new_[1627]_  = \new_[56176]_  & \new_[56163]_ ;
  assign \new_[1628]_  = \new_[56152]_  & \new_[56139]_ ;
  assign \new_[1629]_  = \new_[56128]_  & \new_[56115]_ ;
  assign \new_[1630]_  = \new_[56104]_  & \new_[56091]_ ;
  assign \new_[1631]_  = \new_[56080]_  & \new_[56067]_ ;
  assign \new_[1632]_  = \new_[56056]_  & \new_[56043]_ ;
  assign \new_[1633]_  = \new_[56032]_  & \new_[56019]_ ;
  assign \new_[1634]_  = \new_[56008]_  & \new_[55995]_ ;
  assign \new_[1635]_  = \new_[55984]_  & \new_[55971]_ ;
  assign \new_[1636]_  = \new_[55960]_  & \new_[55947]_ ;
  assign \new_[1637]_  = \new_[55936]_  & \new_[55923]_ ;
  assign \new_[1638]_  = \new_[55912]_  & \new_[55899]_ ;
  assign \new_[1639]_  = \new_[55888]_  & \new_[55875]_ ;
  assign \new_[1640]_  = \new_[55864]_  & \new_[55851]_ ;
  assign \new_[1641]_  = \new_[55840]_  & \new_[55827]_ ;
  assign \new_[1642]_  = \new_[55816]_  & \new_[55803]_ ;
  assign \new_[1643]_  = \new_[55792]_  & \new_[55779]_ ;
  assign \new_[1644]_  = \new_[55768]_  & \new_[55755]_ ;
  assign \new_[1645]_  = \new_[55744]_  & \new_[55731]_ ;
  assign \new_[1646]_  = \new_[55720]_  & \new_[55707]_ ;
  assign \new_[1647]_  = \new_[55696]_  & \new_[55683]_ ;
  assign \new_[1648]_  = \new_[55672]_  & \new_[55659]_ ;
  assign \new_[1649]_  = \new_[55648]_  & \new_[55635]_ ;
  assign \new_[1650]_  = \new_[55624]_  & \new_[55611]_ ;
  assign \new_[1651]_  = \new_[55600]_  & \new_[55587]_ ;
  assign \new_[1652]_  = \new_[55576]_  & \new_[55563]_ ;
  assign \new_[1653]_  = \new_[55552]_  & \new_[55539]_ ;
  assign \new_[1654]_  = \new_[55528]_  & \new_[55515]_ ;
  assign \new_[1655]_  = \new_[55504]_  & \new_[55491]_ ;
  assign \new_[1656]_  = \new_[55480]_  & \new_[55467]_ ;
  assign \new_[1657]_  = \new_[55456]_  & \new_[55443]_ ;
  assign \new_[1658]_  = \new_[55432]_  & \new_[55419]_ ;
  assign \new_[1659]_  = \new_[55408]_  & \new_[55395]_ ;
  assign \new_[1660]_  = \new_[55384]_  & \new_[55371]_ ;
  assign \new_[1661]_  = \new_[55360]_  & \new_[55347]_ ;
  assign \new_[1662]_  = \new_[55336]_  & \new_[55323]_ ;
  assign \new_[1663]_  = \new_[55312]_  & \new_[55299]_ ;
  assign \new_[1664]_  = \new_[55288]_  & \new_[55275]_ ;
  assign \new_[1665]_  = \new_[55264]_  & \new_[55251]_ ;
  assign \new_[1666]_  = \new_[55240]_  & \new_[55227]_ ;
  assign \new_[1667]_  = \new_[55216]_  & \new_[55203]_ ;
  assign \new_[1668]_  = \new_[55192]_  & \new_[55179]_ ;
  assign \new_[1669]_  = \new_[55168]_  & \new_[55155]_ ;
  assign \new_[1670]_  = \new_[55144]_  & \new_[55131]_ ;
  assign \new_[1671]_  = \new_[55120]_  & \new_[55107]_ ;
  assign \new_[1672]_  = \new_[55096]_  & \new_[55083]_ ;
  assign \new_[1673]_  = \new_[55072]_  & \new_[55059]_ ;
  assign \new_[1674]_  = \new_[55048]_  & \new_[55035]_ ;
  assign \new_[1675]_  = \new_[55024]_  & \new_[55011]_ ;
  assign \new_[1676]_  = \new_[55000]_  & \new_[54987]_ ;
  assign \new_[1677]_  = \new_[54976]_  & \new_[54963]_ ;
  assign \new_[1678]_  = \new_[54952]_  & \new_[54939]_ ;
  assign \new_[1679]_  = \new_[54928]_  & \new_[54915]_ ;
  assign \new_[1680]_  = \new_[54904]_  & \new_[54891]_ ;
  assign \new_[1681]_  = \new_[54880]_  & \new_[54867]_ ;
  assign \new_[1682]_  = \new_[54856]_  & \new_[54843]_ ;
  assign \new_[1683]_  = \new_[54832]_  & \new_[54819]_ ;
  assign \new_[1684]_  = \new_[54808]_  & \new_[54795]_ ;
  assign \new_[1685]_  = \new_[54784]_  & \new_[54771]_ ;
  assign \new_[1686]_  = \new_[54760]_  & \new_[54747]_ ;
  assign \new_[1687]_  = \new_[54736]_  & \new_[54723]_ ;
  assign \new_[1688]_  = \new_[54712]_  & \new_[54699]_ ;
  assign \new_[1689]_  = \new_[54688]_  & \new_[54675]_ ;
  assign \new_[1690]_  = \new_[54664]_  & \new_[54651]_ ;
  assign \new_[1691]_  = \new_[54640]_  & \new_[54627]_ ;
  assign \new_[1692]_  = \new_[54616]_  & \new_[54603]_ ;
  assign \new_[1693]_  = \new_[54592]_  & \new_[54579]_ ;
  assign \new_[1694]_  = \new_[54568]_  & \new_[54555]_ ;
  assign \new_[1695]_  = \new_[54544]_  & \new_[54531]_ ;
  assign \new_[1696]_  = \new_[54520]_  & \new_[54507]_ ;
  assign \new_[1697]_  = \new_[54496]_  & \new_[54483]_ ;
  assign \new_[1698]_  = \new_[54472]_  & \new_[54459]_ ;
  assign \new_[1699]_  = \new_[54448]_  & \new_[54435]_ ;
  assign \new_[1700]_  = \new_[54424]_  & \new_[54411]_ ;
  assign \new_[1701]_  = \new_[54400]_  & \new_[54387]_ ;
  assign \new_[1702]_  = \new_[54376]_  & \new_[54363]_ ;
  assign \new_[1703]_  = \new_[54352]_  & \new_[54339]_ ;
  assign \new_[1704]_  = \new_[54328]_  & \new_[54315]_ ;
  assign \new_[1705]_  = \new_[54304]_  & \new_[54291]_ ;
  assign \new_[1706]_  = \new_[54280]_  & \new_[54267]_ ;
  assign \new_[1707]_  = \new_[54256]_  & \new_[54243]_ ;
  assign \new_[1708]_  = \new_[54232]_  & \new_[54219]_ ;
  assign \new_[1709]_  = \new_[54208]_  & \new_[54195]_ ;
  assign \new_[1710]_  = \new_[54184]_  & \new_[54171]_ ;
  assign \new_[1711]_  = \new_[54160]_  & \new_[54147]_ ;
  assign \new_[1712]_  = \new_[54136]_  & \new_[54123]_ ;
  assign \new_[1713]_  = \new_[54112]_  & \new_[54099]_ ;
  assign \new_[1714]_  = \new_[54088]_  & \new_[54075]_ ;
  assign \new_[1715]_  = \new_[54064]_  & \new_[54051]_ ;
  assign \new_[1716]_  = \new_[54040]_  & \new_[54027]_ ;
  assign \new_[1717]_  = \new_[54016]_  & \new_[54003]_ ;
  assign \new_[1718]_  = \new_[53992]_  & \new_[53979]_ ;
  assign \new_[1719]_  = \new_[53968]_  & \new_[53955]_ ;
  assign \new_[1720]_  = \new_[53944]_  & \new_[53931]_ ;
  assign \new_[1721]_  = \new_[53920]_  & \new_[53907]_ ;
  assign \new_[1722]_  = \new_[53896]_  & \new_[53883]_ ;
  assign \new_[1723]_  = \new_[53872]_  & \new_[53859]_ ;
  assign \new_[1724]_  = \new_[53848]_  & \new_[53835]_ ;
  assign \new_[1725]_  = \new_[53824]_  & \new_[53811]_ ;
  assign \new_[1726]_  = \new_[53800]_  & \new_[53787]_ ;
  assign \new_[1727]_  = \new_[53776]_  & \new_[53763]_ ;
  assign \new_[1728]_  = \new_[53752]_  & \new_[53739]_ ;
  assign \new_[1729]_  = \new_[53728]_  & \new_[53715]_ ;
  assign \new_[1730]_  = \new_[53704]_  & \new_[53691]_ ;
  assign \new_[1731]_  = \new_[53680]_  & \new_[53667]_ ;
  assign \new_[1732]_  = \new_[53656]_  & \new_[53643]_ ;
  assign \new_[1733]_  = \new_[53632]_  & \new_[53619]_ ;
  assign \new_[1734]_  = \new_[53608]_  & \new_[53595]_ ;
  assign \new_[1735]_  = \new_[53584]_  & \new_[53571]_ ;
  assign \new_[1736]_  = \new_[53560]_  & \new_[53547]_ ;
  assign \new_[1737]_  = \new_[53536]_  & \new_[53523]_ ;
  assign \new_[1738]_  = \new_[53512]_  & \new_[53499]_ ;
  assign \new_[1739]_  = \new_[53488]_  & \new_[53475]_ ;
  assign \new_[1740]_  = \new_[53464]_  & \new_[53451]_ ;
  assign \new_[1741]_  = \new_[53440]_  & \new_[53427]_ ;
  assign \new_[1742]_  = \new_[53416]_  & \new_[53403]_ ;
  assign \new_[1743]_  = \new_[53392]_  & \new_[53379]_ ;
  assign \new_[1744]_  = \new_[53368]_  & \new_[53355]_ ;
  assign \new_[1745]_  = \new_[53344]_  & \new_[53331]_ ;
  assign \new_[1746]_  = \new_[53320]_  & \new_[53307]_ ;
  assign \new_[1747]_  = \new_[53296]_  & \new_[53283]_ ;
  assign \new_[1748]_  = \new_[53272]_  & \new_[53259]_ ;
  assign \new_[1749]_  = \new_[53248]_  & \new_[53235]_ ;
  assign \new_[1750]_  = \new_[53224]_  & \new_[53211]_ ;
  assign \new_[1751]_  = \new_[53200]_  & \new_[53187]_ ;
  assign \new_[1752]_  = \new_[53176]_  & \new_[53163]_ ;
  assign \new_[1753]_  = \new_[53152]_  & \new_[53139]_ ;
  assign \new_[1754]_  = \new_[53128]_  & \new_[53115]_ ;
  assign \new_[1755]_  = \new_[53104]_  & \new_[53091]_ ;
  assign \new_[1756]_  = \new_[53080]_  & \new_[53067]_ ;
  assign \new_[1757]_  = \new_[53056]_  & \new_[53043]_ ;
  assign \new_[1758]_  = \new_[53032]_  & \new_[53019]_ ;
  assign \new_[1759]_  = \new_[53008]_  & \new_[52995]_ ;
  assign \new_[1760]_  = \new_[52984]_  & \new_[52971]_ ;
  assign \new_[1761]_  = \new_[52960]_  & \new_[52947]_ ;
  assign \new_[1762]_  = \new_[52936]_  & \new_[52923]_ ;
  assign \new_[1763]_  = \new_[52912]_  & \new_[52899]_ ;
  assign \new_[1764]_  = \new_[52888]_  & \new_[52875]_ ;
  assign \new_[1765]_  = \new_[52864]_  & \new_[52851]_ ;
  assign \new_[1766]_  = \new_[52840]_  & \new_[52827]_ ;
  assign \new_[1767]_  = \new_[52816]_  & \new_[52803]_ ;
  assign \new_[1768]_  = \new_[52792]_  & \new_[52779]_ ;
  assign \new_[1769]_  = \new_[52768]_  & \new_[52755]_ ;
  assign \new_[1770]_  = \new_[52744]_  & \new_[52731]_ ;
  assign \new_[1771]_  = \new_[52720]_  & \new_[52707]_ ;
  assign \new_[1772]_  = \new_[52696]_  & \new_[52683]_ ;
  assign \new_[1773]_  = \new_[52672]_  & \new_[52659]_ ;
  assign \new_[1774]_  = \new_[52648]_  & \new_[52635]_ ;
  assign \new_[1775]_  = \new_[52624]_  & \new_[52611]_ ;
  assign \new_[1776]_  = \new_[52600]_  & \new_[52587]_ ;
  assign \new_[1777]_  = \new_[52576]_  & \new_[52563]_ ;
  assign \new_[1778]_  = \new_[52552]_  & \new_[52539]_ ;
  assign \new_[1779]_  = \new_[52528]_  & \new_[52515]_ ;
  assign \new_[1780]_  = \new_[52504]_  & \new_[52491]_ ;
  assign \new_[1781]_  = \new_[52480]_  & \new_[52467]_ ;
  assign \new_[1782]_  = \new_[52456]_  & \new_[52443]_ ;
  assign \new_[1783]_  = \new_[52432]_  & \new_[52419]_ ;
  assign \new_[1784]_  = \new_[52408]_  & \new_[52395]_ ;
  assign \new_[1785]_  = \new_[52384]_  & \new_[52371]_ ;
  assign \new_[1786]_  = \new_[52360]_  & \new_[52347]_ ;
  assign \new_[1787]_  = \new_[52336]_  & \new_[52323]_ ;
  assign \new_[1788]_  = \new_[52312]_  & \new_[52299]_ ;
  assign \new_[1789]_  = \new_[52288]_  & \new_[52275]_ ;
  assign \new_[1790]_  = \new_[52264]_  & \new_[52251]_ ;
  assign \new_[1791]_  = \new_[52240]_  & \new_[52227]_ ;
  assign \new_[1792]_  = \new_[52216]_  & \new_[52203]_ ;
  assign \new_[1793]_  = \new_[52192]_  & \new_[52179]_ ;
  assign \new_[1794]_  = \new_[52168]_  & \new_[52155]_ ;
  assign \new_[1795]_  = \new_[52144]_  & \new_[52131]_ ;
  assign \new_[1796]_  = \new_[52120]_  & \new_[52107]_ ;
  assign \new_[1797]_  = \new_[52096]_  & \new_[52083]_ ;
  assign \new_[1798]_  = \new_[52072]_  & \new_[52059]_ ;
  assign \new_[1799]_  = \new_[52048]_  & \new_[52035]_ ;
  assign \new_[1800]_  = \new_[52024]_  & \new_[52011]_ ;
  assign \new_[1801]_  = \new_[52000]_  & \new_[51987]_ ;
  assign \new_[1802]_  = \new_[51976]_  & \new_[51963]_ ;
  assign \new_[1803]_  = \new_[51952]_  & \new_[51939]_ ;
  assign \new_[1804]_  = \new_[51928]_  & \new_[51915]_ ;
  assign \new_[1805]_  = \new_[51904]_  & \new_[51891]_ ;
  assign \new_[1806]_  = \new_[51880]_  & \new_[51867]_ ;
  assign \new_[1807]_  = \new_[51856]_  & \new_[51843]_ ;
  assign \new_[1808]_  = \new_[51832]_  & \new_[51819]_ ;
  assign \new_[1809]_  = \new_[51808]_  & \new_[51795]_ ;
  assign \new_[1810]_  = \new_[51784]_  & \new_[51771]_ ;
  assign \new_[1811]_  = \new_[51760]_  & \new_[51747]_ ;
  assign \new_[1812]_  = \new_[51736]_  & \new_[51723]_ ;
  assign \new_[1813]_  = \new_[51712]_  & \new_[51699]_ ;
  assign \new_[1814]_  = \new_[51688]_  & \new_[51675]_ ;
  assign \new_[1815]_  = \new_[51664]_  & \new_[51651]_ ;
  assign \new_[1816]_  = \new_[51640]_  & \new_[51627]_ ;
  assign \new_[1817]_  = \new_[51616]_  & \new_[51603]_ ;
  assign \new_[1818]_  = \new_[51592]_  & \new_[51579]_ ;
  assign \new_[1819]_  = \new_[51568]_  & \new_[51555]_ ;
  assign \new_[1820]_  = \new_[51544]_  & \new_[51531]_ ;
  assign \new_[1821]_  = \new_[51520]_  & \new_[51507]_ ;
  assign \new_[1822]_  = \new_[51496]_  & \new_[51483]_ ;
  assign \new_[1823]_  = \new_[51472]_  & \new_[51459]_ ;
  assign \new_[1824]_  = \new_[51448]_  & \new_[51435]_ ;
  assign \new_[1825]_  = \new_[51424]_  & \new_[51411]_ ;
  assign \new_[1826]_  = \new_[51400]_  & \new_[51387]_ ;
  assign \new_[1827]_  = \new_[51376]_  & \new_[51363]_ ;
  assign \new_[1828]_  = \new_[51352]_  & \new_[51339]_ ;
  assign \new_[1829]_  = \new_[51328]_  & \new_[51315]_ ;
  assign \new_[1830]_  = \new_[51304]_  & \new_[51291]_ ;
  assign \new_[1831]_  = \new_[51280]_  & \new_[51267]_ ;
  assign \new_[1832]_  = \new_[51256]_  & \new_[51243]_ ;
  assign \new_[1833]_  = \new_[51232]_  & \new_[51219]_ ;
  assign \new_[1834]_  = \new_[51208]_  & \new_[51195]_ ;
  assign \new_[1835]_  = \new_[51184]_  & \new_[51171]_ ;
  assign \new_[1836]_  = \new_[51160]_  & \new_[51147]_ ;
  assign \new_[1837]_  = \new_[51136]_  & \new_[51123]_ ;
  assign \new_[1838]_  = \new_[51112]_  & \new_[51099]_ ;
  assign \new_[1839]_  = \new_[51088]_  & \new_[51075]_ ;
  assign \new_[1840]_  = \new_[51064]_  & \new_[51051]_ ;
  assign \new_[1841]_  = \new_[51040]_  & \new_[51027]_ ;
  assign \new_[1842]_  = \new_[51016]_  & \new_[51003]_ ;
  assign \new_[1843]_  = \new_[50992]_  & \new_[50979]_ ;
  assign \new_[1844]_  = \new_[50968]_  & \new_[50955]_ ;
  assign \new_[1845]_  = \new_[50944]_  & \new_[50931]_ ;
  assign \new_[1846]_  = \new_[50920]_  & \new_[50907]_ ;
  assign \new_[1847]_  = \new_[50896]_  & \new_[50883]_ ;
  assign \new_[1848]_  = \new_[50872]_  & \new_[50859]_ ;
  assign \new_[1849]_  = \new_[50848]_  & \new_[50835]_ ;
  assign \new_[1850]_  = \new_[50824]_  & \new_[50811]_ ;
  assign \new_[1851]_  = \new_[50800]_  & \new_[50787]_ ;
  assign \new_[1852]_  = \new_[50776]_  & \new_[50763]_ ;
  assign \new_[1853]_  = \new_[50752]_  & \new_[50739]_ ;
  assign \new_[1854]_  = \new_[50728]_  & \new_[50715]_ ;
  assign \new_[1855]_  = \new_[50704]_  & \new_[50691]_ ;
  assign \new_[1856]_  = \new_[50680]_  & \new_[50667]_ ;
  assign \new_[1857]_  = \new_[50656]_  & \new_[50643]_ ;
  assign \new_[1858]_  = \new_[50632]_  & \new_[50619]_ ;
  assign \new_[1859]_  = \new_[50608]_  & \new_[50595]_ ;
  assign \new_[1860]_  = \new_[50584]_  & \new_[50571]_ ;
  assign \new_[1861]_  = \new_[50560]_  & \new_[50547]_ ;
  assign \new_[1862]_  = \new_[50536]_  & \new_[50523]_ ;
  assign \new_[1863]_  = \new_[50512]_  & \new_[50499]_ ;
  assign \new_[1864]_  = \new_[50488]_  & \new_[50475]_ ;
  assign \new_[1865]_  = \new_[50464]_  & \new_[50451]_ ;
  assign \new_[1866]_  = \new_[50440]_  & \new_[50427]_ ;
  assign \new_[1867]_  = \new_[50416]_  & \new_[50403]_ ;
  assign \new_[1868]_  = \new_[50392]_  & \new_[50379]_ ;
  assign \new_[1869]_  = \new_[50368]_  & \new_[50355]_ ;
  assign \new_[1870]_  = \new_[50344]_  & \new_[50331]_ ;
  assign \new_[1871]_  = \new_[50320]_  & \new_[50307]_ ;
  assign \new_[1872]_  = \new_[50296]_  & \new_[50283]_ ;
  assign \new_[1873]_  = \new_[50272]_  & \new_[50259]_ ;
  assign \new_[1874]_  = \new_[50248]_  & \new_[50235]_ ;
  assign \new_[1875]_  = \new_[50224]_  & \new_[50211]_ ;
  assign \new_[1876]_  = \new_[50200]_  & \new_[50187]_ ;
  assign \new_[1877]_  = \new_[50176]_  & \new_[50163]_ ;
  assign \new_[1878]_  = \new_[50152]_  & \new_[50139]_ ;
  assign \new_[1879]_  = \new_[50128]_  & \new_[50115]_ ;
  assign \new_[1880]_  = \new_[50104]_  & \new_[50091]_ ;
  assign \new_[1881]_  = \new_[50080]_  & \new_[50067]_ ;
  assign \new_[1882]_  = \new_[50056]_  & \new_[50043]_ ;
  assign \new_[1883]_  = \new_[50032]_  & \new_[50019]_ ;
  assign \new_[1884]_  = \new_[50008]_  & \new_[49995]_ ;
  assign \new_[1885]_  = \new_[49984]_  & \new_[49971]_ ;
  assign \new_[1886]_  = \new_[49960]_  & \new_[49947]_ ;
  assign \new_[1887]_  = \new_[49936]_  & \new_[49923]_ ;
  assign \new_[1888]_  = \new_[49912]_  & \new_[49899]_ ;
  assign \new_[1889]_  = \new_[49888]_  & \new_[49875]_ ;
  assign \new_[1890]_  = \new_[49864]_  & \new_[49851]_ ;
  assign \new_[1891]_  = \new_[49840]_  & \new_[49827]_ ;
  assign \new_[1892]_  = \new_[49816]_  & \new_[49803]_ ;
  assign \new_[1893]_  = \new_[49792]_  & \new_[49779]_ ;
  assign \new_[1894]_  = \new_[49768]_  & \new_[49755]_ ;
  assign \new_[1895]_  = \new_[49744]_  & \new_[49731]_ ;
  assign \new_[1896]_  = \new_[49720]_  & \new_[49707]_ ;
  assign \new_[1897]_  = \new_[49696]_  & \new_[49683]_ ;
  assign \new_[1898]_  = \new_[49672]_  & \new_[49659]_ ;
  assign \new_[1899]_  = \new_[49648]_  & \new_[49635]_ ;
  assign \new_[1900]_  = \new_[49624]_  & \new_[49611]_ ;
  assign \new_[1901]_  = \new_[49600]_  & \new_[49587]_ ;
  assign \new_[1902]_  = \new_[49576]_  & \new_[49563]_ ;
  assign \new_[1903]_  = \new_[49552]_  & \new_[49539]_ ;
  assign \new_[1904]_  = \new_[49528]_  & \new_[49515]_ ;
  assign \new_[1905]_  = \new_[49504]_  & \new_[49491]_ ;
  assign \new_[1906]_  = \new_[49480]_  & \new_[49467]_ ;
  assign \new_[1907]_  = \new_[49456]_  & \new_[49443]_ ;
  assign \new_[1908]_  = \new_[49432]_  & \new_[49419]_ ;
  assign \new_[1909]_  = \new_[49408]_  & \new_[49395]_ ;
  assign \new_[1910]_  = \new_[49384]_  & \new_[49371]_ ;
  assign \new_[1911]_  = \new_[49360]_  & \new_[49347]_ ;
  assign \new_[1912]_  = \new_[49336]_  & \new_[49323]_ ;
  assign \new_[1913]_  = \new_[49312]_  & \new_[49299]_ ;
  assign \new_[1914]_  = \new_[49288]_  & \new_[49275]_ ;
  assign \new_[1915]_  = \new_[49264]_  & \new_[49251]_ ;
  assign \new_[1916]_  = \new_[49240]_  & \new_[49227]_ ;
  assign \new_[1917]_  = \new_[49216]_  & \new_[49203]_ ;
  assign \new_[1918]_  = \new_[49192]_  & \new_[49179]_ ;
  assign \new_[1919]_  = \new_[49168]_  & \new_[49155]_ ;
  assign \new_[1920]_  = \new_[49144]_  & \new_[49131]_ ;
  assign \new_[1921]_  = \new_[49120]_  & \new_[49107]_ ;
  assign \new_[1922]_  = \new_[49096]_  & \new_[49083]_ ;
  assign \new_[1923]_  = \new_[49072]_  & \new_[49059]_ ;
  assign \new_[1924]_  = \new_[49048]_  & \new_[49035]_ ;
  assign \new_[1925]_  = \new_[49024]_  & \new_[49011]_ ;
  assign \new_[1926]_  = \new_[49000]_  & \new_[48987]_ ;
  assign \new_[1927]_  = \new_[48976]_  & \new_[48963]_ ;
  assign \new_[1928]_  = \new_[48952]_  & \new_[48939]_ ;
  assign \new_[1929]_  = \new_[48928]_  & \new_[48915]_ ;
  assign \new_[1930]_  = \new_[48904]_  & \new_[48891]_ ;
  assign \new_[1931]_  = \new_[48880]_  & \new_[48867]_ ;
  assign \new_[1932]_  = \new_[48856]_  & \new_[48843]_ ;
  assign \new_[1933]_  = \new_[48832]_  & \new_[48819]_ ;
  assign \new_[1934]_  = \new_[48808]_  & \new_[48795]_ ;
  assign \new_[1935]_  = \new_[48784]_  & \new_[48771]_ ;
  assign \new_[1936]_  = \new_[48760]_  & \new_[48747]_ ;
  assign \new_[1937]_  = \new_[48736]_  & \new_[48723]_ ;
  assign \new_[1938]_  = \new_[48712]_  & \new_[48699]_ ;
  assign \new_[1939]_  = \new_[48688]_  & \new_[48675]_ ;
  assign \new_[1940]_  = \new_[48664]_  & \new_[48651]_ ;
  assign \new_[1941]_  = \new_[48640]_  & \new_[48627]_ ;
  assign \new_[1942]_  = \new_[48616]_  & \new_[48603]_ ;
  assign \new_[1943]_  = \new_[48592]_  & \new_[48579]_ ;
  assign \new_[1944]_  = \new_[48568]_  & \new_[48555]_ ;
  assign \new_[1945]_  = \new_[48544]_  & \new_[48531]_ ;
  assign \new_[1946]_  = \new_[48520]_  & \new_[48507]_ ;
  assign \new_[1947]_  = \new_[48496]_  & \new_[48483]_ ;
  assign \new_[1948]_  = \new_[48472]_  & \new_[48459]_ ;
  assign \new_[1949]_  = \new_[48448]_  & \new_[48435]_ ;
  assign \new_[1950]_  = \new_[48424]_  & \new_[48411]_ ;
  assign \new_[1951]_  = \new_[48400]_  & \new_[48387]_ ;
  assign \new_[1952]_  = \new_[48376]_  & \new_[48363]_ ;
  assign \new_[1953]_  = \new_[48352]_  & \new_[48339]_ ;
  assign \new_[1954]_  = \new_[48328]_  & \new_[48315]_ ;
  assign \new_[1955]_  = \new_[48304]_  & \new_[48291]_ ;
  assign \new_[1956]_  = \new_[48280]_  & \new_[48267]_ ;
  assign \new_[1957]_  = \new_[48256]_  & \new_[48243]_ ;
  assign \new_[1958]_  = \new_[48232]_  & \new_[48219]_ ;
  assign \new_[1959]_  = \new_[48208]_  & \new_[48195]_ ;
  assign \new_[1960]_  = \new_[48184]_  & \new_[48171]_ ;
  assign \new_[1961]_  = \new_[48160]_  & \new_[48147]_ ;
  assign \new_[1962]_  = \new_[48136]_  & \new_[48123]_ ;
  assign \new_[1963]_  = \new_[48112]_  & \new_[48099]_ ;
  assign \new_[1964]_  = \new_[48088]_  & \new_[48075]_ ;
  assign \new_[1965]_  = \new_[48064]_  & \new_[48051]_ ;
  assign \new_[1966]_  = \new_[48040]_  & \new_[48027]_ ;
  assign \new_[1967]_  = \new_[48016]_  & \new_[48003]_ ;
  assign \new_[1968]_  = \new_[47992]_  & \new_[47979]_ ;
  assign \new_[1969]_  = \new_[47968]_  & \new_[47955]_ ;
  assign \new_[1970]_  = \new_[47944]_  & \new_[47931]_ ;
  assign \new_[1971]_  = \new_[47920]_  & \new_[47907]_ ;
  assign \new_[1972]_  = \new_[47896]_  & \new_[47883]_ ;
  assign \new_[1973]_  = \new_[47872]_  & \new_[47859]_ ;
  assign \new_[1974]_  = \new_[47848]_  & \new_[47835]_ ;
  assign \new_[1975]_  = \new_[47824]_  & \new_[47811]_ ;
  assign \new_[1976]_  = \new_[47800]_  & \new_[47787]_ ;
  assign \new_[1977]_  = \new_[47776]_  & \new_[47763]_ ;
  assign \new_[1978]_  = \new_[47752]_  & \new_[47739]_ ;
  assign \new_[1979]_  = \new_[47728]_  & \new_[47715]_ ;
  assign \new_[1980]_  = \new_[47704]_  & \new_[47691]_ ;
  assign \new_[1981]_  = \new_[47680]_  & \new_[47667]_ ;
  assign \new_[1982]_  = \new_[47656]_  & \new_[47643]_ ;
  assign \new_[1983]_  = \new_[47632]_  & \new_[47619]_ ;
  assign \new_[1984]_  = \new_[47608]_  & \new_[47595]_ ;
  assign \new_[1985]_  = \new_[47584]_  & \new_[47571]_ ;
  assign \new_[1986]_  = \new_[47560]_  & \new_[47547]_ ;
  assign \new_[1987]_  = \new_[47536]_  & \new_[47523]_ ;
  assign \new_[1988]_  = \new_[47512]_  & \new_[47499]_ ;
  assign \new_[1989]_  = \new_[47488]_  & \new_[47475]_ ;
  assign \new_[1990]_  = \new_[47464]_  & \new_[47451]_ ;
  assign \new_[1991]_  = \new_[47440]_  & \new_[47427]_ ;
  assign \new_[1992]_  = \new_[47416]_  & \new_[47403]_ ;
  assign \new_[1993]_  = \new_[47392]_  & \new_[47379]_ ;
  assign \new_[1994]_  = \new_[47368]_  & \new_[47355]_ ;
  assign \new_[1995]_  = \new_[47344]_  & \new_[47331]_ ;
  assign \new_[1996]_  = \new_[47320]_  & \new_[47307]_ ;
  assign \new_[1997]_  = \new_[47296]_  & \new_[47283]_ ;
  assign \new_[1998]_  = \new_[47272]_  & \new_[47259]_ ;
  assign \new_[1999]_  = \new_[47248]_  & \new_[47235]_ ;
  assign \new_[2000]_  = \new_[47224]_  & \new_[47211]_ ;
  assign \new_[2001]_  = \new_[47200]_  & \new_[47187]_ ;
  assign \new_[2002]_  = \new_[47176]_  & \new_[47163]_ ;
  assign \new_[2003]_  = \new_[47152]_  & \new_[47139]_ ;
  assign \new_[2004]_  = \new_[47128]_  & \new_[47115]_ ;
  assign \new_[2005]_  = \new_[47104]_  & \new_[47091]_ ;
  assign \new_[2006]_  = \new_[47080]_  & \new_[47067]_ ;
  assign \new_[2007]_  = \new_[47056]_  & \new_[47043]_ ;
  assign \new_[2008]_  = \new_[47032]_  & \new_[47019]_ ;
  assign \new_[2009]_  = \new_[47008]_  & \new_[46995]_ ;
  assign \new_[2010]_  = \new_[46984]_  & \new_[46971]_ ;
  assign \new_[2011]_  = \new_[46960]_  & \new_[46947]_ ;
  assign \new_[2012]_  = \new_[46936]_  & \new_[46923]_ ;
  assign \new_[2013]_  = \new_[46912]_  & \new_[46899]_ ;
  assign \new_[2014]_  = \new_[46888]_  & \new_[46875]_ ;
  assign \new_[2015]_  = \new_[46864]_  & \new_[46851]_ ;
  assign \new_[2016]_  = \new_[46840]_  & \new_[46827]_ ;
  assign \new_[2017]_  = \new_[46816]_  & \new_[46803]_ ;
  assign \new_[2018]_  = \new_[46792]_  & \new_[46779]_ ;
  assign \new_[2019]_  = \new_[46768]_  & \new_[46755]_ ;
  assign \new_[2020]_  = \new_[46744]_  & \new_[46731]_ ;
  assign \new_[2021]_  = \new_[46720]_  & \new_[46707]_ ;
  assign \new_[2022]_  = \new_[46696]_  & \new_[46683]_ ;
  assign \new_[2023]_  = \new_[46672]_  & \new_[46659]_ ;
  assign \new_[2024]_  = \new_[46648]_  & \new_[46635]_ ;
  assign \new_[2025]_  = \new_[46624]_  & \new_[46611]_ ;
  assign \new_[2026]_  = \new_[46600]_  & \new_[46587]_ ;
  assign \new_[2027]_  = \new_[46576]_  & \new_[46563]_ ;
  assign \new_[2028]_  = \new_[46552]_  & \new_[46539]_ ;
  assign \new_[2029]_  = \new_[46528]_  & \new_[46515]_ ;
  assign \new_[2030]_  = \new_[46504]_  & \new_[46491]_ ;
  assign \new_[2031]_  = \new_[46480]_  & \new_[46467]_ ;
  assign \new_[2032]_  = \new_[46456]_  & \new_[46443]_ ;
  assign \new_[2033]_  = \new_[46432]_  & \new_[46419]_ ;
  assign \new_[2034]_  = \new_[46408]_  & \new_[46395]_ ;
  assign \new_[2035]_  = \new_[46384]_  & \new_[46371]_ ;
  assign \new_[2036]_  = \new_[46360]_  & \new_[46347]_ ;
  assign \new_[2037]_  = \new_[46336]_  & \new_[46323]_ ;
  assign \new_[2038]_  = \new_[46312]_  & \new_[46299]_ ;
  assign \new_[2039]_  = \new_[46288]_  & \new_[46275]_ ;
  assign \new_[2040]_  = \new_[46264]_  & \new_[46251]_ ;
  assign \new_[2041]_  = \new_[46240]_  & \new_[46227]_ ;
  assign \new_[2042]_  = \new_[46216]_  & \new_[46203]_ ;
  assign \new_[2043]_  = \new_[46192]_  & \new_[46179]_ ;
  assign \new_[2044]_  = \new_[46168]_  & \new_[46155]_ ;
  assign \new_[2045]_  = \new_[46144]_  & \new_[46131]_ ;
  assign \new_[2046]_  = \new_[46120]_  & \new_[46107]_ ;
  assign \new_[2047]_  = \new_[46096]_  & \new_[46083]_ ;
  assign \new_[2048]_  = \new_[46072]_  & \new_[46059]_ ;
  assign \new_[2049]_  = \new_[46048]_  & \new_[46035]_ ;
  assign \new_[2050]_  = \new_[46024]_  & \new_[46011]_ ;
  assign \new_[2051]_  = \new_[46000]_  & \new_[45987]_ ;
  assign \new_[2052]_  = \new_[45976]_  & \new_[45963]_ ;
  assign \new_[2053]_  = \new_[45952]_  & \new_[45939]_ ;
  assign \new_[2054]_  = \new_[45928]_  & \new_[45915]_ ;
  assign \new_[2055]_  = \new_[45904]_  & \new_[45891]_ ;
  assign \new_[2056]_  = \new_[45880]_  & \new_[45867]_ ;
  assign \new_[2057]_  = \new_[45856]_  & \new_[45843]_ ;
  assign \new_[2058]_  = \new_[45832]_  & \new_[45819]_ ;
  assign \new_[2059]_  = \new_[45808]_  & \new_[45795]_ ;
  assign \new_[2060]_  = \new_[45784]_  & \new_[45771]_ ;
  assign \new_[2061]_  = \new_[45760]_  & \new_[45747]_ ;
  assign \new_[2062]_  = \new_[45736]_  & \new_[45723]_ ;
  assign \new_[2063]_  = \new_[45712]_  & \new_[45699]_ ;
  assign \new_[2064]_  = \new_[45688]_  & \new_[45675]_ ;
  assign \new_[2065]_  = \new_[45664]_  & \new_[45651]_ ;
  assign \new_[2066]_  = \new_[45640]_  & \new_[45627]_ ;
  assign \new_[2067]_  = \new_[45616]_  & \new_[45603]_ ;
  assign \new_[2068]_  = \new_[45592]_  & \new_[45579]_ ;
  assign \new_[2069]_  = \new_[45568]_  & \new_[45555]_ ;
  assign \new_[2070]_  = \new_[45544]_  & \new_[45531]_ ;
  assign \new_[2071]_  = \new_[45520]_  & \new_[45507]_ ;
  assign \new_[2072]_  = \new_[45496]_  & \new_[45483]_ ;
  assign \new_[2073]_  = \new_[45472]_  & \new_[45459]_ ;
  assign \new_[2074]_  = \new_[45448]_  & \new_[45435]_ ;
  assign \new_[2075]_  = \new_[45424]_  & \new_[45411]_ ;
  assign \new_[2076]_  = \new_[45400]_  & \new_[45387]_ ;
  assign \new_[2077]_  = \new_[45376]_  & \new_[45363]_ ;
  assign \new_[2078]_  = \new_[45352]_  & \new_[45339]_ ;
  assign \new_[2079]_  = \new_[45328]_  & \new_[45315]_ ;
  assign \new_[2080]_  = \new_[45304]_  & \new_[45291]_ ;
  assign \new_[2081]_  = \new_[45280]_  & \new_[45267]_ ;
  assign \new_[2082]_  = \new_[45256]_  & \new_[45243]_ ;
  assign \new_[2083]_  = \new_[45232]_  & \new_[45219]_ ;
  assign \new_[2084]_  = \new_[45208]_  & \new_[45195]_ ;
  assign \new_[2085]_  = \new_[45184]_  & \new_[45171]_ ;
  assign \new_[2086]_  = \new_[45160]_  & \new_[45147]_ ;
  assign \new_[2087]_  = \new_[45136]_  & \new_[45123]_ ;
  assign \new_[2088]_  = \new_[45112]_  & \new_[45099]_ ;
  assign \new_[2089]_  = \new_[45088]_  & \new_[45075]_ ;
  assign \new_[2090]_  = \new_[45064]_  & \new_[45051]_ ;
  assign \new_[2091]_  = \new_[45040]_  & \new_[45027]_ ;
  assign \new_[2092]_  = \new_[45016]_  & \new_[45003]_ ;
  assign \new_[2093]_  = \new_[44992]_  & \new_[44979]_ ;
  assign \new_[2094]_  = \new_[44968]_  & \new_[44955]_ ;
  assign \new_[2095]_  = \new_[44944]_  & \new_[44931]_ ;
  assign \new_[2096]_  = \new_[44920]_  & \new_[44907]_ ;
  assign \new_[2097]_  = \new_[44896]_  & \new_[44883]_ ;
  assign \new_[2098]_  = \new_[44872]_  & \new_[44859]_ ;
  assign \new_[2099]_  = \new_[44848]_  & \new_[44835]_ ;
  assign \new_[2100]_  = \new_[44824]_  & \new_[44811]_ ;
  assign \new_[2101]_  = \new_[44800]_  & \new_[44787]_ ;
  assign \new_[2102]_  = \new_[44776]_  & \new_[44763]_ ;
  assign \new_[2103]_  = \new_[44752]_  & \new_[44739]_ ;
  assign \new_[2104]_  = \new_[44728]_  & \new_[44715]_ ;
  assign \new_[2105]_  = \new_[44704]_  & \new_[44691]_ ;
  assign \new_[2106]_  = \new_[44680]_  & \new_[44667]_ ;
  assign \new_[2107]_  = \new_[44656]_  & \new_[44643]_ ;
  assign \new_[2108]_  = \new_[44632]_  & \new_[44619]_ ;
  assign \new_[2109]_  = \new_[44608]_  & \new_[44595]_ ;
  assign \new_[2110]_  = \new_[44584]_  & \new_[44571]_ ;
  assign \new_[2111]_  = \new_[44560]_  & \new_[44547]_ ;
  assign \new_[2112]_  = \new_[44536]_  & \new_[44523]_ ;
  assign \new_[2113]_  = \new_[44512]_  & \new_[44499]_ ;
  assign \new_[2114]_  = \new_[44488]_  & \new_[44475]_ ;
  assign \new_[2115]_  = \new_[44464]_  & \new_[44451]_ ;
  assign \new_[2116]_  = \new_[44440]_  & \new_[44427]_ ;
  assign \new_[2117]_  = \new_[44416]_  & \new_[44403]_ ;
  assign \new_[2118]_  = \new_[44392]_  & \new_[44379]_ ;
  assign \new_[2119]_  = \new_[44368]_  & \new_[44355]_ ;
  assign \new_[2120]_  = \new_[44344]_  & \new_[44331]_ ;
  assign \new_[2121]_  = \new_[44320]_  & \new_[44307]_ ;
  assign \new_[2122]_  = \new_[44296]_  & \new_[44283]_ ;
  assign \new_[2123]_  = \new_[44272]_  & \new_[44259]_ ;
  assign \new_[2124]_  = \new_[44248]_  & \new_[44235]_ ;
  assign \new_[2125]_  = \new_[44224]_  & \new_[44211]_ ;
  assign \new_[2126]_  = \new_[44200]_  & \new_[44187]_ ;
  assign \new_[2127]_  = \new_[44176]_  & \new_[44163]_ ;
  assign \new_[2128]_  = \new_[44152]_  & \new_[44139]_ ;
  assign \new_[2129]_  = \new_[44128]_  & \new_[44115]_ ;
  assign \new_[2130]_  = \new_[44104]_  & \new_[44091]_ ;
  assign \new_[2131]_  = \new_[44080]_  & \new_[44067]_ ;
  assign \new_[2132]_  = \new_[44056]_  & \new_[44043]_ ;
  assign \new_[2133]_  = \new_[44032]_  & \new_[44019]_ ;
  assign \new_[2134]_  = \new_[44008]_  & \new_[43995]_ ;
  assign \new_[2135]_  = \new_[43984]_  & \new_[43971]_ ;
  assign \new_[2136]_  = \new_[43960]_  & \new_[43947]_ ;
  assign \new_[2137]_  = \new_[43936]_  & \new_[43923]_ ;
  assign \new_[2138]_  = \new_[43912]_  & \new_[43899]_ ;
  assign \new_[2139]_  = \new_[43888]_  & \new_[43875]_ ;
  assign \new_[2140]_  = \new_[43864]_  & \new_[43851]_ ;
  assign \new_[2141]_  = \new_[43840]_  & \new_[43827]_ ;
  assign \new_[2142]_  = \new_[43816]_  & \new_[43803]_ ;
  assign \new_[2143]_  = \new_[43792]_  & \new_[43779]_ ;
  assign \new_[2144]_  = \new_[43768]_  & \new_[43755]_ ;
  assign \new_[2145]_  = \new_[43744]_  & \new_[43731]_ ;
  assign \new_[2146]_  = \new_[43720]_  & \new_[43707]_ ;
  assign \new_[2147]_  = \new_[43696]_  & \new_[43683]_ ;
  assign \new_[2148]_  = \new_[43672]_  & \new_[43659]_ ;
  assign \new_[2149]_  = \new_[43648]_  & \new_[43635]_ ;
  assign \new_[2150]_  = \new_[43624]_  & \new_[43611]_ ;
  assign \new_[2151]_  = \new_[43600]_  & \new_[43587]_ ;
  assign \new_[2152]_  = \new_[43576]_  & \new_[43563]_ ;
  assign \new_[2153]_  = \new_[43552]_  & \new_[43539]_ ;
  assign \new_[2154]_  = \new_[43528]_  & \new_[43515]_ ;
  assign \new_[2155]_  = \new_[43504]_  & \new_[43491]_ ;
  assign \new_[2156]_  = \new_[43480]_  & \new_[43467]_ ;
  assign \new_[2157]_  = \new_[43456]_  & \new_[43443]_ ;
  assign \new_[2158]_  = \new_[43432]_  & \new_[43419]_ ;
  assign \new_[2159]_  = \new_[43408]_  & \new_[43395]_ ;
  assign \new_[2160]_  = \new_[43384]_  & \new_[43371]_ ;
  assign \new_[2161]_  = \new_[43360]_  & \new_[43347]_ ;
  assign \new_[2162]_  = \new_[43336]_  & \new_[43323]_ ;
  assign \new_[2163]_  = \new_[43312]_  & \new_[43299]_ ;
  assign \new_[2164]_  = \new_[43288]_  & \new_[43275]_ ;
  assign \new_[2165]_  = \new_[43264]_  & \new_[43251]_ ;
  assign \new_[2166]_  = \new_[43240]_  & \new_[43227]_ ;
  assign \new_[2167]_  = \new_[43216]_  & \new_[43203]_ ;
  assign \new_[2168]_  = \new_[43192]_  & \new_[43179]_ ;
  assign \new_[2169]_  = \new_[43168]_  & \new_[43155]_ ;
  assign \new_[2170]_  = \new_[43144]_  & \new_[43131]_ ;
  assign \new_[2171]_  = \new_[43120]_  & \new_[43107]_ ;
  assign \new_[2172]_  = \new_[43096]_  & \new_[43083]_ ;
  assign \new_[2173]_  = \new_[43072]_  & \new_[43059]_ ;
  assign \new_[2174]_  = \new_[43048]_  & \new_[43035]_ ;
  assign \new_[2175]_  = \new_[43024]_  & \new_[43011]_ ;
  assign \new_[2176]_  = \new_[43000]_  & \new_[42987]_ ;
  assign \new_[2177]_  = \new_[42976]_  & \new_[42963]_ ;
  assign \new_[2178]_  = \new_[42952]_  & \new_[42939]_ ;
  assign \new_[2179]_  = \new_[42928]_  & \new_[42915]_ ;
  assign \new_[2180]_  = \new_[42904]_  & \new_[42891]_ ;
  assign \new_[2181]_  = \new_[42880]_  & \new_[42867]_ ;
  assign \new_[2182]_  = \new_[42856]_  & \new_[42843]_ ;
  assign \new_[2183]_  = \new_[42832]_  & \new_[42819]_ ;
  assign \new_[2184]_  = \new_[42808]_  & \new_[42795]_ ;
  assign \new_[2185]_  = \new_[42784]_  & \new_[42771]_ ;
  assign \new_[2186]_  = \new_[42760]_  & \new_[42747]_ ;
  assign \new_[2187]_  = \new_[42736]_  & \new_[42723]_ ;
  assign \new_[2188]_  = \new_[42712]_  & \new_[42699]_ ;
  assign \new_[2189]_  = \new_[42688]_  & \new_[42675]_ ;
  assign \new_[2190]_  = \new_[42664]_  & \new_[42651]_ ;
  assign \new_[2191]_  = \new_[42640]_  & \new_[42627]_ ;
  assign \new_[2192]_  = \new_[42616]_  & \new_[42603]_ ;
  assign \new_[2193]_  = \new_[42592]_  & \new_[42579]_ ;
  assign \new_[2194]_  = \new_[42568]_  & \new_[42555]_ ;
  assign \new_[2195]_  = \new_[42544]_  & \new_[42531]_ ;
  assign \new_[2196]_  = \new_[42520]_  & \new_[42507]_ ;
  assign \new_[2197]_  = \new_[42496]_  & \new_[42483]_ ;
  assign \new_[2198]_  = \new_[42472]_  & \new_[42459]_ ;
  assign \new_[2199]_  = \new_[42448]_  & \new_[42435]_ ;
  assign \new_[2200]_  = \new_[42424]_  & \new_[42411]_ ;
  assign \new_[2201]_  = \new_[42400]_  & \new_[42387]_ ;
  assign \new_[2202]_  = \new_[42376]_  & \new_[42363]_ ;
  assign \new_[2203]_  = \new_[42352]_  & \new_[42339]_ ;
  assign \new_[2204]_  = \new_[42328]_  & \new_[42315]_ ;
  assign \new_[2205]_  = \new_[42304]_  & \new_[42291]_ ;
  assign \new_[2206]_  = \new_[42280]_  & \new_[42267]_ ;
  assign \new_[2207]_  = \new_[42256]_  & \new_[42243]_ ;
  assign \new_[2208]_  = \new_[42232]_  & \new_[42219]_ ;
  assign \new_[2209]_  = \new_[42208]_  & \new_[42195]_ ;
  assign \new_[2210]_  = \new_[42184]_  & \new_[42171]_ ;
  assign \new_[2211]_  = \new_[42160]_  & \new_[42147]_ ;
  assign \new_[2212]_  = \new_[42136]_  & \new_[42123]_ ;
  assign \new_[2213]_  = \new_[42112]_  & \new_[42099]_ ;
  assign \new_[2214]_  = \new_[42088]_  & \new_[42075]_ ;
  assign \new_[2215]_  = \new_[42064]_  & \new_[42051]_ ;
  assign \new_[2216]_  = \new_[42040]_  & \new_[42027]_ ;
  assign \new_[2217]_  = \new_[42016]_  & \new_[42003]_ ;
  assign \new_[2218]_  = \new_[41992]_  & \new_[41979]_ ;
  assign \new_[2219]_  = \new_[41968]_  & \new_[41955]_ ;
  assign \new_[2220]_  = \new_[41944]_  & \new_[41931]_ ;
  assign \new_[2221]_  = \new_[41920]_  & \new_[41907]_ ;
  assign \new_[2222]_  = \new_[41896]_  & \new_[41883]_ ;
  assign \new_[2223]_  = \new_[41872]_  & \new_[41859]_ ;
  assign \new_[2224]_  = \new_[41848]_  & \new_[41835]_ ;
  assign \new_[2225]_  = \new_[41824]_  & \new_[41811]_ ;
  assign \new_[2226]_  = \new_[41800]_  & \new_[41787]_ ;
  assign \new_[2227]_  = \new_[41776]_  & \new_[41763]_ ;
  assign \new_[2228]_  = \new_[41752]_  & \new_[41739]_ ;
  assign \new_[2229]_  = \new_[41728]_  & \new_[41715]_ ;
  assign \new_[2230]_  = \new_[41704]_  & \new_[41691]_ ;
  assign \new_[2231]_  = \new_[41680]_  & \new_[41667]_ ;
  assign \new_[2232]_  = \new_[41656]_  & \new_[41643]_ ;
  assign \new_[2233]_  = \new_[41632]_  & \new_[41619]_ ;
  assign \new_[2234]_  = \new_[41608]_  & \new_[41595]_ ;
  assign \new_[2235]_  = \new_[41584]_  & \new_[41571]_ ;
  assign \new_[2236]_  = \new_[41560]_  & \new_[41547]_ ;
  assign \new_[2237]_  = \new_[41536]_  & \new_[41523]_ ;
  assign \new_[2238]_  = \new_[41512]_  & \new_[41499]_ ;
  assign \new_[2239]_  = \new_[41488]_  & \new_[41475]_ ;
  assign \new_[2240]_  = \new_[41464]_  & \new_[41451]_ ;
  assign \new_[2241]_  = \new_[41440]_  & \new_[41427]_ ;
  assign \new_[2242]_  = \new_[41416]_  & \new_[41403]_ ;
  assign \new_[2243]_  = \new_[41392]_  & \new_[41379]_ ;
  assign \new_[2244]_  = \new_[41368]_  & \new_[41355]_ ;
  assign \new_[2245]_  = \new_[41344]_  & \new_[41331]_ ;
  assign \new_[2246]_  = \new_[41320]_  & \new_[41307]_ ;
  assign \new_[2247]_  = \new_[41296]_  & \new_[41283]_ ;
  assign \new_[2248]_  = \new_[41272]_  & \new_[41259]_ ;
  assign \new_[2249]_  = \new_[41248]_  & \new_[41235]_ ;
  assign \new_[2250]_  = \new_[41224]_  & \new_[41211]_ ;
  assign \new_[2251]_  = \new_[41200]_  & \new_[41187]_ ;
  assign \new_[2252]_  = \new_[41176]_  & \new_[41163]_ ;
  assign \new_[2253]_  = \new_[41152]_  & \new_[41139]_ ;
  assign \new_[2254]_  = \new_[41128]_  & \new_[41115]_ ;
  assign \new_[2255]_  = \new_[41104]_  & \new_[41091]_ ;
  assign \new_[2256]_  = \new_[41080]_  & \new_[41067]_ ;
  assign \new_[2257]_  = \new_[41056]_  & \new_[41043]_ ;
  assign \new_[2258]_  = \new_[41032]_  & \new_[41019]_ ;
  assign \new_[2259]_  = \new_[41008]_  & \new_[40995]_ ;
  assign \new_[2260]_  = \new_[40984]_  & \new_[40971]_ ;
  assign \new_[2261]_  = \new_[40960]_  & \new_[40947]_ ;
  assign \new_[2262]_  = \new_[40936]_  & \new_[40923]_ ;
  assign \new_[2263]_  = \new_[40912]_  & \new_[40899]_ ;
  assign \new_[2264]_  = \new_[40888]_  & \new_[40875]_ ;
  assign \new_[2265]_  = \new_[40864]_  & \new_[40851]_ ;
  assign \new_[2266]_  = \new_[40840]_  & \new_[40827]_ ;
  assign \new_[2267]_  = \new_[40816]_  & \new_[40803]_ ;
  assign \new_[2268]_  = \new_[40792]_  & \new_[40779]_ ;
  assign \new_[2269]_  = \new_[40768]_  & \new_[40755]_ ;
  assign \new_[2270]_  = \new_[40744]_  & \new_[40731]_ ;
  assign \new_[2271]_  = \new_[40720]_  & \new_[40707]_ ;
  assign \new_[2272]_  = \new_[40696]_  & \new_[40683]_ ;
  assign \new_[2273]_  = \new_[40672]_  & \new_[40659]_ ;
  assign \new_[2274]_  = \new_[40648]_  & \new_[40635]_ ;
  assign \new_[2275]_  = \new_[40624]_  & \new_[40611]_ ;
  assign \new_[2276]_  = \new_[40600]_  & \new_[40587]_ ;
  assign \new_[2277]_  = \new_[40576]_  & \new_[40563]_ ;
  assign \new_[2278]_  = \new_[40552]_  & \new_[40539]_ ;
  assign \new_[2279]_  = \new_[40528]_  & \new_[40515]_ ;
  assign \new_[2280]_  = \new_[40504]_  & \new_[40491]_ ;
  assign \new_[2281]_  = \new_[40480]_  & \new_[40467]_ ;
  assign \new_[2282]_  = \new_[40456]_  & \new_[40443]_ ;
  assign \new_[2283]_  = \new_[40432]_  & \new_[40419]_ ;
  assign \new_[2284]_  = \new_[40408]_  & \new_[40395]_ ;
  assign \new_[2285]_  = \new_[40384]_  & \new_[40371]_ ;
  assign \new_[2286]_  = \new_[40360]_  & \new_[40347]_ ;
  assign \new_[2287]_  = \new_[40336]_  & \new_[40323]_ ;
  assign \new_[2288]_  = \new_[40312]_  & \new_[40299]_ ;
  assign \new_[2289]_  = \new_[40288]_  & \new_[40275]_ ;
  assign \new_[2290]_  = \new_[40264]_  & \new_[40251]_ ;
  assign \new_[2291]_  = \new_[40240]_  & \new_[40227]_ ;
  assign \new_[2292]_  = \new_[40216]_  & \new_[40203]_ ;
  assign \new_[2293]_  = \new_[40192]_  & \new_[40179]_ ;
  assign \new_[2294]_  = \new_[40168]_  & \new_[40155]_ ;
  assign \new_[2295]_  = \new_[40144]_  & \new_[40131]_ ;
  assign \new_[2296]_  = \new_[40120]_  & \new_[40107]_ ;
  assign \new_[2297]_  = \new_[40096]_  & \new_[40083]_ ;
  assign \new_[2298]_  = \new_[40072]_  & \new_[40059]_ ;
  assign \new_[2299]_  = \new_[40048]_  & \new_[40035]_ ;
  assign \new_[2300]_  = \new_[40024]_  & \new_[40011]_ ;
  assign \new_[2301]_  = \new_[40000]_  & \new_[39987]_ ;
  assign \new_[2302]_  = \new_[39976]_  & \new_[39963]_ ;
  assign \new_[2303]_  = \new_[39952]_  & \new_[39939]_ ;
  assign \new_[2304]_  = \new_[39928]_  & \new_[39915]_ ;
  assign \new_[2305]_  = \new_[39904]_  & \new_[39891]_ ;
  assign \new_[2306]_  = \new_[39880]_  & \new_[39867]_ ;
  assign \new_[2307]_  = \new_[39856]_  & \new_[39843]_ ;
  assign \new_[2308]_  = \new_[39832]_  & \new_[39819]_ ;
  assign \new_[2309]_  = \new_[39808]_  & \new_[39795]_ ;
  assign \new_[2310]_  = \new_[39784]_  & \new_[39771]_ ;
  assign \new_[2311]_  = \new_[39760]_  & \new_[39747]_ ;
  assign \new_[2312]_  = \new_[39736]_  & \new_[39723]_ ;
  assign \new_[2313]_  = \new_[39712]_  & \new_[39699]_ ;
  assign \new_[2314]_  = \new_[39688]_  & \new_[39675]_ ;
  assign \new_[2315]_  = \new_[39664]_  & \new_[39651]_ ;
  assign \new_[2316]_  = \new_[39640]_  & \new_[39627]_ ;
  assign \new_[2317]_  = \new_[39616]_  & \new_[39603]_ ;
  assign \new_[2318]_  = \new_[39592]_  & \new_[39579]_ ;
  assign \new_[2319]_  = \new_[39568]_  & \new_[39555]_ ;
  assign \new_[2320]_  = \new_[39544]_  & \new_[39531]_ ;
  assign \new_[2321]_  = \new_[39520]_  & \new_[39507]_ ;
  assign \new_[2322]_  = \new_[39496]_  & \new_[39483]_ ;
  assign \new_[2323]_  = \new_[39472]_  & \new_[39459]_ ;
  assign \new_[2324]_  = \new_[39448]_  & \new_[39435]_ ;
  assign \new_[2325]_  = \new_[39424]_  & \new_[39411]_ ;
  assign \new_[2326]_  = \new_[39400]_  & \new_[39387]_ ;
  assign \new_[2327]_  = \new_[39376]_  & \new_[39363]_ ;
  assign \new_[2328]_  = \new_[39352]_  & \new_[39339]_ ;
  assign \new_[2329]_  = \new_[39328]_  & \new_[39315]_ ;
  assign \new_[2330]_  = \new_[39304]_  & \new_[39291]_ ;
  assign \new_[2331]_  = \new_[39280]_  & \new_[39267]_ ;
  assign \new_[2332]_  = \new_[39256]_  & \new_[39243]_ ;
  assign \new_[2333]_  = \new_[39232]_  & \new_[39219]_ ;
  assign \new_[2334]_  = \new_[39208]_  & \new_[39195]_ ;
  assign \new_[2335]_  = \new_[39184]_  & \new_[39171]_ ;
  assign \new_[2336]_  = \new_[39160]_  & \new_[39147]_ ;
  assign \new_[2337]_  = \new_[39136]_  & \new_[39123]_ ;
  assign \new_[2338]_  = \new_[39112]_  & \new_[39099]_ ;
  assign \new_[2339]_  = \new_[39088]_  & \new_[39075]_ ;
  assign \new_[2340]_  = \new_[39064]_  & \new_[39051]_ ;
  assign \new_[2341]_  = \new_[39040]_  & \new_[39027]_ ;
  assign \new_[2342]_  = \new_[39016]_  & \new_[39003]_ ;
  assign \new_[2343]_  = \new_[38992]_  & \new_[38979]_ ;
  assign \new_[2344]_  = \new_[38968]_  & \new_[38955]_ ;
  assign \new_[2345]_  = \new_[38944]_  & \new_[38931]_ ;
  assign \new_[2346]_  = \new_[38920]_  & \new_[38907]_ ;
  assign \new_[2347]_  = \new_[38896]_  & \new_[38883]_ ;
  assign \new_[2348]_  = \new_[38872]_  & \new_[38859]_ ;
  assign \new_[2349]_  = \new_[38848]_  & \new_[38835]_ ;
  assign \new_[2350]_  = \new_[38824]_  & \new_[38811]_ ;
  assign \new_[2351]_  = \new_[38800]_  & \new_[38787]_ ;
  assign \new_[2352]_  = \new_[38776]_  & \new_[38763]_ ;
  assign \new_[2353]_  = \new_[38752]_  & \new_[38739]_ ;
  assign \new_[2354]_  = \new_[38728]_  & \new_[38715]_ ;
  assign \new_[2355]_  = \new_[38704]_  & \new_[38691]_ ;
  assign \new_[2356]_  = \new_[38680]_  & \new_[38667]_ ;
  assign \new_[2357]_  = \new_[38656]_  & \new_[38643]_ ;
  assign \new_[2358]_  = \new_[38632]_  & \new_[38619]_ ;
  assign \new_[2359]_  = \new_[38608]_  & \new_[38595]_ ;
  assign \new_[2360]_  = \new_[38584]_  & \new_[38571]_ ;
  assign \new_[2361]_  = \new_[38560]_  & \new_[38547]_ ;
  assign \new_[2362]_  = \new_[38536]_  & \new_[38523]_ ;
  assign \new_[2363]_  = \new_[38512]_  & \new_[38499]_ ;
  assign \new_[2364]_  = \new_[38488]_  & \new_[38475]_ ;
  assign \new_[2365]_  = \new_[38464]_  & \new_[38451]_ ;
  assign \new_[2366]_  = \new_[38440]_  & \new_[38427]_ ;
  assign \new_[2367]_  = \new_[38416]_  & \new_[38403]_ ;
  assign \new_[2368]_  = \new_[38392]_  & \new_[38379]_ ;
  assign \new_[2369]_  = \new_[38368]_  & \new_[38355]_ ;
  assign \new_[2370]_  = \new_[38344]_  & \new_[38331]_ ;
  assign \new_[2371]_  = \new_[38320]_  & \new_[38307]_ ;
  assign \new_[2372]_  = \new_[38296]_  & \new_[38283]_ ;
  assign \new_[2373]_  = \new_[38272]_  & \new_[38259]_ ;
  assign \new_[2374]_  = \new_[38248]_  & \new_[38235]_ ;
  assign \new_[2375]_  = \new_[38224]_  & \new_[38211]_ ;
  assign \new_[2376]_  = \new_[38200]_  & \new_[38187]_ ;
  assign \new_[2377]_  = \new_[38176]_  & \new_[38163]_ ;
  assign \new_[2378]_  = \new_[38152]_  & \new_[38139]_ ;
  assign \new_[2379]_  = \new_[38128]_  & \new_[38115]_ ;
  assign \new_[2380]_  = \new_[38104]_  & \new_[38091]_ ;
  assign \new_[2381]_  = \new_[38080]_  & \new_[38067]_ ;
  assign \new_[2382]_  = \new_[38056]_  & \new_[38043]_ ;
  assign \new_[2383]_  = \new_[38032]_  & \new_[38019]_ ;
  assign \new_[2384]_  = \new_[38008]_  & \new_[37995]_ ;
  assign \new_[2385]_  = \new_[37984]_  & \new_[37971]_ ;
  assign \new_[2386]_  = \new_[37960]_  & \new_[37947]_ ;
  assign \new_[2387]_  = \new_[37936]_  & \new_[37923]_ ;
  assign \new_[2388]_  = \new_[37912]_  & \new_[37899]_ ;
  assign \new_[2389]_  = \new_[37888]_  & \new_[37875]_ ;
  assign \new_[2390]_  = \new_[37864]_  & \new_[37851]_ ;
  assign \new_[2391]_  = \new_[37840]_  & \new_[37827]_ ;
  assign \new_[2392]_  = \new_[37816]_  & \new_[37803]_ ;
  assign \new_[2393]_  = \new_[37792]_  & \new_[37779]_ ;
  assign \new_[2394]_  = \new_[37768]_  & \new_[37755]_ ;
  assign \new_[2395]_  = \new_[37744]_  & \new_[37731]_ ;
  assign \new_[2396]_  = \new_[37720]_  & \new_[37707]_ ;
  assign \new_[2397]_  = \new_[37696]_  & \new_[37683]_ ;
  assign \new_[2398]_  = \new_[37672]_  & \new_[37659]_ ;
  assign \new_[2399]_  = \new_[37648]_  & \new_[37637]_ ;
  assign \new_[2400]_  = \new_[37626]_  & \new_[37615]_ ;
  assign \new_[2401]_  = \new_[37604]_  & \new_[37593]_ ;
  assign \new_[2402]_  = \new_[37582]_  & \new_[37571]_ ;
  assign \new_[2403]_  = \new_[37560]_  & \new_[37549]_ ;
  assign \new_[2404]_  = \new_[37538]_  & \new_[37527]_ ;
  assign \new_[2405]_  = \new_[37516]_  & \new_[37505]_ ;
  assign \new_[2406]_  = \new_[37494]_  & \new_[37483]_ ;
  assign \new_[2407]_  = \new_[37472]_  & \new_[37461]_ ;
  assign \new_[2408]_  = \new_[37450]_  & \new_[37439]_ ;
  assign \new_[2409]_  = \new_[37428]_  & \new_[37417]_ ;
  assign \new_[2410]_  = \new_[37406]_  & \new_[37395]_ ;
  assign \new_[2411]_  = \new_[37384]_  & \new_[37373]_ ;
  assign \new_[2412]_  = \new_[37362]_  & \new_[37351]_ ;
  assign \new_[2413]_  = \new_[37340]_  & \new_[37329]_ ;
  assign \new_[2414]_  = \new_[37318]_  & \new_[37307]_ ;
  assign \new_[2415]_  = \new_[37296]_  & \new_[37285]_ ;
  assign \new_[2416]_  = \new_[37274]_  & \new_[37263]_ ;
  assign \new_[2417]_  = \new_[37252]_  & \new_[37241]_ ;
  assign \new_[2418]_  = \new_[37230]_  & \new_[37219]_ ;
  assign \new_[2419]_  = \new_[37208]_  & \new_[37197]_ ;
  assign \new_[2420]_  = \new_[37186]_  & \new_[37175]_ ;
  assign \new_[2421]_  = \new_[37164]_  & \new_[37153]_ ;
  assign \new_[2422]_  = \new_[37142]_  & \new_[37131]_ ;
  assign \new_[2423]_  = \new_[37120]_  & \new_[37109]_ ;
  assign \new_[2424]_  = \new_[37098]_  & \new_[37087]_ ;
  assign \new_[2425]_  = \new_[37076]_  & \new_[37065]_ ;
  assign \new_[2426]_  = \new_[37054]_  & \new_[37043]_ ;
  assign \new_[2427]_  = \new_[37032]_  & \new_[37021]_ ;
  assign \new_[2428]_  = \new_[37010]_  & \new_[36999]_ ;
  assign \new_[2429]_  = \new_[36988]_  & \new_[36977]_ ;
  assign \new_[2430]_  = \new_[36966]_  & \new_[36955]_ ;
  assign \new_[2431]_  = \new_[36944]_  & \new_[36933]_ ;
  assign \new_[2432]_  = \new_[36922]_  & \new_[36911]_ ;
  assign \new_[2433]_  = \new_[36900]_  & \new_[36889]_ ;
  assign \new_[2434]_  = \new_[36878]_  & \new_[36867]_ ;
  assign \new_[2435]_  = \new_[36856]_  & \new_[36845]_ ;
  assign \new_[2436]_  = \new_[36834]_  & \new_[36823]_ ;
  assign \new_[2437]_  = \new_[36812]_  & \new_[36801]_ ;
  assign \new_[2438]_  = \new_[36790]_  & \new_[36779]_ ;
  assign \new_[2439]_  = \new_[36768]_  & \new_[36757]_ ;
  assign \new_[2440]_  = \new_[36746]_  & \new_[36735]_ ;
  assign \new_[2441]_  = \new_[36724]_  & \new_[36713]_ ;
  assign \new_[2442]_  = \new_[36702]_  & \new_[36691]_ ;
  assign \new_[2443]_  = \new_[36680]_  & \new_[36669]_ ;
  assign \new_[2444]_  = \new_[36658]_  & \new_[36647]_ ;
  assign \new_[2445]_  = \new_[36636]_  & \new_[36625]_ ;
  assign \new_[2446]_  = \new_[36614]_  & \new_[36603]_ ;
  assign \new_[2447]_  = \new_[36592]_  & \new_[36581]_ ;
  assign \new_[2448]_  = \new_[36570]_  & \new_[36559]_ ;
  assign \new_[2449]_  = \new_[36548]_  & \new_[36537]_ ;
  assign \new_[2450]_  = \new_[36526]_  & \new_[36515]_ ;
  assign \new_[2451]_  = \new_[36504]_  & \new_[36493]_ ;
  assign \new_[2452]_  = \new_[36482]_  & \new_[36471]_ ;
  assign \new_[2453]_  = \new_[36460]_  & \new_[36449]_ ;
  assign \new_[2454]_  = \new_[36438]_  & \new_[36427]_ ;
  assign \new_[2455]_  = \new_[36416]_  & \new_[36405]_ ;
  assign \new_[2456]_  = \new_[36394]_  & \new_[36383]_ ;
  assign \new_[2457]_  = \new_[36372]_  & \new_[36361]_ ;
  assign \new_[2458]_  = \new_[36350]_  & \new_[36339]_ ;
  assign \new_[2459]_  = \new_[36328]_  & \new_[36317]_ ;
  assign \new_[2460]_  = \new_[36306]_  & \new_[36295]_ ;
  assign \new_[2461]_  = \new_[36284]_  & \new_[36273]_ ;
  assign \new_[2462]_  = \new_[36262]_  & \new_[36251]_ ;
  assign \new_[2463]_  = \new_[36240]_  & \new_[36229]_ ;
  assign \new_[2464]_  = \new_[36218]_  & \new_[36207]_ ;
  assign \new_[2465]_  = \new_[36196]_  & \new_[36185]_ ;
  assign \new_[2466]_  = \new_[36174]_  & \new_[36163]_ ;
  assign \new_[2467]_  = \new_[36152]_  & \new_[36141]_ ;
  assign \new_[2468]_  = \new_[36130]_  & \new_[36119]_ ;
  assign \new_[2469]_  = \new_[36108]_  & \new_[36097]_ ;
  assign \new_[2470]_  = \new_[36086]_  & \new_[36075]_ ;
  assign \new_[2471]_  = \new_[36064]_  & \new_[36053]_ ;
  assign \new_[2472]_  = \new_[36042]_  & \new_[36031]_ ;
  assign \new_[2473]_  = \new_[36020]_  & \new_[36009]_ ;
  assign \new_[2474]_  = \new_[35998]_  & \new_[35987]_ ;
  assign \new_[2475]_  = \new_[35976]_  & \new_[35965]_ ;
  assign \new_[2476]_  = \new_[35954]_  & \new_[35943]_ ;
  assign \new_[2477]_  = \new_[35932]_  & \new_[35921]_ ;
  assign \new_[2478]_  = \new_[35910]_  & \new_[35899]_ ;
  assign \new_[2479]_  = \new_[35888]_  & \new_[35877]_ ;
  assign \new_[2480]_  = \new_[35866]_  & \new_[35855]_ ;
  assign \new_[2481]_  = \new_[35844]_  & \new_[35833]_ ;
  assign \new_[2482]_  = \new_[35822]_  & \new_[35811]_ ;
  assign \new_[2483]_  = \new_[35800]_  & \new_[35789]_ ;
  assign \new_[2484]_  = \new_[35778]_  & \new_[35767]_ ;
  assign \new_[2485]_  = \new_[35756]_  & \new_[35745]_ ;
  assign \new_[2486]_  = \new_[35734]_  & \new_[35723]_ ;
  assign \new_[2487]_  = \new_[35712]_  & \new_[35701]_ ;
  assign \new_[2488]_  = \new_[35690]_  & \new_[35679]_ ;
  assign \new_[2489]_  = \new_[35668]_  & \new_[35657]_ ;
  assign \new_[2490]_  = \new_[35646]_  & \new_[35635]_ ;
  assign \new_[2491]_  = \new_[35624]_  & \new_[35613]_ ;
  assign \new_[2492]_  = \new_[35602]_  & \new_[35591]_ ;
  assign \new_[2493]_  = \new_[35580]_  & \new_[35569]_ ;
  assign \new_[2494]_  = \new_[35558]_  & \new_[35547]_ ;
  assign \new_[2495]_  = \new_[35536]_  & \new_[35525]_ ;
  assign \new_[2496]_  = \new_[35514]_  & \new_[35503]_ ;
  assign \new_[2497]_  = \new_[35492]_  & \new_[35481]_ ;
  assign \new_[2498]_  = \new_[35470]_  & \new_[35459]_ ;
  assign \new_[2499]_  = \new_[35448]_  & \new_[35437]_ ;
  assign \new_[2500]_  = \new_[35426]_  & \new_[35415]_ ;
  assign \new_[2501]_  = \new_[35404]_  & \new_[35393]_ ;
  assign \new_[2502]_  = \new_[35382]_  & \new_[35371]_ ;
  assign \new_[2503]_  = \new_[35360]_  & \new_[35349]_ ;
  assign \new_[2504]_  = \new_[35338]_  & \new_[35327]_ ;
  assign \new_[2505]_  = \new_[35316]_  & \new_[35305]_ ;
  assign \new_[2506]_  = \new_[35294]_  & \new_[35283]_ ;
  assign \new_[2507]_  = \new_[35272]_  & \new_[35261]_ ;
  assign \new_[2508]_  = \new_[35250]_  & \new_[35239]_ ;
  assign \new_[2509]_  = \new_[35228]_  & \new_[35217]_ ;
  assign \new_[2510]_  = \new_[35206]_  & \new_[35195]_ ;
  assign \new_[2511]_  = \new_[35184]_  & \new_[35173]_ ;
  assign \new_[2512]_  = \new_[35162]_  & \new_[35151]_ ;
  assign \new_[2513]_  = \new_[35140]_  & \new_[35129]_ ;
  assign \new_[2514]_  = \new_[35118]_  & \new_[35107]_ ;
  assign \new_[2515]_  = \new_[35096]_  & \new_[35085]_ ;
  assign \new_[2516]_  = \new_[35074]_  & \new_[35063]_ ;
  assign \new_[2517]_  = \new_[35052]_  & \new_[35041]_ ;
  assign \new_[2518]_  = \new_[35030]_  & \new_[35019]_ ;
  assign \new_[2519]_  = \new_[35008]_  & \new_[34997]_ ;
  assign \new_[2520]_  = \new_[34986]_  & \new_[34975]_ ;
  assign \new_[2521]_  = \new_[34964]_  & \new_[34953]_ ;
  assign \new_[2522]_  = \new_[34942]_  & \new_[34931]_ ;
  assign \new_[2523]_  = \new_[34920]_  & \new_[34909]_ ;
  assign \new_[2524]_  = \new_[34898]_  & \new_[34887]_ ;
  assign \new_[2525]_  = \new_[34876]_  & \new_[34865]_ ;
  assign \new_[2526]_  = \new_[34854]_  & \new_[34843]_ ;
  assign \new_[2527]_  = \new_[34832]_  & \new_[34821]_ ;
  assign \new_[2528]_  = \new_[34810]_  & \new_[34799]_ ;
  assign \new_[2529]_  = \new_[34788]_  & \new_[34777]_ ;
  assign \new_[2530]_  = \new_[34766]_  & \new_[34755]_ ;
  assign \new_[2531]_  = \new_[34744]_  & \new_[34733]_ ;
  assign \new_[2532]_  = \new_[34722]_  & \new_[34711]_ ;
  assign \new_[2533]_  = \new_[34700]_  & \new_[34689]_ ;
  assign \new_[2534]_  = \new_[34678]_  & \new_[34667]_ ;
  assign \new_[2535]_  = \new_[34656]_  & \new_[34645]_ ;
  assign \new_[2536]_  = \new_[34634]_  & \new_[34623]_ ;
  assign \new_[2537]_  = \new_[34612]_  & \new_[34601]_ ;
  assign \new_[2538]_  = \new_[34590]_  & \new_[34579]_ ;
  assign \new_[2539]_  = \new_[34568]_  & \new_[34557]_ ;
  assign \new_[2540]_  = \new_[34546]_  & \new_[34535]_ ;
  assign \new_[2541]_  = \new_[34524]_  & \new_[34513]_ ;
  assign \new_[2542]_  = \new_[34502]_  & \new_[34491]_ ;
  assign \new_[2543]_  = \new_[34480]_  & \new_[34469]_ ;
  assign \new_[2544]_  = \new_[34458]_  & \new_[34447]_ ;
  assign \new_[2545]_  = \new_[34436]_  & \new_[34425]_ ;
  assign \new_[2546]_  = \new_[34414]_  & \new_[34403]_ ;
  assign \new_[2547]_  = \new_[34392]_  & \new_[34381]_ ;
  assign \new_[2548]_  = \new_[34370]_  & \new_[34359]_ ;
  assign \new_[2549]_  = \new_[34348]_  & \new_[34337]_ ;
  assign \new_[2550]_  = \new_[34326]_  & \new_[34315]_ ;
  assign \new_[2551]_  = \new_[34304]_  & \new_[34293]_ ;
  assign \new_[2552]_  = \new_[34282]_  & \new_[34271]_ ;
  assign \new_[2553]_  = \new_[34260]_  & \new_[34249]_ ;
  assign \new_[2554]_  = \new_[34238]_  & \new_[34227]_ ;
  assign \new_[2555]_  = \new_[34216]_  & \new_[34205]_ ;
  assign \new_[2556]_  = \new_[34194]_  & \new_[34183]_ ;
  assign \new_[2557]_  = \new_[34172]_  & \new_[34161]_ ;
  assign \new_[2558]_  = \new_[34150]_  & \new_[34139]_ ;
  assign \new_[2559]_  = \new_[34128]_  & \new_[34117]_ ;
  assign \new_[2560]_  = \new_[34106]_  & \new_[34095]_ ;
  assign \new_[2561]_  = \new_[34084]_  & \new_[34073]_ ;
  assign \new_[2562]_  = \new_[34062]_  & \new_[34051]_ ;
  assign \new_[2563]_  = \new_[34040]_  & \new_[34029]_ ;
  assign \new_[2564]_  = \new_[34018]_  & \new_[34007]_ ;
  assign \new_[2565]_  = \new_[33996]_  & \new_[33985]_ ;
  assign \new_[2566]_  = \new_[33974]_  & \new_[33963]_ ;
  assign \new_[2567]_  = \new_[33952]_  & \new_[33941]_ ;
  assign \new_[2568]_  = \new_[33930]_  & \new_[33919]_ ;
  assign \new_[2569]_  = \new_[33908]_  & \new_[33897]_ ;
  assign \new_[2570]_  = \new_[33886]_  & \new_[33875]_ ;
  assign \new_[2571]_  = \new_[33864]_  & \new_[33853]_ ;
  assign \new_[2572]_  = \new_[33842]_  & \new_[33831]_ ;
  assign \new_[2573]_  = \new_[33820]_  & \new_[33809]_ ;
  assign \new_[2574]_  = \new_[33798]_  & \new_[33787]_ ;
  assign \new_[2575]_  = \new_[33776]_  & \new_[33765]_ ;
  assign \new_[2576]_  = \new_[33754]_  & \new_[33743]_ ;
  assign \new_[2577]_  = \new_[33732]_  & \new_[33721]_ ;
  assign \new_[2578]_  = \new_[33710]_  & \new_[33699]_ ;
  assign \new_[2579]_  = \new_[33688]_  & \new_[33677]_ ;
  assign \new_[2580]_  = \new_[33666]_  & \new_[33655]_ ;
  assign \new_[2581]_  = \new_[33644]_  & \new_[33633]_ ;
  assign \new_[2582]_  = \new_[33622]_  & \new_[33611]_ ;
  assign \new_[2583]_  = \new_[33600]_  & \new_[33589]_ ;
  assign \new_[2584]_  = \new_[33578]_  & \new_[33567]_ ;
  assign \new_[2585]_  = \new_[33556]_  & \new_[33545]_ ;
  assign \new_[2586]_  = \new_[33534]_  & \new_[33523]_ ;
  assign \new_[2587]_  = \new_[33512]_  & \new_[33501]_ ;
  assign \new_[2588]_  = \new_[33490]_  & \new_[33479]_ ;
  assign \new_[2589]_  = \new_[33468]_  & \new_[33457]_ ;
  assign \new_[2590]_  = \new_[33446]_  & \new_[33435]_ ;
  assign \new_[2591]_  = \new_[33424]_  & \new_[33413]_ ;
  assign \new_[2592]_  = \new_[33402]_  & \new_[33391]_ ;
  assign \new_[2593]_  = \new_[33380]_  & \new_[33369]_ ;
  assign \new_[2594]_  = \new_[33358]_  & \new_[33347]_ ;
  assign \new_[2595]_  = \new_[33336]_  & \new_[33325]_ ;
  assign \new_[2596]_  = \new_[33314]_  & \new_[33303]_ ;
  assign \new_[2597]_  = \new_[33292]_  & \new_[33281]_ ;
  assign \new_[2598]_  = \new_[33270]_  & \new_[33259]_ ;
  assign \new_[2599]_  = \new_[33248]_  & \new_[33237]_ ;
  assign \new_[2600]_  = \new_[33226]_  & \new_[33215]_ ;
  assign \new_[2601]_  = \new_[33204]_  & \new_[33193]_ ;
  assign \new_[2602]_  = \new_[33182]_  & \new_[33171]_ ;
  assign \new_[2603]_  = \new_[33160]_  & \new_[33149]_ ;
  assign \new_[2604]_  = \new_[33138]_  & \new_[33127]_ ;
  assign \new_[2605]_  = \new_[33116]_  & \new_[33105]_ ;
  assign \new_[2606]_  = \new_[33094]_  & \new_[33083]_ ;
  assign \new_[2607]_  = \new_[33072]_  & \new_[33061]_ ;
  assign \new_[2608]_  = \new_[33050]_  & \new_[33039]_ ;
  assign \new_[2609]_  = \new_[33028]_  & \new_[33017]_ ;
  assign \new_[2610]_  = \new_[33006]_  & \new_[32995]_ ;
  assign \new_[2611]_  = \new_[32984]_  & \new_[32973]_ ;
  assign \new_[2612]_  = \new_[32962]_  & \new_[32951]_ ;
  assign \new_[2613]_  = \new_[32940]_  & \new_[32929]_ ;
  assign \new_[2614]_  = \new_[32918]_  & \new_[32907]_ ;
  assign \new_[2615]_  = \new_[32896]_  & \new_[32885]_ ;
  assign \new_[2616]_  = \new_[32874]_  & \new_[32863]_ ;
  assign \new_[2617]_  = \new_[32852]_  & \new_[32841]_ ;
  assign \new_[2618]_  = \new_[32830]_  & \new_[32819]_ ;
  assign \new_[2619]_  = \new_[32808]_  & \new_[32797]_ ;
  assign \new_[2620]_  = \new_[32786]_  & \new_[32775]_ ;
  assign \new_[2621]_  = \new_[32764]_  & \new_[32753]_ ;
  assign \new_[2622]_  = \new_[32742]_  & \new_[32731]_ ;
  assign \new_[2623]_  = \new_[32720]_  & \new_[32709]_ ;
  assign \new_[2624]_  = \new_[32698]_  & \new_[32687]_ ;
  assign \new_[2625]_  = \new_[32676]_  & \new_[32665]_ ;
  assign \new_[2626]_  = \new_[32654]_  & \new_[32643]_ ;
  assign \new_[2627]_  = \new_[32632]_  & \new_[32621]_ ;
  assign \new_[2628]_  = \new_[32610]_  & \new_[32599]_ ;
  assign \new_[2629]_  = \new_[32588]_  & \new_[32577]_ ;
  assign \new_[2630]_  = \new_[32566]_  & \new_[32555]_ ;
  assign \new_[2631]_  = \new_[32544]_  & \new_[32533]_ ;
  assign \new_[2632]_  = \new_[32522]_  & \new_[32511]_ ;
  assign \new_[2633]_  = \new_[32500]_  & \new_[32489]_ ;
  assign \new_[2634]_  = \new_[32478]_  & \new_[32467]_ ;
  assign \new_[2635]_  = \new_[32456]_  & \new_[32445]_ ;
  assign \new_[2636]_  = \new_[32434]_  & \new_[32423]_ ;
  assign \new_[2637]_  = \new_[32412]_  & \new_[32401]_ ;
  assign \new_[2638]_  = \new_[32390]_  & \new_[32379]_ ;
  assign \new_[2639]_  = \new_[32368]_  & \new_[32357]_ ;
  assign \new_[2640]_  = \new_[32346]_  & \new_[32335]_ ;
  assign \new_[2641]_  = \new_[32324]_  & \new_[32313]_ ;
  assign \new_[2642]_  = \new_[32302]_  & \new_[32291]_ ;
  assign \new_[2643]_  = \new_[32280]_  & \new_[32269]_ ;
  assign \new_[2644]_  = \new_[32258]_  & \new_[32247]_ ;
  assign \new_[2645]_  = \new_[32236]_  & \new_[32225]_ ;
  assign \new_[2646]_  = \new_[32214]_  & \new_[32203]_ ;
  assign \new_[2647]_  = \new_[32192]_  & \new_[32181]_ ;
  assign \new_[2648]_  = \new_[32170]_  & \new_[32159]_ ;
  assign \new_[2649]_  = \new_[32148]_  & \new_[32137]_ ;
  assign \new_[2650]_  = \new_[32126]_  & \new_[32115]_ ;
  assign \new_[2651]_  = \new_[32104]_  & \new_[32093]_ ;
  assign \new_[2652]_  = \new_[32082]_  & \new_[32071]_ ;
  assign \new_[2653]_  = \new_[32060]_  & \new_[32049]_ ;
  assign \new_[2654]_  = \new_[32038]_  & \new_[32027]_ ;
  assign \new_[2655]_  = \new_[32016]_  & \new_[32005]_ ;
  assign \new_[2656]_  = \new_[31994]_  & \new_[31983]_ ;
  assign \new_[2657]_  = \new_[31972]_  & \new_[31961]_ ;
  assign \new_[2658]_  = \new_[31950]_  & \new_[31939]_ ;
  assign \new_[2659]_  = \new_[31928]_  & \new_[31917]_ ;
  assign \new_[2660]_  = \new_[31906]_  & \new_[31895]_ ;
  assign \new_[2661]_  = \new_[31884]_  & \new_[31873]_ ;
  assign \new_[2662]_  = \new_[31862]_  & \new_[31851]_ ;
  assign \new_[2663]_  = \new_[31840]_  & \new_[31829]_ ;
  assign \new_[2664]_  = \new_[31818]_  & \new_[31807]_ ;
  assign \new_[2665]_  = \new_[31796]_  & \new_[31785]_ ;
  assign \new_[2666]_  = \new_[31774]_  & \new_[31763]_ ;
  assign \new_[2667]_  = \new_[31752]_  & \new_[31741]_ ;
  assign \new_[2668]_  = \new_[31730]_  & \new_[31719]_ ;
  assign \new_[2669]_  = \new_[31708]_  & \new_[31697]_ ;
  assign \new_[2670]_  = \new_[31686]_  & \new_[31675]_ ;
  assign \new_[2671]_  = \new_[31664]_  & \new_[31653]_ ;
  assign \new_[2672]_  = \new_[31642]_  & \new_[31631]_ ;
  assign \new_[2673]_  = \new_[31620]_  & \new_[31609]_ ;
  assign \new_[2674]_  = \new_[31598]_  & \new_[31587]_ ;
  assign \new_[2675]_  = \new_[31576]_  & \new_[31565]_ ;
  assign \new_[2676]_  = \new_[31554]_  & \new_[31543]_ ;
  assign \new_[2677]_  = \new_[31532]_  & \new_[31521]_ ;
  assign \new_[2678]_  = \new_[31510]_  & \new_[31499]_ ;
  assign \new_[2679]_  = \new_[31488]_  & \new_[31477]_ ;
  assign \new_[2680]_  = \new_[31466]_  & \new_[31455]_ ;
  assign \new_[2681]_  = \new_[31444]_  & \new_[31433]_ ;
  assign \new_[2682]_  = \new_[31422]_  & \new_[31411]_ ;
  assign \new_[2683]_  = \new_[31400]_  & \new_[31389]_ ;
  assign \new_[2684]_  = \new_[31378]_  & \new_[31367]_ ;
  assign \new_[2685]_  = \new_[31356]_  & \new_[31345]_ ;
  assign \new_[2686]_  = \new_[31334]_  & \new_[31323]_ ;
  assign \new_[2687]_  = \new_[31312]_  & \new_[31301]_ ;
  assign \new_[2688]_  = \new_[31290]_  & \new_[31279]_ ;
  assign \new_[2689]_  = \new_[31268]_  & \new_[31257]_ ;
  assign \new_[2690]_  = \new_[31246]_  & \new_[31235]_ ;
  assign \new_[2691]_  = \new_[31224]_  & \new_[31213]_ ;
  assign \new_[2692]_  = \new_[31202]_  & \new_[31191]_ ;
  assign \new_[2693]_  = \new_[31180]_  & \new_[31169]_ ;
  assign \new_[2694]_  = \new_[31158]_  & \new_[31147]_ ;
  assign \new_[2695]_  = \new_[31136]_  & \new_[31125]_ ;
  assign \new_[2696]_  = \new_[31114]_  & \new_[31103]_ ;
  assign \new_[2697]_  = \new_[31092]_  & \new_[31081]_ ;
  assign \new_[2698]_  = \new_[31070]_  & \new_[31059]_ ;
  assign \new_[2699]_  = \new_[31048]_  & \new_[31037]_ ;
  assign \new_[2700]_  = \new_[31026]_  & \new_[31015]_ ;
  assign \new_[2701]_  = \new_[31004]_  & \new_[30993]_ ;
  assign \new_[2702]_  = \new_[30982]_  & \new_[30971]_ ;
  assign \new_[2703]_  = \new_[30960]_  & \new_[30949]_ ;
  assign \new_[2704]_  = \new_[30938]_  & \new_[30927]_ ;
  assign \new_[2705]_  = \new_[30916]_  & \new_[30905]_ ;
  assign \new_[2706]_  = \new_[30894]_  & \new_[30883]_ ;
  assign \new_[2707]_  = \new_[30872]_  & \new_[30861]_ ;
  assign \new_[2708]_  = \new_[30850]_  & \new_[30839]_ ;
  assign \new_[2709]_  = \new_[30828]_  & \new_[30817]_ ;
  assign \new_[2710]_  = \new_[30806]_  & \new_[30795]_ ;
  assign \new_[2711]_  = \new_[30784]_  & \new_[30773]_ ;
  assign \new_[2712]_  = \new_[30762]_  & \new_[30751]_ ;
  assign \new_[2713]_  = \new_[30740]_  & \new_[30729]_ ;
  assign \new_[2714]_  = \new_[30718]_  & \new_[30707]_ ;
  assign \new_[2715]_  = \new_[30696]_  & \new_[30685]_ ;
  assign \new_[2716]_  = \new_[30674]_  & \new_[30663]_ ;
  assign \new_[2717]_  = \new_[30652]_  & \new_[30641]_ ;
  assign \new_[2718]_  = \new_[30630]_  & \new_[30619]_ ;
  assign \new_[2719]_  = \new_[30608]_  & \new_[30597]_ ;
  assign \new_[2720]_  = \new_[30586]_  & \new_[30575]_ ;
  assign \new_[2721]_  = \new_[30564]_  & \new_[30553]_ ;
  assign \new_[2722]_  = \new_[30542]_  & \new_[30531]_ ;
  assign \new_[2723]_  = \new_[30520]_  & \new_[30509]_ ;
  assign \new_[2724]_  = \new_[30498]_  & \new_[30487]_ ;
  assign \new_[2725]_  = \new_[30476]_  & \new_[30465]_ ;
  assign \new_[2726]_  = \new_[30454]_  & \new_[30443]_ ;
  assign \new_[2727]_  = \new_[30432]_  & \new_[30421]_ ;
  assign \new_[2728]_  = \new_[30410]_  & \new_[30399]_ ;
  assign \new_[2729]_  = \new_[30388]_  & \new_[30377]_ ;
  assign \new_[2730]_  = \new_[30366]_  & \new_[30355]_ ;
  assign \new_[2731]_  = \new_[30344]_  & \new_[30333]_ ;
  assign \new_[2732]_  = \new_[30322]_  & \new_[30311]_ ;
  assign \new_[2733]_  = \new_[30300]_  & \new_[30289]_ ;
  assign \new_[2734]_  = \new_[30278]_  & \new_[30267]_ ;
  assign \new_[2735]_  = \new_[30256]_  & \new_[30245]_ ;
  assign \new_[2736]_  = \new_[30234]_  & \new_[30223]_ ;
  assign \new_[2737]_  = \new_[30212]_  & \new_[30201]_ ;
  assign \new_[2738]_  = \new_[30190]_  & \new_[30179]_ ;
  assign \new_[2739]_  = \new_[30168]_  & \new_[30157]_ ;
  assign \new_[2740]_  = \new_[30146]_  & \new_[30135]_ ;
  assign \new_[2741]_  = \new_[30124]_  & \new_[30113]_ ;
  assign \new_[2742]_  = \new_[30102]_  & \new_[30091]_ ;
  assign \new_[2743]_  = \new_[30080]_  & \new_[30069]_ ;
  assign \new_[2744]_  = \new_[30058]_  & \new_[30047]_ ;
  assign \new_[2745]_  = \new_[30036]_  & \new_[30025]_ ;
  assign \new_[2746]_  = \new_[30014]_  & \new_[30003]_ ;
  assign \new_[2747]_  = \new_[29992]_  & \new_[29981]_ ;
  assign \new_[2748]_  = \new_[29970]_  & \new_[29959]_ ;
  assign \new_[2749]_  = \new_[29948]_  & \new_[29937]_ ;
  assign \new_[2750]_  = \new_[29926]_  & \new_[29915]_ ;
  assign \new_[2751]_  = \new_[29904]_  & \new_[29893]_ ;
  assign \new_[2752]_  = \new_[29882]_  & \new_[29871]_ ;
  assign \new_[2753]_  = \new_[29860]_  & \new_[29849]_ ;
  assign \new_[2754]_  = \new_[29838]_  & \new_[29827]_ ;
  assign \new_[2755]_  = \new_[29816]_  & \new_[29805]_ ;
  assign \new_[2756]_  = \new_[29794]_  & \new_[29783]_ ;
  assign \new_[2757]_  = \new_[29772]_  & \new_[29761]_ ;
  assign \new_[2758]_  = \new_[29750]_  & \new_[29739]_ ;
  assign \new_[2759]_  = \new_[29728]_  & \new_[29717]_ ;
  assign \new_[2760]_  = \new_[29706]_  & \new_[29695]_ ;
  assign \new_[2761]_  = \new_[29684]_  & \new_[29673]_ ;
  assign \new_[2762]_  = \new_[29662]_  & \new_[29651]_ ;
  assign \new_[2763]_  = \new_[29640]_  & \new_[29629]_ ;
  assign \new_[2764]_  = \new_[29618]_  & \new_[29607]_ ;
  assign \new_[2765]_  = \new_[29596]_  & \new_[29585]_ ;
  assign \new_[2766]_  = \new_[29574]_  & \new_[29563]_ ;
  assign \new_[2767]_  = \new_[29552]_  & \new_[29541]_ ;
  assign \new_[2768]_  = \new_[29530]_  & \new_[29519]_ ;
  assign \new_[2769]_  = \new_[29508]_  & \new_[29497]_ ;
  assign \new_[2770]_  = \new_[29486]_  & \new_[29475]_ ;
  assign \new_[2771]_  = \new_[29464]_  & \new_[29453]_ ;
  assign \new_[2772]_  = \new_[29442]_  & \new_[29431]_ ;
  assign \new_[2773]_  = \new_[29420]_  & \new_[29409]_ ;
  assign \new_[2774]_  = \new_[29398]_  & \new_[29387]_ ;
  assign \new_[2775]_  = \new_[29376]_  & \new_[29365]_ ;
  assign \new_[2776]_  = \new_[29354]_  & \new_[29343]_ ;
  assign \new_[2777]_  = \new_[29332]_  & \new_[29321]_ ;
  assign \new_[2778]_  = \new_[29310]_  & \new_[29299]_ ;
  assign \new_[2779]_  = \new_[29288]_  & \new_[29277]_ ;
  assign \new_[2780]_  = \new_[29266]_  & \new_[29255]_ ;
  assign \new_[2781]_  = \new_[29244]_  & \new_[29233]_ ;
  assign \new_[2782]_  = \new_[29222]_  & \new_[29211]_ ;
  assign \new_[2783]_  = \new_[29200]_  & \new_[29189]_ ;
  assign \new_[2784]_  = \new_[29178]_  & \new_[29167]_ ;
  assign \new_[2785]_  = \new_[29156]_  & \new_[29145]_ ;
  assign \new_[2786]_  = \new_[29134]_  & \new_[29123]_ ;
  assign \new_[2787]_  = \new_[29112]_  & \new_[29101]_ ;
  assign \new_[2788]_  = \new_[29090]_  & \new_[29079]_ ;
  assign \new_[2789]_  = \new_[29068]_  & \new_[29057]_ ;
  assign \new_[2790]_  = \new_[29046]_  & \new_[29035]_ ;
  assign \new_[2791]_  = \new_[29024]_  & \new_[29013]_ ;
  assign \new_[2792]_  = \new_[29002]_  & \new_[28991]_ ;
  assign \new_[2793]_  = \new_[28980]_  & \new_[28969]_ ;
  assign \new_[2794]_  = \new_[28958]_  & \new_[28947]_ ;
  assign \new_[2795]_  = \new_[28936]_  & \new_[28925]_ ;
  assign \new_[2796]_  = \new_[28914]_  & \new_[28903]_ ;
  assign \new_[2797]_  = \new_[28892]_  & \new_[28881]_ ;
  assign \new_[2798]_  = \new_[28870]_  & \new_[28859]_ ;
  assign \new_[2799]_  = \new_[28848]_  & \new_[28837]_ ;
  assign \new_[2800]_  = \new_[28826]_  & \new_[28815]_ ;
  assign \new_[2801]_  = \new_[28804]_  & \new_[28793]_ ;
  assign \new_[2802]_  = \new_[28782]_  & \new_[28771]_ ;
  assign \new_[2803]_  = \new_[28760]_  & \new_[28749]_ ;
  assign \new_[2804]_  = \new_[28738]_  & \new_[28727]_ ;
  assign \new_[2805]_  = \new_[28716]_  & \new_[28705]_ ;
  assign \new_[2806]_  = \new_[28694]_  & \new_[28683]_ ;
  assign \new_[2807]_  = \new_[28672]_  & \new_[28661]_ ;
  assign \new_[2808]_  = \new_[28650]_  & \new_[28639]_ ;
  assign \new_[2809]_  = \new_[28628]_  & \new_[28617]_ ;
  assign \new_[2810]_  = \new_[28606]_  & \new_[28595]_ ;
  assign \new_[2811]_  = \new_[28584]_  & \new_[28573]_ ;
  assign \new_[2812]_  = \new_[28562]_  & \new_[28551]_ ;
  assign \new_[2813]_  = \new_[28540]_  & \new_[28529]_ ;
  assign \new_[2814]_  = \new_[28518]_  & \new_[28507]_ ;
  assign \new_[2815]_  = \new_[28496]_  & \new_[28485]_ ;
  assign \new_[2816]_  = \new_[28474]_  & \new_[28463]_ ;
  assign \new_[2817]_  = \new_[28452]_  & \new_[28441]_ ;
  assign \new_[2818]_  = \new_[28430]_  & \new_[28419]_ ;
  assign \new_[2819]_  = \new_[28408]_  & \new_[28397]_ ;
  assign \new_[2820]_  = \new_[28386]_  & \new_[28375]_ ;
  assign \new_[2821]_  = \new_[28364]_  & \new_[28353]_ ;
  assign \new_[2822]_  = \new_[28342]_  & \new_[28331]_ ;
  assign \new_[2823]_  = \new_[28320]_  & \new_[28309]_ ;
  assign \new_[2824]_  = \new_[28298]_  & \new_[28287]_ ;
  assign \new_[2825]_  = \new_[28276]_  & \new_[28265]_ ;
  assign \new_[2826]_  = \new_[28254]_  & \new_[28243]_ ;
  assign \new_[2827]_  = \new_[28232]_  & \new_[28221]_ ;
  assign \new_[2828]_  = \new_[28210]_  & \new_[28199]_ ;
  assign \new_[2829]_  = \new_[28188]_  & \new_[28177]_ ;
  assign \new_[2830]_  = \new_[28166]_  & \new_[28155]_ ;
  assign \new_[2831]_  = \new_[28144]_  & \new_[28133]_ ;
  assign \new_[2832]_  = \new_[28122]_  & \new_[28111]_ ;
  assign \new_[2833]_  = \new_[28100]_  & \new_[28089]_ ;
  assign \new_[2834]_  = \new_[28078]_  & \new_[28067]_ ;
  assign \new_[2835]_  = \new_[28056]_  & \new_[28045]_ ;
  assign \new_[2836]_  = \new_[28034]_  & \new_[28023]_ ;
  assign \new_[2837]_  = \new_[28012]_  & \new_[28001]_ ;
  assign \new_[2838]_  = \new_[27990]_  & \new_[27979]_ ;
  assign \new_[2839]_  = \new_[27968]_  & \new_[27957]_ ;
  assign \new_[2840]_  = \new_[27946]_  & \new_[27935]_ ;
  assign \new_[2841]_  = \new_[27924]_  & \new_[27913]_ ;
  assign \new_[2842]_  = \new_[27902]_  & \new_[27891]_ ;
  assign \new_[2843]_  = \new_[27880]_  & \new_[27869]_ ;
  assign \new_[2844]_  = \new_[27858]_  & \new_[27847]_ ;
  assign \new_[2845]_  = \new_[27836]_  & \new_[27825]_ ;
  assign \new_[2846]_  = \new_[27814]_  & \new_[27803]_ ;
  assign \new_[2847]_  = \new_[27792]_  & \new_[27781]_ ;
  assign \new_[2848]_  = \new_[27770]_  & \new_[27759]_ ;
  assign \new_[2849]_  = \new_[27748]_  & \new_[27737]_ ;
  assign \new_[2850]_  = \new_[27726]_  & \new_[27715]_ ;
  assign \new_[2851]_  = \new_[27704]_  & \new_[27693]_ ;
  assign \new_[2852]_  = \new_[27682]_  & \new_[27671]_ ;
  assign \new_[2853]_  = \new_[27660]_  & \new_[27649]_ ;
  assign \new_[2854]_  = \new_[27638]_  & \new_[27627]_ ;
  assign \new_[2855]_  = \new_[27616]_  & \new_[27605]_ ;
  assign \new_[2856]_  = \new_[27594]_  & \new_[27583]_ ;
  assign \new_[2857]_  = \new_[27572]_  & \new_[27561]_ ;
  assign \new_[2858]_  = \new_[27550]_  & \new_[27539]_ ;
  assign \new_[2859]_  = \new_[27528]_  & \new_[27517]_ ;
  assign \new_[2860]_  = \new_[27506]_  & \new_[27495]_ ;
  assign \new_[2861]_  = \new_[27484]_  & \new_[27473]_ ;
  assign \new_[2862]_  = \new_[27462]_  & \new_[27451]_ ;
  assign \new_[2863]_  = \new_[27440]_  & \new_[27429]_ ;
  assign \new_[2864]_  = \new_[27418]_  & \new_[27407]_ ;
  assign \new_[2865]_  = \new_[27396]_  & \new_[27385]_ ;
  assign \new_[2866]_  = \new_[27374]_  & \new_[27363]_ ;
  assign \new_[2867]_  = \new_[27352]_  & \new_[27341]_ ;
  assign \new_[2868]_  = \new_[27330]_  & \new_[27319]_ ;
  assign \new_[2869]_  = \new_[27308]_  & \new_[27297]_ ;
  assign \new_[2870]_  = \new_[27286]_  & \new_[27275]_ ;
  assign \new_[2871]_  = \new_[27264]_  & \new_[27253]_ ;
  assign \new_[2872]_  = \new_[27242]_  & \new_[27231]_ ;
  assign \new_[2873]_  = \new_[27220]_  & \new_[27209]_ ;
  assign \new_[2874]_  = \new_[27198]_  & \new_[27187]_ ;
  assign \new_[2875]_  = \new_[27176]_  & \new_[27165]_ ;
  assign \new_[2876]_  = \new_[27154]_  & \new_[27143]_ ;
  assign \new_[2877]_  = \new_[27132]_  & \new_[27121]_ ;
  assign \new_[2878]_  = \new_[27110]_  & \new_[27099]_ ;
  assign \new_[2879]_  = \new_[27088]_  & \new_[27077]_ ;
  assign \new_[2880]_  = \new_[27066]_  & \new_[27055]_ ;
  assign \new_[2881]_  = \new_[27044]_  & \new_[27033]_ ;
  assign \new_[2882]_  = \new_[27022]_  & \new_[27011]_ ;
  assign \new_[2883]_  = \new_[27000]_  & \new_[26989]_ ;
  assign \new_[2884]_  = \new_[26978]_  & \new_[26967]_ ;
  assign \new_[2885]_  = \new_[26956]_  & \new_[26945]_ ;
  assign \new_[2886]_  = \new_[26934]_  & \new_[26923]_ ;
  assign \new_[2887]_  = \new_[26912]_  & \new_[26901]_ ;
  assign \new_[2888]_  = \new_[26890]_  & \new_[26879]_ ;
  assign \new_[2889]_  = \new_[26868]_  & \new_[26857]_ ;
  assign \new_[2890]_  = \new_[26846]_  & \new_[26835]_ ;
  assign \new_[2891]_  = \new_[26824]_  & \new_[26813]_ ;
  assign \new_[2892]_  = \new_[26802]_  & \new_[26791]_ ;
  assign \new_[2893]_  = \new_[26780]_  & \new_[26769]_ ;
  assign \new_[2894]_  = \new_[26758]_  & \new_[26747]_ ;
  assign \new_[2895]_  = \new_[26736]_  & \new_[26725]_ ;
  assign \new_[2896]_  = \new_[26714]_  & \new_[26703]_ ;
  assign \new_[2897]_  = \new_[26692]_  & \new_[26681]_ ;
  assign \new_[2898]_  = \new_[26670]_  & \new_[26659]_ ;
  assign \new_[2899]_  = \new_[26648]_  & \new_[26637]_ ;
  assign \new_[2900]_  = \new_[26626]_  & \new_[26615]_ ;
  assign \new_[2901]_  = \new_[26604]_  & \new_[26593]_ ;
  assign \new_[2902]_  = \new_[26582]_  & \new_[26571]_ ;
  assign \new_[2903]_  = \new_[26560]_  & \new_[26549]_ ;
  assign \new_[2904]_  = \new_[26538]_  & \new_[26527]_ ;
  assign \new_[2905]_  = \new_[26516]_  & \new_[26505]_ ;
  assign \new_[2906]_  = \new_[26494]_  & \new_[26483]_ ;
  assign \new_[2907]_  = \new_[26472]_  & \new_[26461]_ ;
  assign \new_[2908]_  = \new_[26450]_  & \new_[26439]_ ;
  assign \new_[2909]_  = \new_[26428]_  & \new_[26417]_ ;
  assign \new_[2910]_  = \new_[26406]_  & \new_[26395]_ ;
  assign \new_[2911]_  = \new_[26384]_  & \new_[26373]_ ;
  assign \new_[2912]_  = \new_[26362]_  & \new_[26351]_ ;
  assign \new_[2913]_  = \new_[26340]_  & \new_[26329]_ ;
  assign \new_[2914]_  = \new_[26318]_  & \new_[26307]_ ;
  assign \new_[2915]_  = \new_[26296]_  & \new_[26285]_ ;
  assign \new_[2916]_  = \new_[26274]_  & \new_[26263]_ ;
  assign \new_[2917]_  = \new_[26252]_  & \new_[26241]_ ;
  assign \new_[2918]_  = \new_[26230]_  & \new_[26219]_ ;
  assign \new_[2919]_  = \new_[26208]_  & \new_[26197]_ ;
  assign \new_[2920]_  = \new_[26186]_  & \new_[26175]_ ;
  assign \new_[2921]_  = \new_[26164]_  & \new_[26153]_ ;
  assign \new_[2922]_  = \new_[26142]_  & \new_[26131]_ ;
  assign \new_[2923]_  = \new_[26120]_  & \new_[26109]_ ;
  assign \new_[2924]_  = \new_[26098]_  & \new_[26087]_ ;
  assign \new_[2925]_  = \new_[26076]_  & \new_[26065]_ ;
  assign \new_[2926]_  = \new_[26054]_  & \new_[26043]_ ;
  assign \new_[2927]_  = \new_[26032]_  & \new_[26021]_ ;
  assign \new_[2928]_  = \new_[26010]_  & \new_[25999]_ ;
  assign \new_[2929]_  = \new_[25988]_  & \new_[25977]_ ;
  assign \new_[2930]_  = \new_[25966]_  & \new_[25955]_ ;
  assign \new_[2931]_  = \new_[25944]_  & \new_[25933]_ ;
  assign \new_[2932]_  = \new_[25922]_  & \new_[25911]_ ;
  assign \new_[2933]_  = \new_[25900]_  & \new_[25889]_ ;
  assign \new_[2934]_  = \new_[25878]_  & \new_[25867]_ ;
  assign \new_[2935]_  = \new_[25856]_  & \new_[25845]_ ;
  assign \new_[2936]_  = \new_[25834]_  & \new_[25823]_ ;
  assign \new_[2937]_  = \new_[25812]_  & \new_[25801]_ ;
  assign \new_[2938]_  = \new_[25790]_  & \new_[25779]_ ;
  assign \new_[2939]_  = \new_[25768]_  & \new_[25757]_ ;
  assign \new_[2940]_  = \new_[25746]_  & \new_[25735]_ ;
  assign \new_[2941]_  = \new_[25724]_  & \new_[25713]_ ;
  assign \new_[2942]_  = \new_[25702]_  & \new_[25691]_ ;
  assign \new_[2943]_  = \new_[25680]_  & \new_[25669]_ ;
  assign \new_[2944]_  = \new_[25658]_  & \new_[25647]_ ;
  assign \new_[2945]_  = \new_[25636]_  & \new_[25625]_ ;
  assign \new_[2946]_  = \new_[25614]_  & \new_[25603]_ ;
  assign \new_[2947]_  = \new_[25592]_  & \new_[25581]_ ;
  assign \new_[2948]_  = \new_[25570]_  & \new_[25559]_ ;
  assign \new_[2949]_  = \new_[25548]_  & \new_[25537]_ ;
  assign \new_[2950]_  = \new_[25526]_  & \new_[25515]_ ;
  assign \new_[2951]_  = \new_[25504]_  & \new_[25493]_ ;
  assign \new_[2952]_  = \new_[25482]_  & \new_[25471]_ ;
  assign \new_[2953]_  = \new_[25460]_  & \new_[25449]_ ;
  assign \new_[2954]_  = \new_[25438]_  & \new_[25427]_ ;
  assign \new_[2955]_  = \new_[25416]_  & \new_[25405]_ ;
  assign \new_[2956]_  = \new_[25394]_  & \new_[25383]_ ;
  assign \new_[2957]_  = \new_[25372]_  & \new_[25361]_ ;
  assign \new_[2958]_  = \new_[25350]_  & \new_[25339]_ ;
  assign \new_[2959]_  = \new_[25328]_  & \new_[25317]_ ;
  assign \new_[2960]_  = \new_[25306]_  & \new_[25295]_ ;
  assign \new_[2961]_  = \new_[25284]_  & \new_[25273]_ ;
  assign \new_[2962]_  = \new_[25262]_  & \new_[25251]_ ;
  assign \new_[2963]_  = \new_[25240]_  & \new_[25229]_ ;
  assign \new_[2964]_  = \new_[25218]_  & \new_[25207]_ ;
  assign \new_[2965]_  = \new_[25196]_  & \new_[25185]_ ;
  assign \new_[2966]_  = \new_[25174]_  & \new_[25163]_ ;
  assign \new_[2967]_  = \new_[25152]_  & \new_[25141]_ ;
  assign \new_[2968]_  = \new_[25130]_  & \new_[25119]_ ;
  assign \new_[2969]_  = \new_[25108]_  & \new_[25097]_ ;
  assign \new_[2970]_  = \new_[25086]_  & \new_[25075]_ ;
  assign \new_[2971]_  = \new_[25064]_  & \new_[25053]_ ;
  assign \new_[2972]_  = \new_[25042]_  & \new_[25031]_ ;
  assign \new_[2973]_  = \new_[25020]_  & \new_[25009]_ ;
  assign \new_[2974]_  = \new_[24998]_  & \new_[24987]_ ;
  assign \new_[2975]_  = \new_[24976]_  & \new_[24965]_ ;
  assign \new_[2976]_  = \new_[24954]_  & \new_[24943]_ ;
  assign \new_[2977]_  = \new_[24932]_  & \new_[24921]_ ;
  assign \new_[2978]_  = \new_[24910]_  & \new_[24899]_ ;
  assign \new_[2979]_  = \new_[24888]_  & \new_[24877]_ ;
  assign \new_[2980]_  = \new_[24866]_  & \new_[24855]_ ;
  assign \new_[2981]_  = \new_[24844]_  & \new_[24833]_ ;
  assign \new_[2982]_  = \new_[24822]_  & \new_[24811]_ ;
  assign \new_[2983]_  = \new_[24800]_  & \new_[24789]_ ;
  assign \new_[2984]_  = \new_[24778]_  & \new_[24767]_ ;
  assign \new_[2985]_  = \new_[24756]_  & \new_[24745]_ ;
  assign \new_[2986]_  = \new_[24734]_  & \new_[24723]_ ;
  assign \new_[2987]_  = \new_[24712]_  & \new_[24701]_ ;
  assign \new_[2988]_  = \new_[24690]_  & \new_[24679]_ ;
  assign \new_[2989]_  = \new_[24668]_  & \new_[24657]_ ;
  assign \new_[2990]_  = \new_[24646]_  & \new_[24635]_ ;
  assign \new_[2991]_  = \new_[24624]_  & \new_[24613]_ ;
  assign \new_[2992]_  = \new_[24602]_  & \new_[24591]_ ;
  assign \new_[2993]_  = \new_[24580]_  & \new_[24569]_ ;
  assign \new_[2994]_  = \new_[24558]_  & \new_[24547]_ ;
  assign \new_[2995]_  = \new_[24536]_  & \new_[24525]_ ;
  assign \new_[2996]_  = \new_[24514]_  & \new_[24503]_ ;
  assign \new_[2997]_  = \new_[24492]_  & \new_[24481]_ ;
  assign \new_[2998]_  = \new_[24470]_  & \new_[24459]_ ;
  assign \new_[2999]_  = \new_[24448]_  & \new_[24437]_ ;
  assign \new_[3000]_  = \new_[24426]_  & \new_[24415]_ ;
  assign \new_[3001]_  = \new_[24404]_  & \new_[24393]_ ;
  assign \new_[3002]_  = \new_[24382]_  & \new_[24371]_ ;
  assign \new_[3003]_  = \new_[24360]_  & \new_[24349]_ ;
  assign \new_[3004]_  = \new_[24338]_  & \new_[24327]_ ;
  assign \new_[3005]_  = \new_[24316]_  & \new_[24305]_ ;
  assign \new_[3006]_  = \new_[24294]_  & \new_[24283]_ ;
  assign \new_[3007]_  = \new_[24272]_  & \new_[24261]_ ;
  assign \new_[3008]_  = \new_[24250]_  & \new_[24239]_ ;
  assign \new_[3009]_  = \new_[24228]_  & \new_[24217]_ ;
  assign \new_[3010]_  = \new_[24206]_  & \new_[24195]_ ;
  assign \new_[3011]_  = \new_[24184]_  & \new_[24173]_ ;
  assign \new_[3012]_  = \new_[24162]_  & \new_[24151]_ ;
  assign \new_[3013]_  = \new_[24140]_  & \new_[24129]_ ;
  assign \new_[3014]_  = \new_[24118]_  & \new_[24107]_ ;
  assign \new_[3015]_  = \new_[24096]_  & \new_[24085]_ ;
  assign \new_[3016]_  = \new_[24074]_  & \new_[24063]_ ;
  assign \new_[3017]_  = \new_[24052]_  & \new_[24041]_ ;
  assign \new_[3018]_  = \new_[24030]_  & \new_[24019]_ ;
  assign \new_[3019]_  = \new_[24008]_  & \new_[23997]_ ;
  assign \new_[3020]_  = \new_[23986]_  & \new_[23975]_ ;
  assign \new_[3021]_  = \new_[23964]_  & \new_[23953]_ ;
  assign \new_[3022]_  = \new_[23942]_  & \new_[23931]_ ;
  assign \new_[3023]_  = \new_[23920]_  & \new_[23909]_ ;
  assign \new_[3024]_  = \new_[23898]_  & \new_[23887]_ ;
  assign \new_[3025]_  = \new_[23876]_  & \new_[23865]_ ;
  assign \new_[3026]_  = \new_[23854]_  & \new_[23843]_ ;
  assign \new_[3027]_  = \new_[23832]_  & \new_[23821]_ ;
  assign \new_[3028]_  = \new_[23810]_  & \new_[23799]_ ;
  assign \new_[3029]_  = \new_[23788]_  & \new_[23777]_ ;
  assign \new_[3030]_  = \new_[23766]_  & \new_[23755]_ ;
  assign \new_[3031]_  = \new_[23744]_  & \new_[23733]_ ;
  assign \new_[3032]_  = \new_[23722]_  & \new_[23711]_ ;
  assign \new_[3033]_  = \new_[23700]_  & \new_[23689]_ ;
  assign \new_[3034]_  = \new_[23678]_  & \new_[23667]_ ;
  assign \new_[3035]_  = \new_[23656]_  & \new_[23645]_ ;
  assign \new_[3036]_  = \new_[23634]_  & \new_[23623]_ ;
  assign \new_[3037]_  = \new_[23612]_  & \new_[23601]_ ;
  assign \new_[3038]_  = \new_[23590]_  & \new_[23579]_ ;
  assign \new_[3039]_  = \new_[23568]_  & \new_[23557]_ ;
  assign \new_[3040]_  = \new_[23546]_  & \new_[23535]_ ;
  assign \new_[3041]_  = \new_[23524]_  & \new_[23513]_ ;
  assign \new_[3042]_  = \new_[23502]_  & \new_[23491]_ ;
  assign \new_[3043]_  = \new_[23480]_  & \new_[23469]_ ;
  assign \new_[3044]_  = \new_[23458]_  & \new_[23447]_ ;
  assign \new_[3045]_  = \new_[23436]_  & \new_[23425]_ ;
  assign \new_[3046]_  = \new_[23414]_  & \new_[23403]_ ;
  assign \new_[3047]_  = \new_[23392]_  & \new_[23381]_ ;
  assign \new_[3048]_  = \new_[23370]_  & \new_[23359]_ ;
  assign \new_[3049]_  = \new_[23348]_  & \new_[23337]_ ;
  assign \new_[3050]_  = \new_[23326]_  & \new_[23315]_ ;
  assign \new_[3051]_  = \new_[23304]_  & \new_[23293]_ ;
  assign \new_[3052]_  = \new_[23282]_  & \new_[23271]_ ;
  assign \new_[3053]_  = \new_[23260]_  & \new_[23249]_ ;
  assign \new_[3054]_  = \new_[23238]_  & \new_[23227]_ ;
  assign \new_[3055]_  = \new_[23216]_  & \new_[23205]_ ;
  assign \new_[3056]_  = \new_[23196]_  & \new_[23185]_ ;
  assign \new_[3057]_  = \new_[23176]_  & \new_[23165]_ ;
  assign \new_[3058]_  = \new_[23156]_  & \new_[23145]_ ;
  assign \new_[3059]_  = \new_[23136]_  & \new_[23125]_ ;
  assign \new_[3060]_  = \new_[23116]_  & \new_[23105]_ ;
  assign \new_[3061]_  = \new_[23096]_  & \new_[23085]_ ;
  assign \new_[3062]_  = \new_[23076]_  & \new_[23065]_ ;
  assign \new_[3063]_  = \new_[23056]_  & \new_[23045]_ ;
  assign \new_[3064]_  = \new_[23036]_  & \new_[23025]_ ;
  assign \new_[3065]_  = \new_[23016]_  & \new_[23005]_ ;
  assign \new_[3066]_  = \new_[22996]_  & \new_[22985]_ ;
  assign \new_[3067]_  = \new_[22976]_  & \new_[22965]_ ;
  assign \new_[3068]_  = \new_[22956]_  & \new_[22945]_ ;
  assign \new_[3069]_  = \new_[22936]_  & \new_[22925]_ ;
  assign \new_[3070]_  = \new_[22916]_  & \new_[22905]_ ;
  assign \new_[3071]_  = \new_[22896]_  & \new_[22885]_ ;
  assign \new_[3072]_  = \new_[22876]_  & \new_[22865]_ ;
  assign \new_[3073]_  = \new_[22856]_  & \new_[22845]_ ;
  assign \new_[3074]_  = \new_[22836]_  & \new_[22825]_ ;
  assign \new_[3075]_  = \new_[22816]_  & \new_[22805]_ ;
  assign \new_[3076]_  = \new_[22796]_  & \new_[22785]_ ;
  assign \new_[3077]_  = \new_[22776]_  & \new_[22765]_ ;
  assign \new_[3078]_  = \new_[22756]_  & \new_[22745]_ ;
  assign \new_[3079]_  = \new_[22736]_  & \new_[22725]_ ;
  assign \new_[3080]_  = \new_[22716]_  & \new_[22705]_ ;
  assign \new_[3081]_  = \new_[22696]_  & \new_[22685]_ ;
  assign \new_[3082]_  = \new_[22676]_  & \new_[22665]_ ;
  assign \new_[3083]_  = \new_[22656]_  & \new_[22645]_ ;
  assign \new_[3084]_  = \new_[22636]_  & \new_[22625]_ ;
  assign \new_[3085]_  = \new_[22616]_  & \new_[22605]_ ;
  assign \new_[3086]_  = \new_[22596]_  & \new_[22585]_ ;
  assign \new_[3087]_  = \new_[22576]_  & \new_[22565]_ ;
  assign \new_[3088]_  = \new_[22556]_  & \new_[22545]_ ;
  assign \new_[3089]_  = \new_[22536]_  & \new_[22525]_ ;
  assign \new_[3090]_  = \new_[22516]_  & \new_[22505]_ ;
  assign \new_[3091]_  = \new_[22496]_  & \new_[22485]_ ;
  assign \new_[3092]_  = \new_[22476]_  & \new_[22465]_ ;
  assign \new_[3093]_  = \new_[22456]_  & \new_[22445]_ ;
  assign \new_[3094]_  = \new_[22436]_  & \new_[22425]_ ;
  assign \new_[3095]_  = \new_[22416]_  & \new_[22405]_ ;
  assign \new_[3096]_  = \new_[22396]_  & \new_[22385]_ ;
  assign \new_[3097]_  = \new_[22376]_  & \new_[22365]_ ;
  assign \new_[3098]_  = \new_[22356]_  & \new_[22345]_ ;
  assign \new_[3099]_  = \new_[22336]_  & \new_[22325]_ ;
  assign \new_[3100]_  = \new_[22316]_  & \new_[22305]_ ;
  assign \new_[3101]_  = \new_[22296]_  & \new_[22285]_ ;
  assign \new_[3102]_  = \new_[22276]_  & \new_[22265]_ ;
  assign \new_[3103]_  = \new_[22256]_  & \new_[22245]_ ;
  assign \new_[3104]_  = \new_[22236]_  & \new_[22225]_ ;
  assign \new_[3105]_  = \new_[22216]_  & \new_[22205]_ ;
  assign \new_[3106]_  = \new_[22196]_  & \new_[22185]_ ;
  assign \new_[3107]_  = \new_[22176]_  & \new_[22165]_ ;
  assign \new_[3108]_  = \new_[22156]_  & \new_[22145]_ ;
  assign \new_[3109]_  = \new_[22136]_  & \new_[22125]_ ;
  assign \new_[3110]_  = \new_[22116]_  & \new_[22105]_ ;
  assign \new_[3111]_  = \new_[22096]_  & \new_[22085]_ ;
  assign \new_[3112]_  = \new_[22076]_  & \new_[22065]_ ;
  assign \new_[3113]_  = \new_[22056]_  & \new_[22045]_ ;
  assign \new_[3114]_  = \new_[22036]_  & \new_[22025]_ ;
  assign \new_[3115]_  = \new_[22016]_  & \new_[22005]_ ;
  assign \new_[3116]_  = \new_[21996]_  & \new_[21985]_ ;
  assign \new_[3117]_  = \new_[21976]_  & \new_[21965]_ ;
  assign \new_[3118]_  = \new_[21956]_  & \new_[21945]_ ;
  assign \new_[3119]_  = \new_[21936]_  & \new_[21925]_ ;
  assign \new_[3120]_  = \new_[21916]_  & \new_[21905]_ ;
  assign \new_[3121]_  = \new_[21896]_  & \new_[21885]_ ;
  assign \new_[3122]_  = \new_[21876]_  & \new_[21865]_ ;
  assign \new_[3123]_  = \new_[21856]_  & \new_[21845]_ ;
  assign \new_[3124]_  = \new_[21836]_  & \new_[21825]_ ;
  assign \new_[3125]_  = \new_[21816]_  & \new_[21805]_ ;
  assign \new_[3126]_  = \new_[21796]_  & \new_[21785]_ ;
  assign \new_[3127]_  = \new_[21776]_  & \new_[21765]_ ;
  assign \new_[3128]_  = \new_[21756]_  & \new_[21745]_ ;
  assign \new_[3129]_  = \new_[21736]_  & \new_[21725]_ ;
  assign \new_[3130]_  = \new_[21716]_  & \new_[21705]_ ;
  assign \new_[3131]_  = \new_[21696]_  & \new_[21685]_ ;
  assign \new_[3132]_  = \new_[21676]_  & \new_[21665]_ ;
  assign \new_[3133]_  = \new_[21656]_  & \new_[21645]_ ;
  assign \new_[3134]_  = \new_[21636]_  & \new_[21625]_ ;
  assign \new_[3135]_  = \new_[21616]_  & \new_[21605]_ ;
  assign \new_[3136]_  = \new_[21596]_  & \new_[21585]_ ;
  assign \new_[3137]_  = \new_[21576]_  & \new_[21565]_ ;
  assign \new_[3138]_  = \new_[21556]_  & \new_[21545]_ ;
  assign \new_[3139]_  = \new_[21536]_  & \new_[21525]_ ;
  assign \new_[3140]_  = \new_[21516]_  & \new_[21505]_ ;
  assign \new_[3141]_  = \new_[21496]_  & \new_[21485]_ ;
  assign \new_[3142]_  = \new_[21476]_  & \new_[21465]_ ;
  assign \new_[3143]_  = \new_[21456]_  & \new_[21445]_ ;
  assign \new_[3144]_  = \new_[21436]_  & \new_[21425]_ ;
  assign \new_[3145]_  = \new_[21416]_  & \new_[21405]_ ;
  assign \new_[3146]_  = \new_[21396]_  & \new_[21385]_ ;
  assign \new_[3147]_  = \new_[21376]_  & \new_[21365]_ ;
  assign \new_[3148]_  = \new_[21356]_  & \new_[21345]_ ;
  assign \new_[3149]_  = \new_[21336]_  & \new_[21325]_ ;
  assign \new_[3150]_  = \new_[21316]_  & \new_[21305]_ ;
  assign \new_[3151]_  = \new_[21296]_  & \new_[21285]_ ;
  assign \new_[3152]_  = \new_[21276]_  & \new_[21265]_ ;
  assign \new_[3153]_  = \new_[21256]_  & \new_[21245]_ ;
  assign \new_[3154]_  = \new_[21236]_  & \new_[21225]_ ;
  assign \new_[3155]_  = \new_[21216]_  & \new_[21205]_ ;
  assign \new_[3156]_  = \new_[21196]_  & \new_[21185]_ ;
  assign \new_[3157]_  = \new_[21176]_  & \new_[21165]_ ;
  assign \new_[3158]_  = \new_[21156]_  & \new_[21145]_ ;
  assign \new_[3159]_  = \new_[21136]_  & \new_[21125]_ ;
  assign \new_[3160]_  = \new_[21116]_  & \new_[21105]_ ;
  assign \new_[3161]_  = \new_[21096]_  & \new_[21085]_ ;
  assign \new_[3162]_  = \new_[21076]_  & \new_[21065]_ ;
  assign \new_[3163]_  = \new_[21056]_  & \new_[21045]_ ;
  assign \new_[3164]_  = \new_[21036]_  & \new_[21025]_ ;
  assign \new_[3165]_  = \new_[21016]_  & \new_[21005]_ ;
  assign \new_[3166]_  = \new_[20996]_  & \new_[20985]_ ;
  assign \new_[3167]_  = \new_[20976]_  & \new_[20965]_ ;
  assign \new_[3168]_  = \new_[20956]_  & \new_[20945]_ ;
  assign \new_[3169]_  = \new_[20936]_  & \new_[20925]_ ;
  assign \new_[3170]_  = \new_[20916]_  & \new_[20905]_ ;
  assign \new_[3171]_  = \new_[20896]_  & \new_[20885]_ ;
  assign \new_[3172]_  = \new_[20876]_  & \new_[20865]_ ;
  assign \new_[3173]_  = \new_[20856]_  & \new_[20845]_ ;
  assign \new_[3174]_  = \new_[20836]_  & \new_[20825]_ ;
  assign \new_[3175]_  = \new_[20816]_  & \new_[20805]_ ;
  assign \new_[3176]_  = \new_[20796]_  & \new_[20785]_ ;
  assign \new_[3177]_  = \new_[20776]_  & \new_[20765]_ ;
  assign \new_[3178]_  = \new_[20756]_  & \new_[20745]_ ;
  assign \new_[3179]_  = \new_[20736]_  & \new_[20725]_ ;
  assign \new_[3180]_  = \new_[20716]_  & \new_[20705]_ ;
  assign \new_[3181]_  = \new_[20696]_  & \new_[20685]_ ;
  assign \new_[3182]_  = \new_[20676]_  & \new_[20665]_ ;
  assign \new_[3183]_  = \new_[20656]_  & \new_[20645]_ ;
  assign \new_[3184]_  = \new_[20636]_  & \new_[20625]_ ;
  assign \new_[3185]_  = \new_[20616]_  & \new_[20605]_ ;
  assign \new_[3186]_  = \new_[20596]_  & \new_[20585]_ ;
  assign \new_[3187]_  = \new_[20576]_  & \new_[20565]_ ;
  assign \new_[3188]_  = \new_[20556]_  & \new_[20545]_ ;
  assign \new_[3189]_  = \new_[20536]_  & \new_[20525]_ ;
  assign \new_[3190]_  = \new_[20516]_  & \new_[20505]_ ;
  assign \new_[3191]_  = \new_[20496]_  & \new_[20485]_ ;
  assign \new_[3192]_  = \new_[20476]_  & \new_[20465]_ ;
  assign \new_[3193]_  = \new_[20456]_  & \new_[20445]_ ;
  assign \new_[3194]_  = \new_[20436]_  & \new_[20425]_ ;
  assign \new_[3195]_  = \new_[20416]_  & \new_[20405]_ ;
  assign \new_[3196]_  = \new_[20396]_  & \new_[20385]_ ;
  assign \new_[3197]_  = \new_[20376]_  & \new_[20365]_ ;
  assign \new_[3198]_  = \new_[20356]_  & \new_[20345]_ ;
  assign \new_[3199]_  = \new_[20336]_  & \new_[20325]_ ;
  assign \new_[3200]_  = \new_[20316]_  & \new_[20305]_ ;
  assign \new_[3201]_  = \new_[20296]_  & \new_[20285]_ ;
  assign \new_[3202]_  = \new_[20276]_  & \new_[20265]_ ;
  assign \new_[3203]_  = \new_[20256]_  & \new_[20245]_ ;
  assign \new_[3204]_  = \new_[20236]_  & \new_[20225]_ ;
  assign \new_[3205]_  = \new_[20216]_  & \new_[20205]_ ;
  assign \new_[3206]_  = \new_[20196]_  & \new_[20185]_ ;
  assign \new_[3207]_  = \new_[20176]_  & \new_[20165]_ ;
  assign \new_[3208]_  = \new_[20156]_  & \new_[20145]_ ;
  assign \new_[3209]_  = \new_[20136]_  & \new_[20125]_ ;
  assign \new_[3210]_  = \new_[20116]_  & \new_[20105]_ ;
  assign \new_[3211]_  = \new_[20096]_  & \new_[20085]_ ;
  assign \new_[3212]_  = \new_[20076]_  & \new_[20065]_ ;
  assign \new_[3213]_  = \new_[20056]_  & \new_[20045]_ ;
  assign \new_[3214]_  = \new_[20036]_  & \new_[20025]_ ;
  assign \new_[3215]_  = \new_[20016]_  & \new_[20005]_ ;
  assign \new_[3216]_  = \new_[19996]_  & \new_[19985]_ ;
  assign \new_[3217]_  = \new_[19976]_  & \new_[19965]_ ;
  assign \new_[3218]_  = \new_[19956]_  & \new_[19945]_ ;
  assign \new_[3219]_  = \new_[19936]_  & \new_[19925]_ ;
  assign \new_[3220]_  = \new_[19916]_  & \new_[19905]_ ;
  assign \new_[3221]_  = \new_[19896]_  & \new_[19885]_ ;
  assign \new_[3222]_  = \new_[19876]_  & \new_[19865]_ ;
  assign \new_[3223]_  = \new_[19856]_  & \new_[19845]_ ;
  assign \new_[3224]_  = \new_[19836]_  & \new_[19825]_ ;
  assign \new_[3225]_  = \new_[19816]_  & \new_[19805]_ ;
  assign \new_[3226]_  = \new_[19796]_  & \new_[19785]_ ;
  assign \new_[3227]_  = \new_[19776]_  & \new_[19765]_ ;
  assign \new_[3228]_  = \new_[19756]_  & \new_[19745]_ ;
  assign \new_[3229]_  = \new_[19736]_  & \new_[19725]_ ;
  assign \new_[3230]_  = \new_[19716]_  & \new_[19705]_ ;
  assign \new_[3231]_  = \new_[19696]_  & \new_[19685]_ ;
  assign \new_[3232]_  = \new_[19676]_  & \new_[19665]_ ;
  assign \new_[3233]_  = \new_[19656]_  & \new_[19645]_ ;
  assign \new_[3234]_  = \new_[19636]_  & \new_[19625]_ ;
  assign \new_[3235]_  = \new_[19616]_  & \new_[19605]_ ;
  assign \new_[3236]_  = \new_[19596]_  & \new_[19585]_ ;
  assign \new_[3237]_  = \new_[19576]_  & \new_[19565]_ ;
  assign \new_[3238]_  = \new_[19556]_  & \new_[19545]_ ;
  assign \new_[3239]_  = \new_[19536]_  & \new_[19525]_ ;
  assign \new_[3240]_  = \new_[19516]_  & \new_[19505]_ ;
  assign \new_[3241]_  = \new_[19496]_  & \new_[19485]_ ;
  assign \new_[3242]_  = \new_[19476]_  & \new_[19465]_ ;
  assign \new_[3243]_  = \new_[19456]_  & \new_[19445]_ ;
  assign \new_[3244]_  = \new_[19436]_  & \new_[19425]_ ;
  assign \new_[3245]_  = \new_[19416]_  & \new_[19405]_ ;
  assign \new_[3246]_  = \new_[19396]_  & \new_[19385]_ ;
  assign \new_[3247]_  = \new_[19376]_  & \new_[19365]_ ;
  assign \new_[3248]_  = \new_[19356]_  & \new_[19345]_ ;
  assign \new_[3249]_  = \new_[19336]_  & \new_[19325]_ ;
  assign \new_[3250]_  = \new_[19316]_  & \new_[19305]_ ;
  assign \new_[3251]_  = \new_[19296]_  & \new_[19285]_ ;
  assign \new_[3252]_  = \new_[19276]_  & \new_[19265]_ ;
  assign \new_[3253]_  = \new_[19256]_  & \new_[19245]_ ;
  assign \new_[3254]_  = \new_[19236]_  & \new_[19225]_ ;
  assign \new_[3255]_  = \new_[19216]_  & \new_[19205]_ ;
  assign \new_[3256]_  = \new_[19196]_  & \new_[19185]_ ;
  assign \new_[3257]_  = \new_[19176]_  & \new_[19165]_ ;
  assign \new_[3258]_  = \new_[19156]_  & \new_[19145]_ ;
  assign \new_[3259]_  = \new_[19136]_  & \new_[19125]_ ;
  assign \new_[3260]_  = \new_[19116]_  & \new_[19105]_ ;
  assign \new_[3261]_  = \new_[19096]_  & \new_[19085]_ ;
  assign \new_[3262]_  = \new_[19076]_  & \new_[19065]_ ;
  assign \new_[3263]_  = \new_[19056]_  & \new_[19045]_ ;
  assign \new_[3264]_  = \new_[19036]_  & \new_[19025]_ ;
  assign \new_[3265]_  = \new_[19016]_  & \new_[19005]_ ;
  assign \new_[3266]_  = \new_[18996]_  & \new_[18985]_ ;
  assign \new_[3267]_  = \new_[18976]_  & \new_[18965]_ ;
  assign \new_[3268]_  = \new_[18956]_  & \new_[18945]_ ;
  assign \new_[3269]_  = \new_[18936]_  & \new_[18925]_ ;
  assign \new_[3270]_  = \new_[18916]_  & \new_[18905]_ ;
  assign \new_[3271]_  = \new_[18896]_  & \new_[18885]_ ;
  assign \new_[3272]_  = \new_[18876]_  & \new_[18865]_ ;
  assign \new_[3273]_  = \new_[18856]_  & \new_[18845]_ ;
  assign \new_[3274]_  = \new_[18836]_  & \new_[18825]_ ;
  assign \new_[3275]_  = \new_[18816]_  & \new_[18805]_ ;
  assign \new_[3276]_  = \new_[18796]_  & \new_[18785]_ ;
  assign \new_[3277]_  = \new_[18776]_  & \new_[18765]_ ;
  assign \new_[3278]_  = \new_[18756]_  & \new_[18745]_ ;
  assign \new_[3279]_  = \new_[18736]_  & \new_[18725]_ ;
  assign \new_[3280]_  = \new_[18716]_  & \new_[18705]_ ;
  assign \new_[3281]_  = \new_[18696]_  & \new_[18685]_ ;
  assign \new_[3282]_  = \new_[18676]_  & \new_[18665]_ ;
  assign \new_[3283]_  = \new_[18656]_  & \new_[18645]_ ;
  assign \new_[3284]_  = \new_[18636]_  & \new_[18625]_ ;
  assign \new_[3285]_  = \new_[18616]_  & \new_[18605]_ ;
  assign \new_[3286]_  = \new_[18596]_  & \new_[18585]_ ;
  assign \new_[3287]_  = \new_[18576]_  & \new_[18565]_ ;
  assign \new_[3288]_  = \new_[18556]_  & \new_[18545]_ ;
  assign \new_[3289]_  = \new_[18536]_  & \new_[18525]_ ;
  assign \new_[3290]_  = \new_[18516]_  & \new_[18505]_ ;
  assign \new_[3291]_  = \new_[18496]_  & \new_[18485]_ ;
  assign \new_[3292]_  = \new_[18476]_  & \new_[18465]_ ;
  assign \new_[3293]_  = \new_[18456]_  & \new_[18445]_ ;
  assign \new_[3294]_  = \new_[18436]_  & \new_[18425]_ ;
  assign \new_[3295]_  = \new_[18416]_  & \new_[18405]_ ;
  assign \new_[3296]_  = \new_[18396]_  & \new_[18385]_ ;
  assign \new_[3297]_  = \new_[18376]_  & \new_[18365]_ ;
  assign \new_[3298]_  = \new_[18356]_  & \new_[18345]_ ;
  assign \new_[3299]_  = \new_[18336]_  & \new_[18325]_ ;
  assign \new_[3300]_  = \new_[18316]_  & \new_[18305]_ ;
  assign \new_[3301]_  = \new_[18296]_  & \new_[18285]_ ;
  assign \new_[3302]_  = \new_[18276]_  & \new_[18265]_ ;
  assign \new_[3303]_  = \new_[18256]_  & \new_[18245]_ ;
  assign \new_[3304]_  = \new_[18236]_  & \new_[18225]_ ;
  assign \new_[3305]_  = \new_[18216]_  & \new_[18205]_ ;
  assign \new_[3306]_  = \new_[18196]_  & \new_[18185]_ ;
  assign \new_[3307]_  = \new_[18176]_  & \new_[18165]_ ;
  assign \new_[3308]_  = \new_[18156]_  & \new_[18145]_ ;
  assign \new_[3309]_  = \new_[18136]_  & \new_[18125]_ ;
  assign \new_[3310]_  = \new_[18116]_  & \new_[18105]_ ;
  assign \new_[3311]_  = \new_[18096]_  & \new_[18085]_ ;
  assign \new_[3312]_  = \new_[18076]_  & \new_[18065]_ ;
  assign \new_[3313]_  = \new_[18056]_  & \new_[18045]_ ;
  assign \new_[3314]_  = \new_[18036]_  & \new_[18025]_ ;
  assign \new_[3315]_  = \new_[18016]_  & \new_[18005]_ ;
  assign \new_[3316]_  = \new_[17996]_  & \new_[17985]_ ;
  assign \new_[3317]_  = \new_[17976]_  & \new_[17965]_ ;
  assign \new_[3318]_  = \new_[17956]_  & \new_[17945]_ ;
  assign \new_[3319]_  = \new_[17936]_  & \new_[17925]_ ;
  assign \new_[3320]_  = \new_[17916]_  & \new_[17905]_ ;
  assign \new_[3321]_  = \new_[17896]_  & \new_[17885]_ ;
  assign \new_[3322]_  = \new_[17876]_  & \new_[17865]_ ;
  assign \new_[3323]_  = \new_[17856]_  & \new_[17845]_ ;
  assign \new_[3324]_  = \new_[17836]_  & \new_[17825]_ ;
  assign \new_[3325]_  = \new_[17816]_  & \new_[17805]_ ;
  assign \new_[3326]_  = \new_[17796]_  & \new_[17785]_ ;
  assign \new_[3327]_  = \new_[17776]_  & \new_[17765]_ ;
  assign \new_[3328]_  = \new_[17756]_  & \new_[17745]_ ;
  assign \new_[3329]_  = \new_[17736]_  & \new_[17725]_ ;
  assign \new_[3330]_  = \new_[17716]_  & \new_[17705]_ ;
  assign \new_[3331]_  = \new_[17696]_  & \new_[17685]_ ;
  assign \new_[3332]_  = \new_[17676]_  & \new_[17665]_ ;
  assign \new_[3333]_  = \new_[17656]_  & \new_[17645]_ ;
  assign \new_[3334]_  = \new_[17636]_  & \new_[17625]_ ;
  assign \new_[3335]_  = \new_[17616]_  & \new_[17605]_ ;
  assign \new_[3336]_  = \new_[17596]_  & \new_[17585]_ ;
  assign \new_[3337]_  = \new_[17576]_  & \new_[17565]_ ;
  assign \new_[3338]_  = \new_[17556]_  & \new_[17545]_ ;
  assign \new_[3339]_  = \new_[17536]_  & \new_[17525]_ ;
  assign \new_[3340]_  = \new_[17516]_  & \new_[17505]_ ;
  assign \new_[3341]_  = \new_[17496]_  & \new_[17485]_ ;
  assign \new_[3342]_  = \new_[17476]_  & \new_[17465]_ ;
  assign \new_[3343]_  = \new_[17456]_  & \new_[17445]_ ;
  assign \new_[3344]_  = \new_[17436]_  & \new_[17425]_ ;
  assign \new_[3345]_  = \new_[17416]_  & \new_[17405]_ ;
  assign \new_[3346]_  = \new_[17396]_  & \new_[17385]_ ;
  assign \new_[3347]_  = \new_[17376]_  & \new_[17365]_ ;
  assign \new_[3348]_  = \new_[17356]_  & \new_[17345]_ ;
  assign \new_[3349]_  = \new_[17336]_  & \new_[17325]_ ;
  assign \new_[3350]_  = \new_[17316]_  & \new_[17305]_ ;
  assign \new_[3351]_  = \new_[17296]_  & \new_[17285]_ ;
  assign \new_[3352]_  = \new_[17276]_  & \new_[17265]_ ;
  assign \new_[3353]_  = \new_[17256]_  & \new_[17245]_ ;
  assign \new_[3354]_  = \new_[17236]_  & \new_[17225]_ ;
  assign \new_[3355]_  = \new_[17216]_  & \new_[17205]_ ;
  assign \new_[3356]_  = \new_[17196]_  & \new_[17185]_ ;
  assign \new_[3357]_  = \new_[17176]_  & \new_[17165]_ ;
  assign \new_[3358]_  = \new_[17156]_  & \new_[17145]_ ;
  assign \new_[3359]_  = \new_[17136]_  & \new_[17125]_ ;
  assign \new_[3360]_  = \new_[17116]_  & \new_[17105]_ ;
  assign \new_[3361]_  = \new_[17096]_  & \new_[17085]_ ;
  assign \new_[3362]_  = \new_[17076]_  & \new_[17065]_ ;
  assign \new_[3363]_  = \new_[17056]_  & \new_[17045]_ ;
  assign \new_[3364]_  = \new_[17036]_  & \new_[17025]_ ;
  assign \new_[3365]_  = \new_[17016]_  & \new_[17005]_ ;
  assign \new_[3366]_  = \new_[16996]_  & \new_[16985]_ ;
  assign \new_[3367]_  = \new_[16976]_  & \new_[16965]_ ;
  assign \new_[3368]_  = \new_[16956]_  & \new_[16945]_ ;
  assign \new_[3369]_  = \new_[16936]_  & \new_[16925]_ ;
  assign \new_[3370]_  = \new_[16916]_  & \new_[16905]_ ;
  assign \new_[3371]_  = \new_[16896]_  & \new_[16885]_ ;
  assign \new_[3372]_  = \new_[16876]_  & \new_[16865]_ ;
  assign \new_[3373]_  = \new_[16856]_  & \new_[16845]_ ;
  assign \new_[3374]_  = \new_[16836]_  & \new_[16825]_ ;
  assign \new_[3375]_  = \new_[16816]_  & \new_[16807]_ ;
  assign \new_[3376]_  = \new_[16798]_  & \new_[16789]_ ;
  assign \new_[3377]_  = \new_[16780]_  & \new_[16771]_ ;
  assign \new_[3378]_  = \new_[16762]_  & \new_[16753]_ ;
  assign \new_[3379]_  = \new_[16744]_  & \new_[16735]_ ;
  assign \new_[3380]_  = \new_[16726]_  & \new_[16717]_ ;
  assign \new_[3381]_  = \new_[16708]_  & \new_[16699]_ ;
  assign \new_[3382]_  = \new_[16690]_  & \new_[16681]_ ;
  assign \new_[3383]_  = \new_[16672]_  & \new_[16663]_ ;
  assign \new_[3384]_  = \new_[16654]_  & \new_[16645]_ ;
  assign \new_[3385]_  = \new_[16636]_  & \new_[16627]_ ;
  assign \new_[3386]_  = \new_[16618]_  & \new_[16609]_ ;
  assign \new_[3387]_  = \new_[16600]_  & \new_[16591]_ ;
  assign \new_[3388]_  = \new_[16582]_  & \new_[16573]_ ;
  assign \new_[3389]_  = \new_[16564]_  & \new_[16555]_ ;
  assign \new_[3390]_  = \new_[16546]_  & \new_[16537]_ ;
  assign \new_[3391]_  = \new_[16528]_  & \new_[16519]_ ;
  assign \new_[3392]_  = \new_[16510]_  & \new_[16501]_ ;
  assign \new_[3393]_  = \new_[16492]_  & \new_[16483]_ ;
  assign \new_[3394]_  = \new_[16474]_  & \new_[16465]_ ;
  assign \new_[3395]_  = \new_[16456]_  & \new_[16447]_ ;
  assign \new_[3396]_  = \new_[16438]_  & \new_[16429]_ ;
  assign \new_[3397]_  = \new_[16420]_  & \new_[16411]_ ;
  assign \new_[3398]_  = \new_[16402]_  & \new_[16393]_ ;
  assign \new_[3399]_  = \new_[16384]_  & \new_[16375]_ ;
  assign \new_[3400]_  = \new_[16366]_  & \new_[16357]_ ;
  assign \new_[3401]_  = \new_[16348]_  & \new_[16339]_ ;
  assign \new_[3402]_  = \new_[16330]_  & \new_[16321]_ ;
  assign \new_[3403]_  = \new_[16312]_  & \new_[16303]_ ;
  assign \new_[3404]_  = \new_[16294]_  & \new_[16285]_ ;
  assign \new_[3405]_  = \new_[16276]_  & \new_[16267]_ ;
  assign \new_[3406]_  = \new_[16258]_  & \new_[16249]_ ;
  assign \new_[3407]_  = \new_[16240]_  & \new_[16231]_ ;
  assign \new_[3408]_  = \new_[16222]_  & \new_[16213]_ ;
  assign \new_[3409]_  = \new_[16204]_  & \new_[16195]_ ;
  assign \new_[3410]_  = \new_[16186]_  & \new_[16177]_ ;
  assign \new_[3411]_  = \new_[16168]_  & \new_[16159]_ ;
  assign \new_[3412]_  = \new_[16150]_  & \new_[16141]_ ;
  assign \new_[3413]_  = \new_[16132]_  & \new_[16123]_ ;
  assign \new_[3414]_  = \new_[16114]_  & \new_[16105]_ ;
  assign \new_[3415]_  = \new_[16096]_  & \new_[16087]_ ;
  assign \new_[3416]_  = \new_[16078]_  & \new_[16069]_ ;
  assign \new_[3417]_  = \new_[16060]_  & \new_[16051]_ ;
  assign \new_[3418]_  = \new_[16042]_  & \new_[16033]_ ;
  assign \new_[3419]_  = \new_[16024]_  & \new_[16015]_ ;
  assign \new_[3420]_  = \new_[16006]_  & \new_[15997]_ ;
  assign \new_[3421]_  = \new_[15988]_  & \new_[15979]_ ;
  assign \new_[3422]_  = \new_[15970]_  & \new_[15961]_ ;
  assign \new_[3423]_  = \new_[15952]_  & \new_[15943]_ ;
  assign \new_[3424]_  = \new_[15934]_  & \new_[15925]_ ;
  assign \new_[3425]_  = \new_[15916]_  & \new_[15907]_ ;
  assign \new_[3426]_  = \new_[15898]_  & \new_[15889]_ ;
  assign \new_[3427]_  = \new_[15880]_  & \new_[15871]_ ;
  assign \new_[3428]_  = \new_[15862]_  & \new_[15853]_ ;
  assign \new_[3429]_  = \new_[15844]_  & \new_[15835]_ ;
  assign \new_[3430]_  = \new_[15826]_  & \new_[15817]_ ;
  assign \new_[3431]_  = \new_[15808]_  & \new_[15799]_ ;
  assign \new_[3432]_  = \new_[15790]_  & \new_[15781]_ ;
  assign \new_[3433]_  = \new_[15772]_  & \new_[15763]_ ;
  assign \new_[3434]_  = \new_[15754]_  & \new_[15745]_ ;
  assign \new_[3435]_  = \new_[15736]_  & \new_[15727]_ ;
  assign \new_[3436]_  = \new_[15718]_  & \new_[15709]_ ;
  assign \new_[3437]_  = \new_[15700]_  & \new_[15691]_ ;
  assign \new_[3438]_  = \new_[15682]_  & \new_[15673]_ ;
  assign \new_[3439]_  = \new_[15664]_  & \new_[15655]_ ;
  assign \new_[3440]_  = \new_[15646]_  & \new_[15637]_ ;
  assign \new_[3441]_  = \new_[15628]_  & \new_[15619]_ ;
  assign \new_[3442]_  = \new_[15610]_  & \new_[15601]_ ;
  assign \new_[3443]_  = \new_[15592]_  & \new_[15583]_ ;
  assign \new_[3444]_  = \new_[15574]_  & \new_[15565]_ ;
  assign \new_[3445]_  = \new_[15556]_  & \new_[15547]_ ;
  assign \new_[3446]_  = \new_[15538]_  & \new_[15529]_ ;
  assign \new_[3447]_  = \new_[15520]_  & \new_[15511]_ ;
  assign \new_[3448]_  = \new_[15502]_  & \new_[15493]_ ;
  assign \new_[3449]_  = \new_[15484]_  & \new_[15475]_ ;
  assign \new_[3450]_  = \new_[15466]_  & \new_[15457]_ ;
  assign \new_[3451]_  = \new_[15448]_  & \new_[15439]_ ;
  assign \new_[3452]_  = \new_[15430]_  & \new_[15421]_ ;
  assign \new_[3453]_  = \new_[15412]_  & \new_[15403]_ ;
  assign \new_[3454]_  = \new_[15394]_  & \new_[15385]_ ;
  assign \new_[3455]_  = \new_[15376]_  & \new_[15367]_ ;
  assign \new_[3456]_  = \new_[15358]_  & \new_[15349]_ ;
  assign \new_[3457]_  = \new_[15340]_  & \new_[15331]_ ;
  assign \new_[3458]_  = \new_[15322]_  & \new_[15313]_ ;
  assign \new_[3459]_  = \new_[15304]_  & \new_[15295]_ ;
  assign \new_[3460]_  = \new_[15286]_  & \new_[15277]_ ;
  assign \new_[3461]_  = \new_[15268]_  & \new_[15259]_ ;
  assign \new_[3462]_  = \new_[15250]_  & \new_[15241]_ ;
  assign \new_[3463]_  = \new_[15232]_  & \new_[15223]_ ;
  assign \new_[3464]_  = \new_[15214]_  & \new_[15205]_ ;
  assign \new_[3465]_  = \new_[15196]_  & \new_[15187]_ ;
  assign \new_[3466]_  = \new_[15178]_  & \new_[15169]_ ;
  assign \new_[3467]_  = \new_[15160]_  & \new_[15151]_ ;
  assign \new_[3468]_  = \new_[15142]_  & \new_[15133]_ ;
  assign \new_[3469]_  = \new_[15124]_  & \new_[15115]_ ;
  assign \new_[3470]_  = \new_[15106]_  & \new_[15097]_ ;
  assign \new_[3471]_  = \new_[15088]_  & \new_[15079]_ ;
  assign \new_[3472]_  = \new_[15070]_  & \new_[15061]_ ;
  assign \new_[3473]_  = \new_[15052]_  & \new_[15043]_ ;
  assign \new_[3474]_  = \new_[15034]_  & \new_[15025]_ ;
  assign \new_[3475]_  = \new_[15016]_  & \new_[15007]_ ;
  assign \new_[3476]_  = \new_[14998]_  & \new_[14989]_ ;
  assign \new_[3477]_  = \new_[14980]_  & \new_[14971]_ ;
  assign \new_[3478]_  = \new_[14962]_  & \new_[14953]_ ;
  assign \new_[3479]_  = \new_[14944]_  & \new_[14935]_ ;
  assign \new_[3480]_  = \new_[14926]_  & \new_[14917]_ ;
  assign \new_[3481]_  = \new_[14908]_  & \new_[14899]_ ;
  assign \new_[3482]_  = \new_[14890]_  & \new_[14881]_ ;
  assign \new_[3483]_  = \new_[14872]_  & \new_[14863]_ ;
  assign \new_[3484]_  = \new_[14854]_  & \new_[14845]_ ;
  assign \new_[3485]_  = \new_[14836]_  & \new_[14827]_ ;
  assign \new_[3486]_  = \new_[14818]_  & \new_[14809]_ ;
  assign \new_[3487]_  = \new_[14800]_  & \new_[14791]_ ;
  assign \new_[3488]_  = \new_[14782]_  & \new_[14773]_ ;
  assign \new_[3489]_  = \new_[14764]_  & \new_[14755]_ ;
  assign \new_[3490]_  = \new_[14746]_  & \new_[14737]_ ;
  assign \new_[3491]_  = \new_[14728]_  & \new_[14719]_ ;
  assign \new_[3492]_  = \new_[14710]_  & \new_[14701]_ ;
  assign \new_[3493]_  = \new_[14692]_  & \new_[14683]_ ;
  assign \new_[3494]_  = \new_[14674]_  & \new_[14665]_ ;
  assign \new_[3495]_  = \new_[14656]_  & \new_[14647]_ ;
  assign \new_[3496]_  = \new_[14638]_  & \new_[14629]_ ;
  assign \new_[3497]_  = \new_[14620]_  & \new_[14611]_ ;
  assign \new_[3498]_  = \new_[14602]_  & \new_[14593]_ ;
  assign \new_[3499]_  = \new_[14584]_  & \new_[14575]_ ;
  assign \new_[3500]_  = \new_[14566]_  & \new_[14557]_ ;
  assign \new_[3501]_  = \new_[14548]_  & \new_[14539]_ ;
  assign \new_[3502]_  = \new_[14530]_  & \new_[14521]_ ;
  assign \new_[3503]_  = \new_[14512]_  & \new_[14503]_ ;
  assign \new_[3504]_  = \new_[14494]_  & \new_[14485]_ ;
  assign \new_[3505]_  = \new_[14476]_  & \new_[14467]_ ;
  assign \new_[3506]_  = \new_[14458]_  & \new_[14449]_ ;
  assign \new_[3507]_  = \new_[14440]_  & \new_[14431]_ ;
  assign \new_[3508]_  = \new_[14422]_  & \new_[14413]_ ;
  assign \new_[3509]_  = \new_[14404]_  & \new_[14395]_ ;
  assign \new_[3510]_  = \new_[14386]_  & \new_[14377]_ ;
  assign \new_[3511]_  = \new_[14368]_  & \new_[14359]_ ;
  assign \new_[3512]_  = \new_[14350]_  & \new_[14341]_ ;
  assign \new_[3513]_  = \new_[14332]_  & \new_[14323]_ ;
  assign \new_[3514]_  = \new_[14314]_  & \new_[14305]_ ;
  assign \new_[3515]_  = \new_[14296]_  & \new_[14287]_ ;
  assign \new_[3516]_  = \new_[14278]_  & \new_[14269]_ ;
  assign \new_[3517]_  = \new_[14260]_  & \new_[14251]_ ;
  assign \new_[3518]_  = \new_[14242]_  & \new_[14233]_ ;
  assign \new_[3519]_  = \new_[14224]_  & \new_[14215]_ ;
  assign \new_[3520]_  = \new_[14206]_  & \new_[14197]_ ;
  assign \new_[3521]_  = \new_[14188]_  & \new_[14179]_ ;
  assign \new_[3522]_  = \new_[14170]_  & \new_[14161]_ ;
  assign \new_[3523]_  = \new_[14152]_  & \new_[14143]_ ;
  assign \new_[3524]_  = \new_[14134]_  & \new_[14125]_ ;
  assign \new_[3525]_  = \new_[14116]_  & \new_[14107]_ ;
  assign \new_[3526]_  = \new_[14098]_  & \new_[14089]_ ;
  assign \new_[3527]_  = \new_[14080]_  & \new_[14071]_ ;
  assign \new_[3528]_  = \new_[14062]_  & \new_[14053]_ ;
  assign \new_[3529]_  = \new_[14044]_  & \new_[14035]_ ;
  assign \new_[3530]_  = \new_[14026]_  & \new_[14017]_ ;
  assign \new_[3531]_  = \new_[14008]_  & \new_[13999]_ ;
  assign \new_[3532]_  = \new_[13990]_  & \new_[13981]_ ;
  assign \new_[3533]_  = \new_[13972]_  & \new_[13963]_ ;
  assign \new_[3534]_  = \new_[13954]_  & \new_[13945]_ ;
  assign \new_[3535]_  = \new_[13936]_  & \new_[13927]_ ;
  assign \new_[3536]_  = \new_[13918]_  & \new_[13909]_ ;
  assign \new_[3537]_  = \new_[13900]_  & \new_[13891]_ ;
  assign \new_[3538]_  = \new_[13882]_  & \new_[13873]_ ;
  assign \new_[3539]_  = \new_[13864]_  & \new_[13855]_ ;
  assign \new_[3540]_  = \new_[13846]_  & \new_[13837]_ ;
  assign \new_[3541]_  = \new_[13828]_  & \new_[13819]_ ;
  assign \new_[3542]_  = \new_[13810]_  & \new_[13801]_ ;
  assign \new_[3543]_  = \new_[13792]_  & \new_[13783]_ ;
  assign \new_[3544]_  = \new_[13774]_  & \new_[13765]_ ;
  assign \new_[3545]_  = \new_[13756]_  & \new_[13747]_ ;
  assign \new_[3546]_  = \new_[13738]_  & \new_[13729]_ ;
  assign \new_[3547]_  = \new_[13720]_  & \new_[13711]_ ;
  assign \new_[3548]_  = \new_[13702]_  & \new_[13693]_ ;
  assign \new_[3549]_  = \new_[13684]_  & \new_[13675]_ ;
  assign \new_[3550]_  = \new_[13666]_  & \new_[13657]_ ;
  assign \new_[3551]_  = \new_[13648]_  & \new_[13639]_ ;
  assign \new_[3552]_  = \new_[13630]_  & \new_[13621]_ ;
  assign \new_[3553]_  = \new_[13612]_  & \new_[13603]_ ;
  assign \new_[3554]_  = \new_[13594]_  & \new_[13585]_ ;
  assign \new_[3555]_  = \new_[13576]_  & \new_[13567]_ ;
  assign \new_[3556]_  = \new_[13558]_  & \new_[13549]_ ;
  assign \new_[3557]_  = \new_[13540]_  & \new_[13531]_ ;
  assign \new_[3558]_  = \new_[13522]_  & \new_[13513]_ ;
  assign \new_[3559]_  = \new_[13504]_  & \new_[13495]_ ;
  assign \new_[3560]_  = \new_[13486]_  & \new_[13477]_ ;
  assign \new_[3561]_  = \new_[13468]_  & \new_[13459]_ ;
  assign \new_[3562]_  = \new_[13450]_  & \new_[13441]_ ;
  assign \new_[3563]_  = \new_[13432]_  & \new_[13423]_ ;
  assign \new_[3564]_  = \new_[13414]_  & \new_[13405]_ ;
  assign \new_[3565]_  = \new_[13396]_  & \new_[13387]_ ;
  assign \new_[3566]_  = \new_[13378]_  & \new_[13369]_ ;
  assign \new_[3567]_  = \new_[13360]_  & \new_[13351]_ ;
  assign \new_[3568]_  = \new_[13342]_  & \new_[13333]_ ;
  assign \new_[3569]_  = \new_[13324]_  & \new_[13315]_ ;
  assign \new_[3570]_  = \new_[13306]_  & \new_[13297]_ ;
  assign \new_[3571]_  = \new_[13288]_  & \new_[13279]_ ;
  assign \new_[3572]_  = \new_[13270]_  & \new_[13261]_ ;
  assign \new_[3573]_  = \new_[13252]_  & \new_[13243]_ ;
  assign \new_[3574]_  = \new_[13234]_  & \new_[13225]_ ;
  assign \new_[3575]_  = \new_[13216]_  & \new_[13207]_ ;
  assign \new_[3576]_  = \new_[13198]_  & \new_[13189]_ ;
  assign \new_[3577]_  = \new_[13180]_  & \new_[13171]_ ;
  assign \new_[3578]_  = \new_[13162]_  & \new_[13153]_ ;
  assign \new_[3579]_  = \new_[13144]_  & \new_[13135]_ ;
  assign \new_[3580]_  = \new_[13126]_  & \new_[13117]_ ;
  assign \new_[3581]_  = \new_[13108]_  & \new_[13099]_ ;
  assign \new_[3582]_  = \new_[13090]_  & \new_[13081]_ ;
  assign \new_[3583]_  = \new_[13072]_  & \new_[13063]_ ;
  assign \new_[3584]_  = \new_[13054]_  & \new_[13045]_ ;
  assign \new_[3585]_  = \new_[13036]_  & \new_[13027]_ ;
  assign \new_[3586]_  = \new_[13018]_  & \new_[13009]_ ;
  assign \new_[3587]_  = \new_[13000]_  & \new_[12991]_ ;
  assign \new_[3588]_  = \new_[12982]_  & \new_[12973]_ ;
  assign \new_[3589]_  = \new_[12964]_  & \new_[12955]_ ;
  assign \new_[3590]_  = \new_[12946]_  & \new_[12937]_ ;
  assign \new_[3591]_  = \new_[12928]_  & \new_[12919]_ ;
  assign \new_[3592]_  = \new_[12910]_  & \new_[12901]_ ;
  assign \new_[3593]_  = \new_[12892]_  & \new_[12883]_ ;
  assign \new_[3594]_  = \new_[12874]_  & \new_[12865]_ ;
  assign \new_[3595]_  = \new_[12856]_  & \new_[12847]_ ;
  assign \new_[3596]_  = \new_[12838]_  & \new_[12829]_ ;
  assign \new_[3597]_  = \new_[12820]_  & \new_[12811]_ ;
  assign \new_[3598]_  = \new_[12802]_  & \new_[12793]_ ;
  assign \new_[3599]_  = \new_[12784]_  & \new_[12775]_ ;
  assign \new_[3600]_  = \new_[12766]_  & \new_[12757]_ ;
  assign \new_[3601]_  = \new_[12748]_  & \new_[12739]_ ;
  assign \new_[3602]_  = \new_[12730]_  & \new_[12721]_ ;
  assign \new_[3603]_  = \new_[12712]_  & \new_[12703]_ ;
  assign \new_[3604]_  = \new_[12694]_  & \new_[12685]_ ;
  assign \new_[3605]_  = \new_[12676]_  & \new_[12667]_ ;
  assign \new_[3606]_  = \new_[12658]_  & \new_[12649]_ ;
  assign \new_[3607]_  = \new_[12640]_  & \new_[12631]_ ;
  assign \new_[3608]_  = \new_[12622]_  & \new_[12613]_ ;
  assign \new_[3609]_  = \new_[12604]_  & \new_[12595]_ ;
  assign \new_[3610]_  = \new_[12586]_  & \new_[12577]_ ;
  assign \new_[3611]_  = \new_[12568]_  & \new_[12559]_ ;
  assign \new_[3612]_  = \new_[12550]_  & \new_[12541]_ ;
  assign \new_[3613]_  = \new_[12532]_  & \new_[12523]_ ;
  assign \new_[3614]_  = \new_[12514]_  & \new_[12505]_ ;
  assign \new_[3615]_  = \new_[12496]_  & \new_[12487]_ ;
  assign \new_[3616]_  = \new_[12478]_  & \new_[12469]_ ;
  assign \new_[3617]_  = \new_[12460]_  & \new_[12451]_ ;
  assign \new_[3618]_  = \new_[12442]_  & \new_[12433]_ ;
  assign \new_[3619]_  = \new_[12424]_  & \new_[12415]_ ;
  assign \new_[3620]_  = \new_[12406]_  & \new_[12397]_ ;
  assign \new_[3621]_  = \new_[12388]_  & \new_[12379]_ ;
  assign \new_[3622]_  = \new_[12370]_  & \new_[12361]_ ;
  assign \new_[3623]_  = \new_[12352]_  & \new_[12343]_ ;
  assign \new_[3624]_  = \new_[12334]_  & \new_[12325]_ ;
  assign \new_[3625]_  = \new_[12316]_  & \new_[12307]_ ;
  assign \new_[3626]_  = \new_[12298]_  & \new_[12289]_ ;
  assign \new_[3627]_  = \new_[12280]_  & \new_[12271]_ ;
  assign \new_[3628]_  = \new_[12262]_  & \new_[12253]_ ;
  assign \new_[3629]_  = \new_[12244]_  & \new_[12235]_ ;
  assign \new_[3630]_  = \new_[12226]_  & \new_[12217]_ ;
  assign \new_[3631]_  = \new_[12208]_  & \new_[12199]_ ;
  assign \new_[3632]_  = \new_[12190]_  & \new_[12181]_ ;
  assign \new_[3633]_  = \new_[12172]_  & \new_[12163]_ ;
  assign \new_[3634]_  = \new_[12154]_  & \new_[12145]_ ;
  assign \new_[3635]_  = \new_[12136]_  & \new_[12127]_ ;
  assign \new_[3636]_  = \new_[12118]_  & \new_[12109]_ ;
  assign \new_[3637]_  = \new_[12100]_  & \new_[12091]_ ;
  assign \new_[3638]_  = \new_[12082]_  & \new_[12073]_ ;
  assign \new_[3639]_  = \new_[12064]_  & \new_[12055]_ ;
  assign \new_[3640]_  = \new_[12048]_  & \new_[12039]_ ;
  assign \new_[3641]_  = \new_[12032]_  & \new_[12023]_ ;
  assign \new_[3642]_  = \new_[12016]_  & \new_[12007]_ ;
  assign \new_[3643]_  = \new_[12000]_  & \new_[11991]_ ;
  assign \new_[3644]_  = \new_[11984]_  & \new_[11975]_ ;
  assign \new_[3645]_  = \new_[11968]_  & \new_[11959]_ ;
  assign \new_[3646]_  = \new_[11952]_  & \new_[11943]_ ;
  assign \new_[3647]_  = \new_[11936]_  & \new_[11927]_ ;
  assign \new_[3648]_  = \new_[11920]_  & \new_[11911]_ ;
  assign \new_[3649]_  = \new_[11904]_  & \new_[11895]_ ;
  assign \new_[3650]_  = \new_[11888]_  & \new_[11879]_ ;
  assign \new_[3651]_  = \new_[11872]_  & \new_[11863]_ ;
  assign \new_[3652]_  = \new_[11856]_  & \new_[11847]_ ;
  assign \new_[3653]_  = \new_[11840]_  & \new_[11831]_ ;
  assign \new_[3654]_  = \new_[11824]_  & \new_[11815]_ ;
  assign \new_[3655]_  = \new_[11808]_  & \new_[11799]_ ;
  assign \new_[3656]_  = \new_[11792]_  & \new_[11783]_ ;
  assign \new_[3657]_  = \new_[11776]_  & \new_[11767]_ ;
  assign \new_[3658]_  = \new_[11760]_  & \new_[11751]_ ;
  assign \new_[3659]_  = \new_[11744]_  & \new_[11735]_ ;
  assign \new_[3660]_  = \new_[11728]_  & \new_[11719]_ ;
  assign \new_[3661]_  = \new_[11712]_  & \new_[11703]_ ;
  assign \new_[3662]_  = \new_[11696]_  & \new_[11687]_ ;
  assign \new_[3663]_  = \new_[11680]_  & \new_[11671]_ ;
  assign \new_[3664]_  = \new_[11664]_  & \new_[11655]_ ;
  assign \new_[3665]_  = \new_[11648]_  & \new_[11639]_ ;
  assign \new_[3666]_  = \new_[11632]_  & \new_[11623]_ ;
  assign \new_[3667]_  = \new_[11616]_  & \new_[11607]_ ;
  assign \new_[3668]_  = \new_[11600]_  & \new_[11591]_ ;
  assign \new_[3669]_  = \new_[11584]_  & \new_[11575]_ ;
  assign \new_[3670]_  = \new_[11568]_  & \new_[11559]_ ;
  assign \new_[3671]_  = \new_[11552]_  & \new_[11545]_ ;
  assign \new_[3672]_  = \new_[11538]_  & \new_[11531]_ ;
  assign \new_[3673]_  = \new_[11524]_  & \new_[11517]_ ;
  assign \new_[3674]_  = \new_[11510]_  & \new_[11503]_ ;
  assign \new_[3675]_  = \new_[11496]_  & \new_[11489]_ ;
  assign \new_[3676]_  = \new_[11482]_  & \new_[11475]_ ;
  assign \new_[3677]_  = \new_[11468]_  & \new_[11461]_ ;
  assign \new_[3678]_  = \new_[11454]_  & \new_[11447]_ ;
  assign \new_[3679]_  = \new_[11440]_  & \new_[11433]_ ;
  assign \new_[3680]_  = \new_[11426]_  & \new_[11419]_ ;
  assign \new_[3681]_  = \new_[11412]_  & \new_[11405]_ ;
  assign \new_[3682]_  = \new_[11398]_  & \new_[11391]_ ;
  assign \new_[3683]_  = \new_[11384]_  & \new_[11377]_ ;
  assign \new_[3684]_  = \new_[11370]_  & \new_[11363]_ ;
  assign \new_[3685]_  = \new_[11356]_  & \new_[11349]_ ;
  assign \new_[3686]_  = \new_[11342]_  & \new_[11335]_ ;
  assign \new_[3687]_  = \new_[11328]_  & \new_[11321]_ ;
  assign \new_[3688]_  = \new_[11314]_  & \new_[11307]_ ;
  assign \new_[3689]_  = \new_[11300]_  & \new_[11293]_ ;
  assign \new_[3690]_  = \new_[11286]_  & \new_[11279]_ ;
  assign \new_[3691]_  = \new_[11272]_  & \new_[11265]_ ;
  assign \new_[3692]_  = \new_[11258]_  & \new_[11251]_ ;
  assign \new_[3693]_  = \new_[11244]_  & \new_[11237]_ ;
  assign \new_[3694]_  = \new_[11230]_  & \new_[11223]_ ;
  assign \new_[3695]_  = \new_[11216]_  & \new_[11209]_ ;
  assign \new_[3696]_  = \new_[11202]_  & \new_[11195]_ ;
  assign \new_[3697]_  = \new_[11188]_  & \new_[11181]_ ;
  assign \new_[3698]_  = \new_[11174]_  & \new_[11167]_ ;
  assign \new_[3699]_  = \new_[11160]_  & \new_[11153]_ ;
  assign \new_[3700]_  = \new_[11146]_  & \new_[11139]_ ;
  assign \new_[3701]_  = \new_[11132]_  & \new_[11125]_ ;
  assign \new_[3702]_  = \new_[11118]_  & \new_[11111]_ ;
  assign \new_[3706]_  = \new_[3700]_  | \new_[3701]_ ;
  assign \new_[3707]_  = \new_[3702]_  | \new_[3706]_ ;
  assign \new_[3710]_  = \new_[3698]_  | \new_[3699]_ ;
  assign \new_[3713]_  = \new_[3696]_  | \new_[3697]_ ;
  assign \new_[3714]_  = \new_[3713]_  | \new_[3710]_ ;
  assign \new_[3715]_  = \new_[3714]_  | \new_[3707]_ ;
  assign \new_[3719]_  = \new_[3693]_  | \new_[3694]_ ;
  assign \new_[3720]_  = \new_[3695]_  | \new_[3719]_ ;
  assign \new_[3723]_  = \new_[3691]_  | \new_[3692]_ ;
  assign \new_[3726]_  = \new_[3689]_  | \new_[3690]_ ;
  assign \new_[3727]_  = \new_[3726]_  | \new_[3723]_ ;
  assign \new_[3728]_  = \new_[3727]_  | \new_[3720]_ ;
  assign \new_[3729]_  = \new_[3728]_  | \new_[3715]_ ;
  assign \new_[3733]_  = \new_[3686]_  | \new_[3687]_ ;
  assign \new_[3734]_  = \new_[3688]_  | \new_[3733]_ ;
  assign \new_[3737]_  = \new_[3684]_  | \new_[3685]_ ;
  assign \new_[3740]_  = \new_[3682]_  | \new_[3683]_ ;
  assign \new_[3741]_  = \new_[3740]_  | \new_[3737]_ ;
  assign \new_[3742]_  = \new_[3741]_  | \new_[3734]_ ;
  assign \new_[3746]_  = \new_[3679]_  | \new_[3680]_ ;
  assign \new_[3747]_  = \new_[3681]_  | \new_[3746]_ ;
  assign \new_[3750]_  = \new_[3677]_  | \new_[3678]_ ;
  assign \new_[3753]_  = \new_[3675]_  | \new_[3676]_ ;
  assign \new_[3754]_  = \new_[3753]_  | \new_[3750]_ ;
  assign \new_[3755]_  = \new_[3754]_  | \new_[3747]_ ;
  assign \new_[3756]_  = \new_[3755]_  | \new_[3742]_ ;
  assign \new_[3757]_  = \new_[3756]_  | \new_[3729]_ ;
  assign \new_[3761]_  = \new_[3672]_  | \new_[3673]_ ;
  assign \new_[3762]_  = \new_[3674]_  | \new_[3761]_ ;
  assign \new_[3765]_  = \new_[3670]_  | \new_[3671]_ ;
  assign \new_[3768]_  = \new_[3668]_  | \new_[3669]_ ;
  assign \new_[3769]_  = \new_[3768]_  | \new_[3765]_ ;
  assign \new_[3770]_  = \new_[3769]_  | \new_[3762]_ ;
  assign \new_[3774]_  = \new_[3665]_  | \new_[3666]_ ;
  assign \new_[3775]_  = \new_[3667]_  | \new_[3774]_ ;
  assign \new_[3778]_  = \new_[3663]_  | \new_[3664]_ ;
  assign \new_[3781]_  = \new_[3661]_  | \new_[3662]_ ;
  assign \new_[3782]_  = \new_[3781]_  | \new_[3778]_ ;
  assign \new_[3783]_  = \new_[3782]_  | \new_[3775]_ ;
  assign \new_[3784]_  = \new_[3783]_  | \new_[3770]_ ;
  assign \new_[3788]_  = \new_[3658]_  | \new_[3659]_ ;
  assign \new_[3789]_  = \new_[3660]_  | \new_[3788]_ ;
  assign \new_[3792]_  = \new_[3656]_  | \new_[3657]_ ;
  assign \new_[3795]_  = \new_[3654]_  | \new_[3655]_ ;
  assign \new_[3796]_  = \new_[3795]_  | \new_[3792]_ ;
  assign \new_[3797]_  = \new_[3796]_  | \new_[3789]_ ;
  assign \new_[3800]_  = \new_[3652]_  | \new_[3653]_ ;
  assign \new_[3803]_  = \new_[3650]_  | \new_[3651]_ ;
  assign \new_[3804]_  = \new_[3803]_  | \new_[3800]_ ;
  assign \new_[3807]_  = \new_[3648]_  | \new_[3649]_ ;
  assign \new_[3810]_  = \new_[3646]_  | \new_[3647]_ ;
  assign \new_[3811]_  = \new_[3810]_  | \new_[3807]_ ;
  assign \new_[3812]_  = \new_[3811]_  | \new_[3804]_ ;
  assign \new_[3813]_  = \new_[3812]_  | \new_[3797]_ ;
  assign \new_[3814]_  = \new_[3813]_  | \new_[3784]_ ;
  assign \new_[3815]_  = \new_[3814]_  | \new_[3757]_ ;
  assign \new_[3819]_  = \new_[3643]_  | \new_[3644]_ ;
  assign \new_[3820]_  = \new_[3645]_  | \new_[3819]_ ;
  assign \new_[3823]_  = \new_[3641]_  | \new_[3642]_ ;
  assign \new_[3826]_  = \new_[3639]_  | \new_[3640]_ ;
  assign \new_[3827]_  = \new_[3826]_  | \new_[3823]_ ;
  assign \new_[3828]_  = \new_[3827]_  | \new_[3820]_ ;
  assign \new_[3832]_  = \new_[3636]_  | \new_[3637]_ ;
  assign \new_[3833]_  = \new_[3638]_  | \new_[3832]_ ;
  assign \new_[3836]_  = \new_[3634]_  | \new_[3635]_ ;
  assign \new_[3839]_  = \new_[3632]_  | \new_[3633]_ ;
  assign \new_[3840]_  = \new_[3839]_  | \new_[3836]_ ;
  assign \new_[3841]_  = \new_[3840]_  | \new_[3833]_ ;
  assign \new_[3842]_  = \new_[3841]_  | \new_[3828]_ ;
  assign \new_[3846]_  = \new_[3629]_  | \new_[3630]_ ;
  assign \new_[3847]_  = \new_[3631]_  | \new_[3846]_ ;
  assign \new_[3850]_  = \new_[3627]_  | \new_[3628]_ ;
  assign \new_[3853]_  = \new_[3625]_  | \new_[3626]_ ;
  assign \new_[3854]_  = \new_[3853]_  | \new_[3850]_ ;
  assign \new_[3855]_  = \new_[3854]_  | \new_[3847]_ ;
  assign \new_[3858]_  = \new_[3623]_  | \new_[3624]_ ;
  assign \new_[3861]_  = \new_[3621]_  | \new_[3622]_ ;
  assign \new_[3862]_  = \new_[3861]_  | \new_[3858]_ ;
  assign \new_[3865]_  = \new_[3619]_  | \new_[3620]_ ;
  assign \new_[3868]_  = \new_[3617]_  | \new_[3618]_ ;
  assign \new_[3869]_  = \new_[3868]_  | \new_[3865]_ ;
  assign \new_[3870]_  = \new_[3869]_  | \new_[3862]_ ;
  assign \new_[3871]_  = \new_[3870]_  | \new_[3855]_ ;
  assign \new_[3872]_  = \new_[3871]_  | \new_[3842]_ ;
  assign \new_[3876]_  = \new_[3614]_  | \new_[3615]_ ;
  assign \new_[3877]_  = \new_[3616]_  | \new_[3876]_ ;
  assign \new_[3880]_  = \new_[3612]_  | \new_[3613]_ ;
  assign \new_[3883]_  = \new_[3610]_  | \new_[3611]_ ;
  assign \new_[3884]_  = \new_[3883]_  | \new_[3880]_ ;
  assign \new_[3885]_  = \new_[3884]_  | \new_[3877]_ ;
  assign \new_[3889]_  = \new_[3607]_  | \new_[3608]_ ;
  assign \new_[3890]_  = \new_[3609]_  | \new_[3889]_ ;
  assign \new_[3893]_  = \new_[3605]_  | \new_[3606]_ ;
  assign \new_[3896]_  = \new_[3603]_  | \new_[3604]_ ;
  assign \new_[3897]_  = \new_[3896]_  | \new_[3893]_ ;
  assign \new_[3898]_  = \new_[3897]_  | \new_[3890]_ ;
  assign \new_[3899]_  = \new_[3898]_  | \new_[3885]_ ;
  assign \new_[3903]_  = \new_[3600]_  | \new_[3601]_ ;
  assign \new_[3904]_  = \new_[3602]_  | \new_[3903]_ ;
  assign \new_[3907]_  = \new_[3598]_  | \new_[3599]_ ;
  assign \new_[3910]_  = \new_[3596]_  | \new_[3597]_ ;
  assign \new_[3911]_  = \new_[3910]_  | \new_[3907]_ ;
  assign \new_[3912]_  = \new_[3911]_  | \new_[3904]_ ;
  assign \new_[3915]_  = \new_[3594]_  | \new_[3595]_ ;
  assign \new_[3918]_  = \new_[3592]_  | \new_[3593]_ ;
  assign \new_[3919]_  = \new_[3918]_  | \new_[3915]_ ;
  assign \new_[3922]_  = \new_[3590]_  | \new_[3591]_ ;
  assign \new_[3925]_  = \new_[3588]_  | \new_[3589]_ ;
  assign \new_[3926]_  = \new_[3925]_  | \new_[3922]_ ;
  assign \new_[3927]_  = \new_[3926]_  | \new_[3919]_ ;
  assign \new_[3928]_  = \new_[3927]_  | \new_[3912]_ ;
  assign \new_[3929]_  = \new_[3928]_  | \new_[3899]_ ;
  assign \new_[3930]_  = \new_[3929]_  | \new_[3872]_ ;
  assign \new_[3931]_  = \new_[3930]_  | \new_[3815]_ ;
  assign \new_[3935]_  = \new_[3585]_  | \new_[3586]_ ;
  assign \new_[3936]_  = \new_[3587]_  | \new_[3935]_ ;
  assign \new_[3939]_  = \new_[3583]_  | \new_[3584]_ ;
  assign \new_[3942]_  = \new_[3581]_  | \new_[3582]_ ;
  assign \new_[3943]_  = \new_[3942]_  | \new_[3939]_ ;
  assign \new_[3944]_  = \new_[3943]_  | \new_[3936]_ ;
  assign \new_[3948]_  = \new_[3578]_  | \new_[3579]_ ;
  assign \new_[3949]_  = \new_[3580]_  | \new_[3948]_ ;
  assign \new_[3952]_  = \new_[3576]_  | \new_[3577]_ ;
  assign \new_[3955]_  = \new_[3574]_  | \new_[3575]_ ;
  assign \new_[3956]_  = \new_[3955]_  | \new_[3952]_ ;
  assign \new_[3957]_  = \new_[3956]_  | \new_[3949]_ ;
  assign \new_[3958]_  = \new_[3957]_  | \new_[3944]_ ;
  assign \new_[3962]_  = \new_[3571]_  | \new_[3572]_ ;
  assign \new_[3963]_  = \new_[3573]_  | \new_[3962]_ ;
  assign \new_[3966]_  = \new_[3569]_  | \new_[3570]_ ;
  assign \new_[3969]_  = \new_[3567]_  | \new_[3568]_ ;
  assign \new_[3970]_  = \new_[3969]_  | \new_[3966]_ ;
  assign \new_[3971]_  = \new_[3970]_  | \new_[3963]_ ;
  assign \new_[3974]_  = \new_[3565]_  | \new_[3566]_ ;
  assign \new_[3977]_  = \new_[3563]_  | \new_[3564]_ ;
  assign \new_[3978]_  = \new_[3977]_  | \new_[3974]_ ;
  assign \new_[3981]_  = \new_[3561]_  | \new_[3562]_ ;
  assign \new_[3984]_  = \new_[3559]_  | \new_[3560]_ ;
  assign \new_[3985]_  = \new_[3984]_  | \new_[3981]_ ;
  assign \new_[3986]_  = \new_[3985]_  | \new_[3978]_ ;
  assign \new_[3987]_  = \new_[3986]_  | \new_[3971]_ ;
  assign \new_[3988]_  = \new_[3987]_  | \new_[3958]_ ;
  assign \new_[3992]_  = \new_[3556]_  | \new_[3557]_ ;
  assign \new_[3993]_  = \new_[3558]_  | \new_[3992]_ ;
  assign \new_[3996]_  = \new_[3554]_  | \new_[3555]_ ;
  assign \new_[3999]_  = \new_[3552]_  | \new_[3553]_ ;
  assign \new_[4000]_  = \new_[3999]_  | \new_[3996]_ ;
  assign \new_[4001]_  = \new_[4000]_  | \new_[3993]_ ;
  assign \new_[4005]_  = \new_[3549]_  | \new_[3550]_ ;
  assign \new_[4006]_  = \new_[3551]_  | \new_[4005]_ ;
  assign \new_[4009]_  = \new_[3547]_  | \new_[3548]_ ;
  assign \new_[4012]_  = \new_[3545]_  | \new_[3546]_ ;
  assign \new_[4013]_  = \new_[4012]_  | \new_[4009]_ ;
  assign \new_[4014]_  = \new_[4013]_  | \new_[4006]_ ;
  assign \new_[4015]_  = \new_[4014]_  | \new_[4001]_ ;
  assign \new_[4019]_  = \new_[3542]_  | \new_[3543]_ ;
  assign \new_[4020]_  = \new_[3544]_  | \new_[4019]_ ;
  assign \new_[4023]_  = \new_[3540]_  | \new_[3541]_ ;
  assign \new_[4026]_  = \new_[3538]_  | \new_[3539]_ ;
  assign \new_[4027]_  = \new_[4026]_  | \new_[4023]_ ;
  assign \new_[4028]_  = \new_[4027]_  | \new_[4020]_ ;
  assign \new_[4031]_  = \new_[3536]_  | \new_[3537]_ ;
  assign \new_[4034]_  = \new_[3534]_  | \new_[3535]_ ;
  assign \new_[4035]_  = \new_[4034]_  | \new_[4031]_ ;
  assign \new_[4038]_  = \new_[3532]_  | \new_[3533]_ ;
  assign \new_[4041]_  = \new_[3530]_  | \new_[3531]_ ;
  assign \new_[4042]_  = \new_[4041]_  | \new_[4038]_ ;
  assign \new_[4043]_  = \new_[4042]_  | \new_[4035]_ ;
  assign \new_[4044]_  = \new_[4043]_  | \new_[4028]_ ;
  assign \new_[4045]_  = \new_[4044]_  | \new_[4015]_ ;
  assign \new_[4046]_  = \new_[4045]_  | \new_[3988]_ ;
  assign \new_[4050]_  = \new_[3527]_  | \new_[3528]_ ;
  assign \new_[4051]_  = \new_[3529]_  | \new_[4050]_ ;
  assign \new_[4054]_  = \new_[3525]_  | \new_[3526]_ ;
  assign \new_[4057]_  = \new_[3523]_  | \new_[3524]_ ;
  assign \new_[4058]_  = \new_[4057]_  | \new_[4054]_ ;
  assign \new_[4059]_  = \new_[4058]_  | \new_[4051]_ ;
  assign \new_[4063]_  = \new_[3520]_  | \new_[3521]_ ;
  assign \new_[4064]_  = \new_[3522]_  | \new_[4063]_ ;
  assign \new_[4067]_  = \new_[3518]_  | \new_[3519]_ ;
  assign \new_[4070]_  = \new_[3516]_  | \new_[3517]_ ;
  assign \new_[4071]_  = \new_[4070]_  | \new_[4067]_ ;
  assign \new_[4072]_  = \new_[4071]_  | \new_[4064]_ ;
  assign \new_[4073]_  = \new_[4072]_  | \new_[4059]_ ;
  assign \new_[4077]_  = \new_[3513]_  | \new_[3514]_ ;
  assign \new_[4078]_  = \new_[3515]_  | \new_[4077]_ ;
  assign \new_[4081]_  = \new_[3511]_  | \new_[3512]_ ;
  assign \new_[4084]_  = \new_[3509]_  | \new_[3510]_ ;
  assign \new_[4085]_  = \new_[4084]_  | \new_[4081]_ ;
  assign \new_[4086]_  = \new_[4085]_  | \new_[4078]_ ;
  assign \new_[4089]_  = \new_[3507]_  | \new_[3508]_ ;
  assign \new_[4092]_  = \new_[3505]_  | \new_[3506]_ ;
  assign \new_[4093]_  = \new_[4092]_  | \new_[4089]_ ;
  assign \new_[4096]_  = \new_[3503]_  | \new_[3504]_ ;
  assign \new_[4099]_  = \new_[3501]_  | \new_[3502]_ ;
  assign \new_[4100]_  = \new_[4099]_  | \new_[4096]_ ;
  assign \new_[4101]_  = \new_[4100]_  | \new_[4093]_ ;
  assign \new_[4102]_  = \new_[4101]_  | \new_[4086]_ ;
  assign \new_[4103]_  = \new_[4102]_  | \new_[4073]_ ;
  assign \new_[4107]_  = \new_[3498]_  | \new_[3499]_ ;
  assign \new_[4108]_  = \new_[3500]_  | \new_[4107]_ ;
  assign \new_[4111]_  = \new_[3496]_  | \new_[3497]_ ;
  assign \new_[4114]_  = \new_[3494]_  | \new_[3495]_ ;
  assign \new_[4115]_  = \new_[4114]_  | \new_[4111]_ ;
  assign \new_[4116]_  = \new_[4115]_  | \new_[4108]_ ;
  assign \new_[4120]_  = \new_[3491]_  | \new_[3492]_ ;
  assign \new_[4121]_  = \new_[3493]_  | \new_[4120]_ ;
  assign \new_[4124]_  = \new_[3489]_  | \new_[3490]_ ;
  assign \new_[4127]_  = \new_[3487]_  | \new_[3488]_ ;
  assign \new_[4128]_  = \new_[4127]_  | \new_[4124]_ ;
  assign \new_[4129]_  = \new_[4128]_  | \new_[4121]_ ;
  assign \new_[4130]_  = \new_[4129]_  | \new_[4116]_ ;
  assign \new_[4134]_  = \new_[3484]_  | \new_[3485]_ ;
  assign \new_[4135]_  = \new_[3486]_  | \new_[4134]_ ;
  assign \new_[4138]_  = \new_[3482]_  | \new_[3483]_ ;
  assign \new_[4141]_  = \new_[3480]_  | \new_[3481]_ ;
  assign \new_[4142]_  = \new_[4141]_  | \new_[4138]_ ;
  assign \new_[4143]_  = \new_[4142]_  | \new_[4135]_ ;
  assign \new_[4146]_  = \new_[3478]_  | \new_[3479]_ ;
  assign \new_[4149]_  = \new_[3476]_  | \new_[3477]_ ;
  assign \new_[4150]_  = \new_[4149]_  | \new_[4146]_ ;
  assign \new_[4153]_  = \new_[3474]_  | \new_[3475]_ ;
  assign \new_[4156]_  = \new_[3472]_  | \new_[3473]_ ;
  assign \new_[4157]_  = \new_[4156]_  | \new_[4153]_ ;
  assign \new_[4158]_  = \new_[4157]_  | \new_[4150]_ ;
  assign \new_[4159]_  = \new_[4158]_  | \new_[4143]_ ;
  assign \new_[4160]_  = \new_[4159]_  | \new_[4130]_ ;
  assign \new_[4161]_  = \new_[4160]_  | \new_[4103]_ ;
  assign \new_[4162]_  = \new_[4161]_  | \new_[4046]_ ;
  assign \new_[4163]_  = \new_[4162]_  | \new_[3931]_ ;
  assign \new_[4167]_  = \new_[3469]_  | \new_[3470]_ ;
  assign \new_[4168]_  = \new_[3471]_  | \new_[4167]_ ;
  assign \new_[4171]_  = \new_[3467]_  | \new_[3468]_ ;
  assign \new_[4174]_  = \new_[3465]_  | \new_[3466]_ ;
  assign \new_[4175]_  = \new_[4174]_  | \new_[4171]_ ;
  assign \new_[4176]_  = \new_[4175]_  | \new_[4168]_ ;
  assign \new_[4180]_  = \new_[3462]_  | \new_[3463]_ ;
  assign \new_[4181]_  = \new_[3464]_  | \new_[4180]_ ;
  assign \new_[4184]_  = \new_[3460]_  | \new_[3461]_ ;
  assign \new_[4187]_  = \new_[3458]_  | \new_[3459]_ ;
  assign \new_[4188]_  = \new_[4187]_  | \new_[4184]_ ;
  assign \new_[4189]_  = \new_[4188]_  | \new_[4181]_ ;
  assign \new_[4190]_  = \new_[4189]_  | \new_[4176]_ ;
  assign \new_[4194]_  = \new_[3455]_  | \new_[3456]_ ;
  assign \new_[4195]_  = \new_[3457]_  | \new_[4194]_ ;
  assign \new_[4198]_  = \new_[3453]_  | \new_[3454]_ ;
  assign \new_[4201]_  = \new_[3451]_  | \new_[3452]_ ;
  assign \new_[4202]_  = \new_[4201]_  | \new_[4198]_ ;
  assign \new_[4203]_  = \new_[4202]_  | \new_[4195]_ ;
  assign \new_[4207]_  = \new_[3448]_  | \new_[3449]_ ;
  assign \new_[4208]_  = \new_[3450]_  | \new_[4207]_ ;
  assign \new_[4211]_  = \new_[3446]_  | \new_[3447]_ ;
  assign \new_[4214]_  = \new_[3444]_  | \new_[3445]_ ;
  assign \new_[4215]_  = \new_[4214]_  | \new_[4211]_ ;
  assign \new_[4216]_  = \new_[4215]_  | \new_[4208]_ ;
  assign \new_[4217]_  = \new_[4216]_  | \new_[4203]_ ;
  assign \new_[4218]_  = \new_[4217]_  | \new_[4190]_ ;
  assign \new_[4222]_  = \new_[3441]_  | \new_[3442]_ ;
  assign \new_[4223]_  = \new_[3443]_  | \new_[4222]_ ;
  assign \new_[4226]_  = \new_[3439]_  | \new_[3440]_ ;
  assign \new_[4229]_  = \new_[3437]_  | \new_[3438]_ ;
  assign \new_[4230]_  = \new_[4229]_  | \new_[4226]_ ;
  assign \new_[4231]_  = \new_[4230]_  | \new_[4223]_ ;
  assign \new_[4235]_  = \new_[3434]_  | \new_[3435]_ ;
  assign \new_[4236]_  = \new_[3436]_  | \new_[4235]_ ;
  assign \new_[4239]_  = \new_[3432]_  | \new_[3433]_ ;
  assign \new_[4242]_  = \new_[3430]_  | \new_[3431]_ ;
  assign \new_[4243]_  = \new_[4242]_  | \new_[4239]_ ;
  assign \new_[4244]_  = \new_[4243]_  | \new_[4236]_ ;
  assign \new_[4245]_  = \new_[4244]_  | \new_[4231]_ ;
  assign \new_[4249]_  = \new_[3427]_  | \new_[3428]_ ;
  assign \new_[4250]_  = \new_[3429]_  | \new_[4249]_ ;
  assign \new_[4253]_  = \new_[3425]_  | \new_[3426]_ ;
  assign \new_[4256]_  = \new_[3423]_  | \new_[3424]_ ;
  assign \new_[4257]_  = \new_[4256]_  | \new_[4253]_ ;
  assign \new_[4258]_  = \new_[4257]_  | \new_[4250]_ ;
  assign \new_[4261]_  = \new_[3421]_  | \new_[3422]_ ;
  assign \new_[4264]_  = \new_[3419]_  | \new_[3420]_ ;
  assign \new_[4265]_  = \new_[4264]_  | \new_[4261]_ ;
  assign \new_[4268]_  = \new_[3417]_  | \new_[3418]_ ;
  assign \new_[4271]_  = \new_[3415]_  | \new_[3416]_ ;
  assign \new_[4272]_  = \new_[4271]_  | \new_[4268]_ ;
  assign \new_[4273]_  = \new_[4272]_  | \new_[4265]_ ;
  assign \new_[4274]_  = \new_[4273]_  | \new_[4258]_ ;
  assign \new_[4275]_  = \new_[4274]_  | \new_[4245]_ ;
  assign \new_[4276]_  = \new_[4275]_  | \new_[4218]_ ;
  assign \new_[4280]_  = \new_[3412]_  | \new_[3413]_ ;
  assign \new_[4281]_  = \new_[3414]_  | \new_[4280]_ ;
  assign \new_[4284]_  = \new_[3410]_  | \new_[3411]_ ;
  assign \new_[4287]_  = \new_[3408]_  | \new_[3409]_ ;
  assign \new_[4288]_  = \new_[4287]_  | \new_[4284]_ ;
  assign \new_[4289]_  = \new_[4288]_  | \new_[4281]_ ;
  assign \new_[4293]_  = \new_[3405]_  | \new_[3406]_ ;
  assign \new_[4294]_  = \new_[3407]_  | \new_[4293]_ ;
  assign \new_[4297]_  = \new_[3403]_  | \new_[3404]_ ;
  assign \new_[4300]_  = \new_[3401]_  | \new_[3402]_ ;
  assign \new_[4301]_  = \new_[4300]_  | \new_[4297]_ ;
  assign \new_[4302]_  = \new_[4301]_  | \new_[4294]_ ;
  assign \new_[4303]_  = \new_[4302]_  | \new_[4289]_ ;
  assign \new_[4307]_  = \new_[3398]_  | \new_[3399]_ ;
  assign \new_[4308]_  = \new_[3400]_  | \new_[4307]_ ;
  assign \new_[4311]_  = \new_[3396]_  | \new_[3397]_ ;
  assign \new_[4314]_  = \new_[3394]_  | \new_[3395]_ ;
  assign \new_[4315]_  = \new_[4314]_  | \new_[4311]_ ;
  assign \new_[4316]_  = \new_[4315]_  | \new_[4308]_ ;
  assign \new_[4319]_  = \new_[3392]_  | \new_[3393]_ ;
  assign \new_[4322]_  = \new_[3390]_  | \new_[3391]_ ;
  assign \new_[4323]_  = \new_[4322]_  | \new_[4319]_ ;
  assign \new_[4326]_  = \new_[3388]_  | \new_[3389]_ ;
  assign \new_[4329]_  = \new_[3386]_  | \new_[3387]_ ;
  assign \new_[4330]_  = \new_[4329]_  | \new_[4326]_ ;
  assign \new_[4331]_  = \new_[4330]_  | \new_[4323]_ ;
  assign \new_[4332]_  = \new_[4331]_  | \new_[4316]_ ;
  assign \new_[4333]_  = \new_[4332]_  | \new_[4303]_ ;
  assign \new_[4337]_  = \new_[3383]_  | \new_[3384]_ ;
  assign \new_[4338]_  = \new_[3385]_  | \new_[4337]_ ;
  assign \new_[4341]_  = \new_[3381]_  | \new_[3382]_ ;
  assign \new_[4344]_  = \new_[3379]_  | \new_[3380]_ ;
  assign \new_[4345]_  = \new_[4344]_  | \new_[4341]_ ;
  assign \new_[4346]_  = \new_[4345]_  | \new_[4338]_ ;
  assign \new_[4350]_  = \new_[3376]_  | \new_[3377]_ ;
  assign \new_[4351]_  = \new_[3378]_  | \new_[4350]_ ;
  assign \new_[4354]_  = \new_[3374]_  | \new_[3375]_ ;
  assign \new_[4357]_  = \new_[3372]_  | \new_[3373]_ ;
  assign \new_[4358]_  = \new_[4357]_  | \new_[4354]_ ;
  assign \new_[4359]_  = \new_[4358]_  | \new_[4351]_ ;
  assign \new_[4360]_  = \new_[4359]_  | \new_[4346]_ ;
  assign \new_[4364]_  = \new_[3369]_  | \new_[3370]_ ;
  assign \new_[4365]_  = \new_[3371]_  | \new_[4364]_ ;
  assign \new_[4368]_  = \new_[3367]_  | \new_[3368]_ ;
  assign \new_[4371]_  = \new_[3365]_  | \new_[3366]_ ;
  assign \new_[4372]_  = \new_[4371]_  | \new_[4368]_ ;
  assign \new_[4373]_  = \new_[4372]_  | \new_[4365]_ ;
  assign \new_[4376]_  = \new_[3363]_  | \new_[3364]_ ;
  assign \new_[4379]_  = \new_[3361]_  | \new_[3362]_ ;
  assign \new_[4380]_  = \new_[4379]_  | \new_[4376]_ ;
  assign \new_[4383]_  = \new_[3359]_  | \new_[3360]_ ;
  assign \new_[4386]_  = \new_[3357]_  | \new_[3358]_ ;
  assign \new_[4387]_  = \new_[4386]_  | \new_[4383]_ ;
  assign \new_[4388]_  = \new_[4387]_  | \new_[4380]_ ;
  assign \new_[4389]_  = \new_[4388]_  | \new_[4373]_ ;
  assign \new_[4390]_  = \new_[4389]_  | \new_[4360]_ ;
  assign \new_[4391]_  = \new_[4390]_  | \new_[4333]_ ;
  assign \new_[4392]_  = \new_[4391]_  | \new_[4276]_ ;
  assign \new_[4396]_  = \new_[3354]_  | \new_[3355]_ ;
  assign \new_[4397]_  = \new_[3356]_  | \new_[4396]_ ;
  assign \new_[4400]_  = \new_[3352]_  | \new_[3353]_ ;
  assign \new_[4403]_  = \new_[3350]_  | \new_[3351]_ ;
  assign \new_[4404]_  = \new_[4403]_  | \new_[4400]_ ;
  assign \new_[4405]_  = \new_[4404]_  | \new_[4397]_ ;
  assign \new_[4409]_  = \new_[3347]_  | \new_[3348]_ ;
  assign \new_[4410]_  = \new_[3349]_  | \new_[4409]_ ;
  assign \new_[4413]_  = \new_[3345]_  | \new_[3346]_ ;
  assign \new_[4416]_  = \new_[3343]_  | \new_[3344]_ ;
  assign \new_[4417]_  = \new_[4416]_  | \new_[4413]_ ;
  assign \new_[4418]_  = \new_[4417]_  | \new_[4410]_ ;
  assign \new_[4419]_  = \new_[4418]_  | \new_[4405]_ ;
  assign \new_[4423]_  = \new_[3340]_  | \new_[3341]_ ;
  assign \new_[4424]_  = \new_[3342]_  | \new_[4423]_ ;
  assign \new_[4427]_  = \new_[3338]_  | \new_[3339]_ ;
  assign \new_[4430]_  = \new_[3336]_  | \new_[3337]_ ;
  assign \new_[4431]_  = \new_[4430]_  | \new_[4427]_ ;
  assign \new_[4432]_  = \new_[4431]_  | \new_[4424]_ ;
  assign \new_[4435]_  = \new_[3334]_  | \new_[3335]_ ;
  assign \new_[4438]_  = \new_[3332]_  | \new_[3333]_ ;
  assign \new_[4439]_  = \new_[4438]_  | \new_[4435]_ ;
  assign \new_[4442]_  = \new_[3330]_  | \new_[3331]_ ;
  assign \new_[4445]_  = \new_[3328]_  | \new_[3329]_ ;
  assign \new_[4446]_  = \new_[4445]_  | \new_[4442]_ ;
  assign \new_[4447]_  = \new_[4446]_  | \new_[4439]_ ;
  assign \new_[4448]_  = \new_[4447]_  | \new_[4432]_ ;
  assign \new_[4449]_  = \new_[4448]_  | \new_[4419]_ ;
  assign \new_[4453]_  = \new_[3325]_  | \new_[3326]_ ;
  assign \new_[4454]_  = \new_[3327]_  | \new_[4453]_ ;
  assign \new_[4457]_  = \new_[3323]_  | \new_[3324]_ ;
  assign \new_[4460]_  = \new_[3321]_  | \new_[3322]_ ;
  assign \new_[4461]_  = \new_[4460]_  | \new_[4457]_ ;
  assign \new_[4462]_  = \new_[4461]_  | \new_[4454]_ ;
  assign \new_[4466]_  = \new_[3318]_  | \new_[3319]_ ;
  assign \new_[4467]_  = \new_[3320]_  | \new_[4466]_ ;
  assign \new_[4470]_  = \new_[3316]_  | \new_[3317]_ ;
  assign \new_[4473]_  = \new_[3314]_  | \new_[3315]_ ;
  assign \new_[4474]_  = \new_[4473]_  | \new_[4470]_ ;
  assign \new_[4475]_  = \new_[4474]_  | \new_[4467]_ ;
  assign \new_[4476]_  = \new_[4475]_  | \new_[4462]_ ;
  assign \new_[4480]_  = \new_[3311]_  | \new_[3312]_ ;
  assign \new_[4481]_  = \new_[3313]_  | \new_[4480]_ ;
  assign \new_[4484]_  = \new_[3309]_  | \new_[3310]_ ;
  assign \new_[4487]_  = \new_[3307]_  | \new_[3308]_ ;
  assign \new_[4488]_  = \new_[4487]_  | \new_[4484]_ ;
  assign \new_[4489]_  = \new_[4488]_  | \new_[4481]_ ;
  assign \new_[4492]_  = \new_[3305]_  | \new_[3306]_ ;
  assign \new_[4495]_  = \new_[3303]_  | \new_[3304]_ ;
  assign \new_[4496]_  = \new_[4495]_  | \new_[4492]_ ;
  assign \new_[4499]_  = \new_[3301]_  | \new_[3302]_ ;
  assign \new_[4502]_  = \new_[3299]_  | \new_[3300]_ ;
  assign \new_[4503]_  = \new_[4502]_  | \new_[4499]_ ;
  assign \new_[4504]_  = \new_[4503]_  | \new_[4496]_ ;
  assign \new_[4505]_  = \new_[4504]_  | \new_[4489]_ ;
  assign \new_[4506]_  = \new_[4505]_  | \new_[4476]_ ;
  assign \new_[4507]_  = \new_[4506]_  | \new_[4449]_ ;
  assign \new_[4511]_  = \new_[3296]_  | \new_[3297]_ ;
  assign \new_[4512]_  = \new_[3298]_  | \new_[4511]_ ;
  assign \new_[4515]_  = \new_[3294]_  | \new_[3295]_ ;
  assign \new_[4518]_  = \new_[3292]_  | \new_[3293]_ ;
  assign \new_[4519]_  = \new_[4518]_  | \new_[4515]_ ;
  assign \new_[4520]_  = \new_[4519]_  | \new_[4512]_ ;
  assign \new_[4524]_  = \new_[3289]_  | \new_[3290]_ ;
  assign \new_[4525]_  = \new_[3291]_  | \new_[4524]_ ;
  assign \new_[4528]_  = \new_[3287]_  | \new_[3288]_ ;
  assign \new_[4531]_  = \new_[3285]_  | \new_[3286]_ ;
  assign \new_[4532]_  = \new_[4531]_  | \new_[4528]_ ;
  assign \new_[4533]_  = \new_[4532]_  | \new_[4525]_ ;
  assign \new_[4534]_  = \new_[4533]_  | \new_[4520]_ ;
  assign \new_[4538]_  = \new_[3282]_  | \new_[3283]_ ;
  assign \new_[4539]_  = \new_[3284]_  | \new_[4538]_ ;
  assign \new_[4542]_  = \new_[3280]_  | \new_[3281]_ ;
  assign \new_[4545]_  = \new_[3278]_  | \new_[3279]_ ;
  assign \new_[4546]_  = \new_[4545]_  | \new_[4542]_ ;
  assign \new_[4547]_  = \new_[4546]_  | \new_[4539]_ ;
  assign \new_[4550]_  = \new_[3276]_  | \new_[3277]_ ;
  assign \new_[4553]_  = \new_[3274]_  | \new_[3275]_ ;
  assign \new_[4554]_  = \new_[4553]_  | \new_[4550]_ ;
  assign \new_[4557]_  = \new_[3272]_  | \new_[3273]_ ;
  assign \new_[4560]_  = \new_[3270]_  | \new_[3271]_ ;
  assign \new_[4561]_  = \new_[4560]_  | \new_[4557]_ ;
  assign \new_[4562]_  = \new_[4561]_  | \new_[4554]_ ;
  assign \new_[4563]_  = \new_[4562]_  | \new_[4547]_ ;
  assign \new_[4564]_  = \new_[4563]_  | \new_[4534]_ ;
  assign \new_[4568]_  = \new_[3267]_  | \new_[3268]_ ;
  assign \new_[4569]_  = \new_[3269]_  | \new_[4568]_ ;
  assign \new_[4572]_  = \new_[3265]_  | \new_[3266]_ ;
  assign \new_[4575]_  = \new_[3263]_  | \new_[3264]_ ;
  assign \new_[4576]_  = \new_[4575]_  | \new_[4572]_ ;
  assign \new_[4577]_  = \new_[4576]_  | \new_[4569]_ ;
  assign \new_[4581]_  = \new_[3260]_  | \new_[3261]_ ;
  assign \new_[4582]_  = \new_[3262]_  | \new_[4581]_ ;
  assign \new_[4585]_  = \new_[3258]_  | \new_[3259]_ ;
  assign \new_[4588]_  = \new_[3256]_  | \new_[3257]_ ;
  assign \new_[4589]_  = \new_[4588]_  | \new_[4585]_ ;
  assign \new_[4590]_  = \new_[4589]_  | \new_[4582]_ ;
  assign \new_[4591]_  = \new_[4590]_  | \new_[4577]_ ;
  assign \new_[4595]_  = \new_[3253]_  | \new_[3254]_ ;
  assign \new_[4596]_  = \new_[3255]_  | \new_[4595]_ ;
  assign \new_[4599]_  = \new_[3251]_  | \new_[3252]_ ;
  assign \new_[4602]_  = \new_[3249]_  | \new_[3250]_ ;
  assign \new_[4603]_  = \new_[4602]_  | \new_[4599]_ ;
  assign \new_[4604]_  = \new_[4603]_  | \new_[4596]_ ;
  assign \new_[4607]_  = \new_[3247]_  | \new_[3248]_ ;
  assign \new_[4610]_  = \new_[3245]_  | \new_[3246]_ ;
  assign \new_[4611]_  = \new_[4610]_  | \new_[4607]_ ;
  assign \new_[4614]_  = \new_[3243]_  | \new_[3244]_ ;
  assign \new_[4617]_  = \new_[3241]_  | \new_[3242]_ ;
  assign \new_[4618]_  = \new_[4617]_  | \new_[4614]_ ;
  assign \new_[4619]_  = \new_[4618]_  | \new_[4611]_ ;
  assign \new_[4620]_  = \new_[4619]_  | \new_[4604]_ ;
  assign \new_[4621]_  = \new_[4620]_  | \new_[4591]_ ;
  assign \new_[4622]_  = \new_[4621]_  | \new_[4564]_ ;
  assign \new_[4623]_  = \new_[4622]_  | \new_[4507]_ ;
  assign \new_[4624]_  = \new_[4623]_  | \new_[4392]_ ;
  assign \new_[4625]_  = \new_[4624]_  | \new_[4163]_ ;
  assign \new_[4629]_  = \new_[3238]_  | \new_[3239]_ ;
  assign \new_[4630]_  = \new_[3240]_  | \new_[4629]_ ;
  assign \new_[4633]_  = \new_[3236]_  | \new_[3237]_ ;
  assign \new_[4636]_  = \new_[3234]_  | \new_[3235]_ ;
  assign \new_[4637]_  = \new_[4636]_  | \new_[4633]_ ;
  assign \new_[4638]_  = \new_[4637]_  | \new_[4630]_ ;
  assign \new_[4642]_  = \new_[3231]_  | \new_[3232]_ ;
  assign \new_[4643]_  = \new_[3233]_  | \new_[4642]_ ;
  assign \new_[4646]_  = \new_[3229]_  | \new_[3230]_ ;
  assign \new_[4649]_  = \new_[3227]_  | \new_[3228]_ ;
  assign \new_[4650]_  = \new_[4649]_  | \new_[4646]_ ;
  assign \new_[4651]_  = \new_[4650]_  | \new_[4643]_ ;
  assign \new_[4652]_  = \new_[4651]_  | \new_[4638]_ ;
  assign \new_[4656]_  = \new_[3224]_  | \new_[3225]_ ;
  assign \new_[4657]_  = \new_[3226]_  | \new_[4656]_ ;
  assign \new_[4660]_  = \new_[3222]_  | \new_[3223]_ ;
  assign \new_[4663]_  = \new_[3220]_  | \new_[3221]_ ;
  assign \new_[4664]_  = \new_[4663]_  | \new_[4660]_ ;
  assign \new_[4665]_  = \new_[4664]_  | \new_[4657]_ ;
  assign \new_[4669]_  = \new_[3217]_  | \new_[3218]_ ;
  assign \new_[4670]_  = \new_[3219]_  | \new_[4669]_ ;
  assign \new_[4673]_  = \new_[3215]_  | \new_[3216]_ ;
  assign \new_[4676]_  = \new_[3213]_  | \new_[3214]_ ;
  assign \new_[4677]_  = \new_[4676]_  | \new_[4673]_ ;
  assign \new_[4678]_  = \new_[4677]_  | \new_[4670]_ ;
  assign \new_[4679]_  = \new_[4678]_  | \new_[4665]_ ;
  assign \new_[4680]_  = \new_[4679]_  | \new_[4652]_ ;
  assign \new_[4684]_  = \new_[3210]_  | \new_[3211]_ ;
  assign \new_[4685]_  = \new_[3212]_  | \new_[4684]_ ;
  assign \new_[4688]_  = \new_[3208]_  | \new_[3209]_ ;
  assign \new_[4691]_  = \new_[3206]_  | \new_[3207]_ ;
  assign \new_[4692]_  = \new_[4691]_  | \new_[4688]_ ;
  assign \new_[4693]_  = \new_[4692]_  | \new_[4685]_ ;
  assign \new_[4697]_  = \new_[3203]_  | \new_[3204]_ ;
  assign \new_[4698]_  = \new_[3205]_  | \new_[4697]_ ;
  assign \new_[4701]_  = \new_[3201]_  | \new_[3202]_ ;
  assign \new_[4704]_  = \new_[3199]_  | \new_[3200]_ ;
  assign \new_[4705]_  = \new_[4704]_  | \new_[4701]_ ;
  assign \new_[4706]_  = \new_[4705]_  | \new_[4698]_ ;
  assign \new_[4707]_  = \new_[4706]_  | \new_[4693]_ ;
  assign \new_[4711]_  = \new_[3196]_  | \new_[3197]_ ;
  assign \new_[4712]_  = \new_[3198]_  | \new_[4711]_ ;
  assign \new_[4715]_  = \new_[3194]_  | \new_[3195]_ ;
  assign \new_[4718]_  = \new_[3192]_  | \new_[3193]_ ;
  assign \new_[4719]_  = \new_[4718]_  | \new_[4715]_ ;
  assign \new_[4720]_  = \new_[4719]_  | \new_[4712]_ ;
  assign \new_[4723]_  = \new_[3190]_  | \new_[3191]_ ;
  assign \new_[4726]_  = \new_[3188]_  | \new_[3189]_ ;
  assign \new_[4727]_  = \new_[4726]_  | \new_[4723]_ ;
  assign \new_[4730]_  = \new_[3186]_  | \new_[3187]_ ;
  assign \new_[4733]_  = \new_[3184]_  | \new_[3185]_ ;
  assign \new_[4734]_  = \new_[4733]_  | \new_[4730]_ ;
  assign \new_[4735]_  = \new_[4734]_  | \new_[4727]_ ;
  assign \new_[4736]_  = \new_[4735]_  | \new_[4720]_ ;
  assign \new_[4737]_  = \new_[4736]_  | \new_[4707]_ ;
  assign \new_[4738]_  = \new_[4737]_  | \new_[4680]_ ;
  assign \new_[4742]_  = \new_[3181]_  | \new_[3182]_ ;
  assign \new_[4743]_  = \new_[3183]_  | \new_[4742]_ ;
  assign \new_[4746]_  = \new_[3179]_  | \new_[3180]_ ;
  assign \new_[4749]_  = \new_[3177]_  | \new_[3178]_ ;
  assign \new_[4750]_  = \new_[4749]_  | \new_[4746]_ ;
  assign \new_[4751]_  = \new_[4750]_  | \new_[4743]_ ;
  assign \new_[4755]_  = \new_[3174]_  | \new_[3175]_ ;
  assign \new_[4756]_  = \new_[3176]_  | \new_[4755]_ ;
  assign \new_[4759]_  = \new_[3172]_  | \new_[3173]_ ;
  assign \new_[4762]_  = \new_[3170]_  | \new_[3171]_ ;
  assign \new_[4763]_  = \new_[4762]_  | \new_[4759]_ ;
  assign \new_[4764]_  = \new_[4763]_  | \new_[4756]_ ;
  assign \new_[4765]_  = \new_[4764]_  | \new_[4751]_ ;
  assign \new_[4769]_  = \new_[3167]_  | \new_[3168]_ ;
  assign \new_[4770]_  = \new_[3169]_  | \new_[4769]_ ;
  assign \new_[4773]_  = \new_[3165]_  | \new_[3166]_ ;
  assign \new_[4776]_  = \new_[3163]_  | \new_[3164]_ ;
  assign \new_[4777]_  = \new_[4776]_  | \new_[4773]_ ;
  assign \new_[4778]_  = \new_[4777]_  | \new_[4770]_ ;
  assign \new_[4781]_  = \new_[3161]_  | \new_[3162]_ ;
  assign \new_[4784]_  = \new_[3159]_  | \new_[3160]_ ;
  assign \new_[4785]_  = \new_[4784]_  | \new_[4781]_ ;
  assign \new_[4788]_  = \new_[3157]_  | \new_[3158]_ ;
  assign \new_[4791]_  = \new_[3155]_  | \new_[3156]_ ;
  assign \new_[4792]_  = \new_[4791]_  | \new_[4788]_ ;
  assign \new_[4793]_  = \new_[4792]_  | \new_[4785]_ ;
  assign \new_[4794]_  = \new_[4793]_  | \new_[4778]_ ;
  assign \new_[4795]_  = \new_[4794]_  | \new_[4765]_ ;
  assign \new_[4799]_  = \new_[3152]_  | \new_[3153]_ ;
  assign \new_[4800]_  = \new_[3154]_  | \new_[4799]_ ;
  assign \new_[4803]_  = \new_[3150]_  | \new_[3151]_ ;
  assign \new_[4806]_  = \new_[3148]_  | \new_[3149]_ ;
  assign \new_[4807]_  = \new_[4806]_  | \new_[4803]_ ;
  assign \new_[4808]_  = \new_[4807]_  | \new_[4800]_ ;
  assign \new_[4812]_  = \new_[3145]_  | \new_[3146]_ ;
  assign \new_[4813]_  = \new_[3147]_  | \new_[4812]_ ;
  assign \new_[4816]_  = \new_[3143]_  | \new_[3144]_ ;
  assign \new_[4819]_  = \new_[3141]_  | \new_[3142]_ ;
  assign \new_[4820]_  = \new_[4819]_  | \new_[4816]_ ;
  assign \new_[4821]_  = \new_[4820]_  | \new_[4813]_ ;
  assign \new_[4822]_  = \new_[4821]_  | \new_[4808]_ ;
  assign \new_[4826]_  = \new_[3138]_  | \new_[3139]_ ;
  assign \new_[4827]_  = \new_[3140]_  | \new_[4826]_ ;
  assign \new_[4830]_  = \new_[3136]_  | \new_[3137]_ ;
  assign \new_[4833]_  = \new_[3134]_  | \new_[3135]_ ;
  assign \new_[4834]_  = \new_[4833]_  | \new_[4830]_ ;
  assign \new_[4835]_  = \new_[4834]_  | \new_[4827]_ ;
  assign \new_[4838]_  = \new_[3132]_  | \new_[3133]_ ;
  assign \new_[4841]_  = \new_[3130]_  | \new_[3131]_ ;
  assign \new_[4842]_  = \new_[4841]_  | \new_[4838]_ ;
  assign \new_[4845]_  = \new_[3128]_  | \new_[3129]_ ;
  assign \new_[4848]_  = \new_[3126]_  | \new_[3127]_ ;
  assign \new_[4849]_  = \new_[4848]_  | \new_[4845]_ ;
  assign \new_[4850]_  = \new_[4849]_  | \new_[4842]_ ;
  assign \new_[4851]_  = \new_[4850]_  | \new_[4835]_ ;
  assign \new_[4852]_  = \new_[4851]_  | \new_[4822]_ ;
  assign \new_[4853]_  = \new_[4852]_  | \new_[4795]_ ;
  assign \new_[4854]_  = \new_[4853]_  | \new_[4738]_ ;
  assign \new_[4858]_  = \new_[3123]_  | \new_[3124]_ ;
  assign \new_[4859]_  = \new_[3125]_  | \new_[4858]_ ;
  assign \new_[4862]_  = \new_[3121]_  | \new_[3122]_ ;
  assign \new_[4865]_  = \new_[3119]_  | \new_[3120]_ ;
  assign \new_[4866]_  = \new_[4865]_  | \new_[4862]_ ;
  assign \new_[4867]_  = \new_[4866]_  | \new_[4859]_ ;
  assign \new_[4871]_  = \new_[3116]_  | \new_[3117]_ ;
  assign \new_[4872]_  = \new_[3118]_  | \new_[4871]_ ;
  assign \new_[4875]_  = \new_[3114]_  | \new_[3115]_ ;
  assign \new_[4878]_  = \new_[3112]_  | \new_[3113]_ ;
  assign \new_[4879]_  = \new_[4878]_  | \new_[4875]_ ;
  assign \new_[4880]_  = \new_[4879]_  | \new_[4872]_ ;
  assign \new_[4881]_  = \new_[4880]_  | \new_[4867]_ ;
  assign \new_[4885]_  = \new_[3109]_  | \new_[3110]_ ;
  assign \new_[4886]_  = \new_[3111]_  | \new_[4885]_ ;
  assign \new_[4889]_  = \new_[3107]_  | \new_[3108]_ ;
  assign \new_[4892]_  = \new_[3105]_  | \new_[3106]_ ;
  assign \new_[4893]_  = \new_[4892]_  | \new_[4889]_ ;
  assign \new_[4894]_  = \new_[4893]_  | \new_[4886]_ ;
  assign \new_[4897]_  = \new_[3103]_  | \new_[3104]_ ;
  assign \new_[4900]_  = \new_[3101]_  | \new_[3102]_ ;
  assign \new_[4901]_  = \new_[4900]_  | \new_[4897]_ ;
  assign \new_[4904]_  = \new_[3099]_  | \new_[3100]_ ;
  assign \new_[4907]_  = \new_[3097]_  | \new_[3098]_ ;
  assign \new_[4908]_  = \new_[4907]_  | \new_[4904]_ ;
  assign \new_[4909]_  = \new_[4908]_  | \new_[4901]_ ;
  assign \new_[4910]_  = \new_[4909]_  | \new_[4894]_ ;
  assign \new_[4911]_  = \new_[4910]_  | \new_[4881]_ ;
  assign \new_[4915]_  = \new_[3094]_  | \new_[3095]_ ;
  assign \new_[4916]_  = \new_[3096]_  | \new_[4915]_ ;
  assign \new_[4919]_  = \new_[3092]_  | \new_[3093]_ ;
  assign \new_[4922]_  = \new_[3090]_  | \new_[3091]_ ;
  assign \new_[4923]_  = \new_[4922]_  | \new_[4919]_ ;
  assign \new_[4924]_  = \new_[4923]_  | \new_[4916]_ ;
  assign \new_[4928]_  = \new_[3087]_  | \new_[3088]_ ;
  assign \new_[4929]_  = \new_[3089]_  | \new_[4928]_ ;
  assign \new_[4932]_  = \new_[3085]_  | \new_[3086]_ ;
  assign \new_[4935]_  = \new_[3083]_  | \new_[3084]_ ;
  assign \new_[4936]_  = \new_[4935]_  | \new_[4932]_ ;
  assign \new_[4937]_  = \new_[4936]_  | \new_[4929]_ ;
  assign \new_[4938]_  = \new_[4937]_  | \new_[4924]_ ;
  assign \new_[4942]_  = \new_[3080]_  | \new_[3081]_ ;
  assign \new_[4943]_  = \new_[3082]_  | \new_[4942]_ ;
  assign \new_[4946]_  = \new_[3078]_  | \new_[3079]_ ;
  assign \new_[4949]_  = \new_[3076]_  | \new_[3077]_ ;
  assign \new_[4950]_  = \new_[4949]_  | \new_[4946]_ ;
  assign \new_[4951]_  = \new_[4950]_  | \new_[4943]_ ;
  assign \new_[4954]_  = \new_[3074]_  | \new_[3075]_ ;
  assign \new_[4957]_  = \new_[3072]_  | \new_[3073]_ ;
  assign \new_[4958]_  = \new_[4957]_  | \new_[4954]_ ;
  assign \new_[4961]_  = \new_[3070]_  | \new_[3071]_ ;
  assign \new_[4964]_  = \new_[3068]_  | \new_[3069]_ ;
  assign \new_[4965]_  = \new_[4964]_  | \new_[4961]_ ;
  assign \new_[4966]_  = \new_[4965]_  | \new_[4958]_ ;
  assign \new_[4967]_  = \new_[4966]_  | \new_[4951]_ ;
  assign \new_[4968]_  = \new_[4967]_  | \new_[4938]_ ;
  assign \new_[4969]_  = \new_[4968]_  | \new_[4911]_ ;
  assign \new_[4973]_  = \new_[3065]_  | \new_[3066]_ ;
  assign \new_[4974]_  = \new_[3067]_  | \new_[4973]_ ;
  assign \new_[4977]_  = \new_[3063]_  | \new_[3064]_ ;
  assign \new_[4980]_  = \new_[3061]_  | \new_[3062]_ ;
  assign \new_[4981]_  = \new_[4980]_  | \new_[4977]_ ;
  assign \new_[4982]_  = \new_[4981]_  | \new_[4974]_ ;
  assign \new_[4986]_  = \new_[3058]_  | \new_[3059]_ ;
  assign \new_[4987]_  = \new_[3060]_  | \new_[4986]_ ;
  assign \new_[4990]_  = \new_[3056]_  | \new_[3057]_ ;
  assign \new_[4993]_  = \new_[3054]_  | \new_[3055]_ ;
  assign \new_[4994]_  = \new_[4993]_  | \new_[4990]_ ;
  assign \new_[4995]_  = \new_[4994]_  | \new_[4987]_ ;
  assign \new_[4996]_  = \new_[4995]_  | \new_[4982]_ ;
  assign \new_[5000]_  = \new_[3051]_  | \new_[3052]_ ;
  assign \new_[5001]_  = \new_[3053]_  | \new_[5000]_ ;
  assign \new_[5004]_  = \new_[3049]_  | \new_[3050]_ ;
  assign \new_[5007]_  = \new_[3047]_  | \new_[3048]_ ;
  assign \new_[5008]_  = \new_[5007]_  | \new_[5004]_ ;
  assign \new_[5009]_  = \new_[5008]_  | \new_[5001]_ ;
  assign \new_[5012]_  = \new_[3045]_  | \new_[3046]_ ;
  assign \new_[5015]_  = \new_[3043]_  | \new_[3044]_ ;
  assign \new_[5016]_  = \new_[5015]_  | \new_[5012]_ ;
  assign \new_[5019]_  = \new_[3041]_  | \new_[3042]_ ;
  assign \new_[5022]_  = \new_[3039]_  | \new_[3040]_ ;
  assign \new_[5023]_  = \new_[5022]_  | \new_[5019]_ ;
  assign \new_[5024]_  = \new_[5023]_  | \new_[5016]_ ;
  assign \new_[5025]_  = \new_[5024]_  | \new_[5009]_ ;
  assign \new_[5026]_  = \new_[5025]_  | \new_[4996]_ ;
  assign \new_[5030]_  = \new_[3036]_  | \new_[3037]_ ;
  assign \new_[5031]_  = \new_[3038]_  | \new_[5030]_ ;
  assign \new_[5034]_  = \new_[3034]_  | \new_[3035]_ ;
  assign \new_[5037]_  = \new_[3032]_  | \new_[3033]_ ;
  assign \new_[5038]_  = \new_[5037]_  | \new_[5034]_ ;
  assign \new_[5039]_  = \new_[5038]_  | \new_[5031]_ ;
  assign \new_[5043]_  = \new_[3029]_  | \new_[3030]_ ;
  assign \new_[5044]_  = \new_[3031]_  | \new_[5043]_ ;
  assign \new_[5047]_  = \new_[3027]_  | \new_[3028]_ ;
  assign \new_[5050]_  = \new_[3025]_  | \new_[3026]_ ;
  assign \new_[5051]_  = \new_[5050]_  | \new_[5047]_ ;
  assign \new_[5052]_  = \new_[5051]_  | \new_[5044]_ ;
  assign \new_[5053]_  = \new_[5052]_  | \new_[5039]_ ;
  assign \new_[5057]_  = \new_[3022]_  | \new_[3023]_ ;
  assign \new_[5058]_  = \new_[3024]_  | \new_[5057]_ ;
  assign \new_[5061]_  = \new_[3020]_  | \new_[3021]_ ;
  assign \new_[5064]_  = \new_[3018]_  | \new_[3019]_ ;
  assign \new_[5065]_  = \new_[5064]_  | \new_[5061]_ ;
  assign \new_[5066]_  = \new_[5065]_  | \new_[5058]_ ;
  assign \new_[5069]_  = \new_[3016]_  | \new_[3017]_ ;
  assign \new_[5072]_  = \new_[3014]_  | \new_[3015]_ ;
  assign \new_[5073]_  = \new_[5072]_  | \new_[5069]_ ;
  assign \new_[5076]_  = \new_[3012]_  | \new_[3013]_ ;
  assign \new_[5079]_  = \new_[3010]_  | \new_[3011]_ ;
  assign \new_[5080]_  = \new_[5079]_  | \new_[5076]_ ;
  assign \new_[5081]_  = \new_[5080]_  | \new_[5073]_ ;
  assign \new_[5082]_  = \new_[5081]_  | \new_[5066]_ ;
  assign \new_[5083]_  = \new_[5082]_  | \new_[5053]_ ;
  assign \new_[5084]_  = \new_[5083]_  | \new_[5026]_ ;
  assign \new_[5085]_  = \new_[5084]_  | \new_[4969]_ ;
  assign \new_[5086]_  = \new_[5085]_  | \new_[4854]_ ;
  assign \new_[5090]_  = \new_[3007]_  | \new_[3008]_ ;
  assign \new_[5091]_  = \new_[3009]_  | \new_[5090]_ ;
  assign \new_[5094]_  = \new_[3005]_  | \new_[3006]_ ;
  assign \new_[5097]_  = \new_[3003]_  | \new_[3004]_ ;
  assign \new_[5098]_  = \new_[5097]_  | \new_[5094]_ ;
  assign \new_[5099]_  = \new_[5098]_  | \new_[5091]_ ;
  assign \new_[5103]_  = \new_[3000]_  | \new_[3001]_ ;
  assign \new_[5104]_  = \new_[3002]_  | \new_[5103]_ ;
  assign \new_[5107]_  = \new_[2998]_  | \new_[2999]_ ;
  assign \new_[5110]_  = \new_[2996]_  | \new_[2997]_ ;
  assign \new_[5111]_  = \new_[5110]_  | \new_[5107]_ ;
  assign \new_[5112]_  = \new_[5111]_  | \new_[5104]_ ;
  assign \new_[5113]_  = \new_[5112]_  | \new_[5099]_ ;
  assign \new_[5117]_  = \new_[2993]_  | \new_[2994]_ ;
  assign \new_[5118]_  = \new_[2995]_  | \new_[5117]_ ;
  assign \new_[5121]_  = \new_[2991]_  | \new_[2992]_ ;
  assign \new_[5124]_  = \new_[2989]_  | \new_[2990]_ ;
  assign \new_[5125]_  = \new_[5124]_  | \new_[5121]_ ;
  assign \new_[5126]_  = \new_[5125]_  | \new_[5118]_ ;
  assign \new_[5129]_  = \new_[2987]_  | \new_[2988]_ ;
  assign \new_[5132]_  = \new_[2985]_  | \new_[2986]_ ;
  assign \new_[5133]_  = \new_[5132]_  | \new_[5129]_ ;
  assign \new_[5136]_  = \new_[2983]_  | \new_[2984]_ ;
  assign \new_[5139]_  = \new_[2981]_  | \new_[2982]_ ;
  assign \new_[5140]_  = \new_[5139]_  | \new_[5136]_ ;
  assign \new_[5141]_  = \new_[5140]_  | \new_[5133]_ ;
  assign \new_[5142]_  = \new_[5141]_  | \new_[5126]_ ;
  assign \new_[5143]_  = \new_[5142]_  | \new_[5113]_ ;
  assign \new_[5147]_  = \new_[2978]_  | \new_[2979]_ ;
  assign \new_[5148]_  = \new_[2980]_  | \new_[5147]_ ;
  assign \new_[5151]_  = \new_[2976]_  | \new_[2977]_ ;
  assign \new_[5154]_  = \new_[2974]_  | \new_[2975]_ ;
  assign \new_[5155]_  = \new_[5154]_  | \new_[5151]_ ;
  assign \new_[5156]_  = \new_[5155]_  | \new_[5148]_ ;
  assign \new_[5160]_  = \new_[2971]_  | \new_[2972]_ ;
  assign \new_[5161]_  = \new_[2973]_  | \new_[5160]_ ;
  assign \new_[5164]_  = \new_[2969]_  | \new_[2970]_ ;
  assign \new_[5167]_  = \new_[2967]_  | \new_[2968]_ ;
  assign \new_[5168]_  = \new_[5167]_  | \new_[5164]_ ;
  assign \new_[5169]_  = \new_[5168]_  | \new_[5161]_ ;
  assign \new_[5170]_  = \new_[5169]_  | \new_[5156]_ ;
  assign \new_[5174]_  = \new_[2964]_  | \new_[2965]_ ;
  assign \new_[5175]_  = \new_[2966]_  | \new_[5174]_ ;
  assign \new_[5178]_  = \new_[2962]_  | \new_[2963]_ ;
  assign \new_[5181]_  = \new_[2960]_  | \new_[2961]_ ;
  assign \new_[5182]_  = \new_[5181]_  | \new_[5178]_ ;
  assign \new_[5183]_  = \new_[5182]_  | \new_[5175]_ ;
  assign \new_[5186]_  = \new_[2958]_  | \new_[2959]_ ;
  assign \new_[5189]_  = \new_[2956]_  | \new_[2957]_ ;
  assign \new_[5190]_  = \new_[5189]_  | \new_[5186]_ ;
  assign \new_[5193]_  = \new_[2954]_  | \new_[2955]_ ;
  assign \new_[5196]_  = \new_[2952]_  | \new_[2953]_ ;
  assign \new_[5197]_  = \new_[5196]_  | \new_[5193]_ ;
  assign \new_[5198]_  = \new_[5197]_  | \new_[5190]_ ;
  assign \new_[5199]_  = \new_[5198]_  | \new_[5183]_ ;
  assign \new_[5200]_  = \new_[5199]_  | \new_[5170]_ ;
  assign \new_[5201]_  = \new_[5200]_  | \new_[5143]_ ;
  assign \new_[5205]_  = \new_[2949]_  | \new_[2950]_ ;
  assign \new_[5206]_  = \new_[2951]_  | \new_[5205]_ ;
  assign \new_[5209]_  = \new_[2947]_  | \new_[2948]_ ;
  assign \new_[5212]_  = \new_[2945]_  | \new_[2946]_ ;
  assign \new_[5213]_  = \new_[5212]_  | \new_[5209]_ ;
  assign \new_[5214]_  = \new_[5213]_  | \new_[5206]_ ;
  assign \new_[5218]_  = \new_[2942]_  | \new_[2943]_ ;
  assign \new_[5219]_  = \new_[2944]_  | \new_[5218]_ ;
  assign \new_[5222]_  = \new_[2940]_  | \new_[2941]_ ;
  assign \new_[5225]_  = \new_[2938]_  | \new_[2939]_ ;
  assign \new_[5226]_  = \new_[5225]_  | \new_[5222]_ ;
  assign \new_[5227]_  = \new_[5226]_  | \new_[5219]_ ;
  assign \new_[5228]_  = \new_[5227]_  | \new_[5214]_ ;
  assign \new_[5232]_  = \new_[2935]_  | \new_[2936]_ ;
  assign \new_[5233]_  = \new_[2937]_  | \new_[5232]_ ;
  assign \new_[5236]_  = \new_[2933]_  | \new_[2934]_ ;
  assign \new_[5239]_  = \new_[2931]_  | \new_[2932]_ ;
  assign \new_[5240]_  = \new_[5239]_  | \new_[5236]_ ;
  assign \new_[5241]_  = \new_[5240]_  | \new_[5233]_ ;
  assign \new_[5244]_  = \new_[2929]_  | \new_[2930]_ ;
  assign \new_[5247]_  = \new_[2927]_  | \new_[2928]_ ;
  assign \new_[5248]_  = \new_[5247]_  | \new_[5244]_ ;
  assign \new_[5251]_  = \new_[2925]_  | \new_[2926]_ ;
  assign \new_[5254]_  = \new_[2923]_  | \new_[2924]_ ;
  assign \new_[5255]_  = \new_[5254]_  | \new_[5251]_ ;
  assign \new_[5256]_  = \new_[5255]_  | \new_[5248]_ ;
  assign \new_[5257]_  = \new_[5256]_  | \new_[5241]_ ;
  assign \new_[5258]_  = \new_[5257]_  | \new_[5228]_ ;
  assign \new_[5262]_  = \new_[2920]_  | \new_[2921]_ ;
  assign \new_[5263]_  = \new_[2922]_  | \new_[5262]_ ;
  assign \new_[5266]_  = \new_[2918]_  | \new_[2919]_ ;
  assign \new_[5269]_  = \new_[2916]_  | \new_[2917]_ ;
  assign \new_[5270]_  = \new_[5269]_  | \new_[5266]_ ;
  assign \new_[5271]_  = \new_[5270]_  | \new_[5263]_ ;
  assign \new_[5275]_  = \new_[2913]_  | \new_[2914]_ ;
  assign \new_[5276]_  = \new_[2915]_  | \new_[5275]_ ;
  assign \new_[5279]_  = \new_[2911]_  | \new_[2912]_ ;
  assign \new_[5282]_  = \new_[2909]_  | \new_[2910]_ ;
  assign \new_[5283]_  = \new_[5282]_  | \new_[5279]_ ;
  assign \new_[5284]_  = \new_[5283]_  | \new_[5276]_ ;
  assign \new_[5285]_  = \new_[5284]_  | \new_[5271]_ ;
  assign \new_[5289]_  = \new_[2906]_  | \new_[2907]_ ;
  assign \new_[5290]_  = \new_[2908]_  | \new_[5289]_ ;
  assign \new_[5293]_  = \new_[2904]_  | \new_[2905]_ ;
  assign \new_[5296]_  = \new_[2902]_  | \new_[2903]_ ;
  assign \new_[5297]_  = \new_[5296]_  | \new_[5293]_ ;
  assign \new_[5298]_  = \new_[5297]_  | \new_[5290]_ ;
  assign \new_[5301]_  = \new_[2900]_  | \new_[2901]_ ;
  assign \new_[5304]_  = \new_[2898]_  | \new_[2899]_ ;
  assign \new_[5305]_  = \new_[5304]_  | \new_[5301]_ ;
  assign \new_[5308]_  = \new_[2896]_  | \new_[2897]_ ;
  assign \new_[5311]_  = \new_[2894]_  | \new_[2895]_ ;
  assign \new_[5312]_  = \new_[5311]_  | \new_[5308]_ ;
  assign \new_[5313]_  = \new_[5312]_  | \new_[5305]_ ;
  assign \new_[5314]_  = \new_[5313]_  | \new_[5298]_ ;
  assign \new_[5315]_  = \new_[5314]_  | \new_[5285]_ ;
  assign \new_[5316]_  = \new_[5315]_  | \new_[5258]_ ;
  assign \new_[5317]_  = \new_[5316]_  | \new_[5201]_ ;
  assign \new_[5321]_  = \new_[2891]_  | \new_[2892]_ ;
  assign \new_[5322]_  = \new_[2893]_  | \new_[5321]_ ;
  assign \new_[5325]_  = \new_[2889]_  | \new_[2890]_ ;
  assign \new_[5328]_  = \new_[2887]_  | \new_[2888]_ ;
  assign \new_[5329]_  = \new_[5328]_  | \new_[5325]_ ;
  assign \new_[5330]_  = \new_[5329]_  | \new_[5322]_ ;
  assign \new_[5334]_  = \new_[2884]_  | \new_[2885]_ ;
  assign \new_[5335]_  = \new_[2886]_  | \new_[5334]_ ;
  assign \new_[5338]_  = \new_[2882]_  | \new_[2883]_ ;
  assign \new_[5341]_  = \new_[2880]_  | \new_[2881]_ ;
  assign \new_[5342]_  = \new_[5341]_  | \new_[5338]_ ;
  assign \new_[5343]_  = \new_[5342]_  | \new_[5335]_ ;
  assign \new_[5344]_  = \new_[5343]_  | \new_[5330]_ ;
  assign \new_[5348]_  = \new_[2877]_  | \new_[2878]_ ;
  assign \new_[5349]_  = \new_[2879]_  | \new_[5348]_ ;
  assign \new_[5352]_  = \new_[2875]_  | \new_[2876]_ ;
  assign \new_[5355]_  = \new_[2873]_  | \new_[2874]_ ;
  assign \new_[5356]_  = \new_[5355]_  | \new_[5352]_ ;
  assign \new_[5357]_  = \new_[5356]_  | \new_[5349]_ ;
  assign \new_[5360]_  = \new_[2871]_  | \new_[2872]_ ;
  assign \new_[5363]_  = \new_[2869]_  | \new_[2870]_ ;
  assign \new_[5364]_  = \new_[5363]_  | \new_[5360]_ ;
  assign \new_[5367]_  = \new_[2867]_  | \new_[2868]_ ;
  assign \new_[5370]_  = \new_[2865]_  | \new_[2866]_ ;
  assign \new_[5371]_  = \new_[5370]_  | \new_[5367]_ ;
  assign \new_[5372]_  = \new_[5371]_  | \new_[5364]_ ;
  assign \new_[5373]_  = \new_[5372]_  | \new_[5357]_ ;
  assign \new_[5374]_  = \new_[5373]_  | \new_[5344]_ ;
  assign \new_[5378]_  = \new_[2862]_  | \new_[2863]_ ;
  assign \new_[5379]_  = \new_[2864]_  | \new_[5378]_ ;
  assign \new_[5382]_  = \new_[2860]_  | \new_[2861]_ ;
  assign \new_[5385]_  = \new_[2858]_  | \new_[2859]_ ;
  assign \new_[5386]_  = \new_[5385]_  | \new_[5382]_ ;
  assign \new_[5387]_  = \new_[5386]_  | \new_[5379]_ ;
  assign \new_[5391]_  = \new_[2855]_  | \new_[2856]_ ;
  assign \new_[5392]_  = \new_[2857]_  | \new_[5391]_ ;
  assign \new_[5395]_  = \new_[2853]_  | \new_[2854]_ ;
  assign \new_[5398]_  = \new_[2851]_  | \new_[2852]_ ;
  assign \new_[5399]_  = \new_[5398]_  | \new_[5395]_ ;
  assign \new_[5400]_  = \new_[5399]_  | \new_[5392]_ ;
  assign \new_[5401]_  = \new_[5400]_  | \new_[5387]_ ;
  assign \new_[5405]_  = \new_[2848]_  | \new_[2849]_ ;
  assign \new_[5406]_  = \new_[2850]_  | \new_[5405]_ ;
  assign \new_[5409]_  = \new_[2846]_  | \new_[2847]_ ;
  assign \new_[5412]_  = \new_[2844]_  | \new_[2845]_ ;
  assign \new_[5413]_  = \new_[5412]_  | \new_[5409]_ ;
  assign \new_[5414]_  = \new_[5413]_  | \new_[5406]_ ;
  assign \new_[5417]_  = \new_[2842]_  | \new_[2843]_ ;
  assign \new_[5420]_  = \new_[2840]_  | \new_[2841]_ ;
  assign \new_[5421]_  = \new_[5420]_  | \new_[5417]_ ;
  assign \new_[5424]_  = \new_[2838]_  | \new_[2839]_ ;
  assign \new_[5427]_  = \new_[2836]_  | \new_[2837]_ ;
  assign \new_[5428]_  = \new_[5427]_  | \new_[5424]_ ;
  assign \new_[5429]_  = \new_[5428]_  | \new_[5421]_ ;
  assign \new_[5430]_  = \new_[5429]_  | \new_[5414]_ ;
  assign \new_[5431]_  = \new_[5430]_  | \new_[5401]_ ;
  assign \new_[5432]_  = \new_[5431]_  | \new_[5374]_ ;
  assign \new_[5436]_  = \new_[2833]_  | \new_[2834]_ ;
  assign \new_[5437]_  = \new_[2835]_  | \new_[5436]_ ;
  assign \new_[5440]_  = \new_[2831]_  | \new_[2832]_ ;
  assign \new_[5443]_  = \new_[2829]_  | \new_[2830]_ ;
  assign \new_[5444]_  = \new_[5443]_  | \new_[5440]_ ;
  assign \new_[5445]_  = \new_[5444]_  | \new_[5437]_ ;
  assign \new_[5449]_  = \new_[2826]_  | \new_[2827]_ ;
  assign \new_[5450]_  = \new_[2828]_  | \new_[5449]_ ;
  assign \new_[5453]_  = \new_[2824]_  | \new_[2825]_ ;
  assign \new_[5456]_  = \new_[2822]_  | \new_[2823]_ ;
  assign \new_[5457]_  = \new_[5456]_  | \new_[5453]_ ;
  assign \new_[5458]_  = \new_[5457]_  | \new_[5450]_ ;
  assign \new_[5459]_  = \new_[5458]_  | \new_[5445]_ ;
  assign \new_[5463]_  = \new_[2819]_  | \new_[2820]_ ;
  assign \new_[5464]_  = \new_[2821]_  | \new_[5463]_ ;
  assign \new_[5467]_  = \new_[2817]_  | \new_[2818]_ ;
  assign \new_[5470]_  = \new_[2815]_  | \new_[2816]_ ;
  assign \new_[5471]_  = \new_[5470]_  | \new_[5467]_ ;
  assign \new_[5472]_  = \new_[5471]_  | \new_[5464]_ ;
  assign \new_[5475]_  = \new_[2813]_  | \new_[2814]_ ;
  assign \new_[5478]_  = \new_[2811]_  | \new_[2812]_ ;
  assign \new_[5479]_  = \new_[5478]_  | \new_[5475]_ ;
  assign \new_[5482]_  = \new_[2809]_  | \new_[2810]_ ;
  assign \new_[5485]_  = \new_[2807]_  | \new_[2808]_ ;
  assign \new_[5486]_  = \new_[5485]_  | \new_[5482]_ ;
  assign \new_[5487]_  = \new_[5486]_  | \new_[5479]_ ;
  assign \new_[5488]_  = \new_[5487]_  | \new_[5472]_ ;
  assign \new_[5489]_  = \new_[5488]_  | \new_[5459]_ ;
  assign \new_[5493]_  = \new_[2804]_  | \new_[2805]_ ;
  assign \new_[5494]_  = \new_[2806]_  | \new_[5493]_ ;
  assign \new_[5497]_  = \new_[2802]_  | \new_[2803]_ ;
  assign \new_[5500]_  = \new_[2800]_  | \new_[2801]_ ;
  assign \new_[5501]_  = \new_[5500]_  | \new_[5497]_ ;
  assign \new_[5502]_  = \new_[5501]_  | \new_[5494]_ ;
  assign \new_[5506]_  = \new_[2797]_  | \new_[2798]_ ;
  assign \new_[5507]_  = \new_[2799]_  | \new_[5506]_ ;
  assign \new_[5510]_  = \new_[2795]_  | \new_[2796]_ ;
  assign \new_[5513]_  = \new_[2793]_  | \new_[2794]_ ;
  assign \new_[5514]_  = \new_[5513]_  | \new_[5510]_ ;
  assign \new_[5515]_  = \new_[5514]_  | \new_[5507]_ ;
  assign \new_[5516]_  = \new_[5515]_  | \new_[5502]_ ;
  assign \new_[5520]_  = \new_[2790]_  | \new_[2791]_ ;
  assign \new_[5521]_  = \new_[2792]_  | \new_[5520]_ ;
  assign \new_[5524]_  = \new_[2788]_  | \new_[2789]_ ;
  assign \new_[5527]_  = \new_[2786]_  | \new_[2787]_ ;
  assign \new_[5528]_  = \new_[5527]_  | \new_[5524]_ ;
  assign \new_[5529]_  = \new_[5528]_  | \new_[5521]_ ;
  assign \new_[5532]_  = \new_[2784]_  | \new_[2785]_ ;
  assign \new_[5535]_  = \new_[2782]_  | \new_[2783]_ ;
  assign \new_[5536]_  = \new_[5535]_  | \new_[5532]_ ;
  assign \new_[5539]_  = \new_[2780]_  | \new_[2781]_ ;
  assign \new_[5542]_  = \new_[2778]_  | \new_[2779]_ ;
  assign \new_[5543]_  = \new_[5542]_  | \new_[5539]_ ;
  assign \new_[5544]_  = \new_[5543]_  | \new_[5536]_ ;
  assign \new_[5545]_  = \new_[5544]_  | \new_[5529]_ ;
  assign \new_[5546]_  = \new_[5545]_  | \new_[5516]_ ;
  assign \new_[5547]_  = \new_[5546]_  | \new_[5489]_ ;
  assign \new_[5548]_  = \new_[5547]_  | \new_[5432]_ ;
  assign \new_[5549]_  = \new_[5548]_  | \new_[5317]_ ;
  assign \new_[5550]_  = \new_[5549]_  | \new_[5086]_ ;
  assign \new_[5551]_  = \new_[5550]_  | \new_[4625]_ ;
  assign \new_[5555]_  = \new_[2775]_  | \new_[2776]_ ;
  assign \new_[5556]_  = \new_[2777]_  | \new_[5555]_ ;
  assign \new_[5559]_  = \new_[2773]_  | \new_[2774]_ ;
  assign \new_[5562]_  = \new_[2771]_  | \new_[2772]_ ;
  assign \new_[5563]_  = \new_[5562]_  | \new_[5559]_ ;
  assign \new_[5564]_  = \new_[5563]_  | \new_[5556]_ ;
  assign \new_[5568]_  = \new_[2768]_  | \new_[2769]_ ;
  assign \new_[5569]_  = \new_[2770]_  | \new_[5568]_ ;
  assign \new_[5572]_  = \new_[2766]_  | \new_[2767]_ ;
  assign \new_[5575]_  = \new_[2764]_  | \new_[2765]_ ;
  assign \new_[5576]_  = \new_[5575]_  | \new_[5572]_ ;
  assign \new_[5577]_  = \new_[5576]_  | \new_[5569]_ ;
  assign \new_[5578]_  = \new_[5577]_  | \new_[5564]_ ;
  assign \new_[5582]_  = \new_[2761]_  | \new_[2762]_ ;
  assign \new_[5583]_  = \new_[2763]_  | \new_[5582]_ ;
  assign \new_[5586]_  = \new_[2759]_  | \new_[2760]_ ;
  assign \new_[5589]_  = \new_[2757]_  | \new_[2758]_ ;
  assign \new_[5590]_  = \new_[5589]_  | \new_[5586]_ ;
  assign \new_[5591]_  = \new_[5590]_  | \new_[5583]_ ;
  assign \new_[5595]_  = \new_[2754]_  | \new_[2755]_ ;
  assign \new_[5596]_  = \new_[2756]_  | \new_[5595]_ ;
  assign \new_[5599]_  = \new_[2752]_  | \new_[2753]_ ;
  assign \new_[5602]_  = \new_[2750]_  | \new_[2751]_ ;
  assign \new_[5603]_  = \new_[5602]_  | \new_[5599]_ ;
  assign \new_[5604]_  = \new_[5603]_  | \new_[5596]_ ;
  assign \new_[5605]_  = \new_[5604]_  | \new_[5591]_ ;
  assign \new_[5606]_  = \new_[5605]_  | \new_[5578]_ ;
  assign \new_[5610]_  = \new_[2747]_  | \new_[2748]_ ;
  assign \new_[5611]_  = \new_[2749]_  | \new_[5610]_ ;
  assign \new_[5614]_  = \new_[2745]_  | \new_[2746]_ ;
  assign \new_[5617]_  = \new_[2743]_  | \new_[2744]_ ;
  assign \new_[5618]_  = \new_[5617]_  | \new_[5614]_ ;
  assign \new_[5619]_  = \new_[5618]_  | \new_[5611]_ ;
  assign \new_[5623]_  = \new_[2740]_  | \new_[2741]_ ;
  assign \new_[5624]_  = \new_[2742]_  | \new_[5623]_ ;
  assign \new_[5627]_  = \new_[2738]_  | \new_[2739]_ ;
  assign \new_[5630]_  = \new_[2736]_  | \new_[2737]_ ;
  assign \new_[5631]_  = \new_[5630]_  | \new_[5627]_ ;
  assign \new_[5632]_  = \new_[5631]_  | \new_[5624]_ ;
  assign \new_[5633]_  = \new_[5632]_  | \new_[5619]_ ;
  assign \new_[5637]_  = \new_[2733]_  | \new_[2734]_ ;
  assign \new_[5638]_  = \new_[2735]_  | \new_[5637]_ ;
  assign \new_[5641]_  = \new_[2731]_  | \new_[2732]_ ;
  assign \new_[5644]_  = \new_[2729]_  | \new_[2730]_ ;
  assign \new_[5645]_  = \new_[5644]_  | \new_[5641]_ ;
  assign \new_[5646]_  = \new_[5645]_  | \new_[5638]_ ;
  assign \new_[5649]_  = \new_[2727]_  | \new_[2728]_ ;
  assign \new_[5652]_  = \new_[2725]_  | \new_[2726]_ ;
  assign \new_[5653]_  = \new_[5652]_  | \new_[5649]_ ;
  assign \new_[5656]_  = \new_[2723]_  | \new_[2724]_ ;
  assign \new_[5659]_  = \new_[2721]_  | \new_[2722]_ ;
  assign \new_[5660]_  = \new_[5659]_  | \new_[5656]_ ;
  assign \new_[5661]_  = \new_[5660]_  | \new_[5653]_ ;
  assign \new_[5662]_  = \new_[5661]_  | \new_[5646]_ ;
  assign \new_[5663]_  = \new_[5662]_  | \new_[5633]_ ;
  assign \new_[5664]_  = \new_[5663]_  | \new_[5606]_ ;
  assign \new_[5668]_  = \new_[2718]_  | \new_[2719]_ ;
  assign \new_[5669]_  = \new_[2720]_  | \new_[5668]_ ;
  assign \new_[5672]_  = \new_[2716]_  | \new_[2717]_ ;
  assign \new_[5675]_  = \new_[2714]_  | \new_[2715]_ ;
  assign \new_[5676]_  = \new_[5675]_  | \new_[5672]_ ;
  assign \new_[5677]_  = \new_[5676]_  | \new_[5669]_ ;
  assign \new_[5681]_  = \new_[2711]_  | \new_[2712]_ ;
  assign \new_[5682]_  = \new_[2713]_  | \new_[5681]_ ;
  assign \new_[5685]_  = \new_[2709]_  | \new_[2710]_ ;
  assign \new_[5688]_  = \new_[2707]_  | \new_[2708]_ ;
  assign \new_[5689]_  = \new_[5688]_  | \new_[5685]_ ;
  assign \new_[5690]_  = \new_[5689]_  | \new_[5682]_ ;
  assign \new_[5691]_  = \new_[5690]_  | \new_[5677]_ ;
  assign \new_[5695]_  = \new_[2704]_  | \new_[2705]_ ;
  assign \new_[5696]_  = \new_[2706]_  | \new_[5695]_ ;
  assign \new_[5699]_  = \new_[2702]_  | \new_[2703]_ ;
  assign \new_[5702]_  = \new_[2700]_  | \new_[2701]_ ;
  assign \new_[5703]_  = \new_[5702]_  | \new_[5699]_ ;
  assign \new_[5704]_  = \new_[5703]_  | \new_[5696]_ ;
  assign \new_[5707]_  = \new_[2698]_  | \new_[2699]_ ;
  assign \new_[5710]_  = \new_[2696]_  | \new_[2697]_ ;
  assign \new_[5711]_  = \new_[5710]_  | \new_[5707]_ ;
  assign \new_[5714]_  = \new_[2694]_  | \new_[2695]_ ;
  assign \new_[5717]_  = \new_[2692]_  | \new_[2693]_ ;
  assign \new_[5718]_  = \new_[5717]_  | \new_[5714]_ ;
  assign \new_[5719]_  = \new_[5718]_  | \new_[5711]_ ;
  assign \new_[5720]_  = \new_[5719]_  | \new_[5704]_ ;
  assign \new_[5721]_  = \new_[5720]_  | \new_[5691]_ ;
  assign \new_[5725]_  = \new_[2689]_  | \new_[2690]_ ;
  assign \new_[5726]_  = \new_[2691]_  | \new_[5725]_ ;
  assign \new_[5729]_  = \new_[2687]_  | \new_[2688]_ ;
  assign \new_[5732]_  = \new_[2685]_  | \new_[2686]_ ;
  assign \new_[5733]_  = \new_[5732]_  | \new_[5729]_ ;
  assign \new_[5734]_  = \new_[5733]_  | \new_[5726]_ ;
  assign \new_[5738]_  = \new_[2682]_  | \new_[2683]_ ;
  assign \new_[5739]_  = \new_[2684]_  | \new_[5738]_ ;
  assign \new_[5742]_  = \new_[2680]_  | \new_[2681]_ ;
  assign \new_[5745]_  = \new_[2678]_  | \new_[2679]_ ;
  assign \new_[5746]_  = \new_[5745]_  | \new_[5742]_ ;
  assign \new_[5747]_  = \new_[5746]_  | \new_[5739]_ ;
  assign \new_[5748]_  = \new_[5747]_  | \new_[5734]_ ;
  assign \new_[5752]_  = \new_[2675]_  | \new_[2676]_ ;
  assign \new_[5753]_  = \new_[2677]_  | \new_[5752]_ ;
  assign \new_[5756]_  = \new_[2673]_  | \new_[2674]_ ;
  assign \new_[5759]_  = \new_[2671]_  | \new_[2672]_ ;
  assign \new_[5760]_  = \new_[5759]_  | \new_[5756]_ ;
  assign \new_[5761]_  = \new_[5760]_  | \new_[5753]_ ;
  assign \new_[5764]_  = \new_[2669]_  | \new_[2670]_ ;
  assign \new_[5767]_  = \new_[2667]_  | \new_[2668]_ ;
  assign \new_[5768]_  = \new_[5767]_  | \new_[5764]_ ;
  assign \new_[5771]_  = \new_[2665]_  | \new_[2666]_ ;
  assign \new_[5774]_  = \new_[2663]_  | \new_[2664]_ ;
  assign \new_[5775]_  = \new_[5774]_  | \new_[5771]_ ;
  assign \new_[5776]_  = \new_[5775]_  | \new_[5768]_ ;
  assign \new_[5777]_  = \new_[5776]_  | \new_[5761]_ ;
  assign \new_[5778]_  = \new_[5777]_  | \new_[5748]_ ;
  assign \new_[5779]_  = \new_[5778]_  | \new_[5721]_ ;
  assign \new_[5780]_  = \new_[5779]_  | \new_[5664]_ ;
  assign \new_[5784]_  = \new_[2660]_  | \new_[2661]_ ;
  assign \new_[5785]_  = \new_[2662]_  | \new_[5784]_ ;
  assign \new_[5788]_  = \new_[2658]_  | \new_[2659]_ ;
  assign \new_[5791]_  = \new_[2656]_  | \new_[2657]_ ;
  assign \new_[5792]_  = \new_[5791]_  | \new_[5788]_ ;
  assign \new_[5793]_  = \new_[5792]_  | \new_[5785]_ ;
  assign \new_[5797]_  = \new_[2653]_  | \new_[2654]_ ;
  assign \new_[5798]_  = \new_[2655]_  | \new_[5797]_ ;
  assign \new_[5801]_  = \new_[2651]_  | \new_[2652]_ ;
  assign \new_[5804]_  = \new_[2649]_  | \new_[2650]_ ;
  assign \new_[5805]_  = \new_[5804]_  | \new_[5801]_ ;
  assign \new_[5806]_  = \new_[5805]_  | \new_[5798]_ ;
  assign \new_[5807]_  = \new_[5806]_  | \new_[5793]_ ;
  assign \new_[5811]_  = \new_[2646]_  | \new_[2647]_ ;
  assign \new_[5812]_  = \new_[2648]_  | \new_[5811]_ ;
  assign \new_[5815]_  = \new_[2644]_  | \new_[2645]_ ;
  assign \new_[5818]_  = \new_[2642]_  | \new_[2643]_ ;
  assign \new_[5819]_  = \new_[5818]_  | \new_[5815]_ ;
  assign \new_[5820]_  = \new_[5819]_  | \new_[5812]_ ;
  assign \new_[5823]_  = \new_[2640]_  | \new_[2641]_ ;
  assign \new_[5826]_  = \new_[2638]_  | \new_[2639]_ ;
  assign \new_[5827]_  = \new_[5826]_  | \new_[5823]_ ;
  assign \new_[5830]_  = \new_[2636]_  | \new_[2637]_ ;
  assign \new_[5833]_  = \new_[2634]_  | \new_[2635]_ ;
  assign \new_[5834]_  = \new_[5833]_  | \new_[5830]_ ;
  assign \new_[5835]_  = \new_[5834]_  | \new_[5827]_ ;
  assign \new_[5836]_  = \new_[5835]_  | \new_[5820]_ ;
  assign \new_[5837]_  = \new_[5836]_  | \new_[5807]_ ;
  assign \new_[5841]_  = \new_[2631]_  | \new_[2632]_ ;
  assign \new_[5842]_  = \new_[2633]_  | \new_[5841]_ ;
  assign \new_[5845]_  = \new_[2629]_  | \new_[2630]_ ;
  assign \new_[5848]_  = \new_[2627]_  | \new_[2628]_ ;
  assign \new_[5849]_  = \new_[5848]_  | \new_[5845]_ ;
  assign \new_[5850]_  = \new_[5849]_  | \new_[5842]_ ;
  assign \new_[5854]_  = \new_[2624]_  | \new_[2625]_ ;
  assign \new_[5855]_  = \new_[2626]_  | \new_[5854]_ ;
  assign \new_[5858]_  = \new_[2622]_  | \new_[2623]_ ;
  assign \new_[5861]_  = \new_[2620]_  | \new_[2621]_ ;
  assign \new_[5862]_  = \new_[5861]_  | \new_[5858]_ ;
  assign \new_[5863]_  = \new_[5862]_  | \new_[5855]_ ;
  assign \new_[5864]_  = \new_[5863]_  | \new_[5850]_ ;
  assign \new_[5868]_  = \new_[2617]_  | \new_[2618]_ ;
  assign \new_[5869]_  = \new_[2619]_  | \new_[5868]_ ;
  assign \new_[5872]_  = \new_[2615]_  | \new_[2616]_ ;
  assign \new_[5875]_  = \new_[2613]_  | \new_[2614]_ ;
  assign \new_[5876]_  = \new_[5875]_  | \new_[5872]_ ;
  assign \new_[5877]_  = \new_[5876]_  | \new_[5869]_ ;
  assign \new_[5880]_  = \new_[2611]_  | \new_[2612]_ ;
  assign \new_[5883]_  = \new_[2609]_  | \new_[2610]_ ;
  assign \new_[5884]_  = \new_[5883]_  | \new_[5880]_ ;
  assign \new_[5887]_  = \new_[2607]_  | \new_[2608]_ ;
  assign \new_[5890]_  = \new_[2605]_  | \new_[2606]_ ;
  assign \new_[5891]_  = \new_[5890]_  | \new_[5887]_ ;
  assign \new_[5892]_  = \new_[5891]_  | \new_[5884]_ ;
  assign \new_[5893]_  = \new_[5892]_  | \new_[5877]_ ;
  assign \new_[5894]_  = \new_[5893]_  | \new_[5864]_ ;
  assign \new_[5895]_  = \new_[5894]_  | \new_[5837]_ ;
  assign \new_[5899]_  = \new_[2602]_  | \new_[2603]_ ;
  assign \new_[5900]_  = \new_[2604]_  | \new_[5899]_ ;
  assign \new_[5903]_  = \new_[2600]_  | \new_[2601]_ ;
  assign \new_[5906]_  = \new_[2598]_  | \new_[2599]_ ;
  assign \new_[5907]_  = \new_[5906]_  | \new_[5903]_ ;
  assign \new_[5908]_  = \new_[5907]_  | \new_[5900]_ ;
  assign \new_[5912]_  = \new_[2595]_  | \new_[2596]_ ;
  assign \new_[5913]_  = \new_[2597]_  | \new_[5912]_ ;
  assign \new_[5916]_  = \new_[2593]_  | \new_[2594]_ ;
  assign \new_[5919]_  = \new_[2591]_  | \new_[2592]_ ;
  assign \new_[5920]_  = \new_[5919]_  | \new_[5916]_ ;
  assign \new_[5921]_  = \new_[5920]_  | \new_[5913]_ ;
  assign \new_[5922]_  = \new_[5921]_  | \new_[5908]_ ;
  assign \new_[5926]_  = \new_[2588]_  | \new_[2589]_ ;
  assign \new_[5927]_  = \new_[2590]_  | \new_[5926]_ ;
  assign \new_[5930]_  = \new_[2586]_  | \new_[2587]_ ;
  assign \new_[5933]_  = \new_[2584]_  | \new_[2585]_ ;
  assign \new_[5934]_  = \new_[5933]_  | \new_[5930]_ ;
  assign \new_[5935]_  = \new_[5934]_  | \new_[5927]_ ;
  assign \new_[5938]_  = \new_[2582]_  | \new_[2583]_ ;
  assign \new_[5941]_  = \new_[2580]_  | \new_[2581]_ ;
  assign \new_[5942]_  = \new_[5941]_  | \new_[5938]_ ;
  assign \new_[5945]_  = \new_[2578]_  | \new_[2579]_ ;
  assign \new_[5948]_  = \new_[2576]_  | \new_[2577]_ ;
  assign \new_[5949]_  = \new_[5948]_  | \new_[5945]_ ;
  assign \new_[5950]_  = \new_[5949]_  | \new_[5942]_ ;
  assign \new_[5951]_  = \new_[5950]_  | \new_[5935]_ ;
  assign \new_[5952]_  = \new_[5951]_  | \new_[5922]_ ;
  assign \new_[5956]_  = \new_[2573]_  | \new_[2574]_ ;
  assign \new_[5957]_  = \new_[2575]_  | \new_[5956]_ ;
  assign \new_[5960]_  = \new_[2571]_  | \new_[2572]_ ;
  assign \new_[5963]_  = \new_[2569]_  | \new_[2570]_ ;
  assign \new_[5964]_  = \new_[5963]_  | \new_[5960]_ ;
  assign \new_[5965]_  = \new_[5964]_  | \new_[5957]_ ;
  assign \new_[5969]_  = \new_[2566]_  | \new_[2567]_ ;
  assign \new_[5970]_  = \new_[2568]_  | \new_[5969]_ ;
  assign \new_[5973]_  = \new_[2564]_  | \new_[2565]_ ;
  assign \new_[5976]_  = \new_[2562]_  | \new_[2563]_ ;
  assign \new_[5977]_  = \new_[5976]_  | \new_[5973]_ ;
  assign \new_[5978]_  = \new_[5977]_  | \new_[5970]_ ;
  assign \new_[5979]_  = \new_[5978]_  | \new_[5965]_ ;
  assign \new_[5983]_  = \new_[2559]_  | \new_[2560]_ ;
  assign \new_[5984]_  = \new_[2561]_  | \new_[5983]_ ;
  assign \new_[5987]_  = \new_[2557]_  | \new_[2558]_ ;
  assign \new_[5990]_  = \new_[2555]_  | \new_[2556]_ ;
  assign \new_[5991]_  = \new_[5990]_  | \new_[5987]_ ;
  assign \new_[5992]_  = \new_[5991]_  | \new_[5984]_ ;
  assign \new_[5995]_  = \new_[2553]_  | \new_[2554]_ ;
  assign \new_[5998]_  = \new_[2551]_  | \new_[2552]_ ;
  assign \new_[5999]_  = \new_[5998]_  | \new_[5995]_ ;
  assign \new_[6002]_  = \new_[2549]_  | \new_[2550]_ ;
  assign \new_[6005]_  = \new_[2547]_  | \new_[2548]_ ;
  assign \new_[6006]_  = \new_[6005]_  | \new_[6002]_ ;
  assign \new_[6007]_  = \new_[6006]_  | \new_[5999]_ ;
  assign \new_[6008]_  = \new_[6007]_  | \new_[5992]_ ;
  assign \new_[6009]_  = \new_[6008]_  | \new_[5979]_ ;
  assign \new_[6010]_  = \new_[6009]_  | \new_[5952]_ ;
  assign \new_[6011]_  = \new_[6010]_  | \new_[5895]_ ;
  assign \new_[6012]_  = \new_[6011]_  | \new_[5780]_ ;
  assign \new_[6016]_  = \new_[2544]_  | \new_[2545]_ ;
  assign \new_[6017]_  = \new_[2546]_  | \new_[6016]_ ;
  assign \new_[6020]_  = \new_[2542]_  | \new_[2543]_ ;
  assign \new_[6023]_  = \new_[2540]_  | \new_[2541]_ ;
  assign \new_[6024]_  = \new_[6023]_  | \new_[6020]_ ;
  assign \new_[6025]_  = \new_[6024]_  | \new_[6017]_ ;
  assign \new_[6029]_  = \new_[2537]_  | \new_[2538]_ ;
  assign \new_[6030]_  = \new_[2539]_  | \new_[6029]_ ;
  assign \new_[6033]_  = \new_[2535]_  | \new_[2536]_ ;
  assign \new_[6036]_  = \new_[2533]_  | \new_[2534]_ ;
  assign \new_[6037]_  = \new_[6036]_  | \new_[6033]_ ;
  assign \new_[6038]_  = \new_[6037]_  | \new_[6030]_ ;
  assign \new_[6039]_  = \new_[6038]_  | \new_[6025]_ ;
  assign \new_[6043]_  = \new_[2530]_  | \new_[2531]_ ;
  assign \new_[6044]_  = \new_[2532]_  | \new_[6043]_ ;
  assign \new_[6047]_  = \new_[2528]_  | \new_[2529]_ ;
  assign \new_[6050]_  = \new_[2526]_  | \new_[2527]_ ;
  assign \new_[6051]_  = \new_[6050]_  | \new_[6047]_ ;
  assign \new_[6052]_  = \new_[6051]_  | \new_[6044]_ ;
  assign \new_[6055]_  = \new_[2524]_  | \new_[2525]_ ;
  assign \new_[6058]_  = \new_[2522]_  | \new_[2523]_ ;
  assign \new_[6059]_  = \new_[6058]_  | \new_[6055]_ ;
  assign \new_[6062]_  = \new_[2520]_  | \new_[2521]_ ;
  assign \new_[6065]_  = \new_[2518]_  | \new_[2519]_ ;
  assign \new_[6066]_  = \new_[6065]_  | \new_[6062]_ ;
  assign \new_[6067]_  = \new_[6066]_  | \new_[6059]_ ;
  assign \new_[6068]_  = \new_[6067]_  | \new_[6052]_ ;
  assign \new_[6069]_  = \new_[6068]_  | \new_[6039]_ ;
  assign \new_[6073]_  = \new_[2515]_  | \new_[2516]_ ;
  assign \new_[6074]_  = \new_[2517]_  | \new_[6073]_ ;
  assign \new_[6077]_  = \new_[2513]_  | \new_[2514]_ ;
  assign \new_[6080]_  = \new_[2511]_  | \new_[2512]_ ;
  assign \new_[6081]_  = \new_[6080]_  | \new_[6077]_ ;
  assign \new_[6082]_  = \new_[6081]_  | \new_[6074]_ ;
  assign \new_[6086]_  = \new_[2508]_  | \new_[2509]_ ;
  assign \new_[6087]_  = \new_[2510]_  | \new_[6086]_ ;
  assign \new_[6090]_  = \new_[2506]_  | \new_[2507]_ ;
  assign \new_[6093]_  = \new_[2504]_  | \new_[2505]_ ;
  assign \new_[6094]_  = \new_[6093]_  | \new_[6090]_ ;
  assign \new_[6095]_  = \new_[6094]_  | \new_[6087]_ ;
  assign \new_[6096]_  = \new_[6095]_  | \new_[6082]_ ;
  assign \new_[6100]_  = \new_[2501]_  | \new_[2502]_ ;
  assign \new_[6101]_  = \new_[2503]_  | \new_[6100]_ ;
  assign \new_[6104]_  = \new_[2499]_  | \new_[2500]_ ;
  assign \new_[6107]_  = \new_[2497]_  | \new_[2498]_ ;
  assign \new_[6108]_  = \new_[6107]_  | \new_[6104]_ ;
  assign \new_[6109]_  = \new_[6108]_  | \new_[6101]_ ;
  assign \new_[6112]_  = \new_[2495]_  | \new_[2496]_ ;
  assign \new_[6115]_  = \new_[2493]_  | \new_[2494]_ ;
  assign \new_[6116]_  = \new_[6115]_  | \new_[6112]_ ;
  assign \new_[6119]_  = \new_[2491]_  | \new_[2492]_ ;
  assign \new_[6122]_  = \new_[2489]_  | \new_[2490]_ ;
  assign \new_[6123]_  = \new_[6122]_  | \new_[6119]_ ;
  assign \new_[6124]_  = \new_[6123]_  | \new_[6116]_ ;
  assign \new_[6125]_  = \new_[6124]_  | \new_[6109]_ ;
  assign \new_[6126]_  = \new_[6125]_  | \new_[6096]_ ;
  assign \new_[6127]_  = \new_[6126]_  | \new_[6069]_ ;
  assign \new_[6131]_  = \new_[2486]_  | \new_[2487]_ ;
  assign \new_[6132]_  = \new_[2488]_  | \new_[6131]_ ;
  assign \new_[6135]_  = \new_[2484]_  | \new_[2485]_ ;
  assign \new_[6138]_  = \new_[2482]_  | \new_[2483]_ ;
  assign \new_[6139]_  = \new_[6138]_  | \new_[6135]_ ;
  assign \new_[6140]_  = \new_[6139]_  | \new_[6132]_ ;
  assign \new_[6144]_  = \new_[2479]_  | \new_[2480]_ ;
  assign \new_[6145]_  = \new_[2481]_  | \new_[6144]_ ;
  assign \new_[6148]_  = \new_[2477]_  | \new_[2478]_ ;
  assign \new_[6151]_  = \new_[2475]_  | \new_[2476]_ ;
  assign \new_[6152]_  = \new_[6151]_  | \new_[6148]_ ;
  assign \new_[6153]_  = \new_[6152]_  | \new_[6145]_ ;
  assign \new_[6154]_  = \new_[6153]_  | \new_[6140]_ ;
  assign \new_[6158]_  = \new_[2472]_  | \new_[2473]_ ;
  assign \new_[6159]_  = \new_[2474]_  | \new_[6158]_ ;
  assign \new_[6162]_  = \new_[2470]_  | \new_[2471]_ ;
  assign \new_[6165]_  = \new_[2468]_  | \new_[2469]_ ;
  assign \new_[6166]_  = \new_[6165]_  | \new_[6162]_ ;
  assign \new_[6167]_  = \new_[6166]_  | \new_[6159]_ ;
  assign \new_[6170]_  = \new_[2466]_  | \new_[2467]_ ;
  assign \new_[6173]_  = \new_[2464]_  | \new_[2465]_ ;
  assign \new_[6174]_  = \new_[6173]_  | \new_[6170]_ ;
  assign \new_[6177]_  = \new_[2462]_  | \new_[2463]_ ;
  assign \new_[6180]_  = \new_[2460]_  | \new_[2461]_ ;
  assign \new_[6181]_  = \new_[6180]_  | \new_[6177]_ ;
  assign \new_[6182]_  = \new_[6181]_  | \new_[6174]_ ;
  assign \new_[6183]_  = \new_[6182]_  | \new_[6167]_ ;
  assign \new_[6184]_  = \new_[6183]_  | \new_[6154]_ ;
  assign \new_[6188]_  = \new_[2457]_  | \new_[2458]_ ;
  assign \new_[6189]_  = \new_[2459]_  | \new_[6188]_ ;
  assign \new_[6192]_  = \new_[2455]_  | \new_[2456]_ ;
  assign \new_[6195]_  = \new_[2453]_  | \new_[2454]_ ;
  assign \new_[6196]_  = \new_[6195]_  | \new_[6192]_ ;
  assign \new_[6197]_  = \new_[6196]_  | \new_[6189]_ ;
  assign \new_[6201]_  = \new_[2450]_  | \new_[2451]_ ;
  assign \new_[6202]_  = \new_[2452]_  | \new_[6201]_ ;
  assign \new_[6205]_  = \new_[2448]_  | \new_[2449]_ ;
  assign \new_[6208]_  = \new_[2446]_  | \new_[2447]_ ;
  assign \new_[6209]_  = \new_[6208]_  | \new_[6205]_ ;
  assign \new_[6210]_  = \new_[6209]_  | \new_[6202]_ ;
  assign \new_[6211]_  = \new_[6210]_  | \new_[6197]_ ;
  assign \new_[6215]_  = \new_[2443]_  | \new_[2444]_ ;
  assign \new_[6216]_  = \new_[2445]_  | \new_[6215]_ ;
  assign \new_[6219]_  = \new_[2441]_  | \new_[2442]_ ;
  assign \new_[6222]_  = \new_[2439]_  | \new_[2440]_ ;
  assign \new_[6223]_  = \new_[6222]_  | \new_[6219]_ ;
  assign \new_[6224]_  = \new_[6223]_  | \new_[6216]_ ;
  assign \new_[6227]_  = \new_[2437]_  | \new_[2438]_ ;
  assign \new_[6230]_  = \new_[2435]_  | \new_[2436]_ ;
  assign \new_[6231]_  = \new_[6230]_  | \new_[6227]_ ;
  assign \new_[6234]_  = \new_[2433]_  | \new_[2434]_ ;
  assign \new_[6237]_  = \new_[2431]_  | \new_[2432]_ ;
  assign \new_[6238]_  = \new_[6237]_  | \new_[6234]_ ;
  assign \new_[6239]_  = \new_[6238]_  | \new_[6231]_ ;
  assign \new_[6240]_  = \new_[6239]_  | \new_[6224]_ ;
  assign \new_[6241]_  = \new_[6240]_  | \new_[6211]_ ;
  assign \new_[6242]_  = \new_[6241]_  | \new_[6184]_ ;
  assign \new_[6243]_  = \new_[6242]_  | \new_[6127]_ ;
  assign \new_[6247]_  = \new_[2428]_  | \new_[2429]_ ;
  assign \new_[6248]_  = \new_[2430]_  | \new_[6247]_ ;
  assign \new_[6251]_  = \new_[2426]_  | \new_[2427]_ ;
  assign \new_[6254]_  = \new_[2424]_  | \new_[2425]_ ;
  assign \new_[6255]_  = \new_[6254]_  | \new_[6251]_ ;
  assign \new_[6256]_  = \new_[6255]_  | \new_[6248]_ ;
  assign \new_[6260]_  = \new_[2421]_  | \new_[2422]_ ;
  assign \new_[6261]_  = \new_[2423]_  | \new_[6260]_ ;
  assign \new_[6264]_  = \new_[2419]_  | \new_[2420]_ ;
  assign \new_[6267]_  = \new_[2417]_  | \new_[2418]_ ;
  assign \new_[6268]_  = \new_[6267]_  | \new_[6264]_ ;
  assign \new_[6269]_  = \new_[6268]_  | \new_[6261]_ ;
  assign \new_[6270]_  = \new_[6269]_  | \new_[6256]_ ;
  assign \new_[6274]_  = \new_[2414]_  | \new_[2415]_ ;
  assign \new_[6275]_  = \new_[2416]_  | \new_[6274]_ ;
  assign \new_[6278]_  = \new_[2412]_  | \new_[2413]_ ;
  assign \new_[6281]_  = \new_[2410]_  | \new_[2411]_ ;
  assign \new_[6282]_  = \new_[6281]_  | \new_[6278]_ ;
  assign \new_[6283]_  = \new_[6282]_  | \new_[6275]_ ;
  assign \new_[6286]_  = \new_[2408]_  | \new_[2409]_ ;
  assign \new_[6289]_  = \new_[2406]_  | \new_[2407]_ ;
  assign \new_[6290]_  = \new_[6289]_  | \new_[6286]_ ;
  assign \new_[6293]_  = \new_[2404]_  | \new_[2405]_ ;
  assign \new_[6296]_  = \new_[2402]_  | \new_[2403]_ ;
  assign \new_[6297]_  = \new_[6296]_  | \new_[6293]_ ;
  assign \new_[6298]_  = \new_[6297]_  | \new_[6290]_ ;
  assign \new_[6299]_  = \new_[6298]_  | \new_[6283]_ ;
  assign \new_[6300]_  = \new_[6299]_  | \new_[6270]_ ;
  assign \new_[6304]_  = \new_[2399]_  | \new_[2400]_ ;
  assign \new_[6305]_  = \new_[2401]_  | \new_[6304]_ ;
  assign \new_[6308]_  = \new_[2397]_  | \new_[2398]_ ;
  assign \new_[6311]_  = \new_[2395]_  | \new_[2396]_ ;
  assign \new_[6312]_  = \new_[6311]_  | \new_[6308]_ ;
  assign \new_[6313]_  = \new_[6312]_  | \new_[6305]_ ;
  assign \new_[6317]_  = \new_[2392]_  | \new_[2393]_ ;
  assign \new_[6318]_  = \new_[2394]_  | \new_[6317]_ ;
  assign \new_[6321]_  = \new_[2390]_  | \new_[2391]_ ;
  assign \new_[6324]_  = \new_[2388]_  | \new_[2389]_ ;
  assign \new_[6325]_  = \new_[6324]_  | \new_[6321]_ ;
  assign \new_[6326]_  = \new_[6325]_  | \new_[6318]_ ;
  assign \new_[6327]_  = \new_[6326]_  | \new_[6313]_ ;
  assign \new_[6331]_  = \new_[2385]_  | \new_[2386]_ ;
  assign \new_[6332]_  = \new_[2387]_  | \new_[6331]_ ;
  assign \new_[6335]_  = \new_[2383]_  | \new_[2384]_ ;
  assign \new_[6338]_  = \new_[2381]_  | \new_[2382]_ ;
  assign \new_[6339]_  = \new_[6338]_  | \new_[6335]_ ;
  assign \new_[6340]_  = \new_[6339]_  | \new_[6332]_ ;
  assign \new_[6343]_  = \new_[2379]_  | \new_[2380]_ ;
  assign \new_[6346]_  = \new_[2377]_  | \new_[2378]_ ;
  assign \new_[6347]_  = \new_[6346]_  | \new_[6343]_ ;
  assign \new_[6350]_  = \new_[2375]_  | \new_[2376]_ ;
  assign \new_[6353]_  = \new_[2373]_  | \new_[2374]_ ;
  assign \new_[6354]_  = \new_[6353]_  | \new_[6350]_ ;
  assign \new_[6355]_  = \new_[6354]_  | \new_[6347]_ ;
  assign \new_[6356]_  = \new_[6355]_  | \new_[6340]_ ;
  assign \new_[6357]_  = \new_[6356]_  | \new_[6327]_ ;
  assign \new_[6358]_  = \new_[6357]_  | \new_[6300]_ ;
  assign \new_[6362]_  = \new_[2370]_  | \new_[2371]_ ;
  assign \new_[6363]_  = \new_[2372]_  | \new_[6362]_ ;
  assign \new_[6366]_  = \new_[2368]_  | \new_[2369]_ ;
  assign \new_[6369]_  = \new_[2366]_  | \new_[2367]_ ;
  assign \new_[6370]_  = \new_[6369]_  | \new_[6366]_ ;
  assign \new_[6371]_  = \new_[6370]_  | \new_[6363]_ ;
  assign \new_[6375]_  = \new_[2363]_  | \new_[2364]_ ;
  assign \new_[6376]_  = \new_[2365]_  | \new_[6375]_ ;
  assign \new_[6379]_  = \new_[2361]_  | \new_[2362]_ ;
  assign \new_[6382]_  = \new_[2359]_  | \new_[2360]_ ;
  assign \new_[6383]_  = \new_[6382]_  | \new_[6379]_ ;
  assign \new_[6384]_  = \new_[6383]_  | \new_[6376]_ ;
  assign \new_[6385]_  = \new_[6384]_  | \new_[6371]_ ;
  assign \new_[6389]_  = \new_[2356]_  | \new_[2357]_ ;
  assign \new_[6390]_  = \new_[2358]_  | \new_[6389]_ ;
  assign \new_[6393]_  = \new_[2354]_  | \new_[2355]_ ;
  assign \new_[6396]_  = \new_[2352]_  | \new_[2353]_ ;
  assign \new_[6397]_  = \new_[6396]_  | \new_[6393]_ ;
  assign \new_[6398]_  = \new_[6397]_  | \new_[6390]_ ;
  assign \new_[6401]_  = \new_[2350]_  | \new_[2351]_ ;
  assign \new_[6404]_  = \new_[2348]_  | \new_[2349]_ ;
  assign \new_[6405]_  = \new_[6404]_  | \new_[6401]_ ;
  assign \new_[6408]_  = \new_[2346]_  | \new_[2347]_ ;
  assign \new_[6411]_  = \new_[2344]_  | \new_[2345]_ ;
  assign \new_[6412]_  = \new_[6411]_  | \new_[6408]_ ;
  assign \new_[6413]_  = \new_[6412]_  | \new_[6405]_ ;
  assign \new_[6414]_  = \new_[6413]_  | \new_[6398]_ ;
  assign \new_[6415]_  = \new_[6414]_  | \new_[6385]_ ;
  assign \new_[6419]_  = \new_[2341]_  | \new_[2342]_ ;
  assign \new_[6420]_  = \new_[2343]_  | \new_[6419]_ ;
  assign \new_[6423]_  = \new_[2339]_  | \new_[2340]_ ;
  assign \new_[6426]_  = \new_[2337]_  | \new_[2338]_ ;
  assign \new_[6427]_  = \new_[6426]_  | \new_[6423]_ ;
  assign \new_[6428]_  = \new_[6427]_  | \new_[6420]_ ;
  assign \new_[6432]_  = \new_[2334]_  | \new_[2335]_ ;
  assign \new_[6433]_  = \new_[2336]_  | \new_[6432]_ ;
  assign \new_[6436]_  = \new_[2332]_  | \new_[2333]_ ;
  assign \new_[6439]_  = \new_[2330]_  | \new_[2331]_ ;
  assign \new_[6440]_  = \new_[6439]_  | \new_[6436]_ ;
  assign \new_[6441]_  = \new_[6440]_  | \new_[6433]_ ;
  assign \new_[6442]_  = \new_[6441]_  | \new_[6428]_ ;
  assign \new_[6446]_  = \new_[2327]_  | \new_[2328]_ ;
  assign \new_[6447]_  = \new_[2329]_  | \new_[6446]_ ;
  assign \new_[6450]_  = \new_[2325]_  | \new_[2326]_ ;
  assign \new_[6453]_  = \new_[2323]_  | \new_[2324]_ ;
  assign \new_[6454]_  = \new_[6453]_  | \new_[6450]_ ;
  assign \new_[6455]_  = \new_[6454]_  | \new_[6447]_ ;
  assign \new_[6458]_  = \new_[2321]_  | \new_[2322]_ ;
  assign \new_[6461]_  = \new_[2319]_  | \new_[2320]_ ;
  assign \new_[6462]_  = \new_[6461]_  | \new_[6458]_ ;
  assign \new_[6465]_  = \new_[2317]_  | \new_[2318]_ ;
  assign \new_[6468]_  = \new_[2315]_  | \new_[2316]_ ;
  assign \new_[6469]_  = \new_[6468]_  | \new_[6465]_ ;
  assign \new_[6470]_  = \new_[6469]_  | \new_[6462]_ ;
  assign \new_[6471]_  = \new_[6470]_  | \new_[6455]_ ;
  assign \new_[6472]_  = \new_[6471]_  | \new_[6442]_ ;
  assign \new_[6473]_  = \new_[6472]_  | \new_[6415]_ ;
  assign \new_[6474]_  = \new_[6473]_  | \new_[6358]_ ;
  assign \new_[6475]_  = \new_[6474]_  | \new_[6243]_ ;
  assign \new_[6476]_  = \new_[6475]_  | \new_[6012]_ ;
  assign \new_[6480]_  = \new_[2312]_  | \new_[2313]_ ;
  assign \new_[6481]_  = \new_[2314]_  | \new_[6480]_ ;
  assign \new_[6484]_  = \new_[2310]_  | \new_[2311]_ ;
  assign \new_[6487]_  = \new_[2308]_  | \new_[2309]_ ;
  assign \new_[6488]_  = \new_[6487]_  | \new_[6484]_ ;
  assign \new_[6489]_  = \new_[6488]_  | \new_[6481]_ ;
  assign \new_[6493]_  = \new_[2305]_  | \new_[2306]_ ;
  assign \new_[6494]_  = \new_[2307]_  | \new_[6493]_ ;
  assign \new_[6497]_  = \new_[2303]_  | \new_[2304]_ ;
  assign \new_[6500]_  = \new_[2301]_  | \new_[2302]_ ;
  assign \new_[6501]_  = \new_[6500]_  | \new_[6497]_ ;
  assign \new_[6502]_  = \new_[6501]_  | \new_[6494]_ ;
  assign \new_[6503]_  = \new_[6502]_  | \new_[6489]_ ;
  assign \new_[6507]_  = \new_[2298]_  | \new_[2299]_ ;
  assign \new_[6508]_  = \new_[2300]_  | \new_[6507]_ ;
  assign \new_[6511]_  = \new_[2296]_  | \new_[2297]_ ;
  assign \new_[6514]_  = \new_[2294]_  | \new_[2295]_ ;
  assign \new_[6515]_  = \new_[6514]_  | \new_[6511]_ ;
  assign \new_[6516]_  = \new_[6515]_  | \new_[6508]_ ;
  assign \new_[6520]_  = \new_[2291]_  | \new_[2292]_ ;
  assign \new_[6521]_  = \new_[2293]_  | \new_[6520]_ ;
  assign \new_[6524]_  = \new_[2289]_  | \new_[2290]_ ;
  assign \new_[6527]_  = \new_[2287]_  | \new_[2288]_ ;
  assign \new_[6528]_  = \new_[6527]_  | \new_[6524]_ ;
  assign \new_[6529]_  = \new_[6528]_  | \new_[6521]_ ;
  assign \new_[6530]_  = \new_[6529]_  | \new_[6516]_ ;
  assign \new_[6531]_  = \new_[6530]_  | \new_[6503]_ ;
  assign \new_[6535]_  = \new_[2284]_  | \new_[2285]_ ;
  assign \new_[6536]_  = \new_[2286]_  | \new_[6535]_ ;
  assign \new_[6539]_  = \new_[2282]_  | \new_[2283]_ ;
  assign \new_[6542]_  = \new_[2280]_  | \new_[2281]_ ;
  assign \new_[6543]_  = \new_[6542]_  | \new_[6539]_ ;
  assign \new_[6544]_  = \new_[6543]_  | \new_[6536]_ ;
  assign \new_[6548]_  = \new_[2277]_  | \new_[2278]_ ;
  assign \new_[6549]_  = \new_[2279]_  | \new_[6548]_ ;
  assign \new_[6552]_  = \new_[2275]_  | \new_[2276]_ ;
  assign \new_[6555]_  = \new_[2273]_  | \new_[2274]_ ;
  assign \new_[6556]_  = \new_[6555]_  | \new_[6552]_ ;
  assign \new_[6557]_  = \new_[6556]_  | \new_[6549]_ ;
  assign \new_[6558]_  = \new_[6557]_  | \new_[6544]_ ;
  assign \new_[6562]_  = \new_[2270]_  | \new_[2271]_ ;
  assign \new_[6563]_  = \new_[2272]_  | \new_[6562]_ ;
  assign \new_[6566]_  = \new_[2268]_  | \new_[2269]_ ;
  assign \new_[6569]_  = \new_[2266]_  | \new_[2267]_ ;
  assign \new_[6570]_  = \new_[6569]_  | \new_[6566]_ ;
  assign \new_[6571]_  = \new_[6570]_  | \new_[6563]_ ;
  assign \new_[6574]_  = \new_[2264]_  | \new_[2265]_ ;
  assign \new_[6577]_  = \new_[2262]_  | \new_[2263]_ ;
  assign \new_[6578]_  = \new_[6577]_  | \new_[6574]_ ;
  assign \new_[6581]_  = \new_[2260]_  | \new_[2261]_ ;
  assign \new_[6584]_  = \new_[2258]_  | \new_[2259]_ ;
  assign \new_[6585]_  = \new_[6584]_  | \new_[6581]_ ;
  assign \new_[6586]_  = \new_[6585]_  | \new_[6578]_ ;
  assign \new_[6587]_  = \new_[6586]_  | \new_[6571]_ ;
  assign \new_[6588]_  = \new_[6587]_  | \new_[6558]_ ;
  assign \new_[6589]_  = \new_[6588]_  | \new_[6531]_ ;
  assign \new_[6593]_  = \new_[2255]_  | \new_[2256]_ ;
  assign \new_[6594]_  = \new_[2257]_  | \new_[6593]_ ;
  assign \new_[6597]_  = \new_[2253]_  | \new_[2254]_ ;
  assign \new_[6600]_  = \new_[2251]_  | \new_[2252]_ ;
  assign \new_[6601]_  = \new_[6600]_  | \new_[6597]_ ;
  assign \new_[6602]_  = \new_[6601]_  | \new_[6594]_ ;
  assign \new_[6606]_  = \new_[2248]_  | \new_[2249]_ ;
  assign \new_[6607]_  = \new_[2250]_  | \new_[6606]_ ;
  assign \new_[6610]_  = \new_[2246]_  | \new_[2247]_ ;
  assign \new_[6613]_  = \new_[2244]_  | \new_[2245]_ ;
  assign \new_[6614]_  = \new_[6613]_  | \new_[6610]_ ;
  assign \new_[6615]_  = \new_[6614]_  | \new_[6607]_ ;
  assign \new_[6616]_  = \new_[6615]_  | \new_[6602]_ ;
  assign \new_[6620]_  = \new_[2241]_  | \new_[2242]_ ;
  assign \new_[6621]_  = \new_[2243]_  | \new_[6620]_ ;
  assign \new_[6624]_  = \new_[2239]_  | \new_[2240]_ ;
  assign \new_[6627]_  = \new_[2237]_  | \new_[2238]_ ;
  assign \new_[6628]_  = \new_[6627]_  | \new_[6624]_ ;
  assign \new_[6629]_  = \new_[6628]_  | \new_[6621]_ ;
  assign \new_[6632]_  = \new_[2235]_  | \new_[2236]_ ;
  assign \new_[6635]_  = \new_[2233]_  | \new_[2234]_ ;
  assign \new_[6636]_  = \new_[6635]_  | \new_[6632]_ ;
  assign \new_[6639]_  = \new_[2231]_  | \new_[2232]_ ;
  assign \new_[6642]_  = \new_[2229]_  | \new_[2230]_ ;
  assign \new_[6643]_  = \new_[6642]_  | \new_[6639]_ ;
  assign \new_[6644]_  = \new_[6643]_  | \new_[6636]_ ;
  assign \new_[6645]_  = \new_[6644]_  | \new_[6629]_ ;
  assign \new_[6646]_  = \new_[6645]_  | \new_[6616]_ ;
  assign \new_[6650]_  = \new_[2226]_  | \new_[2227]_ ;
  assign \new_[6651]_  = \new_[2228]_  | \new_[6650]_ ;
  assign \new_[6654]_  = \new_[2224]_  | \new_[2225]_ ;
  assign \new_[6657]_  = \new_[2222]_  | \new_[2223]_ ;
  assign \new_[6658]_  = \new_[6657]_  | \new_[6654]_ ;
  assign \new_[6659]_  = \new_[6658]_  | \new_[6651]_ ;
  assign \new_[6663]_  = \new_[2219]_  | \new_[2220]_ ;
  assign \new_[6664]_  = \new_[2221]_  | \new_[6663]_ ;
  assign \new_[6667]_  = \new_[2217]_  | \new_[2218]_ ;
  assign \new_[6670]_  = \new_[2215]_  | \new_[2216]_ ;
  assign \new_[6671]_  = \new_[6670]_  | \new_[6667]_ ;
  assign \new_[6672]_  = \new_[6671]_  | \new_[6664]_ ;
  assign \new_[6673]_  = \new_[6672]_  | \new_[6659]_ ;
  assign \new_[6677]_  = \new_[2212]_  | \new_[2213]_ ;
  assign \new_[6678]_  = \new_[2214]_  | \new_[6677]_ ;
  assign \new_[6681]_  = \new_[2210]_  | \new_[2211]_ ;
  assign \new_[6684]_  = \new_[2208]_  | \new_[2209]_ ;
  assign \new_[6685]_  = \new_[6684]_  | \new_[6681]_ ;
  assign \new_[6686]_  = \new_[6685]_  | \new_[6678]_ ;
  assign \new_[6689]_  = \new_[2206]_  | \new_[2207]_ ;
  assign \new_[6692]_  = \new_[2204]_  | \new_[2205]_ ;
  assign \new_[6693]_  = \new_[6692]_  | \new_[6689]_ ;
  assign \new_[6696]_  = \new_[2202]_  | \new_[2203]_ ;
  assign \new_[6699]_  = \new_[2200]_  | \new_[2201]_ ;
  assign \new_[6700]_  = \new_[6699]_  | \new_[6696]_ ;
  assign \new_[6701]_  = \new_[6700]_  | \new_[6693]_ ;
  assign \new_[6702]_  = \new_[6701]_  | \new_[6686]_ ;
  assign \new_[6703]_  = \new_[6702]_  | \new_[6673]_ ;
  assign \new_[6704]_  = \new_[6703]_  | \new_[6646]_ ;
  assign \new_[6705]_  = \new_[6704]_  | \new_[6589]_ ;
  assign \new_[6709]_  = \new_[2197]_  | \new_[2198]_ ;
  assign \new_[6710]_  = \new_[2199]_  | \new_[6709]_ ;
  assign \new_[6713]_  = \new_[2195]_  | \new_[2196]_ ;
  assign \new_[6716]_  = \new_[2193]_  | \new_[2194]_ ;
  assign \new_[6717]_  = \new_[6716]_  | \new_[6713]_ ;
  assign \new_[6718]_  = \new_[6717]_  | \new_[6710]_ ;
  assign \new_[6722]_  = \new_[2190]_  | \new_[2191]_ ;
  assign \new_[6723]_  = \new_[2192]_  | \new_[6722]_ ;
  assign \new_[6726]_  = \new_[2188]_  | \new_[2189]_ ;
  assign \new_[6729]_  = \new_[2186]_  | \new_[2187]_ ;
  assign \new_[6730]_  = \new_[6729]_  | \new_[6726]_ ;
  assign \new_[6731]_  = \new_[6730]_  | \new_[6723]_ ;
  assign \new_[6732]_  = \new_[6731]_  | \new_[6718]_ ;
  assign \new_[6736]_  = \new_[2183]_  | \new_[2184]_ ;
  assign \new_[6737]_  = \new_[2185]_  | \new_[6736]_ ;
  assign \new_[6740]_  = \new_[2181]_  | \new_[2182]_ ;
  assign \new_[6743]_  = \new_[2179]_  | \new_[2180]_ ;
  assign \new_[6744]_  = \new_[6743]_  | \new_[6740]_ ;
  assign \new_[6745]_  = \new_[6744]_  | \new_[6737]_ ;
  assign \new_[6748]_  = \new_[2177]_  | \new_[2178]_ ;
  assign \new_[6751]_  = \new_[2175]_  | \new_[2176]_ ;
  assign \new_[6752]_  = \new_[6751]_  | \new_[6748]_ ;
  assign \new_[6755]_  = \new_[2173]_  | \new_[2174]_ ;
  assign \new_[6758]_  = \new_[2171]_  | \new_[2172]_ ;
  assign \new_[6759]_  = \new_[6758]_  | \new_[6755]_ ;
  assign \new_[6760]_  = \new_[6759]_  | \new_[6752]_ ;
  assign \new_[6761]_  = \new_[6760]_  | \new_[6745]_ ;
  assign \new_[6762]_  = \new_[6761]_  | \new_[6732]_ ;
  assign \new_[6766]_  = \new_[2168]_  | \new_[2169]_ ;
  assign \new_[6767]_  = \new_[2170]_  | \new_[6766]_ ;
  assign \new_[6770]_  = \new_[2166]_  | \new_[2167]_ ;
  assign \new_[6773]_  = \new_[2164]_  | \new_[2165]_ ;
  assign \new_[6774]_  = \new_[6773]_  | \new_[6770]_ ;
  assign \new_[6775]_  = \new_[6774]_  | \new_[6767]_ ;
  assign \new_[6779]_  = \new_[2161]_  | \new_[2162]_ ;
  assign \new_[6780]_  = \new_[2163]_  | \new_[6779]_ ;
  assign \new_[6783]_  = \new_[2159]_  | \new_[2160]_ ;
  assign \new_[6786]_  = \new_[2157]_  | \new_[2158]_ ;
  assign \new_[6787]_  = \new_[6786]_  | \new_[6783]_ ;
  assign \new_[6788]_  = \new_[6787]_  | \new_[6780]_ ;
  assign \new_[6789]_  = \new_[6788]_  | \new_[6775]_ ;
  assign \new_[6793]_  = \new_[2154]_  | \new_[2155]_ ;
  assign \new_[6794]_  = \new_[2156]_  | \new_[6793]_ ;
  assign \new_[6797]_  = \new_[2152]_  | \new_[2153]_ ;
  assign \new_[6800]_  = \new_[2150]_  | \new_[2151]_ ;
  assign \new_[6801]_  = \new_[6800]_  | \new_[6797]_ ;
  assign \new_[6802]_  = \new_[6801]_  | \new_[6794]_ ;
  assign \new_[6805]_  = \new_[2148]_  | \new_[2149]_ ;
  assign \new_[6808]_  = \new_[2146]_  | \new_[2147]_ ;
  assign \new_[6809]_  = \new_[6808]_  | \new_[6805]_ ;
  assign \new_[6812]_  = \new_[2144]_  | \new_[2145]_ ;
  assign \new_[6815]_  = \new_[2142]_  | \new_[2143]_ ;
  assign \new_[6816]_  = \new_[6815]_  | \new_[6812]_ ;
  assign \new_[6817]_  = \new_[6816]_  | \new_[6809]_ ;
  assign \new_[6818]_  = \new_[6817]_  | \new_[6802]_ ;
  assign \new_[6819]_  = \new_[6818]_  | \new_[6789]_ ;
  assign \new_[6820]_  = \new_[6819]_  | \new_[6762]_ ;
  assign \new_[6824]_  = \new_[2139]_  | \new_[2140]_ ;
  assign \new_[6825]_  = \new_[2141]_  | \new_[6824]_ ;
  assign \new_[6828]_  = \new_[2137]_  | \new_[2138]_ ;
  assign \new_[6831]_  = \new_[2135]_  | \new_[2136]_ ;
  assign \new_[6832]_  = \new_[6831]_  | \new_[6828]_ ;
  assign \new_[6833]_  = \new_[6832]_  | \new_[6825]_ ;
  assign \new_[6837]_  = \new_[2132]_  | \new_[2133]_ ;
  assign \new_[6838]_  = \new_[2134]_  | \new_[6837]_ ;
  assign \new_[6841]_  = \new_[2130]_  | \new_[2131]_ ;
  assign \new_[6844]_  = \new_[2128]_  | \new_[2129]_ ;
  assign \new_[6845]_  = \new_[6844]_  | \new_[6841]_ ;
  assign \new_[6846]_  = \new_[6845]_  | \new_[6838]_ ;
  assign \new_[6847]_  = \new_[6846]_  | \new_[6833]_ ;
  assign \new_[6851]_  = \new_[2125]_  | \new_[2126]_ ;
  assign \new_[6852]_  = \new_[2127]_  | \new_[6851]_ ;
  assign \new_[6855]_  = \new_[2123]_  | \new_[2124]_ ;
  assign \new_[6858]_  = \new_[2121]_  | \new_[2122]_ ;
  assign \new_[6859]_  = \new_[6858]_  | \new_[6855]_ ;
  assign \new_[6860]_  = \new_[6859]_  | \new_[6852]_ ;
  assign \new_[6863]_  = \new_[2119]_  | \new_[2120]_ ;
  assign \new_[6866]_  = \new_[2117]_  | \new_[2118]_ ;
  assign \new_[6867]_  = \new_[6866]_  | \new_[6863]_ ;
  assign \new_[6870]_  = \new_[2115]_  | \new_[2116]_ ;
  assign \new_[6873]_  = \new_[2113]_  | \new_[2114]_ ;
  assign \new_[6874]_  = \new_[6873]_  | \new_[6870]_ ;
  assign \new_[6875]_  = \new_[6874]_  | \new_[6867]_ ;
  assign \new_[6876]_  = \new_[6875]_  | \new_[6860]_ ;
  assign \new_[6877]_  = \new_[6876]_  | \new_[6847]_ ;
  assign \new_[6881]_  = \new_[2110]_  | \new_[2111]_ ;
  assign \new_[6882]_  = \new_[2112]_  | \new_[6881]_ ;
  assign \new_[6885]_  = \new_[2108]_  | \new_[2109]_ ;
  assign \new_[6888]_  = \new_[2106]_  | \new_[2107]_ ;
  assign \new_[6889]_  = \new_[6888]_  | \new_[6885]_ ;
  assign \new_[6890]_  = \new_[6889]_  | \new_[6882]_ ;
  assign \new_[6894]_  = \new_[2103]_  | \new_[2104]_ ;
  assign \new_[6895]_  = \new_[2105]_  | \new_[6894]_ ;
  assign \new_[6898]_  = \new_[2101]_  | \new_[2102]_ ;
  assign \new_[6901]_  = \new_[2099]_  | \new_[2100]_ ;
  assign \new_[6902]_  = \new_[6901]_  | \new_[6898]_ ;
  assign \new_[6903]_  = \new_[6902]_  | \new_[6895]_ ;
  assign \new_[6904]_  = \new_[6903]_  | \new_[6890]_ ;
  assign \new_[6908]_  = \new_[2096]_  | \new_[2097]_ ;
  assign \new_[6909]_  = \new_[2098]_  | \new_[6908]_ ;
  assign \new_[6912]_  = \new_[2094]_  | \new_[2095]_ ;
  assign \new_[6915]_  = \new_[2092]_  | \new_[2093]_ ;
  assign \new_[6916]_  = \new_[6915]_  | \new_[6912]_ ;
  assign \new_[6917]_  = \new_[6916]_  | \new_[6909]_ ;
  assign \new_[6920]_  = \new_[2090]_  | \new_[2091]_ ;
  assign \new_[6923]_  = \new_[2088]_  | \new_[2089]_ ;
  assign \new_[6924]_  = \new_[6923]_  | \new_[6920]_ ;
  assign \new_[6927]_  = \new_[2086]_  | \new_[2087]_ ;
  assign \new_[6930]_  = \new_[2084]_  | \new_[2085]_ ;
  assign \new_[6931]_  = \new_[6930]_  | \new_[6927]_ ;
  assign \new_[6932]_  = \new_[6931]_  | \new_[6924]_ ;
  assign \new_[6933]_  = \new_[6932]_  | \new_[6917]_ ;
  assign \new_[6934]_  = \new_[6933]_  | \new_[6904]_ ;
  assign \new_[6935]_  = \new_[6934]_  | \new_[6877]_ ;
  assign \new_[6936]_  = \new_[6935]_  | \new_[6820]_ ;
  assign \new_[6937]_  = \new_[6936]_  | \new_[6705]_ ;
  assign \new_[6941]_  = \new_[2081]_  | \new_[2082]_ ;
  assign \new_[6942]_  = \new_[2083]_  | \new_[6941]_ ;
  assign \new_[6945]_  = \new_[2079]_  | \new_[2080]_ ;
  assign \new_[6948]_  = \new_[2077]_  | \new_[2078]_ ;
  assign \new_[6949]_  = \new_[6948]_  | \new_[6945]_ ;
  assign \new_[6950]_  = \new_[6949]_  | \new_[6942]_ ;
  assign \new_[6954]_  = \new_[2074]_  | \new_[2075]_ ;
  assign \new_[6955]_  = \new_[2076]_  | \new_[6954]_ ;
  assign \new_[6958]_  = \new_[2072]_  | \new_[2073]_ ;
  assign \new_[6961]_  = \new_[2070]_  | \new_[2071]_ ;
  assign \new_[6962]_  = \new_[6961]_  | \new_[6958]_ ;
  assign \new_[6963]_  = \new_[6962]_  | \new_[6955]_ ;
  assign \new_[6964]_  = \new_[6963]_  | \new_[6950]_ ;
  assign \new_[6968]_  = \new_[2067]_  | \new_[2068]_ ;
  assign \new_[6969]_  = \new_[2069]_  | \new_[6968]_ ;
  assign \new_[6972]_  = \new_[2065]_  | \new_[2066]_ ;
  assign \new_[6975]_  = \new_[2063]_  | \new_[2064]_ ;
  assign \new_[6976]_  = \new_[6975]_  | \new_[6972]_ ;
  assign \new_[6977]_  = \new_[6976]_  | \new_[6969]_ ;
  assign \new_[6980]_  = \new_[2061]_  | \new_[2062]_ ;
  assign \new_[6983]_  = \new_[2059]_  | \new_[2060]_ ;
  assign \new_[6984]_  = \new_[6983]_  | \new_[6980]_ ;
  assign \new_[6987]_  = \new_[2057]_  | \new_[2058]_ ;
  assign \new_[6990]_  = \new_[2055]_  | \new_[2056]_ ;
  assign \new_[6991]_  = \new_[6990]_  | \new_[6987]_ ;
  assign \new_[6992]_  = \new_[6991]_  | \new_[6984]_ ;
  assign \new_[6993]_  = \new_[6992]_  | \new_[6977]_ ;
  assign \new_[6994]_  = \new_[6993]_  | \new_[6964]_ ;
  assign \new_[6998]_  = \new_[2052]_  | \new_[2053]_ ;
  assign \new_[6999]_  = \new_[2054]_  | \new_[6998]_ ;
  assign \new_[7002]_  = \new_[2050]_  | \new_[2051]_ ;
  assign \new_[7005]_  = \new_[2048]_  | \new_[2049]_ ;
  assign \new_[7006]_  = \new_[7005]_  | \new_[7002]_ ;
  assign \new_[7007]_  = \new_[7006]_  | \new_[6999]_ ;
  assign \new_[7011]_  = \new_[2045]_  | \new_[2046]_ ;
  assign \new_[7012]_  = \new_[2047]_  | \new_[7011]_ ;
  assign \new_[7015]_  = \new_[2043]_  | \new_[2044]_ ;
  assign \new_[7018]_  = \new_[2041]_  | \new_[2042]_ ;
  assign \new_[7019]_  = \new_[7018]_  | \new_[7015]_ ;
  assign \new_[7020]_  = \new_[7019]_  | \new_[7012]_ ;
  assign \new_[7021]_  = \new_[7020]_  | \new_[7007]_ ;
  assign \new_[7025]_  = \new_[2038]_  | \new_[2039]_ ;
  assign \new_[7026]_  = \new_[2040]_  | \new_[7025]_ ;
  assign \new_[7029]_  = \new_[2036]_  | \new_[2037]_ ;
  assign \new_[7032]_  = \new_[2034]_  | \new_[2035]_ ;
  assign \new_[7033]_  = \new_[7032]_  | \new_[7029]_ ;
  assign \new_[7034]_  = \new_[7033]_  | \new_[7026]_ ;
  assign \new_[7037]_  = \new_[2032]_  | \new_[2033]_ ;
  assign \new_[7040]_  = \new_[2030]_  | \new_[2031]_ ;
  assign \new_[7041]_  = \new_[7040]_  | \new_[7037]_ ;
  assign \new_[7044]_  = \new_[2028]_  | \new_[2029]_ ;
  assign \new_[7047]_  = \new_[2026]_  | \new_[2027]_ ;
  assign \new_[7048]_  = \new_[7047]_  | \new_[7044]_ ;
  assign \new_[7049]_  = \new_[7048]_  | \new_[7041]_ ;
  assign \new_[7050]_  = \new_[7049]_  | \new_[7034]_ ;
  assign \new_[7051]_  = \new_[7050]_  | \new_[7021]_ ;
  assign \new_[7052]_  = \new_[7051]_  | \new_[6994]_ ;
  assign \new_[7056]_  = \new_[2023]_  | \new_[2024]_ ;
  assign \new_[7057]_  = \new_[2025]_  | \new_[7056]_ ;
  assign \new_[7060]_  = \new_[2021]_  | \new_[2022]_ ;
  assign \new_[7063]_  = \new_[2019]_  | \new_[2020]_ ;
  assign \new_[7064]_  = \new_[7063]_  | \new_[7060]_ ;
  assign \new_[7065]_  = \new_[7064]_  | \new_[7057]_ ;
  assign \new_[7069]_  = \new_[2016]_  | \new_[2017]_ ;
  assign \new_[7070]_  = \new_[2018]_  | \new_[7069]_ ;
  assign \new_[7073]_  = \new_[2014]_  | \new_[2015]_ ;
  assign \new_[7076]_  = \new_[2012]_  | \new_[2013]_ ;
  assign \new_[7077]_  = \new_[7076]_  | \new_[7073]_ ;
  assign \new_[7078]_  = \new_[7077]_  | \new_[7070]_ ;
  assign \new_[7079]_  = \new_[7078]_  | \new_[7065]_ ;
  assign \new_[7083]_  = \new_[2009]_  | \new_[2010]_ ;
  assign \new_[7084]_  = \new_[2011]_  | \new_[7083]_ ;
  assign \new_[7087]_  = \new_[2007]_  | \new_[2008]_ ;
  assign \new_[7090]_  = \new_[2005]_  | \new_[2006]_ ;
  assign \new_[7091]_  = \new_[7090]_  | \new_[7087]_ ;
  assign \new_[7092]_  = \new_[7091]_  | \new_[7084]_ ;
  assign \new_[7095]_  = \new_[2003]_  | \new_[2004]_ ;
  assign \new_[7098]_  = \new_[2001]_  | \new_[2002]_ ;
  assign \new_[7099]_  = \new_[7098]_  | \new_[7095]_ ;
  assign \new_[7102]_  = \new_[1999]_  | \new_[2000]_ ;
  assign \new_[7105]_  = \new_[1997]_  | \new_[1998]_ ;
  assign \new_[7106]_  = \new_[7105]_  | \new_[7102]_ ;
  assign \new_[7107]_  = \new_[7106]_  | \new_[7099]_ ;
  assign \new_[7108]_  = \new_[7107]_  | \new_[7092]_ ;
  assign \new_[7109]_  = \new_[7108]_  | \new_[7079]_ ;
  assign \new_[7113]_  = \new_[1994]_  | \new_[1995]_ ;
  assign \new_[7114]_  = \new_[1996]_  | \new_[7113]_ ;
  assign \new_[7117]_  = \new_[1992]_  | \new_[1993]_ ;
  assign \new_[7120]_  = \new_[1990]_  | \new_[1991]_ ;
  assign \new_[7121]_  = \new_[7120]_  | \new_[7117]_ ;
  assign \new_[7122]_  = \new_[7121]_  | \new_[7114]_ ;
  assign \new_[7126]_  = \new_[1987]_  | \new_[1988]_ ;
  assign \new_[7127]_  = \new_[1989]_  | \new_[7126]_ ;
  assign \new_[7130]_  = \new_[1985]_  | \new_[1986]_ ;
  assign \new_[7133]_  = \new_[1983]_  | \new_[1984]_ ;
  assign \new_[7134]_  = \new_[7133]_  | \new_[7130]_ ;
  assign \new_[7135]_  = \new_[7134]_  | \new_[7127]_ ;
  assign \new_[7136]_  = \new_[7135]_  | \new_[7122]_ ;
  assign \new_[7140]_  = \new_[1980]_  | \new_[1981]_ ;
  assign \new_[7141]_  = \new_[1982]_  | \new_[7140]_ ;
  assign \new_[7144]_  = \new_[1978]_  | \new_[1979]_ ;
  assign \new_[7147]_  = \new_[1976]_  | \new_[1977]_ ;
  assign \new_[7148]_  = \new_[7147]_  | \new_[7144]_ ;
  assign \new_[7149]_  = \new_[7148]_  | \new_[7141]_ ;
  assign \new_[7152]_  = \new_[1974]_  | \new_[1975]_ ;
  assign \new_[7155]_  = \new_[1972]_  | \new_[1973]_ ;
  assign \new_[7156]_  = \new_[7155]_  | \new_[7152]_ ;
  assign \new_[7159]_  = \new_[1970]_  | \new_[1971]_ ;
  assign \new_[7162]_  = \new_[1968]_  | \new_[1969]_ ;
  assign \new_[7163]_  = \new_[7162]_  | \new_[7159]_ ;
  assign \new_[7164]_  = \new_[7163]_  | \new_[7156]_ ;
  assign \new_[7165]_  = \new_[7164]_  | \new_[7149]_ ;
  assign \new_[7166]_  = \new_[7165]_  | \new_[7136]_ ;
  assign \new_[7167]_  = \new_[7166]_  | \new_[7109]_ ;
  assign \new_[7168]_  = \new_[7167]_  | \new_[7052]_ ;
  assign \new_[7172]_  = \new_[1965]_  | \new_[1966]_ ;
  assign \new_[7173]_  = \new_[1967]_  | \new_[7172]_ ;
  assign \new_[7176]_  = \new_[1963]_  | \new_[1964]_ ;
  assign \new_[7179]_  = \new_[1961]_  | \new_[1962]_ ;
  assign \new_[7180]_  = \new_[7179]_  | \new_[7176]_ ;
  assign \new_[7181]_  = \new_[7180]_  | \new_[7173]_ ;
  assign \new_[7185]_  = \new_[1958]_  | \new_[1959]_ ;
  assign \new_[7186]_  = \new_[1960]_  | \new_[7185]_ ;
  assign \new_[7189]_  = \new_[1956]_  | \new_[1957]_ ;
  assign \new_[7192]_  = \new_[1954]_  | \new_[1955]_ ;
  assign \new_[7193]_  = \new_[7192]_  | \new_[7189]_ ;
  assign \new_[7194]_  = \new_[7193]_  | \new_[7186]_ ;
  assign \new_[7195]_  = \new_[7194]_  | \new_[7181]_ ;
  assign \new_[7199]_  = \new_[1951]_  | \new_[1952]_ ;
  assign \new_[7200]_  = \new_[1953]_  | \new_[7199]_ ;
  assign \new_[7203]_  = \new_[1949]_  | \new_[1950]_ ;
  assign \new_[7206]_  = \new_[1947]_  | \new_[1948]_ ;
  assign \new_[7207]_  = \new_[7206]_  | \new_[7203]_ ;
  assign \new_[7208]_  = \new_[7207]_  | \new_[7200]_ ;
  assign \new_[7211]_  = \new_[1945]_  | \new_[1946]_ ;
  assign \new_[7214]_  = \new_[1943]_  | \new_[1944]_ ;
  assign \new_[7215]_  = \new_[7214]_  | \new_[7211]_ ;
  assign \new_[7218]_  = \new_[1941]_  | \new_[1942]_ ;
  assign \new_[7221]_  = \new_[1939]_  | \new_[1940]_ ;
  assign \new_[7222]_  = \new_[7221]_  | \new_[7218]_ ;
  assign \new_[7223]_  = \new_[7222]_  | \new_[7215]_ ;
  assign \new_[7224]_  = \new_[7223]_  | \new_[7208]_ ;
  assign \new_[7225]_  = \new_[7224]_  | \new_[7195]_ ;
  assign \new_[7229]_  = \new_[1936]_  | \new_[1937]_ ;
  assign \new_[7230]_  = \new_[1938]_  | \new_[7229]_ ;
  assign \new_[7233]_  = \new_[1934]_  | \new_[1935]_ ;
  assign \new_[7236]_  = \new_[1932]_  | \new_[1933]_ ;
  assign \new_[7237]_  = \new_[7236]_  | \new_[7233]_ ;
  assign \new_[7238]_  = \new_[7237]_  | \new_[7230]_ ;
  assign \new_[7242]_  = \new_[1929]_  | \new_[1930]_ ;
  assign \new_[7243]_  = \new_[1931]_  | \new_[7242]_ ;
  assign \new_[7246]_  = \new_[1927]_  | \new_[1928]_ ;
  assign \new_[7249]_  = \new_[1925]_  | \new_[1926]_ ;
  assign \new_[7250]_  = \new_[7249]_  | \new_[7246]_ ;
  assign \new_[7251]_  = \new_[7250]_  | \new_[7243]_ ;
  assign \new_[7252]_  = \new_[7251]_  | \new_[7238]_ ;
  assign \new_[7256]_  = \new_[1922]_  | \new_[1923]_ ;
  assign \new_[7257]_  = \new_[1924]_  | \new_[7256]_ ;
  assign \new_[7260]_  = \new_[1920]_  | \new_[1921]_ ;
  assign \new_[7263]_  = \new_[1918]_  | \new_[1919]_ ;
  assign \new_[7264]_  = \new_[7263]_  | \new_[7260]_ ;
  assign \new_[7265]_  = \new_[7264]_  | \new_[7257]_ ;
  assign \new_[7268]_  = \new_[1916]_  | \new_[1917]_ ;
  assign \new_[7271]_  = \new_[1914]_  | \new_[1915]_ ;
  assign \new_[7272]_  = \new_[7271]_  | \new_[7268]_ ;
  assign \new_[7275]_  = \new_[1912]_  | \new_[1913]_ ;
  assign \new_[7278]_  = \new_[1910]_  | \new_[1911]_ ;
  assign \new_[7279]_  = \new_[7278]_  | \new_[7275]_ ;
  assign \new_[7280]_  = \new_[7279]_  | \new_[7272]_ ;
  assign \new_[7281]_  = \new_[7280]_  | \new_[7265]_ ;
  assign \new_[7282]_  = \new_[7281]_  | \new_[7252]_ ;
  assign \new_[7283]_  = \new_[7282]_  | \new_[7225]_ ;
  assign \new_[7287]_  = \new_[1907]_  | \new_[1908]_ ;
  assign \new_[7288]_  = \new_[1909]_  | \new_[7287]_ ;
  assign \new_[7291]_  = \new_[1905]_  | \new_[1906]_ ;
  assign \new_[7294]_  = \new_[1903]_  | \new_[1904]_ ;
  assign \new_[7295]_  = \new_[7294]_  | \new_[7291]_ ;
  assign \new_[7296]_  = \new_[7295]_  | \new_[7288]_ ;
  assign \new_[7300]_  = \new_[1900]_  | \new_[1901]_ ;
  assign \new_[7301]_  = \new_[1902]_  | \new_[7300]_ ;
  assign \new_[7304]_  = \new_[1898]_  | \new_[1899]_ ;
  assign \new_[7307]_  = \new_[1896]_  | \new_[1897]_ ;
  assign \new_[7308]_  = \new_[7307]_  | \new_[7304]_ ;
  assign \new_[7309]_  = \new_[7308]_  | \new_[7301]_ ;
  assign \new_[7310]_  = \new_[7309]_  | \new_[7296]_ ;
  assign \new_[7314]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[7315]_  = \new_[1895]_  | \new_[7314]_ ;
  assign \new_[7318]_  = \new_[1891]_  | \new_[1892]_ ;
  assign \new_[7321]_  = \new_[1889]_  | \new_[1890]_ ;
  assign \new_[7322]_  = \new_[7321]_  | \new_[7318]_ ;
  assign \new_[7323]_  = \new_[7322]_  | \new_[7315]_ ;
  assign \new_[7326]_  = \new_[1887]_  | \new_[1888]_ ;
  assign \new_[7329]_  = \new_[1885]_  | \new_[1886]_ ;
  assign \new_[7330]_  = \new_[7329]_  | \new_[7326]_ ;
  assign \new_[7333]_  = \new_[1883]_  | \new_[1884]_ ;
  assign \new_[7336]_  = \new_[1881]_  | \new_[1882]_ ;
  assign \new_[7337]_  = \new_[7336]_  | \new_[7333]_ ;
  assign \new_[7338]_  = \new_[7337]_  | \new_[7330]_ ;
  assign \new_[7339]_  = \new_[7338]_  | \new_[7323]_ ;
  assign \new_[7340]_  = \new_[7339]_  | \new_[7310]_ ;
  assign \new_[7344]_  = \new_[1878]_  | \new_[1879]_ ;
  assign \new_[7345]_  = \new_[1880]_  | \new_[7344]_ ;
  assign \new_[7348]_  = \new_[1876]_  | \new_[1877]_ ;
  assign \new_[7351]_  = \new_[1874]_  | \new_[1875]_ ;
  assign \new_[7352]_  = \new_[7351]_  | \new_[7348]_ ;
  assign \new_[7353]_  = \new_[7352]_  | \new_[7345]_ ;
  assign \new_[7357]_  = \new_[1871]_  | \new_[1872]_ ;
  assign \new_[7358]_  = \new_[1873]_  | \new_[7357]_ ;
  assign \new_[7361]_  = \new_[1869]_  | \new_[1870]_ ;
  assign \new_[7364]_  = \new_[1867]_  | \new_[1868]_ ;
  assign \new_[7365]_  = \new_[7364]_  | \new_[7361]_ ;
  assign \new_[7366]_  = \new_[7365]_  | \new_[7358]_ ;
  assign \new_[7367]_  = \new_[7366]_  | \new_[7353]_ ;
  assign \new_[7371]_  = \new_[1864]_  | \new_[1865]_ ;
  assign \new_[7372]_  = \new_[1866]_  | \new_[7371]_ ;
  assign \new_[7375]_  = \new_[1862]_  | \new_[1863]_ ;
  assign \new_[7378]_  = \new_[1860]_  | \new_[1861]_ ;
  assign \new_[7379]_  = \new_[7378]_  | \new_[7375]_ ;
  assign \new_[7380]_  = \new_[7379]_  | \new_[7372]_ ;
  assign \new_[7383]_  = \new_[1858]_  | \new_[1859]_ ;
  assign \new_[7386]_  = \new_[1856]_  | \new_[1857]_ ;
  assign \new_[7387]_  = \new_[7386]_  | \new_[7383]_ ;
  assign \new_[7390]_  = \new_[1854]_  | \new_[1855]_ ;
  assign \new_[7393]_  = \new_[1852]_  | \new_[1853]_ ;
  assign \new_[7394]_  = \new_[7393]_  | \new_[7390]_ ;
  assign \new_[7395]_  = \new_[7394]_  | \new_[7387]_ ;
  assign \new_[7396]_  = \new_[7395]_  | \new_[7380]_ ;
  assign \new_[7397]_  = \new_[7396]_  | \new_[7367]_ ;
  assign \new_[7398]_  = \new_[7397]_  | \new_[7340]_ ;
  assign \new_[7399]_  = \new_[7398]_  | \new_[7283]_ ;
  assign \new_[7400]_  = \new_[7399]_  | \new_[7168]_ ;
  assign \new_[7401]_  = \new_[7400]_  | \new_[6937]_ ;
  assign \new_[7402]_  = \new_[7401]_  | \new_[6476]_ ;
  assign \new_[7403]_  = \new_[7402]_  | \new_[5551]_ ;
  assign \new_[7407]_  = \new_[1849]_  | \new_[1850]_ ;
  assign \new_[7408]_  = \new_[1851]_  | \new_[7407]_ ;
  assign \new_[7411]_  = \new_[1847]_  | \new_[1848]_ ;
  assign \new_[7414]_  = \new_[1845]_  | \new_[1846]_ ;
  assign \new_[7415]_  = \new_[7414]_  | \new_[7411]_ ;
  assign \new_[7416]_  = \new_[7415]_  | \new_[7408]_ ;
  assign \new_[7420]_  = \new_[1842]_  | \new_[1843]_ ;
  assign \new_[7421]_  = \new_[1844]_  | \new_[7420]_ ;
  assign \new_[7424]_  = \new_[1840]_  | \new_[1841]_ ;
  assign \new_[7427]_  = \new_[1838]_  | \new_[1839]_ ;
  assign \new_[7428]_  = \new_[7427]_  | \new_[7424]_ ;
  assign \new_[7429]_  = \new_[7428]_  | \new_[7421]_ ;
  assign \new_[7430]_  = \new_[7429]_  | \new_[7416]_ ;
  assign \new_[7434]_  = \new_[1835]_  | \new_[1836]_ ;
  assign \new_[7435]_  = \new_[1837]_  | \new_[7434]_ ;
  assign \new_[7438]_  = \new_[1833]_  | \new_[1834]_ ;
  assign \new_[7441]_  = \new_[1831]_  | \new_[1832]_ ;
  assign \new_[7442]_  = \new_[7441]_  | \new_[7438]_ ;
  assign \new_[7443]_  = \new_[7442]_  | \new_[7435]_ ;
  assign \new_[7447]_  = \new_[1828]_  | \new_[1829]_ ;
  assign \new_[7448]_  = \new_[1830]_  | \new_[7447]_ ;
  assign \new_[7451]_  = \new_[1826]_  | \new_[1827]_ ;
  assign \new_[7454]_  = \new_[1824]_  | \new_[1825]_ ;
  assign \new_[7455]_  = \new_[7454]_  | \new_[7451]_ ;
  assign \new_[7456]_  = \new_[7455]_  | \new_[7448]_ ;
  assign \new_[7457]_  = \new_[7456]_  | \new_[7443]_ ;
  assign \new_[7458]_  = \new_[7457]_  | \new_[7430]_ ;
  assign \new_[7462]_  = \new_[1821]_  | \new_[1822]_ ;
  assign \new_[7463]_  = \new_[1823]_  | \new_[7462]_ ;
  assign \new_[7466]_  = \new_[1819]_  | \new_[1820]_ ;
  assign \new_[7469]_  = \new_[1817]_  | \new_[1818]_ ;
  assign \new_[7470]_  = \new_[7469]_  | \new_[7466]_ ;
  assign \new_[7471]_  = \new_[7470]_  | \new_[7463]_ ;
  assign \new_[7475]_  = \new_[1814]_  | \new_[1815]_ ;
  assign \new_[7476]_  = \new_[1816]_  | \new_[7475]_ ;
  assign \new_[7479]_  = \new_[1812]_  | \new_[1813]_ ;
  assign \new_[7482]_  = \new_[1810]_  | \new_[1811]_ ;
  assign \new_[7483]_  = \new_[7482]_  | \new_[7479]_ ;
  assign \new_[7484]_  = \new_[7483]_  | \new_[7476]_ ;
  assign \new_[7485]_  = \new_[7484]_  | \new_[7471]_ ;
  assign \new_[7489]_  = \new_[1807]_  | \new_[1808]_ ;
  assign \new_[7490]_  = \new_[1809]_  | \new_[7489]_ ;
  assign \new_[7493]_  = \new_[1805]_  | \new_[1806]_ ;
  assign \new_[7496]_  = \new_[1803]_  | \new_[1804]_ ;
  assign \new_[7497]_  = \new_[7496]_  | \new_[7493]_ ;
  assign \new_[7498]_  = \new_[7497]_  | \new_[7490]_ ;
  assign \new_[7501]_  = \new_[1801]_  | \new_[1802]_ ;
  assign \new_[7504]_  = \new_[1799]_  | \new_[1800]_ ;
  assign \new_[7505]_  = \new_[7504]_  | \new_[7501]_ ;
  assign \new_[7508]_  = \new_[1797]_  | \new_[1798]_ ;
  assign \new_[7511]_  = \new_[1795]_  | \new_[1796]_ ;
  assign \new_[7512]_  = \new_[7511]_  | \new_[7508]_ ;
  assign \new_[7513]_  = \new_[7512]_  | \new_[7505]_ ;
  assign \new_[7514]_  = \new_[7513]_  | \new_[7498]_ ;
  assign \new_[7515]_  = \new_[7514]_  | \new_[7485]_ ;
  assign \new_[7516]_  = \new_[7515]_  | \new_[7458]_ ;
  assign \new_[7520]_  = \new_[1792]_  | \new_[1793]_ ;
  assign \new_[7521]_  = \new_[1794]_  | \new_[7520]_ ;
  assign \new_[7524]_  = \new_[1790]_  | \new_[1791]_ ;
  assign \new_[7527]_  = \new_[1788]_  | \new_[1789]_ ;
  assign \new_[7528]_  = \new_[7527]_  | \new_[7524]_ ;
  assign \new_[7529]_  = \new_[7528]_  | \new_[7521]_ ;
  assign \new_[7533]_  = \new_[1785]_  | \new_[1786]_ ;
  assign \new_[7534]_  = \new_[1787]_  | \new_[7533]_ ;
  assign \new_[7537]_  = \new_[1783]_  | \new_[1784]_ ;
  assign \new_[7540]_  = \new_[1781]_  | \new_[1782]_ ;
  assign \new_[7541]_  = \new_[7540]_  | \new_[7537]_ ;
  assign \new_[7542]_  = \new_[7541]_  | \new_[7534]_ ;
  assign \new_[7543]_  = \new_[7542]_  | \new_[7529]_ ;
  assign \new_[7547]_  = \new_[1778]_  | \new_[1779]_ ;
  assign \new_[7548]_  = \new_[1780]_  | \new_[7547]_ ;
  assign \new_[7551]_  = \new_[1776]_  | \new_[1777]_ ;
  assign \new_[7554]_  = \new_[1774]_  | \new_[1775]_ ;
  assign \new_[7555]_  = \new_[7554]_  | \new_[7551]_ ;
  assign \new_[7556]_  = \new_[7555]_  | \new_[7548]_ ;
  assign \new_[7559]_  = \new_[1772]_  | \new_[1773]_ ;
  assign \new_[7562]_  = \new_[1770]_  | \new_[1771]_ ;
  assign \new_[7563]_  = \new_[7562]_  | \new_[7559]_ ;
  assign \new_[7566]_  = \new_[1768]_  | \new_[1769]_ ;
  assign \new_[7569]_  = \new_[1766]_  | \new_[1767]_ ;
  assign \new_[7570]_  = \new_[7569]_  | \new_[7566]_ ;
  assign \new_[7571]_  = \new_[7570]_  | \new_[7563]_ ;
  assign \new_[7572]_  = \new_[7571]_  | \new_[7556]_ ;
  assign \new_[7573]_  = \new_[7572]_  | \new_[7543]_ ;
  assign \new_[7577]_  = \new_[1763]_  | \new_[1764]_ ;
  assign \new_[7578]_  = \new_[1765]_  | \new_[7577]_ ;
  assign \new_[7581]_  = \new_[1761]_  | \new_[1762]_ ;
  assign \new_[7584]_  = \new_[1759]_  | \new_[1760]_ ;
  assign \new_[7585]_  = \new_[7584]_  | \new_[7581]_ ;
  assign \new_[7586]_  = \new_[7585]_  | \new_[7578]_ ;
  assign \new_[7590]_  = \new_[1756]_  | \new_[1757]_ ;
  assign \new_[7591]_  = \new_[1758]_  | \new_[7590]_ ;
  assign \new_[7594]_  = \new_[1754]_  | \new_[1755]_ ;
  assign \new_[7597]_  = \new_[1752]_  | \new_[1753]_ ;
  assign \new_[7598]_  = \new_[7597]_  | \new_[7594]_ ;
  assign \new_[7599]_  = \new_[7598]_  | \new_[7591]_ ;
  assign \new_[7600]_  = \new_[7599]_  | \new_[7586]_ ;
  assign \new_[7604]_  = \new_[1749]_  | \new_[1750]_ ;
  assign \new_[7605]_  = \new_[1751]_  | \new_[7604]_ ;
  assign \new_[7608]_  = \new_[1747]_  | \new_[1748]_ ;
  assign \new_[7611]_  = \new_[1745]_  | \new_[1746]_ ;
  assign \new_[7612]_  = \new_[7611]_  | \new_[7608]_ ;
  assign \new_[7613]_  = \new_[7612]_  | \new_[7605]_ ;
  assign \new_[7616]_  = \new_[1743]_  | \new_[1744]_ ;
  assign \new_[7619]_  = \new_[1741]_  | \new_[1742]_ ;
  assign \new_[7620]_  = \new_[7619]_  | \new_[7616]_ ;
  assign \new_[7623]_  = \new_[1739]_  | \new_[1740]_ ;
  assign \new_[7626]_  = \new_[1737]_  | \new_[1738]_ ;
  assign \new_[7627]_  = \new_[7626]_  | \new_[7623]_ ;
  assign \new_[7628]_  = \new_[7627]_  | \new_[7620]_ ;
  assign \new_[7629]_  = \new_[7628]_  | \new_[7613]_ ;
  assign \new_[7630]_  = \new_[7629]_  | \new_[7600]_ ;
  assign \new_[7631]_  = \new_[7630]_  | \new_[7573]_ ;
  assign \new_[7632]_  = \new_[7631]_  | \new_[7516]_ ;
  assign \new_[7636]_  = \new_[1734]_  | \new_[1735]_ ;
  assign \new_[7637]_  = \new_[1736]_  | \new_[7636]_ ;
  assign \new_[7640]_  = \new_[1732]_  | \new_[1733]_ ;
  assign \new_[7643]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[7644]_  = \new_[7643]_  | \new_[7640]_ ;
  assign \new_[7645]_  = \new_[7644]_  | \new_[7637]_ ;
  assign \new_[7649]_  = \new_[1727]_  | \new_[1728]_ ;
  assign \new_[7650]_  = \new_[1729]_  | \new_[7649]_ ;
  assign \new_[7653]_  = \new_[1725]_  | \new_[1726]_ ;
  assign \new_[7656]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[7657]_  = \new_[7656]_  | \new_[7653]_ ;
  assign \new_[7658]_  = \new_[7657]_  | \new_[7650]_ ;
  assign \new_[7659]_  = \new_[7658]_  | \new_[7645]_ ;
  assign \new_[7663]_  = \new_[1720]_  | \new_[1721]_ ;
  assign \new_[7664]_  = \new_[1722]_  | \new_[7663]_ ;
  assign \new_[7667]_  = \new_[1718]_  | \new_[1719]_ ;
  assign \new_[7670]_  = \new_[1716]_  | \new_[1717]_ ;
  assign \new_[7671]_  = \new_[7670]_  | \new_[7667]_ ;
  assign \new_[7672]_  = \new_[7671]_  | \new_[7664]_ ;
  assign \new_[7675]_  = \new_[1714]_  | \new_[1715]_ ;
  assign \new_[7678]_  = \new_[1712]_  | \new_[1713]_ ;
  assign \new_[7679]_  = \new_[7678]_  | \new_[7675]_ ;
  assign \new_[7682]_  = \new_[1710]_  | \new_[1711]_ ;
  assign \new_[7685]_  = \new_[1708]_  | \new_[1709]_ ;
  assign \new_[7686]_  = \new_[7685]_  | \new_[7682]_ ;
  assign \new_[7687]_  = \new_[7686]_  | \new_[7679]_ ;
  assign \new_[7688]_  = \new_[7687]_  | \new_[7672]_ ;
  assign \new_[7689]_  = \new_[7688]_  | \new_[7659]_ ;
  assign \new_[7693]_  = \new_[1705]_  | \new_[1706]_ ;
  assign \new_[7694]_  = \new_[1707]_  | \new_[7693]_ ;
  assign \new_[7697]_  = \new_[1703]_  | \new_[1704]_ ;
  assign \new_[7700]_  = \new_[1701]_  | \new_[1702]_ ;
  assign \new_[7701]_  = \new_[7700]_  | \new_[7697]_ ;
  assign \new_[7702]_  = \new_[7701]_  | \new_[7694]_ ;
  assign \new_[7706]_  = \new_[1698]_  | \new_[1699]_ ;
  assign \new_[7707]_  = \new_[1700]_  | \new_[7706]_ ;
  assign \new_[7710]_  = \new_[1696]_  | \new_[1697]_ ;
  assign \new_[7713]_  = \new_[1694]_  | \new_[1695]_ ;
  assign \new_[7714]_  = \new_[7713]_  | \new_[7710]_ ;
  assign \new_[7715]_  = \new_[7714]_  | \new_[7707]_ ;
  assign \new_[7716]_  = \new_[7715]_  | \new_[7702]_ ;
  assign \new_[7720]_  = \new_[1691]_  | \new_[1692]_ ;
  assign \new_[7721]_  = \new_[1693]_  | \new_[7720]_ ;
  assign \new_[7724]_  = \new_[1689]_  | \new_[1690]_ ;
  assign \new_[7727]_  = \new_[1687]_  | \new_[1688]_ ;
  assign \new_[7728]_  = \new_[7727]_  | \new_[7724]_ ;
  assign \new_[7729]_  = \new_[7728]_  | \new_[7721]_ ;
  assign \new_[7732]_  = \new_[1685]_  | \new_[1686]_ ;
  assign \new_[7735]_  = \new_[1683]_  | \new_[1684]_ ;
  assign \new_[7736]_  = \new_[7735]_  | \new_[7732]_ ;
  assign \new_[7739]_  = \new_[1681]_  | \new_[1682]_ ;
  assign \new_[7742]_  = \new_[1679]_  | \new_[1680]_ ;
  assign \new_[7743]_  = \new_[7742]_  | \new_[7739]_ ;
  assign \new_[7744]_  = \new_[7743]_  | \new_[7736]_ ;
  assign \new_[7745]_  = \new_[7744]_  | \new_[7729]_ ;
  assign \new_[7746]_  = \new_[7745]_  | \new_[7716]_ ;
  assign \new_[7747]_  = \new_[7746]_  | \new_[7689]_ ;
  assign \new_[7751]_  = \new_[1676]_  | \new_[1677]_ ;
  assign \new_[7752]_  = \new_[1678]_  | \new_[7751]_ ;
  assign \new_[7755]_  = \new_[1674]_  | \new_[1675]_ ;
  assign \new_[7758]_  = \new_[1672]_  | \new_[1673]_ ;
  assign \new_[7759]_  = \new_[7758]_  | \new_[7755]_ ;
  assign \new_[7760]_  = \new_[7759]_  | \new_[7752]_ ;
  assign \new_[7764]_  = \new_[1669]_  | \new_[1670]_ ;
  assign \new_[7765]_  = \new_[1671]_  | \new_[7764]_ ;
  assign \new_[7768]_  = \new_[1667]_  | \new_[1668]_ ;
  assign \new_[7771]_  = \new_[1665]_  | \new_[1666]_ ;
  assign \new_[7772]_  = \new_[7771]_  | \new_[7768]_ ;
  assign \new_[7773]_  = \new_[7772]_  | \new_[7765]_ ;
  assign \new_[7774]_  = \new_[7773]_  | \new_[7760]_ ;
  assign \new_[7778]_  = \new_[1662]_  | \new_[1663]_ ;
  assign \new_[7779]_  = \new_[1664]_  | \new_[7778]_ ;
  assign \new_[7782]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[7785]_  = \new_[1658]_  | \new_[1659]_ ;
  assign \new_[7786]_  = \new_[7785]_  | \new_[7782]_ ;
  assign \new_[7787]_  = \new_[7786]_  | \new_[7779]_ ;
  assign \new_[7790]_  = \new_[1656]_  | \new_[1657]_ ;
  assign \new_[7793]_  = \new_[1654]_  | \new_[1655]_ ;
  assign \new_[7794]_  = \new_[7793]_  | \new_[7790]_ ;
  assign \new_[7797]_  = \new_[1652]_  | \new_[1653]_ ;
  assign \new_[7800]_  = \new_[1650]_  | \new_[1651]_ ;
  assign \new_[7801]_  = \new_[7800]_  | \new_[7797]_ ;
  assign \new_[7802]_  = \new_[7801]_  | \new_[7794]_ ;
  assign \new_[7803]_  = \new_[7802]_  | \new_[7787]_ ;
  assign \new_[7804]_  = \new_[7803]_  | \new_[7774]_ ;
  assign \new_[7808]_  = \new_[1647]_  | \new_[1648]_ ;
  assign \new_[7809]_  = \new_[1649]_  | \new_[7808]_ ;
  assign \new_[7812]_  = \new_[1645]_  | \new_[1646]_ ;
  assign \new_[7815]_  = \new_[1643]_  | \new_[1644]_ ;
  assign \new_[7816]_  = \new_[7815]_  | \new_[7812]_ ;
  assign \new_[7817]_  = \new_[7816]_  | \new_[7809]_ ;
  assign \new_[7821]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[7822]_  = \new_[1642]_  | \new_[7821]_ ;
  assign \new_[7825]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[7828]_  = \new_[1636]_  | \new_[1637]_ ;
  assign \new_[7829]_  = \new_[7828]_  | \new_[7825]_ ;
  assign \new_[7830]_  = \new_[7829]_  | \new_[7822]_ ;
  assign \new_[7831]_  = \new_[7830]_  | \new_[7817]_ ;
  assign \new_[7835]_  = \new_[1633]_  | \new_[1634]_ ;
  assign \new_[7836]_  = \new_[1635]_  | \new_[7835]_ ;
  assign \new_[7839]_  = \new_[1631]_  | \new_[1632]_ ;
  assign \new_[7842]_  = \new_[1629]_  | \new_[1630]_ ;
  assign \new_[7843]_  = \new_[7842]_  | \new_[7839]_ ;
  assign \new_[7844]_  = \new_[7843]_  | \new_[7836]_ ;
  assign \new_[7847]_  = \new_[1627]_  | \new_[1628]_ ;
  assign \new_[7850]_  = \new_[1625]_  | \new_[1626]_ ;
  assign \new_[7851]_  = \new_[7850]_  | \new_[7847]_ ;
  assign \new_[7854]_  = \new_[1623]_  | \new_[1624]_ ;
  assign \new_[7857]_  = \new_[1621]_  | \new_[1622]_ ;
  assign \new_[7858]_  = \new_[7857]_  | \new_[7854]_ ;
  assign \new_[7859]_  = \new_[7858]_  | \new_[7851]_ ;
  assign \new_[7860]_  = \new_[7859]_  | \new_[7844]_ ;
  assign \new_[7861]_  = \new_[7860]_  | \new_[7831]_ ;
  assign \new_[7862]_  = \new_[7861]_  | \new_[7804]_ ;
  assign \new_[7863]_  = \new_[7862]_  | \new_[7747]_ ;
  assign \new_[7864]_  = \new_[7863]_  | \new_[7632]_ ;
  assign \new_[7868]_  = \new_[1618]_  | \new_[1619]_ ;
  assign \new_[7869]_  = \new_[1620]_  | \new_[7868]_ ;
  assign \new_[7872]_  = \new_[1616]_  | \new_[1617]_ ;
  assign \new_[7875]_  = \new_[1614]_  | \new_[1615]_ ;
  assign \new_[7876]_  = \new_[7875]_  | \new_[7872]_ ;
  assign \new_[7877]_  = \new_[7876]_  | \new_[7869]_ ;
  assign \new_[7881]_  = \new_[1611]_  | \new_[1612]_ ;
  assign \new_[7882]_  = \new_[1613]_  | \new_[7881]_ ;
  assign \new_[7885]_  = \new_[1609]_  | \new_[1610]_ ;
  assign \new_[7888]_  = \new_[1607]_  | \new_[1608]_ ;
  assign \new_[7889]_  = \new_[7888]_  | \new_[7885]_ ;
  assign \new_[7890]_  = \new_[7889]_  | \new_[7882]_ ;
  assign \new_[7891]_  = \new_[7890]_  | \new_[7877]_ ;
  assign \new_[7895]_  = \new_[1604]_  | \new_[1605]_ ;
  assign \new_[7896]_  = \new_[1606]_  | \new_[7895]_ ;
  assign \new_[7899]_  = \new_[1602]_  | \new_[1603]_ ;
  assign \new_[7902]_  = \new_[1600]_  | \new_[1601]_ ;
  assign \new_[7903]_  = \new_[7902]_  | \new_[7899]_ ;
  assign \new_[7904]_  = \new_[7903]_  | \new_[7896]_ ;
  assign \new_[7908]_  = \new_[1597]_  | \new_[1598]_ ;
  assign \new_[7909]_  = \new_[1599]_  | \new_[7908]_ ;
  assign \new_[7912]_  = \new_[1595]_  | \new_[1596]_ ;
  assign \new_[7915]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[7916]_  = \new_[7915]_  | \new_[7912]_ ;
  assign \new_[7917]_  = \new_[7916]_  | \new_[7909]_ ;
  assign \new_[7918]_  = \new_[7917]_  | \new_[7904]_ ;
  assign \new_[7919]_  = \new_[7918]_  | \new_[7891]_ ;
  assign \new_[7923]_  = \new_[1590]_  | \new_[1591]_ ;
  assign \new_[7924]_  = \new_[1592]_  | \new_[7923]_ ;
  assign \new_[7927]_  = \new_[1588]_  | \new_[1589]_ ;
  assign \new_[7930]_  = \new_[1586]_  | \new_[1587]_ ;
  assign \new_[7931]_  = \new_[7930]_  | \new_[7927]_ ;
  assign \new_[7932]_  = \new_[7931]_  | \new_[7924]_ ;
  assign \new_[7936]_  = \new_[1583]_  | \new_[1584]_ ;
  assign \new_[7937]_  = \new_[1585]_  | \new_[7936]_ ;
  assign \new_[7940]_  = \new_[1581]_  | \new_[1582]_ ;
  assign \new_[7943]_  = \new_[1579]_  | \new_[1580]_ ;
  assign \new_[7944]_  = \new_[7943]_  | \new_[7940]_ ;
  assign \new_[7945]_  = \new_[7944]_  | \new_[7937]_ ;
  assign \new_[7946]_  = \new_[7945]_  | \new_[7932]_ ;
  assign \new_[7950]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[7951]_  = \new_[1578]_  | \new_[7950]_ ;
  assign \new_[7954]_  = \new_[1574]_  | \new_[1575]_ ;
  assign \new_[7957]_  = \new_[1572]_  | \new_[1573]_ ;
  assign \new_[7958]_  = \new_[7957]_  | \new_[7954]_ ;
  assign \new_[7959]_  = \new_[7958]_  | \new_[7951]_ ;
  assign \new_[7962]_  = \new_[1570]_  | \new_[1571]_ ;
  assign \new_[7965]_  = \new_[1568]_  | \new_[1569]_ ;
  assign \new_[7966]_  = \new_[7965]_  | \new_[7962]_ ;
  assign \new_[7969]_  = \new_[1566]_  | \new_[1567]_ ;
  assign \new_[7972]_  = \new_[1564]_  | \new_[1565]_ ;
  assign \new_[7973]_  = \new_[7972]_  | \new_[7969]_ ;
  assign \new_[7974]_  = \new_[7973]_  | \new_[7966]_ ;
  assign \new_[7975]_  = \new_[7974]_  | \new_[7959]_ ;
  assign \new_[7976]_  = \new_[7975]_  | \new_[7946]_ ;
  assign \new_[7977]_  = \new_[7976]_  | \new_[7919]_ ;
  assign \new_[7981]_  = \new_[1561]_  | \new_[1562]_ ;
  assign \new_[7982]_  = \new_[1563]_  | \new_[7981]_ ;
  assign \new_[7985]_  = \new_[1559]_  | \new_[1560]_ ;
  assign \new_[7988]_  = \new_[1557]_  | \new_[1558]_ ;
  assign \new_[7989]_  = \new_[7988]_  | \new_[7985]_ ;
  assign \new_[7990]_  = \new_[7989]_  | \new_[7982]_ ;
  assign \new_[7994]_  = \new_[1554]_  | \new_[1555]_ ;
  assign \new_[7995]_  = \new_[1556]_  | \new_[7994]_ ;
  assign \new_[7998]_  = \new_[1552]_  | \new_[1553]_ ;
  assign \new_[8001]_  = \new_[1550]_  | \new_[1551]_ ;
  assign \new_[8002]_  = \new_[8001]_  | \new_[7998]_ ;
  assign \new_[8003]_  = \new_[8002]_  | \new_[7995]_ ;
  assign \new_[8004]_  = \new_[8003]_  | \new_[7990]_ ;
  assign \new_[8008]_  = \new_[1547]_  | \new_[1548]_ ;
  assign \new_[8009]_  = \new_[1549]_  | \new_[8008]_ ;
  assign \new_[8012]_  = \new_[1545]_  | \new_[1546]_ ;
  assign \new_[8015]_  = \new_[1543]_  | \new_[1544]_ ;
  assign \new_[8016]_  = \new_[8015]_  | \new_[8012]_ ;
  assign \new_[8017]_  = \new_[8016]_  | \new_[8009]_ ;
  assign \new_[8020]_  = \new_[1541]_  | \new_[1542]_ ;
  assign \new_[8023]_  = \new_[1539]_  | \new_[1540]_ ;
  assign \new_[8024]_  = \new_[8023]_  | \new_[8020]_ ;
  assign \new_[8027]_  = \new_[1537]_  | \new_[1538]_ ;
  assign \new_[8030]_  = \new_[1535]_  | \new_[1536]_ ;
  assign \new_[8031]_  = \new_[8030]_  | \new_[8027]_ ;
  assign \new_[8032]_  = \new_[8031]_  | \new_[8024]_ ;
  assign \new_[8033]_  = \new_[8032]_  | \new_[8017]_ ;
  assign \new_[8034]_  = \new_[8033]_  | \new_[8004]_ ;
  assign \new_[8038]_  = \new_[1532]_  | \new_[1533]_ ;
  assign \new_[8039]_  = \new_[1534]_  | \new_[8038]_ ;
  assign \new_[8042]_  = \new_[1530]_  | \new_[1531]_ ;
  assign \new_[8045]_  = \new_[1528]_  | \new_[1529]_ ;
  assign \new_[8046]_  = \new_[8045]_  | \new_[8042]_ ;
  assign \new_[8047]_  = \new_[8046]_  | \new_[8039]_ ;
  assign \new_[8051]_  = \new_[1525]_  | \new_[1526]_ ;
  assign \new_[8052]_  = \new_[1527]_  | \new_[8051]_ ;
  assign \new_[8055]_  = \new_[1523]_  | \new_[1524]_ ;
  assign \new_[8058]_  = \new_[1521]_  | \new_[1522]_ ;
  assign \new_[8059]_  = \new_[8058]_  | \new_[8055]_ ;
  assign \new_[8060]_  = \new_[8059]_  | \new_[8052]_ ;
  assign \new_[8061]_  = \new_[8060]_  | \new_[8047]_ ;
  assign \new_[8065]_  = \new_[1518]_  | \new_[1519]_ ;
  assign \new_[8066]_  = \new_[1520]_  | \new_[8065]_ ;
  assign \new_[8069]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[8072]_  = \new_[1514]_  | \new_[1515]_ ;
  assign \new_[8073]_  = \new_[8072]_  | \new_[8069]_ ;
  assign \new_[8074]_  = \new_[8073]_  | \new_[8066]_ ;
  assign \new_[8077]_  = \new_[1512]_  | \new_[1513]_ ;
  assign \new_[8080]_  = \new_[1510]_  | \new_[1511]_ ;
  assign \new_[8081]_  = \new_[8080]_  | \new_[8077]_ ;
  assign \new_[8084]_  = \new_[1508]_  | \new_[1509]_ ;
  assign \new_[8087]_  = \new_[1506]_  | \new_[1507]_ ;
  assign \new_[8088]_  = \new_[8087]_  | \new_[8084]_ ;
  assign \new_[8089]_  = \new_[8088]_  | \new_[8081]_ ;
  assign \new_[8090]_  = \new_[8089]_  | \new_[8074]_ ;
  assign \new_[8091]_  = \new_[8090]_  | \new_[8061]_ ;
  assign \new_[8092]_  = \new_[8091]_  | \new_[8034]_ ;
  assign \new_[8093]_  = \new_[8092]_  | \new_[7977]_ ;
  assign \new_[8097]_  = \new_[1503]_  | \new_[1504]_ ;
  assign \new_[8098]_  = \new_[1505]_  | \new_[8097]_ ;
  assign \new_[8101]_  = \new_[1501]_  | \new_[1502]_ ;
  assign \new_[8104]_  = \new_[1499]_  | \new_[1500]_ ;
  assign \new_[8105]_  = \new_[8104]_  | \new_[8101]_ ;
  assign \new_[8106]_  = \new_[8105]_  | \new_[8098]_ ;
  assign \new_[8110]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[8111]_  = \new_[1498]_  | \new_[8110]_ ;
  assign \new_[8114]_  = \new_[1494]_  | \new_[1495]_ ;
  assign \new_[8117]_  = \new_[1492]_  | \new_[1493]_ ;
  assign \new_[8118]_  = \new_[8117]_  | \new_[8114]_ ;
  assign \new_[8119]_  = \new_[8118]_  | \new_[8111]_ ;
  assign \new_[8120]_  = \new_[8119]_  | \new_[8106]_ ;
  assign \new_[8124]_  = \new_[1489]_  | \new_[1490]_ ;
  assign \new_[8125]_  = \new_[1491]_  | \new_[8124]_ ;
  assign \new_[8128]_  = \new_[1487]_  | \new_[1488]_ ;
  assign \new_[8131]_  = \new_[1485]_  | \new_[1486]_ ;
  assign \new_[8132]_  = \new_[8131]_  | \new_[8128]_ ;
  assign \new_[8133]_  = \new_[8132]_  | \new_[8125]_ ;
  assign \new_[8136]_  = \new_[1483]_  | \new_[1484]_ ;
  assign \new_[8139]_  = \new_[1481]_  | \new_[1482]_ ;
  assign \new_[8140]_  = \new_[8139]_  | \new_[8136]_ ;
  assign \new_[8143]_  = \new_[1479]_  | \new_[1480]_ ;
  assign \new_[8146]_  = \new_[1477]_  | \new_[1478]_ ;
  assign \new_[8147]_  = \new_[8146]_  | \new_[8143]_ ;
  assign \new_[8148]_  = \new_[8147]_  | \new_[8140]_ ;
  assign \new_[8149]_  = \new_[8148]_  | \new_[8133]_ ;
  assign \new_[8150]_  = \new_[8149]_  | \new_[8120]_ ;
  assign \new_[8154]_  = \new_[1474]_  | \new_[1475]_ ;
  assign \new_[8155]_  = \new_[1476]_  | \new_[8154]_ ;
  assign \new_[8158]_  = \new_[1472]_  | \new_[1473]_ ;
  assign \new_[8161]_  = \new_[1470]_  | \new_[1471]_ ;
  assign \new_[8162]_  = \new_[8161]_  | \new_[8158]_ ;
  assign \new_[8163]_  = \new_[8162]_  | \new_[8155]_ ;
  assign \new_[8167]_  = \new_[1467]_  | \new_[1468]_ ;
  assign \new_[8168]_  = \new_[1469]_  | \new_[8167]_ ;
  assign \new_[8171]_  = \new_[1465]_  | \new_[1466]_ ;
  assign \new_[8174]_  = \new_[1463]_  | \new_[1464]_ ;
  assign \new_[8175]_  = \new_[8174]_  | \new_[8171]_ ;
  assign \new_[8176]_  = \new_[8175]_  | \new_[8168]_ ;
  assign \new_[8177]_  = \new_[8176]_  | \new_[8163]_ ;
  assign \new_[8181]_  = \new_[1460]_  | \new_[1461]_ ;
  assign \new_[8182]_  = \new_[1462]_  | \new_[8181]_ ;
  assign \new_[8185]_  = \new_[1458]_  | \new_[1459]_ ;
  assign \new_[8188]_  = \new_[1456]_  | \new_[1457]_ ;
  assign \new_[8189]_  = \new_[8188]_  | \new_[8185]_ ;
  assign \new_[8190]_  = \new_[8189]_  | \new_[8182]_ ;
  assign \new_[8193]_  = \new_[1454]_  | \new_[1455]_ ;
  assign \new_[8196]_  = \new_[1452]_  | \new_[1453]_ ;
  assign \new_[8197]_  = \new_[8196]_  | \new_[8193]_ ;
  assign \new_[8200]_  = \new_[1450]_  | \new_[1451]_ ;
  assign \new_[8203]_  = \new_[1448]_  | \new_[1449]_ ;
  assign \new_[8204]_  = \new_[8203]_  | \new_[8200]_ ;
  assign \new_[8205]_  = \new_[8204]_  | \new_[8197]_ ;
  assign \new_[8206]_  = \new_[8205]_  | \new_[8190]_ ;
  assign \new_[8207]_  = \new_[8206]_  | \new_[8177]_ ;
  assign \new_[8208]_  = \new_[8207]_  | \new_[8150]_ ;
  assign \new_[8212]_  = \new_[1445]_  | \new_[1446]_ ;
  assign \new_[8213]_  = \new_[1447]_  | \new_[8212]_ ;
  assign \new_[8216]_  = \new_[1443]_  | \new_[1444]_ ;
  assign \new_[8219]_  = \new_[1441]_  | \new_[1442]_ ;
  assign \new_[8220]_  = \new_[8219]_  | \new_[8216]_ ;
  assign \new_[8221]_  = \new_[8220]_  | \new_[8213]_ ;
  assign \new_[8225]_  = \new_[1438]_  | \new_[1439]_ ;
  assign \new_[8226]_  = \new_[1440]_  | \new_[8225]_ ;
  assign \new_[8229]_  = \new_[1436]_  | \new_[1437]_ ;
  assign \new_[8232]_  = \new_[1434]_  | \new_[1435]_ ;
  assign \new_[8233]_  = \new_[8232]_  | \new_[8229]_ ;
  assign \new_[8234]_  = \new_[8233]_  | \new_[8226]_ ;
  assign \new_[8235]_  = \new_[8234]_  | \new_[8221]_ ;
  assign \new_[8239]_  = \new_[1431]_  | \new_[1432]_ ;
  assign \new_[8240]_  = \new_[1433]_  | \new_[8239]_ ;
  assign \new_[8243]_  = \new_[1429]_  | \new_[1430]_ ;
  assign \new_[8246]_  = \new_[1427]_  | \new_[1428]_ ;
  assign \new_[8247]_  = \new_[8246]_  | \new_[8243]_ ;
  assign \new_[8248]_  = \new_[8247]_  | \new_[8240]_ ;
  assign \new_[8251]_  = \new_[1425]_  | \new_[1426]_ ;
  assign \new_[8254]_  = \new_[1423]_  | \new_[1424]_ ;
  assign \new_[8255]_  = \new_[8254]_  | \new_[8251]_ ;
  assign \new_[8258]_  = \new_[1421]_  | \new_[1422]_ ;
  assign \new_[8261]_  = \new_[1419]_  | \new_[1420]_ ;
  assign \new_[8262]_  = \new_[8261]_  | \new_[8258]_ ;
  assign \new_[8263]_  = \new_[8262]_  | \new_[8255]_ ;
  assign \new_[8264]_  = \new_[8263]_  | \new_[8248]_ ;
  assign \new_[8265]_  = \new_[8264]_  | \new_[8235]_ ;
  assign \new_[8269]_  = \new_[1416]_  | \new_[1417]_ ;
  assign \new_[8270]_  = \new_[1418]_  | \new_[8269]_ ;
  assign \new_[8273]_  = \new_[1414]_  | \new_[1415]_ ;
  assign \new_[8276]_  = \new_[1412]_  | \new_[1413]_ ;
  assign \new_[8277]_  = \new_[8276]_  | \new_[8273]_ ;
  assign \new_[8278]_  = \new_[8277]_  | \new_[8270]_ ;
  assign \new_[8282]_  = \new_[1409]_  | \new_[1410]_ ;
  assign \new_[8283]_  = \new_[1411]_  | \new_[8282]_ ;
  assign \new_[8286]_  = \new_[1407]_  | \new_[1408]_ ;
  assign \new_[8289]_  = \new_[1405]_  | \new_[1406]_ ;
  assign \new_[8290]_  = \new_[8289]_  | \new_[8286]_ ;
  assign \new_[8291]_  = \new_[8290]_  | \new_[8283]_ ;
  assign \new_[8292]_  = \new_[8291]_  | \new_[8278]_ ;
  assign \new_[8296]_  = \new_[1402]_  | \new_[1403]_ ;
  assign \new_[8297]_  = \new_[1404]_  | \new_[8296]_ ;
  assign \new_[8300]_  = \new_[1400]_  | \new_[1401]_ ;
  assign \new_[8303]_  = \new_[1398]_  | \new_[1399]_ ;
  assign \new_[8304]_  = \new_[8303]_  | \new_[8300]_ ;
  assign \new_[8305]_  = \new_[8304]_  | \new_[8297]_ ;
  assign \new_[8308]_  = \new_[1396]_  | \new_[1397]_ ;
  assign \new_[8311]_  = \new_[1394]_  | \new_[1395]_ ;
  assign \new_[8312]_  = \new_[8311]_  | \new_[8308]_ ;
  assign \new_[8315]_  = \new_[1392]_  | \new_[1393]_ ;
  assign \new_[8318]_  = \new_[1390]_  | \new_[1391]_ ;
  assign \new_[8319]_  = \new_[8318]_  | \new_[8315]_ ;
  assign \new_[8320]_  = \new_[8319]_  | \new_[8312]_ ;
  assign \new_[8321]_  = \new_[8320]_  | \new_[8305]_ ;
  assign \new_[8322]_  = \new_[8321]_  | \new_[8292]_ ;
  assign \new_[8323]_  = \new_[8322]_  | \new_[8265]_ ;
  assign \new_[8324]_  = \new_[8323]_  | \new_[8208]_ ;
  assign \new_[8325]_  = \new_[8324]_  | \new_[8093]_ ;
  assign \new_[8326]_  = \new_[8325]_  | \new_[7864]_ ;
  assign \new_[8330]_  = \new_[1387]_  | \new_[1388]_ ;
  assign \new_[8331]_  = \new_[1389]_  | \new_[8330]_ ;
  assign \new_[8334]_  = \new_[1385]_  | \new_[1386]_ ;
  assign \new_[8337]_  = \new_[1383]_  | \new_[1384]_ ;
  assign \new_[8338]_  = \new_[8337]_  | \new_[8334]_ ;
  assign \new_[8339]_  = \new_[8338]_  | \new_[8331]_ ;
  assign \new_[8343]_  = \new_[1380]_  | \new_[1381]_ ;
  assign \new_[8344]_  = \new_[1382]_  | \new_[8343]_ ;
  assign \new_[8347]_  = \new_[1378]_  | \new_[1379]_ ;
  assign \new_[8350]_  = \new_[1376]_  | \new_[1377]_ ;
  assign \new_[8351]_  = \new_[8350]_  | \new_[8347]_ ;
  assign \new_[8352]_  = \new_[8351]_  | \new_[8344]_ ;
  assign \new_[8353]_  = \new_[8352]_  | \new_[8339]_ ;
  assign \new_[8357]_  = \new_[1373]_  | \new_[1374]_ ;
  assign \new_[8358]_  = \new_[1375]_  | \new_[8357]_ ;
  assign \new_[8361]_  = \new_[1371]_  | \new_[1372]_ ;
  assign \new_[8364]_  = \new_[1369]_  | \new_[1370]_ ;
  assign \new_[8365]_  = \new_[8364]_  | \new_[8361]_ ;
  assign \new_[8366]_  = \new_[8365]_  | \new_[8358]_ ;
  assign \new_[8370]_  = \new_[1366]_  | \new_[1367]_ ;
  assign \new_[8371]_  = \new_[1368]_  | \new_[8370]_ ;
  assign \new_[8374]_  = \new_[1364]_  | \new_[1365]_ ;
  assign \new_[8377]_  = \new_[1362]_  | \new_[1363]_ ;
  assign \new_[8378]_  = \new_[8377]_  | \new_[8374]_ ;
  assign \new_[8379]_  = \new_[8378]_  | \new_[8371]_ ;
  assign \new_[8380]_  = \new_[8379]_  | \new_[8366]_ ;
  assign \new_[8381]_  = \new_[8380]_  | \new_[8353]_ ;
  assign \new_[8385]_  = \new_[1359]_  | \new_[1360]_ ;
  assign \new_[8386]_  = \new_[1361]_  | \new_[8385]_ ;
  assign \new_[8389]_  = \new_[1357]_  | \new_[1358]_ ;
  assign \new_[8392]_  = \new_[1355]_  | \new_[1356]_ ;
  assign \new_[8393]_  = \new_[8392]_  | \new_[8389]_ ;
  assign \new_[8394]_  = \new_[8393]_  | \new_[8386]_ ;
  assign \new_[8398]_  = \new_[1352]_  | \new_[1353]_ ;
  assign \new_[8399]_  = \new_[1354]_  | \new_[8398]_ ;
  assign \new_[8402]_  = \new_[1350]_  | \new_[1351]_ ;
  assign \new_[8405]_  = \new_[1348]_  | \new_[1349]_ ;
  assign \new_[8406]_  = \new_[8405]_  | \new_[8402]_ ;
  assign \new_[8407]_  = \new_[8406]_  | \new_[8399]_ ;
  assign \new_[8408]_  = \new_[8407]_  | \new_[8394]_ ;
  assign \new_[8412]_  = \new_[1345]_  | \new_[1346]_ ;
  assign \new_[8413]_  = \new_[1347]_  | \new_[8412]_ ;
  assign \new_[8416]_  = \new_[1343]_  | \new_[1344]_ ;
  assign \new_[8419]_  = \new_[1341]_  | \new_[1342]_ ;
  assign \new_[8420]_  = \new_[8419]_  | \new_[8416]_ ;
  assign \new_[8421]_  = \new_[8420]_  | \new_[8413]_ ;
  assign \new_[8424]_  = \new_[1339]_  | \new_[1340]_ ;
  assign \new_[8427]_  = \new_[1337]_  | \new_[1338]_ ;
  assign \new_[8428]_  = \new_[8427]_  | \new_[8424]_ ;
  assign \new_[8431]_  = \new_[1335]_  | \new_[1336]_ ;
  assign \new_[8434]_  = \new_[1333]_  | \new_[1334]_ ;
  assign \new_[8435]_  = \new_[8434]_  | \new_[8431]_ ;
  assign \new_[8436]_  = \new_[8435]_  | \new_[8428]_ ;
  assign \new_[8437]_  = \new_[8436]_  | \new_[8421]_ ;
  assign \new_[8438]_  = \new_[8437]_  | \new_[8408]_ ;
  assign \new_[8439]_  = \new_[8438]_  | \new_[8381]_ ;
  assign \new_[8443]_  = \new_[1330]_  | \new_[1331]_ ;
  assign \new_[8444]_  = \new_[1332]_  | \new_[8443]_ ;
  assign \new_[8447]_  = \new_[1328]_  | \new_[1329]_ ;
  assign \new_[8450]_  = \new_[1326]_  | \new_[1327]_ ;
  assign \new_[8451]_  = \new_[8450]_  | \new_[8447]_ ;
  assign \new_[8452]_  = \new_[8451]_  | \new_[8444]_ ;
  assign \new_[8456]_  = \new_[1323]_  | \new_[1324]_ ;
  assign \new_[8457]_  = \new_[1325]_  | \new_[8456]_ ;
  assign \new_[8460]_  = \new_[1321]_  | \new_[1322]_ ;
  assign \new_[8463]_  = \new_[1319]_  | \new_[1320]_ ;
  assign \new_[8464]_  = \new_[8463]_  | \new_[8460]_ ;
  assign \new_[8465]_  = \new_[8464]_  | \new_[8457]_ ;
  assign \new_[8466]_  = \new_[8465]_  | \new_[8452]_ ;
  assign \new_[8470]_  = \new_[1316]_  | \new_[1317]_ ;
  assign \new_[8471]_  = \new_[1318]_  | \new_[8470]_ ;
  assign \new_[8474]_  = \new_[1314]_  | \new_[1315]_ ;
  assign \new_[8477]_  = \new_[1312]_  | \new_[1313]_ ;
  assign \new_[8478]_  = \new_[8477]_  | \new_[8474]_ ;
  assign \new_[8479]_  = \new_[8478]_  | \new_[8471]_ ;
  assign \new_[8482]_  = \new_[1310]_  | \new_[1311]_ ;
  assign \new_[8485]_  = \new_[1308]_  | \new_[1309]_ ;
  assign \new_[8486]_  = \new_[8485]_  | \new_[8482]_ ;
  assign \new_[8489]_  = \new_[1306]_  | \new_[1307]_ ;
  assign \new_[8492]_  = \new_[1304]_  | \new_[1305]_ ;
  assign \new_[8493]_  = \new_[8492]_  | \new_[8489]_ ;
  assign \new_[8494]_  = \new_[8493]_  | \new_[8486]_ ;
  assign \new_[8495]_  = \new_[8494]_  | \new_[8479]_ ;
  assign \new_[8496]_  = \new_[8495]_  | \new_[8466]_ ;
  assign \new_[8500]_  = \new_[1301]_  | \new_[1302]_ ;
  assign \new_[8501]_  = \new_[1303]_  | \new_[8500]_ ;
  assign \new_[8504]_  = \new_[1299]_  | \new_[1300]_ ;
  assign \new_[8507]_  = \new_[1297]_  | \new_[1298]_ ;
  assign \new_[8508]_  = \new_[8507]_  | \new_[8504]_ ;
  assign \new_[8509]_  = \new_[8508]_  | \new_[8501]_ ;
  assign \new_[8513]_  = \new_[1294]_  | \new_[1295]_ ;
  assign \new_[8514]_  = \new_[1296]_  | \new_[8513]_ ;
  assign \new_[8517]_  = \new_[1292]_  | \new_[1293]_ ;
  assign \new_[8520]_  = \new_[1290]_  | \new_[1291]_ ;
  assign \new_[8521]_  = \new_[8520]_  | \new_[8517]_ ;
  assign \new_[8522]_  = \new_[8521]_  | \new_[8514]_ ;
  assign \new_[8523]_  = \new_[8522]_  | \new_[8509]_ ;
  assign \new_[8527]_  = \new_[1287]_  | \new_[1288]_ ;
  assign \new_[8528]_  = \new_[1289]_  | \new_[8527]_ ;
  assign \new_[8531]_  = \new_[1285]_  | \new_[1286]_ ;
  assign \new_[8534]_  = \new_[1283]_  | \new_[1284]_ ;
  assign \new_[8535]_  = \new_[8534]_  | \new_[8531]_ ;
  assign \new_[8536]_  = \new_[8535]_  | \new_[8528]_ ;
  assign \new_[8539]_  = \new_[1281]_  | \new_[1282]_ ;
  assign \new_[8542]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[8543]_  = \new_[8542]_  | \new_[8539]_ ;
  assign \new_[8546]_  = \new_[1277]_  | \new_[1278]_ ;
  assign \new_[8549]_  = \new_[1275]_  | \new_[1276]_ ;
  assign \new_[8550]_  = \new_[8549]_  | \new_[8546]_ ;
  assign \new_[8551]_  = \new_[8550]_  | \new_[8543]_ ;
  assign \new_[8552]_  = \new_[8551]_  | \new_[8536]_ ;
  assign \new_[8553]_  = \new_[8552]_  | \new_[8523]_ ;
  assign \new_[8554]_  = \new_[8553]_  | \new_[8496]_ ;
  assign \new_[8555]_  = \new_[8554]_  | \new_[8439]_ ;
  assign \new_[8559]_  = \new_[1272]_  | \new_[1273]_ ;
  assign \new_[8560]_  = \new_[1274]_  | \new_[8559]_ ;
  assign \new_[8563]_  = \new_[1270]_  | \new_[1271]_ ;
  assign \new_[8566]_  = \new_[1268]_  | \new_[1269]_ ;
  assign \new_[8567]_  = \new_[8566]_  | \new_[8563]_ ;
  assign \new_[8568]_  = \new_[8567]_  | \new_[8560]_ ;
  assign \new_[8572]_  = \new_[1265]_  | \new_[1266]_ ;
  assign \new_[8573]_  = \new_[1267]_  | \new_[8572]_ ;
  assign \new_[8576]_  = \new_[1263]_  | \new_[1264]_ ;
  assign \new_[8579]_  = \new_[1261]_  | \new_[1262]_ ;
  assign \new_[8580]_  = \new_[8579]_  | \new_[8576]_ ;
  assign \new_[8581]_  = \new_[8580]_  | \new_[8573]_ ;
  assign \new_[8582]_  = \new_[8581]_  | \new_[8568]_ ;
  assign \new_[8586]_  = \new_[1258]_  | \new_[1259]_ ;
  assign \new_[8587]_  = \new_[1260]_  | \new_[8586]_ ;
  assign \new_[8590]_  = \new_[1256]_  | \new_[1257]_ ;
  assign \new_[8593]_  = \new_[1254]_  | \new_[1255]_ ;
  assign \new_[8594]_  = \new_[8593]_  | \new_[8590]_ ;
  assign \new_[8595]_  = \new_[8594]_  | \new_[8587]_ ;
  assign \new_[8598]_  = \new_[1252]_  | \new_[1253]_ ;
  assign \new_[8601]_  = \new_[1250]_  | \new_[1251]_ ;
  assign \new_[8602]_  = \new_[8601]_  | \new_[8598]_ ;
  assign \new_[8605]_  = \new_[1248]_  | \new_[1249]_ ;
  assign \new_[8608]_  = \new_[1246]_  | \new_[1247]_ ;
  assign \new_[8609]_  = \new_[8608]_  | \new_[8605]_ ;
  assign \new_[8610]_  = \new_[8609]_  | \new_[8602]_ ;
  assign \new_[8611]_  = \new_[8610]_  | \new_[8595]_ ;
  assign \new_[8612]_  = \new_[8611]_  | \new_[8582]_ ;
  assign \new_[8616]_  = \new_[1243]_  | \new_[1244]_ ;
  assign \new_[8617]_  = \new_[1245]_  | \new_[8616]_ ;
  assign \new_[8620]_  = \new_[1241]_  | \new_[1242]_ ;
  assign \new_[8623]_  = \new_[1239]_  | \new_[1240]_ ;
  assign \new_[8624]_  = \new_[8623]_  | \new_[8620]_ ;
  assign \new_[8625]_  = \new_[8624]_  | \new_[8617]_ ;
  assign \new_[8629]_  = \new_[1236]_  | \new_[1237]_ ;
  assign \new_[8630]_  = \new_[1238]_  | \new_[8629]_ ;
  assign \new_[8633]_  = \new_[1234]_  | \new_[1235]_ ;
  assign \new_[8636]_  = \new_[1232]_  | \new_[1233]_ ;
  assign \new_[8637]_  = \new_[8636]_  | \new_[8633]_ ;
  assign \new_[8638]_  = \new_[8637]_  | \new_[8630]_ ;
  assign \new_[8639]_  = \new_[8638]_  | \new_[8625]_ ;
  assign \new_[8643]_  = \new_[1229]_  | \new_[1230]_ ;
  assign \new_[8644]_  = \new_[1231]_  | \new_[8643]_ ;
  assign \new_[8647]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[8650]_  = \new_[1225]_  | \new_[1226]_ ;
  assign \new_[8651]_  = \new_[8650]_  | \new_[8647]_ ;
  assign \new_[8652]_  = \new_[8651]_  | \new_[8644]_ ;
  assign \new_[8655]_  = \new_[1223]_  | \new_[1224]_ ;
  assign \new_[8658]_  = \new_[1221]_  | \new_[1222]_ ;
  assign \new_[8659]_  = \new_[8658]_  | \new_[8655]_ ;
  assign \new_[8662]_  = \new_[1219]_  | \new_[1220]_ ;
  assign \new_[8665]_  = \new_[1217]_  | \new_[1218]_ ;
  assign \new_[8666]_  = \new_[8665]_  | \new_[8662]_ ;
  assign \new_[8667]_  = \new_[8666]_  | \new_[8659]_ ;
  assign \new_[8668]_  = \new_[8667]_  | \new_[8652]_ ;
  assign \new_[8669]_  = \new_[8668]_  | \new_[8639]_ ;
  assign \new_[8670]_  = \new_[8669]_  | \new_[8612]_ ;
  assign \new_[8674]_  = \new_[1214]_  | \new_[1215]_ ;
  assign \new_[8675]_  = \new_[1216]_  | \new_[8674]_ ;
  assign \new_[8678]_  = \new_[1212]_  | \new_[1213]_ ;
  assign \new_[8681]_  = \new_[1210]_  | \new_[1211]_ ;
  assign \new_[8682]_  = \new_[8681]_  | \new_[8678]_ ;
  assign \new_[8683]_  = \new_[8682]_  | \new_[8675]_ ;
  assign \new_[8687]_  = \new_[1207]_  | \new_[1208]_ ;
  assign \new_[8688]_  = \new_[1209]_  | \new_[8687]_ ;
  assign \new_[8691]_  = \new_[1205]_  | \new_[1206]_ ;
  assign \new_[8694]_  = \new_[1203]_  | \new_[1204]_ ;
  assign \new_[8695]_  = \new_[8694]_  | \new_[8691]_ ;
  assign \new_[8696]_  = \new_[8695]_  | \new_[8688]_ ;
  assign \new_[8697]_  = \new_[8696]_  | \new_[8683]_ ;
  assign \new_[8701]_  = \new_[1200]_  | \new_[1201]_ ;
  assign \new_[8702]_  = \new_[1202]_  | \new_[8701]_ ;
  assign \new_[8705]_  = \new_[1198]_  | \new_[1199]_ ;
  assign \new_[8708]_  = \new_[1196]_  | \new_[1197]_ ;
  assign \new_[8709]_  = \new_[8708]_  | \new_[8705]_ ;
  assign \new_[8710]_  = \new_[8709]_  | \new_[8702]_ ;
  assign \new_[8713]_  = \new_[1194]_  | \new_[1195]_ ;
  assign \new_[8716]_  = \new_[1192]_  | \new_[1193]_ ;
  assign \new_[8717]_  = \new_[8716]_  | \new_[8713]_ ;
  assign \new_[8720]_  = \new_[1190]_  | \new_[1191]_ ;
  assign \new_[8723]_  = \new_[1188]_  | \new_[1189]_ ;
  assign \new_[8724]_  = \new_[8723]_  | \new_[8720]_ ;
  assign \new_[8725]_  = \new_[8724]_  | \new_[8717]_ ;
  assign \new_[8726]_  = \new_[8725]_  | \new_[8710]_ ;
  assign \new_[8727]_  = \new_[8726]_  | \new_[8697]_ ;
  assign \new_[8731]_  = \new_[1185]_  | \new_[1186]_ ;
  assign \new_[8732]_  = \new_[1187]_  | \new_[8731]_ ;
  assign \new_[8735]_  = \new_[1183]_  | \new_[1184]_ ;
  assign \new_[8738]_  = \new_[1181]_  | \new_[1182]_ ;
  assign \new_[8739]_  = \new_[8738]_  | \new_[8735]_ ;
  assign \new_[8740]_  = \new_[8739]_  | \new_[8732]_ ;
  assign \new_[8744]_  = \new_[1178]_  | \new_[1179]_ ;
  assign \new_[8745]_  = \new_[1180]_  | \new_[8744]_ ;
  assign \new_[8748]_  = \new_[1176]_  | \new_[1177]_ ;
  assign \new_[8751]_  = \new_[1174]_  | \new_[1175]_ ;
  assign \new_[8752]_  = \new_[8751]_  | \new_[8748]_ ;
  assign \new_[8753]_  = \new_[8752]_  | \new_[8745]_ ;
  assign \new_[8754]_  = \new_[8753]_  | \new_[8740]_ ;
  assign \new_[8758]_  = \new_[1171]_  | \new_[1172]_ ;
  assign \new_[8759]_  = \new_[1173]_  | \new_[8758]_ ;
  assign \new_[8762]_  = \new_[1169]_  | \new_[1170]_ ;
  assign \new_[8765]_  = \new_[1167]_  | \new_[1168]_ ;
  assign \new_[8766]_  = \new_[8765]_  | \new_[8762]_ ;
  assign \new_[8767]_  = \new_[8766]_  | \new_[8759]_ ;
  assign \new_[8770]_  = \new_[1165]_  | \new_[1166]_ ;
  assign \new_[8773]_  = \new_[1163]_  | \new_[1164]_ ;
  assign \new_[8774]_  = \new_[8773]_  | \new_[8770]_ ;
  assign \new_[8777]_  = \new_[1161]_  | \new_[1162]_ ;
  assign \new_[8780]_  = \new_[1159]_  | \new_[1160]_ ;
  assign \new_[8781]_  = \new_[8780]_  | \new_[8777]_ ;
  assign \new_[8782]_  = \new_[8781]_  | \new_[8774]_ ;
  assign \new_[8783]_  = \new_[8782]_  | \new_[8767]_ ;
  assign \new_[8784]_  = \new_[8783]_  | \new_[8754]_ ;
  assign \new_[8785]_  = \new_[8784]_  | \new_[8727]_ ;
  assign \new_[8786]_  = \new_[8785]_  | \new_[8670]_ ;
  assign \new_[8787]_  = \new_[8786]_  | \new_[8555]_ ;
  assign \new_[8791]_  = \new_[1156]_  | \new_[1157]_ ;
  assign \new_[8792]_  = \new_[1158]_  | \new_[8791]_ ;
  assign \new_[8795]_  = \new_[1154]_  | \new_[1155]_ ;
  assign \new_[8798]_  = \new_[1152]_  | \new_[1153]_ ;
  assign \new_[8799]_  = \new_[8798]_  | \new_[8795]_ ;
  assign \new_[8800]_  = \new_[8799]_  | \new_[8792]_ ;
  assign \new_[8804]_  = \new_[1149]_  | \new_[1150]_ ;
  assign \new_[8805]_  = \new_[1151]_  | \new_[8804]_ ;
  assign \new_[8808]_  = \new_[1147]_  | \new_[1148]_ ;
  assign \new_[8811]_  = \new_[1145]_  | \new_[1146]_ ;
  assign \new_[8812]_  = \new_[8811]_  | \new_[8808]_ ;
  assign \new_[8813]_  = \new_[8812]_  | \new_[8805]_ ;
  assign \new_[8814]_  = \new_[8813]_  | \new_[8800]_ ;
  assign \new_[8818]_  = \new_[1142]_  | \new_[1143]_ ;
  assign \new_[8819]_  = \new_[1144]_  | \new_[8818]_ ;
  assign \new_[8822]_  = \new_[1140]_  | \new_[1141]_ ;
  assign \new_[8825]_  = \new_[1138]_  | \new_[1139]_ ;
  assign \new_[8826]_  = \new_[8825]_  | \new_[8822]_ ;
  assign \new_[8827]_  = \new_[8826]_  | \new_[8819]_ ;
  assign \new_[8830]_  = \new_[1136]_  | \new_[1137]_ ;
  assign \new_[8833]_  = \new_[1134]_  | \new_[1135]_ ;
  assign \new_[8834]_  = \new_[8833]_  | \new_[8830]_ ;
  assign \new_[8837]_  = \new_[1132]_  | \new_[1133]_ ;
  assign \new_[8840]_  = \new_[1130]_  | \new_[1131]_ ;
  assign \new_[8841]_  = \new_[8840]_  | \new_[8837]_ ;
  assign \new_[8842]_  = \new_[8841]_  | \new_[8834]_ ;
  assign \new_[8843]_  = \new_[8842]_  | \new_[8827]_ ;
  assign \new_[8844]_  = \new_[8843]_  | \new_[8814]_ ;
  assign \new_[8848]_  = \new_[1127]_  | \new_[1128]_ ;
  assign \new_[8849]_  = \new_[1129]_  | \new_[8848]_ ;
  assign \new_[8852]_  = \new_[1125]_  | \new_[1126]_ ;
  assign \new_[8855]_  = \new_[1123]_  | \new_[1124]_ ;
  assign \new_[8856]_  = \new_[8855]_  | \new_[8852]_ ;
  assign \new_[8857]_  = \new_[8856]_  | \new_[8849]_ ;
  assign \new_[8861]_  = \new_[1120]_  | \new_[1121]_ ;
  assign \new_[8862]_  = \new_[1122]_  | \new_[8861]_ ;
  assign \new_[8865]_  = \new_[1118]_  | \new_[1119]_ ;
  assign \new_[8868]_  = \new_[1116]_  | \new_[1117]_ ;
  assign \new_[8869]_  = \new_[8868]_  | \new_[8865]_ ;
  assign \new_[8870]_  = \new_[8869]_  | \new_[8862]_ ;
  assign \new_[8871]_  = \new_[8870]_  | \new_[8857]_ ;
  assign \new_[8875]_  = \new_[1113]_  | \new_[1114]_ ;
  assign \new_[8876]_  = \new_[1115]_  | \new_[8875]_ ;
  assign \new_[8879]_  = \new_[1111]_  | \new_[1112]_ ;
  assign \new_[8882]_  = \new_[1109]_  | \new_[1110]_ ;
  assign \new_[8883]_  = \new_[8882]_  | \new_[8879]_ ;
  assign \new_[8884]_  = \new_[8883]_  | \new_[8876]_ ;
  assign \new_[8887]_  = \new_[1107]_  | \new_[1108]_ ;
  assign \new_[8890]_  = \new_[1105]_  | \new_[1106]_ ;
  assign \new_[8891]_  = \new_[8890]_  | \new_[8887]_ ;
  assign \new_[8894]_  = \new_[1103]_  | \new_[1104]_ ;
  assign \new_[8897]_  = \new_[1101]_  | \new_[1102]_ ;
  assign \new_[8898]_  = \new_[8897]_  | \new_[8894]_ ;
  assign \new_[8899]_  = \new_[8898]_  | \new_[8891]_ ;
  assign \new_[8900]_  = \new_[8899]_  | \new_[8884]_ ;
  assign \new_[8901]_  = \new_[8900]_  | \new_[8871]_ ;
  assign \new_[8902]_  = \new_[8901]_  | \new_[8844]_ ;
  assign \new_[8906]_  = \new_[1098]_  | \new_[1099]_ ;
  assign \new_[8907]_  = \new_[1100]_  | \new_[8906]_ ;
  assign \new_[8910]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[8913]_  = \new_[1094]_  | \new_[1095]_ ;
  assign \new_[8914]_  = \new_[8913]_  | \new_[8910]_ ;
  assign \new_[8915]_  = \new_[8914]_  | \new_[8907]_ ;
  assign \new_[8919]_  = \new_[1091]_  | \new_[1092]_ ;
  assign \new_[8920]_  = \new_[1093]_  | \new_[8919]_ ;
  assign \new_[8923]_  = \new_[1089]_  | \new_[1090]_ ;
  assign \new_[8926]_  = \new_[1087]_  | \new_[1088]_ ;
  assign \new_[8927]_  = \new_[8926]_  | \new_[8923]_ ;
  assign \new_[8928]_  = \new_[8927]_  | \new_[8920]_ ;
  assign \new_[8929]_  = \new_[8928]_  | \new_[8915]_ ;
  assign \new_[8933]_  = \new_[1084]_  | \new_[1085]_ ;
  assign \new_[8934]_  = \new_[1086]_  | \new_[8933]_ ;
  assign \new_[8937]_  = \new_[1082]_  | \new_[1083]_ ;
  assign \new_[8940]_  = \new_[1080]_  | \new_[1081]_ ;
  assign \new_[8941]_  = \new_[8940]_  | \new_[8937]_ ;
  assign \new_[8942]_  = \new_[8941]_  | \new_[8934]_ ;
  assign \new_[8945]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[8948]_  = \new_[1076]_  | \new_[1077]_ ;
  assign \new_[8949]_  = \new_[8948]_  | \new_[8945]_ ;
  assign \new_[8952]_  = \new_[1074]_  | \new_[1075]_ ;
  assign \new_[8955]_  = \new_[1072]_  | \new_[1073]_ ;
  assign \new_[8956]_  = \new_[8955]_  | \new_[8952]_ ;
  assign \new_[8957]_  = \new_[8956]_  | \new_[8949]_ ;
  assign \new_[8958]_  = \new_[8957]_  | \new_[8942]_ ;
  assign \new_[8959]_  = \new_[8958]_  | \new_[8929]_ ;
  assign \new_[8963]_  = \new_[1069]_  | \new_[1070]_ ;
  assign \new_[8964]_  = \new_[1071]_  | \new_[8963]_ ;
  assign \new_[8967]_  = \new_[1067]_  | \new_[1068]_ ;
  assign \new_[8970]_  = \new_[1065]_  | \new_[1066]_ ;
  assign \new_[8971]_  = \new_[8970]_  | \new_[8967]_ ;
  assign \new_[8972]_  = \new_[8971]_  | \new_[8964]_ ;
  assign \new_[8976]_  = \new_[1062]_  | \new_[1063]_ ;
  assign \new_[8977]_  = \new_[1064]_  | \new_[8976]_ ;
  assign \new_[8980]_  = \new_[1060]_  | \new_[1061]_ ;
  assign \new_[8983]_  = \new_[1058]_  | \new_[1059]_ ;
  assign \new_[8984]_  = \new_[8983]_  | \new_[8980]_ ;
  assign \new_[8985]_  = \new_[8984]_  | \new_[8977]_ ;
  assign \new_[8986]_  = \new_[8985]_  | \new_[8972]_ ;
  assign \new_[8990]_  = \new_[1055]_  | \new_[1056]_ ;
  assign \new_[8991]_  = \new_[1057]_  | \new_[8990]_ ;
  assign \new_[8994]_  = \new_[1053]_  | \new_[1054]_ ;
  assign \new_[8997]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[8998]_  = \new_[8997]_  | \new_[8994]_ ;
  assign \new_[8999]_  = \new_[8998]_  | \new_[8991]_ ;
  assign \new_[9002]_  = \new_[1049]_  | \new_[1050]_ ;
  assign \new_[9005]_  = \new_[1047]_  | \new_[1048]_ ;
  assign \new_[9006]_  = \new_[9005]_  | \new_[9002]_ ;
  assign \new_[9009]_  = \new_[1045]_  | \new_[1046]_ ;
  assign \new_[9012]_  = \new_[1043]_  | \new_[1044]_ ;
  assign \new_[9013]_  = \new_[9012]_  | \new_[9009]_ ;
  assign \new_[9014]_  = \new_[9013]_  | \new_[9006]_ ;
  assign \new_[9015]_  = \new_[9014]_  | \new_[8999]_ ;
  assign \new_[9016]_  = \new_[9015]_  | \new_[8986]_ ;
  assign \new_[9017]_  = \new_[9016]_  | \new_[8959]_ ;
  assign \new_[9018]_  = \new_[9017]_  | \new_[8902]_ ;
  assign \new_[9022]_  = \new_[1040]_  | \new_[1041]_ ;
  assign \new_[9023]_  = \new_[1042]_  | \new_[9022]_ ;
  assign \new_[9026]_  = \new_[1038]_  | \new_[1039]_ ;
  assign \new_[9029]_  = \new_[1036]_  | \new_[1037]_ ;
  assign \new_[9030]_  = \new_[9029]_  | \new_[9026]_ ;
  assign \new_[9031]_  = \new_[9030]_  | \new_[9023]_ ;
  assign \new_[9035]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[9036]_  = \new_[1035]_  | \new_[9035]_ ;
  assign \new_[9039]_  = \new_[1031]_  | \new_[1032]_ ;
  assign \new_[9042]_  = \new_[1029]_  | \new_[1030]_ ;
  assign \new_[9043]_  = \new_[9042]_  | \new_[9039]_ ;
  assign \new_[9044]_  = \new_[9043]_  | \new_[9036]_ ;
  assign \new_[9045]_  = \new_[9044]_  | \new_[9031]_ ;
  assign \new_[9049]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[9050]_  = \new_[1028]_  | \new_[9049]_ ;
  assign \new_[9053]_  = \new_[1024]_  | \new_[1025]_ ;
  assign \new_[9056]_  = \new_[1022]_  | \new_[1023]_ ;
  assign \new_[9057]_  = \new_[9056]_  | \new_[9053]_ ;
  assign \new_[9058]_  = \new_[9057]_  | \new_[9050]_ ;
  assign \new_[9061]_  = \new_[1020]_  | \new_[1021]_ ;
  assign \new_[9064]_  = \new_[1018]_  | \new_[1019]_ ;
  assign \new_[9065]_  = \new_[9064]_  | \new_[9061]_ ;
  assign \new_[9068]_  = \new_[1016]_  | \new_[1017]_ ;
  assign \new_[9071]_  = \new_[1014]_  | \new_[1015]_ ;
  assign \new_[9072]_  = \new_[9071]_  | \new_[9068]_ ;
  assign \new_[9073]_  = \new_[9072]_  | \new_[9065]_ ;
  assign \new_[9074]_  = \new_[9073]_  | \new_[9058]_ ;
  assign \new_[9075]_  = \new_[9074]_  | \new_[9045]_ ;
  assign \new_[9079]_  = \new_[1011]_  | \new_[1012]_ ;
  assign \new_[9080]_  = \new_[1013]_  | \new_[9079]_ ;
  assign \new_[9083]_  = \new_[1009]_  | \new_[1010]_ ;
  assign \new_[9086]_  = \new_[1007]_  | \new_[1008]_ ;
  assign \new_[9087]_  = \new_[9086]_  | \new_[9083]_ ;
  assign \new_[9088]_  = \new_[9087]_  | \new_[9080]_ ;
  assign \new_[9092]_  = \new_[1004]_  | \new_[1005]_ ;
  assign \new_[9093]_  = \new_[1006]_  | \new_[9092]_ ;
  assign \new_[9096]_  = \new_[1002]_  | \new_[1003]_ ;
  assign \new_[9099]_  = \new_[1000]_  | \new_[1001]_ ;
  assign \new_[9100]_  = \new_[9099]_  | \new_[9096]_ ;
  assign \new_[9101]_  = \new_[9100]_  | \new_[9093]_ ;
  assign \new_[9102]_  = \new_[9101]_  | \new_[9088]_ ;
  assign \new_[9106]_  = \new_[997]_  | \new_[998]_ ;
  assign \new_[9107]_  = \new_[999]_  | \new_[9106]_ ;
  assign \new_[9110]_  = \new_[995]_  | \new_[996]_ ;
  assign \new_[9113]_  = \new_[993]_  | \new_[994]_ ;
  assign \new_[9114]_  = \new_[9113]_  | \new_[9110]_ ;
  assign \new_[9115]_  = \new_[9114]_  | \new_[9107]_ ;
  assign \new_[9118]_  = \new_[991]_  | \new_[992]_ ;
  assign \new_[9121]_  = \new_[989]_  | \new_[990]_ ;
  assign \new_[9122]_  = \new_[9121]_  | \new_[9118]_ ;
  assign \new_[9125]_  = \new_[987]_  | \new_[988]_ ;
  assign \new_[9128]_  = \new_[985]_  | \new_[986]_ ;
  assign \new_[9129]_  = \new_[9128]_  | \new_[9125]_ ;
  assign \new_[9130]_  = \new_[9129]_  | \new_[9122]_ ;
  assign \new_[9131]_  = \new_[9130]_  | \new_[9115]_ ;
  assign \new_[9132]_  = \new_[9131]_  | \new_[9102]_ ;
  assign \new_[9133]_  = \new_[9132]_  | \new_[9075]_ ;
  assign \new_[9137]_  = \new_[982]_  | \new_[983]_ ;
  assign \new_[9138]_  = \new_[984]_  | \new_[9137]_ ;
  assign \new_[9141]_  = \new_[980]_  | \new_[981]_ ;
  assign \new_[9144]_  = \new_[978]_  | \new_[979]_ ;
  assign \new_[9145]_  = \new_[9144]_  | \new_[9141]_ ;
  assign \new_[9146]_  = \new_[9145]_  | \new_[9138]_ ;
  assign \new_[9150]_  = \new_[975]_  | \new_[976]_ ;
  assign \new_[9151]_  = \new_[977]_  | \new_[9150]_ ;
  assign \new_[9154]_  = \new_[973]_  | \new_[974]_ ;
  assign \new_[9157]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[9158]_  = \new_[9157]_  | \new_[9154]_ ;
  assign \new_[9159]_  = \new_[9158]_  | \new_[9151]_ ;
  assign \new_[9160]_  = \new_[9159]_  | \new_[9146]_ ;
  assign \new_[9164]_  = \new_[968]_  | \new_[969]_ ;
  assign \new_[9165]_  = \new_[970]_  | \new_[9164]_ ;
  assign \new_[9168]_  = \new_[966]_  | \new_[967]_ ;
  assign \new_[9171]_  = \new_[964]_  | \new_[965]_ ;
  assign \new_[9172]_  = \new_[9171]_  | \new_[9168]_ ;
  assign \new_[9173]_  = \new_[9172]_  | \new_[9165]_ ;
  assign \new_[9176]_  = \new_[962]_  | \new_[963]_ ;
  assign \new_[9179]_  = \new_[960]_  | \new_[961]_ ;
  assign \new_[9180]_  = \new_[9179]_  | \new_[9176]_ ;
  assign \new_[9183]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[9186]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[9187]_  = \new_[9186]_  | \new_[9183]_ ;
  assign \new_[9188]_  = \new_[9187]_  | \new_[9180]_ ;
  assign \new_[9189]_  = \new_[9188]_  | \new_[9173]_ ;
  assign \new_[9190]_  = \new_[9189]_  | \new_[9160]_ ;
  assign \new_[9194]_  = \new_[953]_  | \new_[954]_ ;
  assign \new_[9195]_  = \new_[955]_  | \new_[9194]_ ;
  assign \new_[9198]_  = \new_[951]_  | \new_[952]_ ;
  assign \new_[9201]_  = \new_[949]_  | \new_[950]_ ;
  assign \new_[9202]_  = \new_[9201]_  | \new_[9198]_ ;
  assign \new_[9203]_  = \new_[9202]_  | \new_[9195]_ ;
  assign \new_[9207]_  = \new_[946]_  | \new_[947]_ ;
  assign \new_[9208]_  = \new_[948]_  | \new_[9207]_ ;
  assign \new_[9211]_  = \new_[944]_  | \new_[945]_ ;
  assign \new_[9214]_  = \new_[942]_  | \new_[943]_ ;
  assign \new_[9215]_  = \new_[9214]_  | \new_[9211]_ ;
  assign \new_[9216]_  = \new_[9215]_  | \new_[9208]_ ;
  assign \new_[9217]_  = \new_[9216]_  | \new_[9203]_ ;
  assign \new_[9221]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[9222]_  = \new_[941]_  | \new_[9221]_ ;
  assign \new_[9225]_  = \new_[937]_  | \new_[938]_ ;
  assign \new_[9228]_  = \new_[935]_  | \new_[936]_ ;
  assign \new_[9229]_  = \new_[9228]_  | \new_[9225]_ ;
  assign \new_[9230]_  = \new_[9229]_  | \new_[9222]_ ;
  assign \new_[9233]_  = \new_[933]_  | \new_[934]_ ;
  assign \new_[9236]_  = \new_[931]_  | \new_[932]_ ;
  assign \new_[9237]_  = \new_[9236]_  | \new_[9233]_ ;
  assign \new_[9240]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[9243]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[9244]_  = \new_[9243]_  | \new_[9240]_ ;
  assign \new_[9245]_  = \new_[9244]_  | \new_[9237]_ ;
  assign \new_[9246]_  = \new_[9245]_  | \new_[9230]_ ;
  assign \new_[9247]_  = \new_[9246]_  | \new_[9217]_ ;
  assign \new_[9248]_  = \new_[9247]_  | \new_[9190]_ ;
  assign \new_[9249]_  = \new_[9248]_  | \new_[9133]_ ;
  assign \new_[9250]_  = \new_[9249]_  | \new_[9018]_ ;
  assign \new_[9251]_  = \new_[9250]_  | \new_[8787]_ ;
  assign \new_[9252]_  = \new_[9251]_  | \new_[8326]_ ;
  assign \new_[9256]_  = \new_[924]_  | \new_[925]_ ;
  assign \new_[9257]_  = \new_[926]_  | \new_[9256]_ ;
  assign \new_[9260]_  = \new_[922]_  | \new_[923]_ ;
  assign \new_[9263]_  = \new_[920]_  | \new_[921]_ ;
  assign \new_[9264]_  = \new_[9263]_  | \new_[9260]_ ;
  assign \new_[9265]_  = \new_[9264]_  | \new_[9257]_ ;
  assign \new_[9269]_  = \new_[917]_  | \new_[918]_ ;
  assign \new_[9270]_  = \new_[919]_  | \new_[9269]_ ;
  assign \new_[9273]_  = \new_[915]_  | \new_[916]_ ;
  assign \new_[9276]_  = \new_[913]_  | \new_[914]_ ;
  assign \new_[9277]_  = \new_[9276]_  | \new_[9273]_ ;
  assign \new_[9278]_  = \new_[9277]_  | \new_[9270]_ ;
  assign \new_[9279]_  = \new_[9278]_  | \new_[9265]_ ;
  assign \new_[9283]_  = \new_[910]_  | \new_[911]_ ;
  assign \new_[9284]_  = \new_[912]_  | \new_[9283]_ ;
  assign \new_[9287]_  = \new_[908]_  | \new_[909]_ ;
  assign \new_[9290]_  = \new_[906]_  | \new_[907]_ ;
  assign \new_[9291]_  = \new_[9290]_  | \new_[9287]_ ;
  assign \new_[9292]_  = \new_[9291]_  | \new_[9284]_ ;
  assign \new_[9296]_  = \new_[903]_  | \new_[904]_ ;
  assign \new_[9297]_  = \new_[905]_  | \new_[9296]_ ;
  assign \new_[9300]_  = \new_[901]_  | \new_[902]_ ;
  assign \new_[9303]_  = \new_[899]_  | \new_[900]_ ;
  assign \new_[9304]_  = \new_[9303]_  | \new_[9300]_ ;
  assign \new_[9305]_  = \new_[9304]_  | \new_[9297]_ ;
  assign \new_[9306]_  = \new_[9305]_  | \new_[9292]_ ;
  assign \new_[9307]_  = \new_[9306]_  | \new_[9279]_ ;
  assign \new_[9311]_  = \new_[896]_  | \new_[897]_ ;
  assign \new_[9312]_  = \new_[898]_  | \new_[9311]_ ;
  assign \new_[9315]_  = \new_[894]_  | \new_[895]_ ;
  assign \new_[9318]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[9319]_  = \new_[9318]_  | \new_[9315]_ ;
  assign \new_[9320]_  = \new_[9319]_  | \new_[9312]_ ;
  assign \new_[9324]_  = \new_[889]_  | \new_[890]_ ;
  assign \new_[9325]_  = \new_[891]_  | \new_[9324]_ ;
  assign \new_[9328]_  = \new_[887]_  | \new_[888]_ ;
  assign \new_[9331]_  = \new_[885]_  | \new_[886]_ ;
  assign \new_[9332]_  = \new_[9331]_  | \new_[9328]_ ;
  assign \new_[9333]_  = \new_[9332]_  | \new_[9325]_ ;
  assign \new_[9334]_  = \new_[9333]_  | \new_[9320]_ ;
  assign \new_[9338]_  = \new_[882]_  | \new_[883]_ ;
  assign \new_[9339]_  = \new_[884]_  | \new_[9338]_ ;
  assign \new_[9342]_  = \new_[880]_  | \new_[881]_ ;
  assign \new_[9345]_  = \new_[878]_  | \new_[879]_ ;
  assign \new_[9346]_  = \new_[9345]_  | \new_[9342]_ ;
  assign \new_[9347]_  = \new_[9346]_  | \new_[9339]_ ;
  assign \new_[9350]_  = \new_[876]_  | \new_[877]_ ;
  assign \new_[9353]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[9354]_  = \new_[9353]_  | \new_[9350]_ ;
  assign \new_[9357]_  = \new_[872]_  | \new_[873]_ ;
  assign \new_[9360]_  = \new_[870]_  | \new_[871]_ ;
  assign \new_[9361]_  = \new_[9360]_  | \new_[9357]_ ;
  assign \new_[9362]_  = \new_[9361]_  | \new_[9354]_ ;
  assign \new_[9363]_  = \new_[9362]_  | \new_[9347]_ ;
  assign \new_[9364]_  = \new_[9363]_  | \new_[9334]_ ;
  assign \new_[9365]_  = \new_[9364]_  | \new_[9307]_ ;
  assign \new_[9369]_  = \new_[867]_  | \new_[868]_ ;
  assign \new_[9370]_  = \new_[869]_  | \new_[9369]_ ;
  assign \new_[9373]_  = \new_[865]_  | \new_[866]_ ;
  assign \new_[9376]_  = \new_[863]_  | \new_[864]_ ;
  assign \new_[9377]_  = \new_[9376]_  | \new_[9373]_ ;
  assign \new_[9378]_  = \new_[9377]_  | \new_[9370]_ ;
  assign \new_[9382]_  = \new_[860]_  | \new_[861]_ ;
  assign \new_[9383]_  = \new_[862]_  | \new_[9382]_ ;
  assign \new_[9386]_  = \new_[858]_  | \new_[859]_ ;
  assign \new_[9389]_  = \new_[856]_  | \new_[857]_ ;
  assign \new_[9390]_  = \new_[9389]_  | \new_[9386]_ ;
  assign \new_[9391]_  = \new_[9390]_  | \new_[9383]_ ;
  assign \new_[9392]_  = \new_[9391]_  | \new_[9378]_ ;
  assign \new_[9396]_  = \new_[853]_  | \new_[854]_ ;
  assign \new_[9397]_  = \new_[855]_  | \new_[9396]_ ;
  assign \new_[9400]_  = \new_[851]_  | \new_[852]_ ;
  assign \new_[9403]_  = \new_[849]_  | \new_[850]_ ;
  assign \new_[9404]_  = \new_[9403]_  | \new_[9400]_ ;
  assign \new_[9405]_  = \new_[9404]_  | \new_[9397]_ ;
  assign \new_[9408]_  = \new_[847]_  | \new_[848]_ ;
  assign \new_[9411]_  = \new_[845]_  | \new_[846]_ ;
  assign \new_[9412]_  = \new_[9411]_  | \new_[9408]_ ;
  assign \new_[9415]_  = \new_[843]_  | \new_[844]_ ;
  assign \new_[9418]_  = \new_[841]_  | \new_[842]_ ;
  assign \new_[9419]_  = \new_[9418]_  | \new_[9415]_ ;
  assign \new_[9420]_  = \new_[9419]_  | \new_[9412]_ ;
  assign \new_[9421]_  = \new_[9420]_  | \new_[9405]_ ;
  assign \new_[9422]_  = \new_[9421]_  | \new_[9392]_ ;
  assign \new_[9426]_  = \new_[838]_  | \new_[839]_ ;
  assign \new_[9427]_  = \new_[840]_  | \new_[9426]_ ;
  assign \new_[9430]_  = \new_[836]_  | \new_[837]_ ;
  assign \new_[9433]_  = \new_[834]_  | \new_[835]_ ;
  assign \new_[9434]_  = \new_[9433]_  | \new_[9430]_ ;
  assign \new_[9435]_  = \new_[9434]_  | \new_[9427]_ ;
  assign \new_[9439]_  = \new_[831]_  | \new_[832]_ ;
  assign \new_[9440]_  = \new_[833]_  | \new_[9439]_ ;
  assign \new_[9443]_  = \new_[829]_  | \new_[830]_ ;
  assign \new_[9446]_  = \new_[827]_  | \new_[828]_ ;
  assign \new_[9447]_  = \new_[9446]_  | \new_[9443]_ ;
  assign \new_[9448]_  = \new_[9447]_  | \new_[9440]_ ;
  assign \new_[9449]_  = \new_[9448]_  | \new_[9435]_ ;
  assign \new_[9453]_  = \new_[824]_  | \new_[825]_ ;
  assign \new_[9454]_  = \new_[826]_  | \new_[9453]_ ;
  assign \new_[9457]_  = \new_[822]_  | \new_[823]_ ;
  assign \new_[9460]_  = \new_[820]_  | \new_[821]_ ;
  assign \new_[9461]_  = \new_[9460]_  | \new_[9457]_ ;
  assign \new_[9462]_  = \new_[9461]_  | \new_[9454]_ ;
  assign \new_[9465]_  = \new_[818]_  | \new_[819]_ ;
  assign \new_[9468]_  = \new_[816]_  | \new_[817]_ ;
  assign \new_[9469]_  = \new_[9468]_  | \new_[9465]_ ;
  assign \new_[9472]_  = \new_[814]_  | \new_[815]_ ;
  assign \new_[9475]_  = \new_[812]_  | \new_[813]_ ;
  assign \new_[9476]_  = \new_[9475]_  | \new_[9472]_ ;
  assign \new_[9477]_  = \new_[9476]_  | \new_[9469]_ ;
  assign \new_[9478]_  = \new_[9477]_  | \new_[9462]_ ;
  assign \new_[9479]_  = \new_[9478]_  | \new_[9449]_ ;
  assign \new_[9480]_  = \new_[9479]_  | \new_[9422]_ ;
  assign \new_[9481]_  = \new_[9480]_  | \new_[9365]_ ;
  assign \new_[9485]_  = \new_[809]_  | \new_[810]_ ;
  assign \new_[9486]_  = \new_[811]_  | \new_[9485]_ ;
  assign \new_[9489]_  = \new_[807]_  | \new_[808]_ ;
  assign \new_[9492]_  = \new_[805]_  | \new_[806]_ ;
  assign \new_[9493]_  = \new_[9492]_  | \new_[9489]_ ;
  assign \new_[9494]_  = \new_[9493]_  | \new_[9486]_ ;
  assign \new_[9498]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[9499]_  = \new_[804]_  | \new_[9498]_ ;
  assign \new_[9502]_  = \new_[800]_  | \new_[801]_ ;
  assign \new_[9505]_  = \new_[798]_  | \new_[799]_ ;
  assign \new_[9506]_  = \new_[9505]_  | \new_[9502]_ ;
  assign \new_[9507]_  = \new_[9506]_  | \new_[9499]_ ;
  assign \new_[9508]_  = \new_[9507]_  | \new_[9494]_ ;
  assign \new_[9512]_  = \new_[795]_  | \new_[796]_ ;
  assign \new_[9513]_  = \new_[797]_  | \new_[9512]_ ;
  assign \new_[9516]_  = \new_[793]_  | \new_[794]_ ;
  assign \new_[9519]_  = \new_[791]_  | \new_[792]_ ;
  assign \new_[9520]_  = \new_[9519]_  | \new_[9516]_ ;
  assign \new_[9521]_  = \new_[9520]_  | \new_[9513]_ ;
  assign \new_[9524]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[9527]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[9528]_  = \new_[9527]_  | \new_[9524]_ ;
  assign \new_[9531]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[9534]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[9535]_  = \new_[9534]_  | \new_[9531]_ ;
  assign \new_[9536]_  = \new_[9535]_  | \new_[9528]_ ;
  assign \new_[9537]_  = \new_[9536]_  | \new_[9521]_ ;
  assign \new_[9538]_  = \new_[9537]_  | \new_[9508]_ ;
  assign \new_[9542]_  = \new_[780]_  | \new_[781]_ ;
  assign \new_[9543]_  = \new_[782]_  | \new_[9542]_ ;
  assign \new_[9546]_  = \new_[778]_  | \new_[779]_ ;
  assign \new_[9549]_  = \new_[776]_  | \new_[777]_ ;
  assign \new_[9550]_  = \new_[9549]_  | \new_[9546]_ ;
  assign \new_[9551]_  = \new_[9550]_  | \new_[9543]_ ;
  assign \new_[9555]_  = \new_[773]_  | \new_[774]_ ;
  assign \new_[9556]_  = \new_[775]_  | \new_[9555]_ ;
  assign \new_[9559]_  = \new_[771]_  | \new_[772]_ ;
  assign \new_[9562]_  = \new_[769]_  | \new_[770]_ ;
  assign \new_[9563]_  = \new_[9562]_  | \new_[9559]_ ;
  assign \new_[9564]_  = \new_[9563]_  | \new_[9556]_ ;
  assign \new_[9565]_  = \new_[9564]_  | \new_[9551]_ ;
  assign \new_[9569]_  = \new_[766]_  | \new_[767]_ ;
  assign \new_[9570]_  = \new_[768]_  | \new_[9569]_ ;
  assign \new_[9573]_  = \new_[764]_  | \new_[765]_ ;
  assign \new_[9576]_  = \new_[762]_  | \new_[763]_ ;
  assign \new_[9577]_  = \new_[9576]_  | \new_[9573]_ ;
  assign \new_[9578]_  = \new_[9577]_  | \new_[9570]_ ;
  assign \new_[9581]_  = \new_[760]_  | \new_[761]_ ;
  assign \new_[9584]_  = \new_[758]_  | \new_[759]_ ;
  assign \new_[9585]_  = \new_[9584]_  | \new_[9581]_ ;
  assign \new_[9588]_  = \new_[756]_  | \new_[757]_ ;
  assign \new_[9591]_  = \new_[754]_  | \new_[755]_ ;
  assign \new_[9592]_  = \new_[9591]_  | \new_[9588]_ ;
  assign \new_[9593]_  = \new_[9592]_  | \new_[9585]_ ;
  assign \new_[9594]_  = \new_[9593]_  | \new_[9578]_ ;
  assign \new_[9595]_  = \new_[9594]_  | \new_[9565]_ ;
  assign \new_[9596]_  = \new_[9595]_  | \new_[9538]_ ;
  assign \new_[9600]_  = \new_[751]_  | \new_[752]_ ;
  assign \new_[9601]_  = \new_[753]_  | \new_[9600]_ ;
  assign \new_[9604]_  = \new_[749]_  | \new_[750]_ ;
  assign \new_[9607]_  = \new_[747]_  | \new_[748]_ ;
  assign \new_[9608]_  = \new_[9607]_  | \new_[9604]_ ;
  assign \new_[9609]_  = \new_[9608]_  | \new_[9601]_ ;
  assign \new_[9613]_  = \new_[744]_  | \new_[745]_ ;
  assign \new_[9614]_  = \new_[746]_  | \new_[9613]_ ;
  assign \new_[9617]_  = \new_[742]_  | \new_[743]_ ;
  assign \new_[9620]_  = \new_[740]_  | \new_[741]_ ;
  assign \new_[9621]_  = \new_[9620]_  | \new_[9617]_ ;
  assign \new_[9622]_  = \new_[9621]_  | \new_[9614]_ ;
  assign \new_[9623]_  = \new_[9622]_  | \new_[9609]_ ;
  assign \new_[9627]_  = \new_[737]_  | \new_[738]_ ;
  assign \new_[9628]_  = \new_[739]_  | \new_[9627]_ ;
  assign \new_[9631]_  = \new_[735]_  | \new_[736]_ ;
  assign \new_[9634]_  = \new_[733]_  | \new_[734]_ ;
  assign \new_[9635]_  = \new_[9634]_  | \new_[9631]_ ;
  assign \new_[9636]_  = \new_[9635]_  | \new_[9628]_ ;
  assign \new_[9639]_  = \new_[731]_  | \new_[732]_ ;
  assign \new_[9642]_  = \new_[729]_  | \new_[730]_ ;
  assign \new_[9643]_  = \new_[9642]_  | \new_[9639]_ ;
  assign \new_[9646]_  = \new_[727]_  | \new_[728]_ ;
  assign \new_[9649]_  = \new_[725]_  | \new_[726]_ ;
  assign \new_[9650]_  = \new_[9649]_  | \new_[9646]_ ;
  assign \new_[9651]_  = \new_[9650]_  | \new_[9643]_ ;
  assign \new_[9652]_  = \new_[9651]_  | \new_[9636]_ ;
  assign \new_[9653]_  = \new_[9652]_  | \new_[9623]_ ;
  assign \new_[9657]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[9658]_  = \new_[724]_  | \new_[9657]_ ;
  assign \new_[9661]_  = \new_[720]_  | \new_[721]_ ;
  assign \new_[9664]_  = \new_[718]_  | \new_[719]_ ;
  assign \new_[9665]_  = \new_[9664]_  | \new_[9661]_ ;
  assign \new_[9666]_  = \new_[9665]_  | \new_[9658]_ ;
  assign \new_[9670]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[9671]_  = \new_[717]_  | \new_[9670]_ ;
  assign \new_[9674]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[9677]_  = \new_[711]_  | \new_[712]_ ;
  assign \new_[9678]_  = \new_[9677]_  | \new_[9674]_ ;
  assign \new_[9679]_  = \new_[9678]_  | \new_[9671]_ ;
  assign \new_[9680]_  = \new_[9679]_  | \new_[9666]_ ;
  assign \new_[9684]_  = \new_[708]_  | \new_[709]_ ;
  assign \new_[9685]_  = \new_[710]_  | \new_[9684]_ ;
  assign \new_[9688]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[9691]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[9692]_  = \new_[9691]_  | \new_[9688]_ ;
  assign \new_[9693]_  = \new_[9692]_  | \new_[9685]_ ;
  assign \new_[9696]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[9699]_  = \new_[700]_  | \new_[701]_ ;
  assign \new_[9700]_  = \new_[9699]_  | \new_[9696]_ ;
  assign \new_[9703]_  = \new_[698]_  | \new_[699]_ ;
  assign \new_[9706]_  = \new_[696]_  | \new_[697]_ ;
  assign \new_[9707]_  = \new_[9706]_  | \new_[9703]_ ;
  assign \new_[9708]_  = \new_[9707]_  | \new_[9700]_ ;
  assign \new_[9709]_  = \new_[9708]_  | \new_[9693]_ ;
  assign \new_[9710]_  = \new_[9709]_  | \new_[9680]_ ;
  assign \new_[9711]_  = \new_[9710]_  | \new_[9653]_ ;
  assign \new_[9712]_  = \new_[9711]_  | \new_[9596]_ ;
  assign \new_[9713]_  = \new_[9712]_  | \new_[9481]_ ;
  assign \new_[9717]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[9718]_  = \new_[695]_  | \new_[9717]_ ;
  assign \new_[9721]_  = \new_[691]_  | \new_[692]_ ;
  assign \new_[9724]_  = \new_[689]_  | \new_[690]_ ;
  assign \new_[9725]_  = \new_[9724]_  | \new_[9721]_ ;
  assign \new_[9726]_  = \new_[9725]_  | \new_[9718]_ ;
  assign \new_[9730]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[9731]_  = \new_[688]_  | \new_[9730]_ ;
  assign \new_[9734]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[9737]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[9738]_  = \new_[9737]_  | \new_[9734]_ ;
  assign \new_[9739]_  = \new_[9738]_  | \new_[9731]_ ;
  assign \new_[9740]_  = \new_[9739]_  | \new_[9726]_ ;
  assign \new_[9744]_  = \new_[679]_  | \new_[680]_ ;
  assign \new_[9745]_  = \new_[681]_  | \new_[9744]_ ;
  assign \new_[9748]_  = \new_[677]_  | \new_[678]_ ;
  assign \new_[9751]_  = \new_[675]_  | \new_[676]_ ;
  assign \new_[9752]_  = \new_[9751]_  | \new_[9748]_ ;
  assign \new_[9753]_  = \new_[9752]_  | \new_[9745]_ ;
  assign \new_[9756]_  = \new_[673]_  | \new_[674]_ ;
  assign \new_[9759]_  = \new_[671]_  | \new_[672]_ ;
  assign \new_[9760]_  = \new_[9759]_  | \new_[9756]_ ;
  assign \new_[9763]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[9766]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[9767]_  = \new_[9766]_  | \new_[9763]_ ;
  assign \new_[9768]_  = \new_[9767]_  | \new_[9760]_ ;
  assign \new_[9769]_  = \new_[9768]_  | \new_[9753]_ ;
  assign \new_[9770]_  = \new_[9769]_  | \new_[9740]_ ;
  assign \new_[9774]_  = \new_[664]_  | \new_[665]_ ;
  assign \new_[9775]_  = \new_[666]_  | \new_[9774]_ ;
  assign \new_[9778]_  = \new_[662]_  | \new_[663]_ ;
  assign \new_[9781]_  = \new_[660]_  | \new_[661]_ ;
  assign \new_[9782]_  = \new_[9781]_  | \new_[9778]_ ;
  assign \new_[9783]_  = \new_[9782]_  | \new_[9775]_ ;
  assign \new_[9787]_  = \new_[657]_  | \new_[658]_ ;
  assign \new_[9788]_  = \new_[659]_  | \new_[9787]_ ;
  assign \new_[9791]_  = \new_[655]_  | \new_[656]_ ;
  assign \new_[9794]_  = \new_[653]_  | \new_[654]_ ;
  assign \new_[9795]_  = \new_[9794]_  | \new_[9791]_ ;
  assign \new_[9796]_  = \new_[9795]_  | \new_[9788]_ ;
  assign \new_[9797]_  = \new_[9796]_  | \new_[9783]_ ;
  assign \new_[9801]_  = \new_[650]_  | \new_[651]_ ;
  assign \new_[9802]_  = \new_[652]_  | \new_[9801]_ ;
  assign \new_[9805]_  = \new_[648]_  | \new_[649]_ ;
  assign \new_[9808]_  = \new_[646]_  | \new_[647]_ ;
  assign \new_[9809]_  = \new_[9808]_  | \new_[9805]_ ;
  assign \new_[9810]_  = \new_[9809]_  | \new_[9802]_ ;
  assign \new_[9813]_  = \new_[644]_  | \new_[645]_ ;
  assign \new_[9816]_  = \new_[642]_  | \new_[643]_ ;
  assign \new_[9817]_  = \new_[9816]_  | \new_[9813]_ ;
  assign \new_[9820]_  = \new_[640]_  | \new_[641]_ ;
  assign \new_[9823]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[9824]_  = \new_[9823]_  | \new_[9820]_ ;
  assign \new_[9825]_  = \new_[9824]_  | \new_[9817]_ ;
  assign \new_[9826]_  = \new_[9825]_  | \new_[9810]_ ;
  assign \new_[9827]_  = \new_[9826]_  | \new_[9797]_ ;
  assign \new_[9828]_  = \new_[9827]_  | \new_[9770]_ ;
  assign \new_[9832]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[9833]_  = \new_[637]_  | \new_[9832]_ ;
  assign \new_[9836]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[9839]_  = \new_[631]_  | \new_[632]_ ;
  assign \new_[9840]_  = \new_[9839]_  | \new_[9836]_ ;
  assign \new_[9841]_  = \new_[9840]_  | \new_[9833]_ ;
  assign \new_[9845]_  = \new_[628]_  | \new_[629]_ ;
  assign \new_[9846]_  = \new_[630]_  | \new_[9845]_ ;
  assign \new_[9849]_  = \new_[626]_  | \new_[627]_ ;
  assign \new_[9852]_  = \new_[624]_  | \new_[625]_ ;
  assign \new_[9853]_  = \new_[9852]_  | \new_[9849]_ ;
  assign \new_[9854]_  = \new_[9853]_  | \new_[9846]_ ;
  assign \new_[9855]_  = \new_[9854]_  | \new_[9841]_ ;
  assign \new_[9859]_  = \new_[621]_  | \new_[622]_ ;
  assign \new_[9860]_  = \new_[623]_  | \new_[9859]_ ;
  assign \new_[9863]_  = \new_[619]_  | \new_[620]_ ;
  assign \new_[9866]_  = \new_[617]_  | \new_[618]_ ;
  assign \new_[9867]_  = \new_[9866]_  | \new_[9863]_ ;
  assign \new_[9868]_  = \new_[9867]_  | \new_[9860]_ ;
  assign \new_[9871]_  = \new_[615]_  | \new_[616]_ ;
  assign \new_[9874]_  = \new_[613]_  | \new_[614]_ ;
  assign \new_[9875]_  = \new_[9874]_  | \new_[9871]_ ;
  assign \new_[9878]_  = \new_[611]_  | \new_[612]_ ;
  assign \new_[9881]_  = \new_[609]_  | \new_[610]_ ;
  assign \new_[9882]_  = \new_[9881]_  | \new_[9878]_ ;
  assign \new_[9883]_  = \new_[9882]_  | \new_[9875]_ ;
  assign \new_[9884]_  = \new_[9883]_  | \new_[9868]_ ;
  assign \new_[9885]_  = \new_[9884]_  | \new_[9855]_ ;
  assign \new_[9889]_  = \new_[606]_  | \new_[607]_ ;
  assign \new_[9890]_  = \new_[608]_  | \new_[9889]_ ;
  assign \new_[9893]_  = \new_[604]_  | \new_[605]_ ;
  assign \new_[9896]_  = \new_[602]_  | \new_[603]_ ;
  assign \new_[9897]_  = \new_[9896]_  | \new_[9893]_ ;
  assign \new_[9898]_  = \new_[9897]_  | \new_[9890]_ ;
  assign \new_[9902]_  = \new_[599]_  | \new_[600]_ ;
  assign \new_[9903]_  = \new_[601]_  | \new_[9902]_ ;
  assign \new_[9906]_  = \new_[597]_  | \new_[598]_ ;
  assign \new_[9909]_  = \new_[595]_  | \new_[596]_ ;
  assign \new_[9910]_  = \new_[9909]_  | \new_[9906]_ ;
  assign \new_[9911]_  = \new_[9910]_  | \new_[9903]_ ;
  assign \new_[9912]_  = \new_[9911]_  | \new_[9898]_ ;
  assign \new_[9916]_  = \new_[592]_  | \new_[593]_ ;
  assign \new_[9917]_  = \new_[594]_  | \new_[9916]_ ;
  assign \new_[9920]_  = \new_[590]_  | \new_[591]_ ;
  assign \new_[9923]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[9924]_  = \new_[9923]_  | \new_[9920]_ ;
  assign \new_[9925]_  = \new_[9924]_  | \new_[9917]_ ;
  assign \new_[9928]_  = \new_[586]_  | \new_[587]_ ;
  assign \new_[9931]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[9932]_  = \new_[9931]_  | \new_[9928]_ ;
  assign \new_[9935]_  = \new_[582]_  | \new_[583]_ ;
  assign \new_[9938]_  = \new_[580]_  | \new_[581]_ ;
  assign \new_[9939]_  = \new_[9938]_  | \new_[9935]_ ;
  assign \new_[9940]_  = \new_[9939]_  | \new_[9932]_ ;
  assign \new_[9941]_  = \new_[9940]_  | \new_[9925]_ ;
  assign \new_[9942]_  = \new_[9941]_  | \new_[9912]_ ;
  assign \new_[9943]_  = \new_[9942]_  | \new_[9885]_ ;
  assign \new_[9944]_  = \new_[9943]_  | \new_[9828]_ ;
  assign \new_[9948]_  = \new_[577]_  | \new_[578]_ ;
  assign \new_[9949]_  = \new_[579]_  | \new_[9948]_ ;
  assign \new_[9952]_  = \new_[575]_  | \new_[576]_ ;
  assign \new_[9955]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[9956]_  = \new_[9955]_  | \new_[9952]_ ;
  assign \new_[9957]_  = \new_[9956]_  | \new_[9949]_ ;
  assign \new_[9961]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[9962]_  = \new_[572]_  | \new_[9961]_ ;
  assign \new_[9965]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[9968]_  = \new_[566]_  | \new_[567]_ ;
  assign \new_[9969]_  = \new_[9968]_  | \new_[9965]_ ;
  assign \new_[9970]_  = \new_[9969]_  | \new_[9962]_ ;
  assign \new_[9971]_  = \new_[9970]_  | \new_[9957]_ ;
  assign \new_[9975]_  = \new_[563]_  | \new_[564]_ ;
  assign \new_[9976]_  = \new_[565]_  | \new_[9975]_ ;
  assign \new_[9979]_  = \new_[561]_  | \new_[562]_ ;
  assign \new_[9982]_  = \new_[559]_  | \new_[560]_ ;
  assign \new_[9983]_  = \new_[9982]_  | \new_[9979]_ ;
  assign \new_[9984]_  = \new_[9983]_  | \new_[9976]_ ;
  assign \new_[9987]_  = \new_[557]_  | \new_[558]_ ;
  assign \new_[9990]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[9991]_  = \new_[9990]_  | \new_[9987]_ ;
  assign \new_[9994]_  = \new_[553]_  | \new_[554]_ ;
  assign \new_[9997]_  = \new_[551]_  | \new_[552]_ ;
  assign \new_[9998]_  = \new_[9997]_  | \new_[9994]_ ;
  assign \new_[9999]_  = \new_[9998]_  | \new_[9991]_ ;
  assign \new_[10000]_  = \new_[9999]_  | \new_[9984]_ ;
  assign \new_[10001]_  = \new_[10000]_  | \new_[9971]_ ;
  assign \new_[10005]_  = \new_[548]_  | \new_[549]_ ;
  assign \new_[10006]_  = \new_[550]_  | \new_[10005]_ ;
  assign \new_[10009]_  = \new_[546]_  | \new_[547]_ ;
  assign \new_[10012]_  = \new_[544]_  | \new_[545]_ ;
  assign \new_[10013]_  = \new_[10012]_  | \new_[10009]_ ;
  assign \new_[10014]_  = \new_[10013]_  | \new_[10006]_ ;
  assign \new_[10018]_  = \new_[541]_  | \new_[542]_ ;
  assign \new_[10019]_  = \new_[543]_  | \new_[10018]_ ;
  assign \new_[10022]_  = \new_[539]_  | \new_[540]_ ;
  assign \new_[10025]_  = \new_[537]_  | \new_[538]_ ;
  assign \new_[10026]_  = \new_[10025]_  | \new_[10022]_ ;
  assign \new_[10027]_  = \new_[10026]_  | \new_[10019]_ ;
  assign \new_[10028]_  = \new_[10027]_  | \new_[10014]_ ;
  assign \new_[10032]_  = \new_[534]_  | \new_[535]_ ;
  assign \new_[10033]_  = \new_[536]_  | \new_[10032]_ ;
  assign \new_[10036]_  = \new_[532]_  | \new_[533]_ ;
  assign \new_[10039]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[10040]_  = \new_[10039]_  | \new_[10036]_ ;
  assign \new_[10041]_  = \new_[10040]_  | \new_[10033]_ ;
  assign \new_[10044]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[10047]_  = \new_[526]_  | \new_[527]_ ;
  assign \new_[10048]_  = \new_[10047]_  | \new_[10044]_ ;
  assign \new_[10051]_  = \new_[524]_  | \new_[525]_ ;
  assign \new_[10054]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[10055]_  = \new_[10054]_  | \new_[10051]_ ;
  assign \new_[10056]_  = \new_[10055]_  | \new_[10048]_ ;
  assign \new_[10057]_  = \new_[10056]_  | \new_[10041]_ ;
  assign \new_[10058]_  = \new_[10057]_  | \new_[10028]_ ;
  assign \new_[10059]_  = \new_[10058]_  | \new_[10001]_ ;
  assign \new_[10063]_  = \new_[519]_  | \new_[520]_ ;
  assign \new_[10064]_  = \new_[521]_  | \new_[10063]_ ;
  assign \new_[10067]_  = \new_[517]_  | \new_[518]_ ;
  assign \new_[10070]_  = \new_[515]_  | \new_[516]_ ;
  assign \new_[10071]_  = \new_[10070]_  | \new_[10067]_ ;
  assign \new_[10072]_  = \new_[10071]_  | \new_[10064]_ ;
  assign \new_[10076]_  = \new_[512]_  | \new_[513]_ ;
  assign \new_[10077]_  = \new_[514]_  | \new_[10076]_ ;
  assign \new_[10080]_  = \new_[510]_  | \new_[511]_ ;
  assign \new_[10083]_  = \new_[508]_  | \new_[509]_ ;
  assign \new_[10084]_  = \new_[10083]_  | \new_[10080]_ ;
  assign \new_[10085]_  = \new_[10084]_  | \new_[10077]_ ;
  assign \new_[10086]_  = \new_[10085]_  | \new_[10072]_ ;
  assign \new_[10090]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[10091]_  = \new_[507]_  | \new_[10090]_ ;
  assign \new_[10094]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[10097]_  = \new_[501]_  | \new_[502]_ ;
  assign \new_[10098]_  = \new_[10097]_  | \new_[10094]_ ;
  assign \new_[10099]_  = \new_[10098]_  | \new_[10091]_ ;
  assign \new_[10102]_  = \new_[499]_  | \new_[500]_ ;
  assign \new_[10105]_  = \new_[497]_  | \new_[498]_ ;
  assign \new_[10106]_  = \new_[10105]_  | \new_[10102]_ ;
  assign \new_[10109]_  = \new_[495]_  | \new_[496]_ ;
  assign \new_[10112]_  = \new_[493]_  | \new_[494]_ ;
  assign \new_[10113]_  = \new_[10112]_  | \new_[10109]_ ;
  assign \new_[10114]_  = \new_[10113]_  | \new_[10106]_ ;
  assign \new_[10115]_  = \new_[10114]_  | \new_[10099]_ ;
  assign \new_[10116]_  = \new_[10115]_  | \new_[10086]_ ;
  assign \new_[10120]_  = \new_[490]_  | \new_[491]_ ;
  assign \new_[10121]_  = \new_[492]_  | \new_[10120]_ ;
  assign \new_[10124]_  = \new_[488]_  | \new_[489]_ ;
  assign \new_[10127]_  = \new_[486]_  | \new_[487]_ ;
  assign \new_[10128]_  = \new_[10127]_  | \new_[10124]_ ;
  assign \new_[10129]_  = \new_[10128]_  | \new_[10121]_ ;
  assign \new_[10133]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[10134]_  = \new_[485]_  | \new_[10133]_ ;
  assign \new_[10137]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[10140]_  = \new_[479]_  | \new_[480]_ ;
  assign \new_[10141]_  = \new_[10140]_  | \new_[10137]_ ;
  assign \new_[10142]_  = \new_[10141]_  | \new_[10134]_ ;
  assign \new_[10143]_  = \new_[10142]_  | \new_[10129]_ ;
  assign \new_[10147]_  = \new_[476]_  | \new_[477]_ ;
  assign \new_[10148]_  = \new_[478]_  | \new_[10147]_ ;
  assign \new_[10151]_  = \new_[474]_  | \new_[475]_ ;
  assign \new_[10154]_  = \new_[472]_  | \new_[473]_ ;
  assign \new_[10155]_  = \new_[10154]_  | \new_[10151]_ ;
  assign \new_[10156]_  = \new_[10155]_  | \new_[10148]_ ;
  assign \new_[10159]_  = \new_[470]_  | \new_[471]_ ;
  assign \new_[10162]_  = \new_[468]_  | \new_[469]_ ;
  assign \new_[10163]_  = \new_[10162]_  | \new_[10159]_ ;
  assign \new_[10166]_  = \new_[466]_  | \new_[467]_ ;
  assign \new_[10169]_  = \new_[464]_  | \new_[465]_ ;
  assign \new_[10170]_  = \new_[10169]_  | \new_[10166]_ ;
  assign \new_[10171]_  = \new_[10170]_  | \new_[10163]_ ;
  assign \new_[10172]_  = \new_[10171]_  | \new_[10156]_ ;
  assign \new_[10173]_  = \new_[10172]_  | \new_[10143]_ ;
  assign \new_[10174]_  = \new_[10173]_  | \new_[10116]_ ;
  assign \new_[10175]_  = \new_[10174]_  | \new_[10059]_ ;
  assign \new_[10176]_  = \new_[10175]_  | \new_[9944]_ ;
  assign \new_[10177]_  = \new_[10176]_  | \new_[9713]_ ;
  assign \new_[10181]_  = \new_[461]_  | \new_[462]_ ;
  assign \new_[10182]_  = \new_[463]_  | \new_[10181]_ ;
  assign \new_[10185]_  = \new_[459]_  | \new_[460]_ ;
  assign \new_[10188]_  = \new_[457]_  | \new_[458]_ ;
  assign \new_[10189]_  = \new_[10188]_  | \new_[10185]_ ;
  assign \new_[10190]_  = \new_[10189]_  | \new_[10182]_ ;
  assign \new_[10194]_  = \new_[454]_  | \new_[455]_ ;
  assign \new_[10195]_  = \new_[456]_  | \new_[10194]_ ;
  assign \new_[10198]_  = \new_[452]_  | \new_[453]_ ;
  assign \new_[10201]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[10202]_  = \new_[10201]_  | \new_[10198]_ ;
  assign \new_[10203]_  = \new_[10202]_  | \new_[10195]_ ;
  assign \new_[10204]_  = \new_[10203]_  | \new_[10190]_ ;
  assign \new_[10208]_  = \new_[447]_  | \new_[448]_ ;
  assign \new_[10209]_  = \new_[449]_  | \new_[10208]_ ;
  assign \new_[10212]_  = \new_[445]_  | \new_[446]_ ;
  assign \new_[10215]_  = \new_[443]_  | \new_[444]_ ;
  assign \new_[10216]_  = \new_[10215]_  | \new_[10212]_ ;
  assign \new_[10217]_  = \new_[10216]_  | \new_[10209]_ ;
  assign \new_[10221]_  = \new_[440]_  | \new_[441]_ ;
  assign \new_[10222]_  = \new_[442]_  | \new_[10221]_ ;
  assign \new_[10225]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[10228]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[10229]_  = \new_[10228]_  | \new_[10225]_ ;
  assign \new_[10230]_  = \new_[10229]_  | \new_[10222]_ ;
  assign \new_[10231]_  = \new_[10230]_  | \new_[10217]_ ;
  assign \new_[10232]_  = \new_[10231]_  | \new_[10204]_ ;
  assign \new_[10236]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[10237]_  = \new_[435]_  | \new_[10236]_ ;
  assign \new_[10240]_  = \new_[431]_  | \new_[432]_ ;
  assign \new_[10243]_  = \new_[429]_  | \new_[430]_ ;
  assign \new_[10244]_  = \new_[10243]_  | \new_[10240]_ ;
  assign \new_[10245]_  = \new_[10244]_  | \new_[10237]_ ;
  assign \new_[10249]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[10250]_  = \new_[428]_  | \new_[10249]_ ;
  assign \new_[10253]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[10256]_  = \new_[422]_  | \new_[423]_ ;
  assign \new_[10257]_  = \new_[10256]_  | \new_[10253]_ ;
  assign \new_[10258]_  = \new_[10257]_  | \new_[10250]_ ;
  assign \new_[10259]_  = \new_[10258]_  | \new_[10245]_ ;
  assign \new_[10263]_  = \new_[419]_  | \new_[420]_ ;
  assign \new_[10264]_  = \new_[421]_  | \new_[10263]_ ;
  assign \new_[10267]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[10270]_  = \new_[415]_  | \new_[416]_ ;
  assign \new_[10271]_  = \new_[10270]_  | \new_[10267]_ ;
  assign \new_[10272]_  = \new_[10271]_  | \new_[10264]_ ;
  assign \new_[10275]_  = \new_[413]_  | \new_[414]_ ;
  assign \new_[10278]_  = \new_[411]_  | \new_[412]_ ;
  assign \new_[10279]_  = \new_[10278]_  | \new_[10275]_ ;
  assign \new_[10282]_  = \new_[409]_  | \new_[410]_ ;
  assign \new_[10285]_  = \new_[407]_  | \new_[408]_ ;
  assign \new_[10286]_  = \new_[10285]_  | \new_[10282]_ ;
  assign \new_[10287]_  = \new_[10286]_  | \new_[10279]_ ;
  assign \new_[10288]_  = \new_[10287]_  | \new_[10272]_ ;
  assign \new_[10289]_  = \new_[10288]_  | \new_[10259]_ ;
  assign \new_[10290]_  = \new_[10289]_  | \new_[10232]_ ;
  assign \new_[10294]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[10295]_  = \new_[406]_  | \new_[10294]_ ;
  assign \new_[10298]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[10301]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[10302]_  = \new_[10301]_  | \new_[10298]_ ;
  assign \new_[10303]_  = \new_[10302]_  | \new_[10295]_ ;
  assign \new_[10307]_  = \new_[397]_  | \new_[398]_ ;
  assign \new_[10308]_  = \new_[399]_  | \new_[10307]_ ;
  assign \new_[10311]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[10314]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[10315]_  = \new_[10314]_  | \new_[10311]_ ;
  assign \new_[10316]_  = \new_[10315]_  | \new_[10308]_ ;
  assign \new_[10317]_  = \new_[10316]_  | \new_[10303]_ ;
  assign \new_[10321]_  = \new_[390]_  | \new_[391]_ ;
  assign \new_[10322]_  = \new_[392]_  | \new_[10321]_ ;
  assign \new_[10325]_  = \new_[388]_  | \new_[389]_ ;
  assign \new_[10328]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[10329]_  = \new_[10328]_  | \new_[10325]_ ;
  assign \new_[10330]_  = \new_[10329]_  | \new_[10322]_ ;
  assign \new_[10333]_  = \new_[384]_  | \new_[385]_ ;
  assign \new_[10336]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[10337]_  = \new_[10336]_  | \new_[10333]_ ;
  assign \new_[10340]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[10343]_  = \new_[378]_  | \new_[379]_ ;
  assign \new_[10344]_  = \new_[10343]_  | \new_[10340]_ ;
  assign \new_[10345]_  = \new_[10344]_  | \new_[10337]_ ;
  assign \new_[10346]_  = \new_[10345]_  | \new_[10330]_ ;
  assign \new_[10347]_  = \new_[10346]_  | \new_[10317]_ ;
  assign \new_[10351]_  = \new_[375]_  | \new_[376]_ ;
  assign \new_[10352]_  = \new_[377]_  | \new_[10351]_ ;
  assign \new_[10355]_  = \new_[373]_  | \new_[374]_ ;
  assign \new_[10358]_  = \new_[371]_  | \new_[372]_ ;
  assign \new_[10359]_  = \new_[10358]_  | \new_[10355]_ ;
  assign \new_[10360]_  = \new_[10359]_  | \new_[10352]_ ;
  assign \new_[10364]_  = \new_[368]_  | \new_[369]_ ;
  assign \new_[10365]_  = \new_[370]_  | \new_[10364]_ ;
  assign \new_[10368]_  = \new_[366]_  | \new_[367]_ ;
  assign \new_[10371]_  = \new_[364]_  | \new_[365]_ ;
  assign \new_[10372]_  = \new_[10371]_  | \new_[10368]_ ;
  assign \new_[10373]_  = \new_[10372]_  | \new_[10365]_ ;
  assign \new_[10374]_  = \new_[10373]_  | \new_[10360]_ ;
  assign \new_[10378]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[10379]_  = \new_[363]_  | \new_[10378]_ ;
  assign \new_[10382]_  = \new_[359]_  | \new_[360]_ ;
  assign \new_[10385]_  = \new_[357]_  | \new_[358]_ ;
  assign \new_[10386]_  = \new_[10385]_  | \new_[10382]_ ;
  assign \new_[10387]_  = \new_[10386]_  | \new_[10379]_ ;
  assign \new_[10390]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[10393]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[10394]_  = \new_[10393]_  | \new_[10390]_ ;
  assign \new_[10397]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[10400]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[10401]_  = \new_[10400]_  | \new_[10397]_ ;
  assign \new_[10402]_  = \new_[10401]_  | \new_[10394]_ ;
  assign \new_[10403]_  = \new_[10402]_  | \new_[10387]_ ;
  assign \new_[10404]_  = \new_[10403]_  | \new_[10374]_ ;
  assign \new_[10405]_  = \new_[10404]_  | \new_[10347]_ ;
  assign \new_[10406]_  = \new_[10405]_  | \new_[10290]_ ;
  assign \new_[10410]_  = \new_[346]_  | \new_[347]_ ;
  assign \new_[10411]_  = \new_[348]_  | \new_[10410]_ ;
  assign \new_[10414]_  = \new_[344]_  | \new_[345]_ ;
  assign \new_[10417]_  = \new_[342]_  | \new_[343]_ ;
  assign \new_[10418]_  = \new_[10417]_  | \new_[10414]_ ;
  assign \new_[10419]_  = \new_[10418]_  | \new_[10411]_ ;
  assign \new_[10423]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[10424]_  = \new_[341]_  | \new_[10423]_ ;
  assign \new_[10427]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[10430]_  = \new_[335]_  | \new_[336]_ ;
  assign \new_[10431]_  = \new_[10430]_  | \new_[10427]_ ;
  assign \new_[10432]_  = \new_[10431]_  | \new_[10424]_ ;
  assign \new_[10433]_  = \new_[10432]_  | \new_[10419]_ ;
  assign \new_[10437]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[10438]_  = \new_[334]_  | \new_[10437]_ ;
  assign \new_[10441]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[10444]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[10445]_  = \new_[10444]_  | \new_[10441]_ ;
  assign \new_[10446]_  = \new_[10445]_  | \new_[10438]_ ;
  assign \new_[10449]_  = \new_[326]_  | \new_[327]_ ;
  assign \new_[10452]_  = \new_[324]_  | \new_[325]_ ;
  assign \new_[10453]_  = \new_[10452]_  | \new_[10449]_ ;
  assign \new_[10456]_  = \new_[322]_  | \new_[323]_ ;
  assign \new_[10459]_  = \new_[320]_  | \new_[321]_ ;
  assign \new_[10460]_  = \new_[10459]_  | \new_[10456]_ ;
  assign \new_[10461]_  = \new_[10460]_  | \new_[10453]_ ;
  assign \new_[10462]_  = \new_[10461]_  | \new_[10446]_ ;
  assign \new_[10463]_  = \new_[10462]_  | \new_[10433]_ ;
  assign \new_[10467]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[10468]_  = \new_[319]_  | \new_[10467]_ ;
  assign \new_[10471]_  = \new_[315]_  | \new_[316]_ ;
  assign \new_[10474]_  = \new_[313]_  | \new_[314]_ ;
  assign \new_[10475]_  = \new_[10474]_  | \new_[10471]_ ;
  assign \new_[10476]_  = \new_[10475]_  | \new_[10468]_ ;
  assign \new_[10480]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[10481]_  = \new_[312]_  | \new_[10480]_ ;
  assign \new_[10484]_  = \new_[308]_  | \new_[309]_ ;
  assign \new_[10487]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[10488]_  = \new_[10487]_  | \new_[10484]_ ;
  assign \new_[10489]_  = \new_[10488]_  | \new_[10481]_ ;
  assign \new_[10490]_  = \new_[10489]_  | \new_[10476]_ ;
  assign \new_[10494]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[10495]_  = \new_[305]_  | \new_[10494]_ ;
  assign \new_[10498]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[10501]_  = \new_[299]_  | \new_[300]_ ;
  assign \new_[10502]_  = \new_[10501]_  | \new_[10498]_ ;
  assign \new_[10503]_  = \new_[10502]_  | \new_[10495]_ ;
  assign \new_[10506]_  = \new_[297]_  | \new_[298]_ ;
  assign \new_[10509]_  = \new_[295]_  | \new_[296]_ ;
  assign \new_[10510]_  = \new_[10509]_  | \new_[10506]_ ;
  assign \new_[10513]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[10516]_  = \new_[291]_  | \new_[292]_ ;
  assign \new_[10517]_  = \new_[10516]_  | \new_[10513]_ ;
  assign \new_[10518]_  = \new_[10517]_  | \new_[10510]_ ;
  assign \new_[10519]_  = \new_[10518]_  | \new_[10503]_ ;
  assign \new_[10520]_  = \new_[10519]_  | \new_[10490]_ ;
  assign \new_[10521]_  = \new_[10520]_  | \new_[10463]_ ;
  assign \new_[10525]_  = \new_[288]_  | \new_[289]_ ;
  assign \new_[10526]_  = \new_[290]_  | \new_[10525]_ ;
  assign \new_[10529]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[10532]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[10533]_  = \new_[10532]_  | \new_[10529]_ ;
  assign \new_[10534]_  = \new_[10533]_  | \new_[10526]_ ;
  assign \new_[10538]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[10539]_  = \new_[283]_  | \new_[10538]_ ;
  assign \new_[10542]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[10545]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[10546]_  = \new_[10545]_  | \new_[10542]_ ;
  assign \new_[10547]_  = \new_[10546]_  | \new_[10539]_ ;
  assign \new_[10548]_  = \new_[10547]_  | \new_[10534]_ ;
  assign \new_[10552]_  = \new_[274]_  | \new_[275]_ ;
  assign \new_[10553]_  = \new_[276]_  | \new_[10552]_ ;
  assign \new_[10556]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[10559]_  = \new_[270]_  | \new_[271]_ ;
  assign \new_[10560]_  = \new_[10559]_  | \new_[10556]_ ;
  assign \new_[10561]_  = \new_[10560]_  | \new_[10553]_ ;
  assign \new_[10564]_  = \new_[268]_  | \new_[269]_ ;
  assign \new_[10567]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[10568]_  = \new_[10567]_  | \new_[10564]_ ;
  assign \new_[10571]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[10574]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[10575]_  = \new_[10574]_  | \new_[10571]_ ;
  assign \new_[10576]_  = \new_[10575]_  | \new_[10568]_ ;
  assign \new_[10577]_  = \new_[10576]_  | \new_[10561]_ ;
  assign \new_[10578]_  = \new_[10577]_  | \new_[10548]_ ;
  assign \new_[10582]_  = \new_[259]_  | \new_[260]_ ;
  assign \new_[10583]_  = \new_[261]_  | \new_[10582]_ ;
  assign \new_[10586]_  = \new_[257]_  | \new_[258]_ ;
  assign \new_[10589]_  = \new_[255]_  | \new_[256]_ ;
  assign \new_[10590]_  = \new_[10589]_  | \new_[10586]_ ;
  assign \new_[10591]_  = \new_[10590]_  | \new_[10583]_ ;
  assign \new_[10595]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[10596]_  = \new_[254]_  | \new_[10595]_ ;
  assign \new_[10599]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[10602]_  = \new_[248]_  | \new_[249]_ ;
  assign \new_[10603]_  = \new_[10602]_  | \new_[10599]_ ;
  assign \new_[10604]_  = \new_[10603]_  | \new_[10596]_ ;
  assign \new_[10605]_  = \new_[10604]_  | \new_[10591]_ ;
  assign \new_[10609]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[10610]_  = \new_[247]_  | \new_[10609]_ ;
  assign \new_[10613]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[10616]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[10617]_  = \new_[10616]_  | \new_[10613]_ ;
  assign \new_[10618]_  = \new_[10617]_  | \new_[10610]_ ;
  assign \new_[10621]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[10624]_  = \new_[237]_  | \new_[238]_ ;
  assign \new_[10625]_  = \new_[10624]_  | \new_[10621]_ ;
  assign \new_[10628]_  = \new_[235]_  | \new_[236]_ ;
  assign \new_[10631]_  = \new_[233]_  | \new_[234]_ ;
  assign \new_[10632]_  = \new_[10631]_  | \new_[10628]_ ;
  assign \new_[10633]_  = \new_[10632]_  | \new_[10625]_ ;
  assign \new_[10634]_  = \new_[10633]_  | \new_[10618]_ ;
  assign \new_[10635]_  = \new_[10634]_  | \new_[10605]_ ;
  assign \new_[10636]_  = \new_[10635]_  | \new_[10578]_ ;
  assign \new_[10637]_  = \new_[10636]_  | \new_[10521]_ ;
  assign \new_[10638]_  = \new_[10637]_  | \new_[10406]_ ;
  assign \new_[10642]_  = \new_[230]_  | \new_[231]_ ;
  assign \new_[10643]_  = \new_[232]_  | \new_[10642]_ ;
  assign \new_[10646]_  = \new_[228]_  | \new_[229]_ ;
  assign \new_[10649]_  = \new_[226]_  | \new_[227]_ ;
  assign \new_[10650]_  = \new_[10649]_  | \new_[10646]_ ;
  assign \new_[10651]_  = \new_[10650]_  | \new_[10643]_ ;
  assign \new_[10655]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[10656]_  = \new_[225]_  | \new_[10655]_ ;
  assign \new_[10659]_  = \new_[221]_  | \new_[222]_ ;
  assign \new_[10662]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[10663]_  = \new_[10662]_  | \new_[10659]_ ;
  assign \new_[10664]_  = \new_[10663]_  | \new_[10656]_ ;
  assign \new_[10665]_  = \new_[10664]_  | \new_[10651]_ ;
  assign \new_[10669]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[10670]_  = \new_[218]_  | \new_[10669]_ ;
  assign \new_[10673]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[10676]_  = \new_[212]_  | \new_[213]_ ;
  assign \new_[10677]_  = \new_[10676]_  | \new_[10673]_ ;
  assign \new_[10678]_  = \new_[10677]_  | \new_[10670]_ ;
  assign \new_[10681]_  = \new_[210]_  | \new_[211]_ ;
  assign \new_[10684]_  = \new_[208]_  | \new_[209]_ ;
  assign \new_[10685]_  = \new_[10684]_  | \new_[10681]_ ;
  assign \new_[10688]_  = \new_[206]_  | \new_[207]_ ;
  assign \new_[10691]_  = \new_[204]_  | \new_[205]_ ;
  assign \new_[10692]_  = \new_[10691]_  | \new_[10688]_ ;
  assign \new_[10693]_  = \new_[10692]_  | \new_[10685]_ ;
  assign \new_[10694]_  = \new_[10693]_  | \new_[10678]_ ;
  assign \new_[10695]_  = \new_[10694]_  | \new_[10665]_ ;
  assign \new_[10699]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[10700]_  = \new_[203]_  | \new_[10699]_ ;
  assign \new_[10703]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[10706]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[10707]_  = \new_[10706]_  | \new_[10703]_ ;
  assign \new_[10708]_  = \new_[10707]_  | \new_[10700]_ ;
  assign \new_[10712]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[10713]_  = \new_[196]_  | \new_[10712]_ ;
  assign \new_[10716]_  = \new_[192]_  | \new_[193]_ ;
  assign \new_[10719]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[10720]_  = \new_[10719]_  | \new_[10716]_ ;
  assign \new_[10721]_  = \new_[10720]_  | \new_[10713]_ ;
  assign \new_[10722]_  = \new_[10721]_  | \new_[10708]_ ;
  assign \new_[10726]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[10727]_  = \new_[189]_  | \new_[10726]_ ;
  assign \new_[10730]_  = \new_[185]_  | \new_[186]_ ;
  assign \new_[10733]_  = \new_[183]_  | \new_[184]_ ;
  assign \new_[10734]_  = \new_[10733]_  | \new_[10730]_ ;
  assign \new_[10735]_  = \new_[10734]_  | \new_[10727]_ ;
  assign \new_[10738]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[10741]_  = \new_[179]_  | \new_[180]_ ;
  assign \new_[10742]_  = \new_[10741]_  | \new_[10738]_ ;
  assign \new_[10745]_  = \new_[177]_  | \new_[178]_ ;
  assign \new_[10748]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[10749]_  = \new_[10748]_  | \new_[10745]_ ;
  assign \new_[10750]_  = \new_[10749]_  | \new_[10742]_ ;
  assign \new_[10751]_  = \new_[10750]_  | \new_[10735]_ ;
  assign \new_[10752]_  = \new_[10751]_  | \new_[10722]_ ;
  assign \new_[10753]_  = \new_[10752]_  | \new_[10695]_ ;
  assign \new_[10757]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[10758]_  = \new_[174]_  | \new_[10757]_ ;
  assign \new_[10761]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[10764]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[10765]_  = \new_[10764]_  | \new_[10761]_ ;
  assign \new_[10766]_  = \new_[10765]_  | \new_[10758]_ ;
  assign \new_[10770]_  = \new_[165]_  | \new_[166]_ ;
  assign \new_[10771]_  = \new_[167]_  | \new_[10770]_ ;
  assign \new_[10774]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[10777]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[10778]_  = \new_[10777]_  | \new_[10774]_ ;
  assign \new_[10779]_  = \new_[10778]_  | \new_[10771]_ ;
  assign \new_[10780]_  = \new_[10779]_  | \new_[10766]_ ;
  assign \new_[10784]_  = \new_[158]_  | \new_[159]_ ;
  assign \new_[10785]_  = \new_[160]_  | \new_[10784]_ ;
  assign \new_[10788]_  = \new_[156]_  | \new_[157]_ ;
  assign \new_[10791]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[10792]_  = \new_[10791]_  | \new_[10788]_ ;
  assign \new_[10793]_  = \new_[10792]_  | \new_[10785]_ ;
  assign \new_[10796]_  = \new_[152]_  | \new_[153]_ ;
  assign \new_[10799]_  = \new_[150]_  | \new_[151]_ ;
  assign \new_[10800]_  = \new_[10799]_  | \new_[10796]_ ;
  assign \new_[10803]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[10806]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[10807]_  = \new_[10806]_  | \new_[10803]_ ;
  assign \new_[10808]_  = \new_[10807]_  | \new_[10800]_ ;
  assign \new_[10809]_  = \new_[10808]_  | \new_[10793]_ ;
  assign \new_[10810]_  = \new_[10809]_  | \new_[10780]_ ;
  assign \new_[10814]_  = \new_[143]_  | \new_[144]_ ;
  assign \new_[10815]_  = \new_[145]_  | \new_[10814]_ ;
  assign \new_[10818]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[10821]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[10822]_  = \new_[10821]_  | \new_[10818]_ ;
  assign \new_[10823]_  = \new_[10822]_  | \new_[10815]_ ;
  assign \new_[10827]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[10828]_  = \new_[138]_  | \new_[10827]_ ;
  assign \new_[10831]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[10834]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[10835]_  = \new_[10834]_  | \new_[10831]_ ;
  assign \new_[10836]_  = \new_[10835]_  | \new_[10828]_ ;
  assign \new_[10837]_  = \new_[10836]_  | \new_[10823]_ ;
  assign \new_[10841]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[10842]_  = \new_[131]_  | \new_[10841]_ ;
  assign \new_[10845]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[10848]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[10849]_  = \new_[10848]_  | \new_[10845]_ ;
  assign \new_[10850]_  = \new_[10849]_  | \new_[10842]_ ;
  assign \new_[10853]_  = \new_[123]_  | \new_[124]_ ;
  assign \new_[10856]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[10857]_  = \new_[10856]_  | \new_[10853]_ ;
  assign \new_[10860]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[10863]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[10864]_  = \new_[10863]_  | \new_[10860]_ ;
  assign \new_[10865]_  = \new_[10864]_  | \new_[10857]_ ;
  assign \new_[10866]_  = \new_[10865]_  | \new_[10850]_ ;
  assign \new_[10867]_  = \new_[10866]_  | \new_[10837]_ ;
  assign \new_[10868]_  = \new_[10867]_  | \new_[10810]_ ;
  assign \new_[10869]_  = \new_[10868]_  | \new_[10753]_ ;
  assign \new_[10873]_  = \new_[114]_  | \new_[115]_ ;
  assign \new_[10874]_  = \new_[116]_  | \new_[10873]_ ;
  assign \new_[10877]_  = \new_[112]_  | \new_[113]_ ;
  assign \new_[10880]_  = \new_[110]_  | \new_[111]_ ;
  assign \new_[10881]_  = \new_[10880]_  | \new_[10877]_ ;
  assign \new_[10882]_  = \new_[10881]_  | \new_[10874]_ ;
  assign \new_[10886]_  = \new_[107]_  | \new_[108]_ ;
  assign \new_[10887]_  = \new_[109]_  | \new_[10886]_ ;
  assign \new_[10890]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[10893]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[10894]_  = \new_[10893]_  | \new_[10890]_ ;
  assign \new_[10895]_  = \new_[10894]_  | \new_[10887]_ ;
  assign \new_[10896]_  = \new_[10895]_  | \new_[10882]_ ;
  assign \new_[10900]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[10901]_  = \new_[102]_  | \new_[10900]_ ;
  assign \new_[10904]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[10907]_  = \new_[96]_  | \new_[97]_ ;
  assign \new_[10908]_  = \new_[10907]_  | \new_[10904]_ ;
  assign \new_[10909]_  = \new_[10908]_  | \new_[10901]_ ;
  assign \new_[10912]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[10915]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[10916]_  = \new_[10915]_  | \new_[10912]_ ;
  assign \new_[10919]_  = \new_[90]_  | \new_[91]_ ;
  assign \new_[10922]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[10923]_  = \new_[10922]_  | \new_[10919]_ ;
  assign \new_[10924]_  = \new_[10923]_  | \new_[10916]_ ;
  assign \new_[10925]_  = \new_[10924]_  | \new_[10909]_ ;
  assign \new_[10926]_  = \new_[10925]_  | \new_[10896]_ ;
  assign \new_[10930]_  = \new_[85]_  | \new_[86]_ ;
  assign \new_[10931]_  = \new_[87]_  | \new_[10930]_ ;
  assign \new_[10934]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[10937]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[10938]_  = \new_[10937]_  | \new_[10934]_ ;
  assign \new_[10939]_  = \new_[10938]_  | \new_[10931]_ ;
  assign \new_[10943]_  = \new_[78]_  | \new_[79]_ ;
  assign \new_[10944]_  = \new_[80]_  | \new_[10943]_ ;
  assign \new_[10947]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[10950]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[10951]_  = \new_[10950]_  | \new_[10947]_ ;
  assign \new_[10952]_  = \new_[10951]_  | \new_[10944]_ ;
  assign \new_[10953]_  = \new_[10952]_  | \new_[10939]_ ;
  assign \new_[10957]_  = \new_[71]_  | \new_[72]_ ;
  assign \new_[10958]_  = \new_[73]_  | \new_[10957]_ ;
  assign \new_[10961]_  = \new_[69]_  | \new_[70]_ ;
  assign \new_[10964]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[10965]_  = \new_[10964]_  | \new_[10961]_ ;
  assign \new_[10966]_  = \new_[10965]_  | \new_[10958]_ ;
  assign \new_[10969]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[10972]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[10973]_  = \new_[10972]_  | \new_[10969]_ ;
  assign \new_[10976]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[10979]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[10980]_  = \new_[10979]_  | \new_[10976]_ ;
  assign \new_[10981]_  = \new_[10980]_  | \new_[10973]_ ;
  assign \new_[10982]_  = \new_[10981]_  | \new_[10966]_ ;
  assign \new_[10983]_  = \new_[10982]_  | \new_[10953]_ ;
  assign \new_[10984]_  = \new_[10983]_  | \new_[10926]_ ;
  assign \new_[10988]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[10989]_  = \new_[58]_  | \new_[10988]_ ;
  assign \new_[10992]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[10995]_  = \new_[52]_  | \new_[53]_ ;
  assign \new_[10996]_  = \new_[10995]_  | \new_[10992]_ ;
  assign \new_[10997]_  = \new_[10996]_  | \new_[10989]_ ;
  assign \new_[11001]_  = \new_[49]_  | \new_[50]_ ;
  assign \new_[11002]_  = \new_[51]_  | \new_[11001]_ ;
  assign \new_[11005]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[11008]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[11009]_  = \new_[11008]_  | \new_[11005]_ ;
  assign \new_[11010]_  = \new_[11009]_  | \new_[11002]_ ;
  assign \new_[11011]_  = \new_[11010]_  | \new_[10997]_ ;
  assign \new_[11015]_  = \new_[42]_  | \new_[43]_ ;
  assign \new_[11016]_  = \new_[44]_  | \new_[11015]_ ;
  assign \new_[11019]_  = \new_[40]_  | \new_[41]_ ;
  assign \new_[11022]_  = \new_[38]_  | \new_[39]_ ;
  assign \new_[11023]_  = \new_[11022]_  | \new_[11019]_ ;
  assign \new_[11024]_  = \new_[11023]_  | \new_[11016]_ ;
  assign \new_[11027]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[11030]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[11031]_  = \new_[11030]_  | \new_[11027]_ ;
  assign \new_[11034]_  = \new_[32]_  | \new_[33]_ ;
  assign \new_[11037]_  = \new_[30]_  | \new_[31]_ ;
  assign \new_[11038]_  = \new_[11037]_  | \new_[11034]_ ;
  assign \new_[11039]_  = \new_[11038]_  | \new_[11031]_ ;
  assign \new_[11040]_  = \new_[11039]_  | \new_[11024]_ ;
  assign \new_[11041]_  = \new_[11040]_  | \new_[11011]_ ;
  assign \new_[11045]_  = \new_[27]_  | \new_[28]_ ;
  assign \new_[11046]_  = \new_[29]_  | \new_[11045]_ ;
  assign \new_[11049]_  = \new_[25]_  | \new_[26]_ ;
  assign \new_[11052]_  = \new_[23]_  | \new_[24]_ ;
  assign \new_[11053]_  = \new_[11052]_  | \new_[11049]_ ;
  assign \new_[11054]_  = \new_[11053]_  | \new_[11046]_ ;
  assign \new_[11058]_  = \new_[20]_  | \new_[21]_ ;
  assign \new_[11059]_  = \new_[22]_  | \new_[11058]_ ;
  assign \new_[11062]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[11065]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[11066]_  = \new_[11065]_  | \new_[11062]_ ;
  assign \new_[11067]_  = \new_[11066]_  | \new_[11059]_ ;
  assign \new_[11068]_  = \new_[11067]_  | \new_[11054]_ ;
  assign \new_[11072]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[11073]_  = \new_[15]_  | \new_[11072]_ ;
  assign \new_[11076]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[11079]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[11080]_  = \new_[11079]_  | \new_[11076]_ ;
  assign \new_[11081]_  = \new_[11080]_  | \new_[11073]_ ;
  assign \new_[11084]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[11087]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[11088]_  = \new_[11087]_  | \new_[11084]_ ;
  assign \new_[11091]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[11094]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[11095]_  = \new_[11094]_  | \new_[11091]_ ;
  assign \new_[11096]_  = \new_[11095]_  | \new_[11088]_ ;
  assign \new_[11097]_  = \new_[11096]_  | \new_[11081]_ ;
  assign \new_[11098]_  = \new_[11097]_  | \new_[11068]_ ;
  assign \new_[11099]_  = \new_[11098]_  | \new_[11041]_ ;
  assign \new_[11100]_  = \new_[11099]_  | \new_[10984]_ ;
  assign \new_[11101]_  = \new_[11100]_  | \new_[10869]_ ;
  assign \new_[11102]_  = \new_[11101]_  | \new_[10638]_ ;
  assign \new_[11103]_  = \new_[11102]_  | \new_[10177]_ ;
  assign \new_[11104]_  = \new_[11103]_  | \new_[9252]_ ;
  assign \new_[11107]_  = A200 & ~A199;
  assign \new_[11110]_  = A202 & A201;
  assign \new_[11111]_  = \new_[11110]_  & \new_[11107]_ ;
  assign \new_[11114]_  = A233 & ~A232;
  assign \new_[11117]_  = A235 & A234;
  assign \new_[11118]_  = \new_[11117]_  & \new_[11114]_ ;
  assign \new_[11121]_  = A200 & ~A199;
  assign \new_[11124]_  = A202 & A201;
  assign \new_[11125]_  = \new_[11124]_  & \new_[11121]_ ;
  assign \new_[11128]_  = A233 & ~A232;
  assign \new_[11131]_  = A236 & A234;
  assign \new_[11132]_  = \new_[11131]_  & \new_[11128]_ ;
  assign \new_[11135]_  = A200 & ~A199;
  assign \new_[11138]_  = A202 & A201;
  assign \new_[11139]_  = \new_[11138]_  & \new_[11135]_ ;
  assign \new_[11142]_  = ~A233 & A232;
  assign \new_[11145]_  = A235 & A234;
  assign \new_[11146]_  = \new_[11145]_  & \new_[11142]_ ;
  assign \new_[11149]_  = A200 & ~A199;
  assign \new_[11152]_  = A202 & A201;
  assign \new_[11153]_  = \new_[11152]_  & \new_[11149]_ ;
  assign \new_[11156]_  = ~A233 & A232;
  assign \new_[11159]_  = A236 & A234;
  assign \new_[11160]_  = \new_[11159]_  & \new_[11156]_ ;
  assign \new_[11163]_  = A200 & ~A199;
  assign \new_[11166]_  = A203 & A201;
  assign \new_[11167]_  = \new_[11166]_  & \new_[11163]_ ;
  assign \new_[11170]_  = A233 & ~A232;
  assign \new_[11173]_  = A235 & A234;
  assign \new_[11174]_  = \new_[11173]_  & \new_[11170]_ ;
  assign \new_[11177]_  = A200 & ~A199;
  assign \new_[11180]_  = A203 & A201;
  assign \new_[11181]_  = \new_[11180]_  & \new_[11177]_ ;
  assign \new_[11184]_  = A233 & ~A232;
  assign \new_[11187]_  = A236 & A234;
  assign \new_[11188]_  = \new_[11187]_  & \new_[11184]_ ;
  assign \new_[11191]_  = A200 & ~A199;
  assign \new_[11194]_  = A203 & A201;
  assign \new_[11195]_  = \new_[11194]_  & \new_[11191]_ ;
  assign \new_[11198]_  = ~A233 & A232;
  assign \new_[11201]_  = A235 & A234;
  assign \new_[11202]_  = \new_[11201]_  & \new_[11198]_ ;
  assign \new_[11205]_  = A200 & ~A199;
  assign \new_[11208]_  = A203 & A201;
  assign \new_[11209]_  = \new_[11208]_  & \new_[11205]_ ;
  assign \new_[11212]_  = ~A233 & A232;
  assign \new_[11215]_  = A236 & A234;
  assign \new_[11216]_  = \new_[11215]_  & \new_[11212]_ ;
  assign \new_[11219]_  = ~A200 & A199;
  assign \new_[11222]_  = A202 & A201;
  assign \new_[11223]_  = \new_[11222]_  & \new_[11219]_ ;
  assign \new_[11226]_  = A233 & ~A232;
  assign \new_[11229]_  = A235 & A234;
  assign \new_[11230]_  = \new_[11229]_  & \new_[11226]_ ;
  assign \new_[11233]_  = ~A200 & A199;
  assign \new_[11236]_  = A202 & A201;
  assign \new_[11237]_  = \new_[11236]_  & \new_[11233]_ ;
  assign \new_[11240]_  = A233 & ~A232;
  assign \new_[11243]_  = A236 & A234;
  assign \new_[11244]_  = \new_[11243]_  & \new_[11240]_ ;
  assign \new_[11247]_  = ~A200 & A199;
  assign \new_[11250]_  = A202 & A201;
  assign \new_[11251]_  = \new_[11250]_  & \new_[11247]_ ;
  assign \new_[11254]_  = ~A233 & A232;
  assign \new_[11257]_  = A235 & A234;
  assign \new_[11258]_  = \new_[11257]_  & \new_[11254]_ ;
  assign \new_[11261]_  = ~A200 & A199;
  assign \new_[11264]_  = A202 & A201;
  assign \new_[11265]_  = \new_[11264]_  & \new_[11261]_ ;
  assign \new_[11268]_  = ~A233 & A232;
  assign \new_[11271]_  = A236 & A234;
  assign \new_[11272]_  = \new_[11271]_  & \new_[11268]_ ;
  assign \new_[11275]_  = ~A200 & A199;
  assign \new_[11278]_  = A203 & A201;
  assign \new_[11279]_  = \new_[11278]_  & \new_[11275]_ ;
  assign \new_[11282]_  = A233 & ~A232;
  assign \new_[11285]_  = A235 & A234;
  assign \new_[11286]_  = \new_[11285]_  & \new_[11282]_ ;
  assign \new_[11289]_  = ~A200 & A199;
  assign \new_[11292]_  = A203 & A201;
  assign \new_[11293]_  = \new_[11292]_  & \new_[11289]_ ;
  assign \new_[11296]_  = A233 & ~A232;
  assign \new_[11299]_  = A236 & A234;
  assign \new_[11300]_  = \new_[11299]_  & \new_[11296]_ ;
  assign \new_[11303]_  = ~A200 & A199;
  assign \new_[11306]_  = A203 & A201;
  assign \new_[11307]_  = \new_[11306]_  & \new_[11303]_ ;
  assign \new_[11310]_  = ~A233 & A232;
  assign \new_[11313]_  = A235 & A234;
  assign \new_[11314]_  = \new_[11313]_  & \new_[11310]_ ;
  assign \new_[11317]_  = ~A200 & A199;
  assign \new_[11320]_  = A203 & A201;
  assign \new_[11321]_  = \new_[11320]_  & \new_[11317]_ ;
  assign \new_[11324]_  = ~A233 & A232;
  assign \new_[11327]_  = A236 & A234;
  assign \new_[11328]_  = \new_[11327]_  & \new_[11324]_ ;
  assign \new_[11331]_  = A168 & ~A170;
  assign \new_[11334]_  = ~A166 & A167;
  assign \new_[11335]_  = \new_[11334]_  & \new_[11331]_ ;
  assign \new_[11338]_  = A233 & ~A232;
  assign \new_[11341]_  = A235 & A234;
  assign \new_[11342]_  = \new_[11341]_  & \new_[11338]_ ;
  assign \new_[11345]_  = A168 & ~A170;
  assign \new_[11348]_  = ~A166 & A167;
  assign \new_[11349]_  = \new_[11348]_  & \new_[11345]_ ;
  assign \new_[11352]_  = A233 & ~A232;
  assign \new_[11355]_  = A236 & A234;
  assign \new_[11356]_  = \new_[11355]_  & \new_[11352]_ ;
  assign \new_[11359]_  = A168 & ~A170;
  assign \new_[11362]_  = ~A166 & A167;
  assign \new_[11363]_  = \new_[11362]_  & \new_[11359]_ ;
  assign \new_[11366]_  = ~A233 & A232;
  assign \new_[11369]_  = A235 & A234;
  assign \new_[11370]_  = \new_[11369]_  & \new_[11366]_ ;
  assign \new_[11373]_  = A168 & ~A170;
  assign \new_[11376]_  = ~A166 & A167;
  assign \new_[11377]_  = \new_[11376]_  & \new_[11373]_ ;
  assign \new_[11380]_  = ~A233 & A232;
  assign \new_[11383]_  = A236 & A234;
  assign \new_[11384]_  = \new_[11383]_  & \new_[11380]_ ;
  assign \new_[11387]_  = A168 & ~A170;
  assign \new_[11390]_  = A166 & ~A167;
  assign \new_[11391]_  = \new_[11390]_  & \new_[11387]_ ;
  assign \new_[11394]_  = A233 & ~A232;
  assign \new_[11397]_  = A235 & A234;
  assign \new_[11398]_  = \new_[11397]_  & \new_[11394]_ ;
  assign \new_[11401]_  = A168 & ~A170;
  assign \new_[11404]_  = A166 & ~A167;
  assign \new_[11405]_  = \new_[11404]_  & \new_[11401]_ ;
  assign \new_[11408]_  = A233 & ~A232;
  assign \new_[11411]_  = A236 & A234;
  assign \new_[11412]_  = \new_[11411]_  & \new_[11408]_ ;
  assign \new_[11415]_  = A168 & ~A170;
  assign \new_[11418]_  = A166 & ~A167;
  assign \new_[11419]_  = \new_[11418]_  & \new_[11415]_ ;
  assign \new_[11422]_  = ~A233 & A232;
  assign \new_[11425]_  = A235 & A234;
  assign \new_[11426]_  = \new_[11425]_  & \new_[11422]_ ;
  assign \new_[11429]_  = A168 & ~A170;
  assign \new_[11432]_  = A166 & ~A167;
  assign \new_[11433]_  = \new_[11432]_  & \new_[11429]_ ;
  assign \new_[11436]_  = ~A233 & A232;
  assign \new_[11439]_  = A236 & A234;
  assign \new_[11440]_  = \new_[11439]_  & \new_[11436]_ ;
  assign \new_[11443]_  = A168 & A169;
  assign \new_[11446]_  = ~A166 & A167;
  assign \new_[11447]_  = \new_[11446]_  & \new_[11443]_ ;
  assign \new_[11450]_  = A233 & ~A232;
  assign \new_[11453]_  = A235 & A234;
  assign \new_[11454]_  = \new_[11453]_  & \new_[11450]_ ;
  assign \new_[11457]_  = A168 & A169;
  assign \new_[11460]_  = ~A166 & A167;
  assign \new_[11461]_  = \new_[11460]_  & \new_[11457]_ ;
  assign \new_[11464]_  = A233 & ~A232;
  assign \new_[11467]_  = A236 & A234;
  assign \new_[11468]_  = \new_[11467]_  & \new_[11464]_ ;
  assign \new_[11471]_  = A168 & A169;
  assign \new_[11474]_  = ~A166 & A167;
  assign \new_[11475]_  = \new_[11474]_  & \new_[11471]_ ;
  assign \new_[11478]_  = ~A233 & A232;
  assign \new_[11481]_  = A235 & A234;
  assign \new_[11482]_  = \new_[11481]_  & \new_[11478]_ ;
  assign \new_[11485]_  = A168 & A169;
  assign \new_[11488]_  = ~A166 & A167;
  assign \new_[11489]_  = \new_[11488]_  & \new_[11485]_ ;
  assign \new_[11492]_  = ~A233 & A232;
  assign \new_[11495]_  = A236 & A234;
  assign \new_[11496]_  = \new_[11495]_  & \new_[11492]_ ;
  assign \new_[11499]_  = A168 & A169;
  assign \new_[11502]_  = A166 & ~A167;
  assign \new_[11503]_  = \new_[11502]_  & \new_[11499]_ ;
  assign \new_[11506]_  = A233 & ~A232;
  assign \new_[11509]_  = A235 & A234;
  assign \new_[11510]_  = \new_[11509]_  & \new_[11506]_ ;
  assign \new_[11513]_  = A168 & A169;
  assign \new_[11516]_  = A166 & ~A167;
  assign \new_[11517]_  = \new_[11516]_  & \new_[11513]_ ;
  assign \new_[11520]_  = A233 & ~A232;
  assign \new_[11523]_  = A236 & A234;
  assign \new_[11524]_  = \new_[11523]_  & \new_[11520]_ ;
  assign \new_[11527]_  = A168 & A169;
  assign \new_[11530]_  = A166 & ~A167;
  assign \new_[11531]_  = \new_[11530]_  & \new_[11527]_ ;
  assign \new_[11534]_  = ~A233 & A232;
  assign \new_[11537]_  = A235 & A234;
  assign \new_[11538]_  = \new_[11537]_  & \new_[11534]_ ;
  assign \new_[11541]_  = A168 & A169;
  assign \new_[11544]_  = A166 & ~A167;
  assign \new_[11545]_  = \new_[11544]_  & \new_[11541]_ ;
  assign \new_[11548]_  = ~A233 & A232;
  assign \new_[11551]_  = A236 & A234;
  assign \new_[11552]_  = \new_[11551]_  & \new_[11548]_ ;
  assign \new_[11555]_  = A200 & ~A199;
  assign \new_[11558]_  = A202 & A201;
  assign \new_[11559]_  = \new_[11558]_  & \new_[11555]_ ;
  assign \new_[11562]_  = A233 & ~A232;
  assign \new_[11566]_  = ~A236 & ~A235;
  assign \new_[11567]_  = ~A234 & \new_[11566]_ ;
  assign \new_[11568]_  = \new_[11567]_  & \new_[11562]_ ;
  assign \new_[11571]_  = A200 & ~A199;
  assign \new_[11574]_  = A202 & A201;
  assign \new_[11575]_  = \new_[11574]_  & \new_[11571]_ ;
  assign \new_[11578]_  = ~A233 & A232;
  assign \new_[11582]_  = ~A236 & ~A235;
  assign \new_[11583]_  = ~A234 & \new_[11582]_ ;
  assign \new_[11584]_  = \new_[11583]_  & \new_[11578]_ ;
  assign \new_[11587]_  = A200 & ~A199;
  assign \new_[11590]_  = A203 & A201;
  assign \new_[11591]_  = \new_[11590]_  & \new_[11587]_ ;
  assign \new_[11594]_  = A233 & ~A232;
  assign \new_[11598]_  = ~A236 & ~A235;
  assign \new_[11599]_  = ~A234 & \new_[11598]_ ;
  assign \new_[11600]_  = \new_[11599]_  & \new_[11594]_ ;
  assign \new_[11603]_  = A200 & ~A199;
  assign \new_[11606]_  = A203 & A201;
  assign \new_[11607]_  = \new_[11606]_  & \new_[11603]_ ;
  assign \new_[11610]_  = ~A233 & A232;
  assign \new_[11614]_  = ~A236 & ~A235;
  assign \new_[11615]_  = ~A234 & \new_[11614]_ ;
  assign \new_[11616]_  = \new_[11615]_  & \new_[11610]_ ;
  assign \new_[11619]_  = A200 & ~A199;
  assign \new_[11622]_  = ~A202 & ~A201;
  assign \new_[11623]_  = \new_[11622]_  & \new_[11619]_ ;
  assign \new_[11626]_  = ~A232 & ~A203;
  assign \new_[11630]_  = A235 & A234;
  assign \new_[11631]_  = A233 & \new_[11630]_ ;
  assign \new_[11632]_  = \new_[11631]_  & \new_[11626]_ ;
  assign \new_[11635]_  = A200 & ~A199;
  assign \new_[11638]_  = ~A202 & ~A201;
  assign \new_[11639]_  = \new_[11638]_  & \new_[11635]_ ;
  assign \new_[11642]_  = ~A232 & ~A203;
  assign \new_[11646]_  = A236 & A234;
  assign \new_[11647]_  = A233 & \new_[11646]_ ;
  assign \new_[11648]_  = \new_[11647]_  & \new_[11642]_ ;
  assign \new_[11651]_  = A200 & ~A199;
  assign \new_[11654]_  = ~A202 & ~A201;
  assign \new_[11655]_  = \new_[11654]_  & \new_[11651]_ ;
  assign \new_[11658]_  = A232 & ~A203;
  assign \new_[11662]_  = A235 & A234;
  assign \new_[11663]_  = ~A233 & \new_[11662]_ ;
  assign \new_[11664]_  = \new_[11663]_  & \new_[11658]_ ;
  assign \new_[11667]_  = A200 & ~A199;
  assign \new_[11670]_  = ~A202 & ~A201;
  assign \new_[11671]_  = \new_[11670]_  & \new_[11667]_ ;
  assign \new_[11674]_  = A232 & ~A203;
  assign \new_[11678]_  = A236 & A234;
  assign \new_[11679]_  = ~A233 & \new_[11678]_ ;
  assign \new_[11680]_  = \new_[11679]_  & \new_[11674]_ ;
  assign \new_[11683]_  = ~A200 & A199;
  assign \new_[11686]_  = A202 & A201;
  assign \new_[11687]_  = \new_[11686]_  & \new_[11683]_ ;
  assign \new_[11690]_  = A233 & ~A232;
  assign \new_[11694]_  = ~A236 & ~A235;
  assign \new_[11695]_  = ~A234 & \new_[11694]_ ;
  assign \new_[11696]_  = \new_[11695]_  & \new_[11690]_ ;
  assign \new_[11699]_  = ~A200 & A199;
  assign \new_[11702]_  = A202 & A201;
  assign \new_[11703]_  = \new_[11702]_  & \new_[11699]_ ;
  assign \new_[11706]_  = ~A233 & A232;
  assign \new_[11710]_  = ~A236 & ~A235;
  assign \new_[11711]_  = ~A234 & \new_[11710]_ ;
  assign \new_[11712]_  = \new_[11711]_  & \new_[11706]_ ;
  assign \new_[11715]_  = ~A200 & A199;
  assign \new_[11718]_  = A203 & A201;
  assign \new_[11719]_  = \new_[11718]_  & \new_[11715]_ ;
  assign \new_[11722]_  = A233 & ~A232;
  assign \new_[11726]_  = ~A236 & ~A235;
  assign \new_[11727]_  = ~A234 & \new_[11726]_ ;
  assign \new_[11728]_  = \new_[11727]_  & \new_[11722]_ ;
  assign \new_[11731]_  = ~A200 & A199;
  assign \new_[11734]_  = A203 & A201;
  assign \new_[11735]_  = \new_[11734]_  & \new_[11731]_ ;
  assign \new_[11738]_  = ~A233 & A232;
  assign \new_[11742]_  = ~A236 & ~A235;
  assign \new_[11743]_  = ~A234 & \new_[11742]_ ;
  assign \new_[11744]_  = \new_[11743]_  & \new_[11738]_ ;
  assign \new_[11747]_  = ~A200 & A199;
  assign \new_[11750]_  = ~A202 & ~A201;
  assign \new_[11751]_  = \new_[11750]_  & \new_[11747]_ ;
  assign \new_[11754]_  = ~A232 & ~A203;
  assign \new_[11758]_  = A235 & A234;
  assign \new_[11759]_  = A233 & \new_[11758]_ ;
  assign \new_[11760]_  = \new_[11759]_  & \new_[11754]_ ;
  assign \new_[11763]_  = ~A200 & A199;
  assign \new_[11766]_  = ~A202 & ~A201;
  assign \new_[11767]_  = \new_[11766]_  & \new_[11763]_ ;
  assign \new_[11770]_  = ~A232 & ~A203;
  assign \new_[11774]_  = A236 & A234;
  assign \new_[11775]_  = A233 & \new_[11774]_ ;
  assign \new_[11776]_  = \new_[11775]_  & \new_[11770]_ ;
  assign \new_[11779]_  = ~A200 & A199;
  assign \new_[11782]_  = ~A202 & ~A201;
  assign \new_[11783]_  = \new_[11782]_  & \new_[11779]_ ;
  assign \new_[11786]_  = A232 & ~A203;
  assign \new_[11790]_  = A235 & A234;
  assign \new_[11791]_  = ~A233 & \new_[11790]_ ;
  assign \new_[11792]_  = \new_[11791]_  & \new_[11786]_ ;
  assign \new_[11795]_  = ~A200 & A199;
  assign \new_[11798]_  = ~A202 & ~A201;
  assign \new_[11799]_  = \new_[11798]_  & \new_[11795]_ ;
  assign \new_[11802]_  = A232 & ~A203;
  assign \new_[11806]_  = A236 & A234;
  assign \new_[11807]_  = ~A233 & \new_[11806]_ ;
  assign \new_[11808]_  = \new_[11807]_  & \new_[11802]_ ;
  assign \new_[11811]_  = A168 & ~A170;
  assign \new_[11814]_  = ~A166 & A167;
  assign \new_[11815]_  = \new_[11814]_  & \new_[11811]_ ;
  assign \new_[11818]_  = A233 & ~A232;
  assign \new_[11822]_  = ~A236 & ~A235;
  assign \new_[11823]_  = ~A234 & \new_[11822]_ ;
  assign \new_[11824]_  = \new_[11823]_  & \new_[11818]_ ;
  assign \new_[11827]_  = A168 & ~A170;
  assign \new_[11830]_  = ~A166 & A167;
  assign \new_[11831]_  = \new_[11830]_  & \new_[11827]_ ;
  assign \new_[11834]_  = ~A233 & A232;
  assign \new_[11838]_  = ~A236 & ~A235;
  assign \new_[11839]_  = ~A234 & \new_[11838]_ ;
  assign \new_[11840]_  = \new_[11839]_  & \new_[11834]_ ;
  assign \new_[11843]_  = A168 & ~A170;
  assign \new_[11846]_  = A166 & ~A167;
  assign \new_[11847]_  = \new_[11846]_  & \new_[11843]_ ;
  assign \new_[11850]_  = A233 & ~A232;
  assign \new_[11854]_  = ~A236 & ~A235;
  assign \new_[11855]_  = ~A234 & \new_[11854]_ ;
  assign \new_[11856]_  = \new_[11855]_  & \new_[11850]_ ;
  assign \new_[11859]_  = A168 & ~A170;
  assign \new_[11862]_  = A166 & ~A167;
  assign \new_[11863]_  = \new_[11862]_  & \new_[11859]_ ;
  assign \new_[11866]_  = ~A233 & A232;
  assign \new_[11870]_  = ~A236 & ~A235;
  assign \new_[11871]_  = ~A234 & \new_[11870]_ ;
  assign \new_[11872]_  = \new_[11871]_  & \new_[11866]_ ;
  assign \new_[11875]_  = A168 & A169;
  assign \new_[11878]_  = ~A166 & A167;
  assign \new_[11879]_  = \new_[11878]_  & \new_[11875]_ ;
  assign \new_[11882]_  = A233 & ~A232;
  assign \new_[11886]_  = ~A236 & ~A235;
  assign \new_[11887]_  = ~A234 & \new_[11886]_ ;
  assign \new_[11888]_  = \new_[11887]_  & \new_[11882]_ ;
  assign \new_[11891]_  = A168 & A169;
  assign \new_[11894]_  = ~A166 & A167;
  assign \new_[11895]_  = \new_[11894]_  & \new_[11891]_ ;
  assign \new_[11898]_  = ~A233 & A232;
  assign \new_[11902]_  = ~A236 & ~A235;
  assign \new_[11903]_  = ~A234 & \new_[11902]_ ;
  assign \new_[11904]_  = \new_[11903]_  & \new_[11898]_ ;
  assign \new_[11907]_  = A168 & A169;
  assign \new_[11910]_  = A166 & ~A167;
  assign \new_[11911]_  = \new_[11910]_  & \new_[11907]_ ;
  assign \new_[11914]_  = A233 & ~A232;
  assign \new_[11918]_  = ~A236 & ~A235;
  assign \new_[11919]_  = ~A234 & \new_[11918]_ ;
  assign \new_[11920]_  = \new_[11919]_  & \new_[11914]_ ;
  assign \new_[11923]_  = A168 & A169;
  assign \new_[11926]_  = A166 & ~A167;
  assign \new_[11927]_  = \new_[11926]_  & \new_[11923]_ ;
  assign \new_[11930]_  = ~A233 & A232;
  assign \new_[11934]_  = ~A236 & ~A235;
  assign \new_[11935]_  = ~A234 & \new_[11934]_ ;
  assign \new_[11936]_  = \new_[11935]_  & \new_[11930]_ ;
  assign \new_[11939]_  = ~A169 & A170;
  assign \new_[11942]_  = A167 & ~A168;
  assign \new_[11943]_  = \new_[11942]_  & \new_[11939]_ ;
  assign \new_[11946]_  = ~A232 & ~A166;
  assign \new_[11950]_  = A235 & A234;
  assign \new_[11951]_  = A233 & \new_[11950]_ ;
  assign \new_[11952]_  = \new_[11951]_  & \new_[11946]_ ;
  assign \new_[11955]_  = ~A169 & A170;
  assign \new_[11958]_  = A167 & ~A168;
  assign \new_[11959]_  = \new_[11958]_  & \new_[11955]_ ;
  assign \new_[11962]_  = ~A232 & ~A166;
  assign \new_[11966]_  = A236 & A234;
  assign \new_[11967]_  = A233 & \new_[11966]_ ;
  assign \new_[11968]_  = \new_[11967]_  & \new_[11962]_ ;
  assign \new_[11971]_  = ~A169 & A170;
  assign \new_[11974]_  = A167 & ~A168;
  assign \new_[11975]_  = \new_[11974]_  & \new_[11971]_ ;
  assign \new_[11978]_  = A232 & ~A166;
  assign \new_[11982]_  = A235 & A234;
  assign \new_[11983]_  = ~A233 & \new_[11982]_ ;
  assign \new_[11984]_  = \new_[11983]_  & \new_[11978]_ ;
  assign \new_[11987]_  = ~A169 & A170;
  assign \new_[11990]_  = A167 & ~A168;
  assign \new_[11991]_  = \new_[11990]_  & \new_[11987]_ ;
  assign \new_[11994]_  = A232 & ~A166;
  assign \new_[11998]_  = A236 & A234;
  assign \new_[11999]_  = ~A233 & \new_[11998]_ ;
  assign \new_[12000]_  = \new_[11999]_  & \new_[11994]_ ;
  assign \new_[12003]_  = ~A169 & A170;
  assign \new_[12006]_  = ~A167 & ~A168;
  assign \new_[12007]_  = \new_[12006]_  & \new_[12003]_ ;
  assign \new_[12010]_  = ~A232 & A166;
  assign \new_[12014]_  = A235 & A234;
  assign \new_[12015]_  = A233 & \new_[12014]_ ;
  assign \new_[12016]_  = \new_[12015]_  & \new_[12010]_ ;
  assign \new_[12019]_  = ~A169 & A170;
  assign \new_[12022]_  = ~A167 & ~A168;
  assign \new_[12023]_  = \new_[12022]_  & \new_[12019]_ ;
  assign \new_[12026]_  = ~A232 & A166;
  assign \new_[12030]_  = A236 & A234;
  assign \new_[12031]_  = A233 & \new_[12030]_ ;
  assign \new_[12032]_  = \new_[12031]_  & \new_[12026]_ ;
  assign \new_[12035]_  = ~A169 & A170;
  assign \new_[12038]_  = ~A167 & ~A168;
  assign \new_[12039]_  = \new_[12038]_  & \new_[12035]_ ;
  assign \new_[12042]_  = A232 & A166;
  assign \new_[12046]_  = A235 & A234;
  assign \new_[12047]_  = ~A233 & \new_[12046]_ ;
  assign \new_[12048]_  = \new_[12047]_  & \new_[12042]_ ;
  assign \new_[12051]_  = ~A169 & A170;
  assign \new_[12054]_  = ~A167 & ~A168;
  assign \new_[12055]_  = \new_[12054]_  & \new_[12051]_ ;
  assign \new_[12058]_  = A232 & A166;
  assign \new_[12062]_  = A236 & A234;
  assign \new_[12063]_  = ~A233 & \new_[12062]_ ;
  assign \new_[12064]_  = \new_[12063]_  & \new_[12058]_ ;
  assign \new_[12067]_  = A200 & ~A199;
  assign \new_[12071]_  = ~A203 & ~A202;
  assign \new_[12072]_  = ~A201 & \new_[12071]_ ;
  assign \new_[12073]_  = \new_[12072]_  & \new_[12067]_ ;
  assign \new_[12076]_  = A233 & ~A232;
  assign \new_[12080]_  = ~A236 & ~A235;
  assign \new_[12081]_  = ~A234 & \new_[12080]_ ;
  assign \new_[12082]_  = \new_[12081]_  & \new_[12076]_ ;
  assign \new_[12085]_  = A200 & ~A199;
  assign \new_[12089]_  = ~A203 & ~A202;
  assign \new_[12090]_  = ~A201 & \new_[12089]_ ;
  assign \new_[12091]_  = \new_[12090]_  & \new_[12085]_ ;
  assign \new_[12094]_  = ~A233 & A232;
  assign \new_[12098]_  = ~A236 & ~A235;
  assign \new_[12099]_  = ~A234 & \new_[12098]_ ;
  assign \new_[12100]_  = \new_[12099]_  & \new_[12094]_ ;
  assign \new_[12103]_  = ~A200 & A199;
  assign \new_[12107]_  = ~A203 & ~A202;
  assign \new_[12108]_  = ~A201 & \new_[12107]_ ;
  assign \new_[12109]_  = \new_[12108]_  & \new_[12103]_ ;
  assign \new_[12112]_  = A233 & ~A232;
  assign \new_[12116]_  = ~A236 & ~A235;
  assign \new_[12117]_  = ~A234 & \new_[12116]_ ;
  assign \new_[12118]_  = \new_[12117]_  & \new_[12112]_ ;
  assign \new_[12121]_  = ~A200 & A199;
  assign \new_[12125]_  = ~A203 & ~A202;
  assign \new_[12126]_  = ~A201 & \new_[12125]_ ;
  assign \new_[12127]_  = \new_[12126]_  & \new_[12121]_ ;
  assign \new_[12130]_  = ~A233 & A232;
  assign \new_[12134]_  = ~A236 & ~A235;
  assign \new_[12135]_  = ~A234 & \new_[12134]_ ;
  assign \new_[12136]_  = \new_[12135]_  & \new_[12130]_ ;
  assign \new_[12139]_  = A166 & A167;
  assign \new_[12143]_  = ~A265 & A202;
  assign \new_[12144]_  = ~A201 & \new_[12143]_ ;
  assign \new_[12145]_  = \new_[12144]_  & \new_[12139]_ ;
  assign \new_[12148]_  = A267 & A266;
  assign \new_[12152]_  = A301 & ~A300;
  assign \new_[12153]_  = A268 & \new_[12152]_ ;
  assign \new_[12154]_  = \new_[12153]_  & \new_[12148]_ ;
  assign \new_[12157]_  = A166 & A167;
  assign \new_[12161]_  = ~A265 & A202;
  assign \new_[12162]_  = ~A201 & \new_[12161]_ ;
  assign \new_[12163]_  = \new_[12162]_  & \new_[12157]_ ;
  assign \new_[12166]_  = A267 & A266;
  assign \new_[12170]_  = A302 & ~A300;
  assign \new_[12171]_  = A268 & \new_[12170]_ ;
  assign \new_[12172]_  = \new_[12171]_  & \new_[12166]_ ;
  assign \new_[12175]_  = A166 & A167;
  assign \new_[12179]_  = ~A265 & A202;
  assign \new_[12180]_  = ~A201 & \new_[12179]_ ;
  assign \new_[12181]_  = \new_[12180]_  & \new_[12175]_ ;
  assign \new_[12184]_  = A267 & A266;
  assign \new_[12188]_  = A299 & A298;
  assign \new_[12189]_  = A268 & \new_[12188]_ ;
  assign \new_[12190]_  = \new_[12189]_  & \new_[12184]_ ;
  assign \new_[12193]_  = A166 & A167;
  assign \new_[12197]_  = ~A265 & A202;
  assign \new_[12198]_  = ~A201 & \new_[12197]_ ;
  assign \new_[12199]_  = \new_[12198]_  & \new_[12193]_ ;
  assign \new_[12202]_  = A267 & A266;
  assign \new_[12206]_  = ~A299 & ~A298;
  assign \new_[12207]_  = A268 & \new_[12206]_ ;
  assign \new_[12208]_  = \new_[12207]_  & \new_[12202]_ ;
  assign \new_[12211]_  = A166 & A167;
  assign \new_[12215]_  = ~A265 & A202;
  assign \new_[12216]_  = ~A201 & \new_[12215]_ ;
  assign \new_[12217]_  = \new_[12216]_  & \new_[12211]_ ;
  assign \new_[12220]_  = A267 & A266;
  assign \new_[12224]_  = A301 & ~A300;
  assign \new_[12225]_  = A269 & \new_[12224]_ ;
  assign \new_[12226]_  = \new_[12225]_  & \new_[12220]_ ;
  assign \new_[12229]_  = A166 & A167;
  assign \new_[12233]_  = ~A265 & A202;
  assign \new_[12234]_  = ~A201 & \new_[12233]_ ;
  assign \new_[12235]_  = \new_[12234]_  & \new_[12229]_ ;
  assign \new_[12238]_  = A267 & A266;
  assign \new_[12242]_  = A302 & ~A300;
  assign \new_[12243]_  = A269 & \new_[12242]_ ;
  assign \new_[12244]_  = \new_[12243]_  & \new_[12238]_ ;
  assign \new_[12247]_  = A166 & A167;
  assign \new_[12251]_  = ~A265 & A202;
  assign \new_[12252]_  = ~A201 & \new_[12251]_ ;
  assign \new_[12253]_  = \new_[12252]_  & \new_[12247]_ ;
  assign \new_[12256]_  = A267 & A266;
  assign \new_[12260]_  = A299 & A298;
  assign \new_[12261]_  = A269 & \new_[12260]_ ;
  assign \new_[12262]_  = \new_[12261]_  & \new_[12256]_ ;
  assign \new_[12265]_  = A166 & A167;
  assign \new_[12269]_  = ~A265 & A202;
  assign \new_[12270]_  = ~A201 & \new_[12269]_ ;
  assign \new_[12271]_  = \new_[12270]_  & \new_[12265]_ ;
  assign \new_[12274]_  = A267 & A266;
  assign \new_[12278]_  = ~A299 & ~A298;
  assign \new_[12279]_  = A269 & \new_[12278]_ ;
  assign \new_[12280]_  = \new_[12279]_  & \new_[12274]_ ;
  assign \new_[12283]_  = A166 & A167;
  assign \new_[12287]_  = A265 & A202;
  assign \new_[12288]_  = ~A201 & \new_[12287]_ ;
  assign \new_[12289]_  = \new_[12288]_  & \new_[12283]_ ;
  assign \new_[12292]_  = A267 & ~A266;
  assign \new_[12296]_  = A301 & ~A300;
  assign \new_[12297]_  = A268 & \new_[12296]_ ;
  assign \new_[12298]_  = \new_[12297]_  & \new_[12292]_ ;
  assign \new_[12301]_  = A166 & A167;
  assign \new_[12305]_  = A265 & A202;
  assign \new_[12306]_  = ~A201 & \new_[12305]_ ;
  assign \new_[12307]_  = \new_[12306]_  & \new_[12301]_ ;
  assign \new_[12310]_  = A267 & ~A266;
  assign \new_[12314]_  = A302 & ~A300;
  assign \new_[12315]_  = A268 & \new_[12314]_ ;
  assign \new_[12316]_  = \new_[12315]_  & \new_[12310]_ ;
  assign \new_[12319]_  = A166 & A167;
  assign \new_[12323]_  = A265 & A202;
  assign \new_[12324]_  = ~A201 & \new_[12323]_ ;
  assign \new_[12325]_  = \new_[12324]_  & \new_[12319]_ ;
  assign \new_[12328]_  = A267 & ~A266;
  assign \new_[12332]_  = A299 & A298;
  assign \new_[12333]_  = A268 & \new_[12332]_ ;
  assign \new_[12334]_  = \new_[12333]_  & \new_[12328]_ ;
  assign \new_[12337]_  = A166 & A167;
  assign \new_[12341]_  = A265 & A202;
  assign \new_[12342]_  = ~A201 & \new_[12341]_ ;
  assign \new_[12343]_  = \new_[12342]_  & \new_[12337]_ ;
  assign \new_[12346]_  = A267 & ~A266;
  assign \new_[12350]_  = ~A299 & ~A298;
  assign \new_[12351]_  = A268 & \new_[12350]_ ;
  assign \new_[12352]_  = \new_[12351]_  & \new_[12346]_ ;
  assign \new_[12355]_  = A166 & A167;
  assign \new_[12359]_  = A265 & A202;
  assign \new_[12360]_  = ~A201 & \new_[12359]_ ;
  assign \new_[12361]_  = \new_[12360]_  & \new_[12355]_ ;
  assign \new_[12364]_  = A267 & ~A266;
  assign \new_[12368]_  = A301 & ~A300;
  assign \new_[12369]_  = A269 & \new_[12368]_ ;
  assign \new_[12370]_  = \new_[12369]_  & \new_[12364]_ ;
  assign \new_[12373]_  = A166 & A167;
  assign \new_[12377]_  = A265 & A202;
  assign \new_[12378]_  = ~A201 & \new_[12377]_ ;
  assign \new_[12379]_  = \new_[12378]_  & \new_[12373]_ ;
  assign \new_[12382]_  = A267 & ~A266;
  assign \new_[12386]_  = A302 & ~A300;
  assign \new_[12387]_  = A269 & \new_[12386]_ ;
  assign \new_[12388]_  = \new_[12387]_  & \new_[12382]_ ;
  assign \new_[12391]_  = A166 & A167;
  assign \new_[12395]_  = A265 & A202;
  assign \new_[12396]_  = ~A201 & \new_[12395]_ ;
  assign \new_[12397]_  = \new_[12396]_  & \new_[12391]_ ;
  assign \new_[12400]_  = A267 & ~A266;
  assign \new_[12404]_  = A299 & A298;
  assign \new_[12405]_  = A269 & \new_[12404]_ ;
  assign \new_[12406]_  = \new_[12405]_  & \new_[12400]_ ;
  assign \new_[12409]_  = A166 & A167;
  assign \new_[12413]_  = A265 & A202;
  assign \new_[12414]_  = ~A201 & \new_[12413]_ ;
  assign \new_[12415]_  = \new_[12414]_  & \new_[12409]_ ;
  assign \new_[12418]_  = A267 & ~A266;
  assign \new_[12422]_  = ~A299 & ~A298;
  assign \new_[12423]_  = A269 & \new_[12422]_ ;
  assign \new_[12424]_  = \new_[12423]_  & \new_[12418]_ ;
  assign \new_[12427]_  = A166 & A167;
  assign \new_[12431]_  = ~A265 & A203;
  assign \new_[12432]_  = ~A201 & \new_[12431]_ ;
  assign \new_[12433]_  = \new_[12432]_  & \new_[12427]_ ;
  assign \new_[12436]_  = A267 & A266;
  assign \new_[12440]_  = A301 & ~A300;
  assign \new_[12441]_  = A268 & \new_[12440]_ ;
  assign \new_[12442]_  = \new_[12441]_  & \new_[12436]_ ;
  assign \new_[12445]_  = A166 & A167;
  assign \new_[12449]_  = ~A265 & A203;
  assign \new_[12450]_  = ~A201 & \new_[12449]_ ;
  assign \new_[12451]_  = \new_[12450]_  & \new_[12445]_ ;
  assign \new_[12454]_  = A267 & A266;
  assign \new_[12458]_  = A302 & ~A300;
  assign \new_[12459]_  = A268 & \new_[12458]_ ;
  assign \new_[12460]_  = \new_[12459]_  & \new_[12454]_ ;
  assign \new_[12463]_  = A166 & A167;
  assign \new_[12467]_  = ~A265 & A203;
  assign \new_[12468]_  = ~A201 & \new_[12467]_ ;
  assign \new_[12469]_  = \new_[12468]_  & \new_[12463]_ ;
  assign \new_[12472]_  = A267 & A266;
  assign \new_[12476]_  = A299 & A298;
  assign \new_[12477]_  = A268 & \new_[12476]_ ;
  assign \new_[12478]_  = \new_[12477]_  & \new_[12472]_ ;
  assign \new_[12481]_  = A166 & A167;
  assign \new_[12485]_  = ~A265 & A203;
  assign \new_[12486]_  = ~A201 & \new_[12485]_ ;
  assign \new_[12487]_  = \new_[12486]_  & \new_[12481]_ ;
  assign \new_[12490]_  = A267 & A266;
  assign \new_[12494]_  = ~A299 & ~A298;
  assign \new_[12495]_  = A268 & \new_[12494]_ ;
  assign \new_[12496]_  = \new_[12495]_  & \new_[12490]_ ;
  assign \new_[12499]_  = A166 & A167;
  assign \new_[12503]_  = ~A265 & A203;
  assign \new_[12504]_  = ~A201 & \new_[12503]_ ;
  assign \new_[12505]_  = \new_[12504]_  & \new_[12499]_ ;
  assign \new_[12508]_  = A267 & A266;
  assign \new_[12512]_  = A301 & ~A300;
  assign \new_[12513]_  = A269 & \new_[12512]_ ;
  assign \new_[12514]_  = \new_[12513]_  & \new_[12508]_ ;
  assign \new_[12517]_  = A166 & A167;
  assign \new_[12521]_  = ~A265 & A203;
  assign \new_[12522]_  = ~A201 & \new_[12521]_ ;
  assign \new_[12523]_  = \new_[12522]_  & \new_[12517]_ ;
  assign \new_[12526]_  = A267 & A266;
  assign \new_[12530]_  = A302 & ~A300;
  assign \new_[12531]_  = A269 & \new_[12530]_ ;
  assign \new_[12532]_  = \new_[12531]_  & \new_[12526]_ ;
  assign \new_[12535]_  = A166 & A167;
  assign \new_[12539]_  = ~A265 & A203;
  assign \new_[12540]_  = ~A201 & \new_[12539]_ ;
  assign \new_[12541]_  = \new_[12540]_  & \new_[12535]_ ;
  assign \new_[12544]_  = A267 & A266;
  assign \new_[12548]_  = A299 & A298;
  assign \new_[12549]_  = A269 & \new_[12548]_ ;
  assign \new_[12550]_  = \new_[12549]_  & \new_[12544]_ ;
  assign \new_[12553]_  = A166 & A167;
  assign \new_[12557]_  = ~A265 & A203;
  assign \new_[12558]_  = ~A201 & \new_[12557]_ ;
  assign \new_[12559]_  = \new_[12558]_  & \new_[12553]_ ;
  assign \new_[12562]_  = A267 & A266;
  assign \new_[12566]_  = ~A299 & ~A298;
  assign \new_[12567]_  = A269 & \new_[12566]_ ;
  assign \new_[12568]_  = \new_[12567]_  & \new_[12562]_ ;
  assign \new_[12571]_  = A166 & A167;
  assign \new_[12575]_  = A265 & A203;
  assign \new_[12576]_  = ~A201 & \new_[12575]_ ;
  assign \new_[12577]_  = \new_[12576]_  & \new_[12571]_ ;
  assign \new_[12580]_  = A267 & ~A266;
  assign \new_[12584]_  = A301 & ~A300;
  assign \new_[12585]_  = A268 & \new_[12584]_ ;
  assign \new_[12586]_  = \new_[12585]_  & \new_[12580]_ ;
  assign \new_[12589]_  = A166 & A167;
  assign \new_[12593]_  = A265 & A203;
  assign \new_[12594]_  = ~A201 & \new_[12593]_ ;
  assign \new_[12595]_  = \new_[12594]_  & \new_[12589]_ ;
  assign \new_[12598]_  = A267 & ~A266;
  assign \new_[12602]_  = A302 & ~A300;
  assign \new_[12603]_  = A268 & \new_[12602]_ ;
  assign \new_[12604]_  = \new_[12603]_  & \new_[12598]_ ;
  assign \new_[12607]_  = A166 & A167;
  assign \new_[12611]_  = A265 & A203;
  assign \new_[12612]_  = ~A201 & \new_[12611]_ ;
  assign \new_[12613]_  = \new_[12612]_  & \new_[12607]_ ;
  assign \new_[12616]_  = A267 & ~A266;
  assign \new_[12620]_  = A299 & A298;
  assign \new_[12621]_  = A268 & \new_[12620]_ ;
  assign \new_[12622]_  = \new_[12621]_  & \new_[12616]_ ;
  assign \new_[12625]_  = A166 & A167;
  assign \new_[12629]_  = A265 & A203;
  assign \new_[12630]_  = ~A201 & \new_[12629]_ ;
  assign \new_[12631]_  = \new_[12630]_  & \new_[12625]_ ;
  assign \new_[12634]_  = A267 & ~A266;
  assign \new_[12638]_  = ~A299 & ~A298;
  assign \new_[12639]_  = A268 & \new_[12638]_ ;
  assign \new_[12640]_  = \new_[12639]_  & \new_[12634]_ ;
  assign \new_[12643]_  = A166 & A167;
  assign \new_[12647]_  = A265 & A203;
  assign \new_[12648]_  = ~A201 & \new_[12647]_ ;
  assign \new_[12649]_  = \new_[12648]_  & \new_[12643]_ ;
  assign \new_[12652]_  = A267 & ~A266;
  assign \new_[12656]_  = A301 & ~A300;
  assign \new_[12657]_  = A269 & \new_[12656]_ ;
  assign \new_[12658]_  = \new_[12657]_  & \new_[12652]_ ;
  assign \new_[12661]_  = A166 & A167;
  assign \new_[12665]_  = A265 & A203;
  assign \new_[12666]_  = ~A201 & \new_[12665]_ ;
  assign \new_[12667]_  = \new_[12666]_  & \new_[12661]_ ;
  assign \new_[12670]_  = A267 & ~A266;
  assign \new_[12674]_  = A302 & ~A300;
  assign \new_[12675]_  = A269 & \new_[12674]_ ;
  assign \new_[12676]_  = \new_[12675]_  & \new_[12670]_ ;
  assign \new_[12679]_  = A166 & A167;
  assign \new_[12683]_  = A265 & A203;
  assign \new_[12684]_  = ~A201 & \new_[12683]_ ;
  assign \new_[12685]_  = \new_[12684]_  & \new_[12679]_ ;
  assign \new_[12688]_  = A267 & ~A266;
  assign \new_[12692]_  = A299 & A298;
  assign \new_[12693]_  = A269 & \new_[12692]_ ;
  assign \new_[12694]_  = \new_[12693]_  & \new_[12688]_ ;
  assign \new_[12697]_  = A166 & A167;
  assign \new_[12701]_  = A265 & A203;
  assign \new_[12702]_  = ~A201 & \new_[12701]_ ;
  assign \new_[12703]_  = \new_[12702]_  & \new_[12697]_ ;
  assign \new_[12706]_  = A267 & ~A266;
  assign \new_[12710]_  = ~A299 & ~A298;
  assign \new_[12711]_  = A269 & \new_[12710]_ ;
  assign \new_[12712]_  = \new_[12711]_  & \new_[12706]_ ;
  assign \new_[12715]_  = A166 & A167;
  assign \new_[12719]_  = ~A265 & A200;
  assign \new_[12720]_  = A199 & \new_[12719]_ ;
  assign \new_[12721]_  = \new_[12720]_  & \new_[12715]_ ;
  assign \new_[12724]_  = A267 & A266;
  assign \new_[12728]_  = A301 & ~A300;
  assign \new_[12729]_  = A268 & \new_[12728]_ ;
  assign \new_[12730]_  = \new_[12729]_  & \new_[12724]_ ;
  assign \new_[12733]_  = A166 & A167;
  assign \new_[12737]_  = ~A265 & A200;
  assign \new_[12738]_  = A199 & \new_[12737]_ ;
  assign \new_[12739]_  = \new_[12738]_  & \new_[12733]_ ;
  assign \new_[12742]_  = A267 & A266;
  assign \new_[12746]_  = A302 & ~A300;
  assign \new_[12747]_  = A268 & \new_[12746]_ ;
  assign \new_[12748]_  = \new_[12747]_  & \new_[12742]_ ;
  assign \new_[12751]_  = A166 & A167;
  assign \new_[12755]_  = ~A265 & A200;
  assign \new_[12756]_  = A199 & \new_[12755]_ ;
  assign \new_[12757]_  = \new_[12756]_  & \new_[12751]_ ;
  assign \new_[12760]_  = A267 & A266;
  assign \new_[12764]_  = A299 & A298;
  assign \new_[12765]_  = A268 & \new_[12764]_ ;
  assign \new_[12766]_  = \new_[12765]_  & \new_[12760]_ ;
  assign \new_[12769]_  = A166 & A167;
  assign \new_[12773]_  = ~A265 & A200;
  assign \new_[12774]_  = A199 & \new_[12773]_ ;
  assign \new_[12775]_  = \new_[12774]_  & \new_[12769]_ ;
  assign \new_[12778]_  = A267 & A266;
  assign \new_[12782]_  = ~A299 & ~A298;
  assign \new_[12783]_  = A268 & \new_[12782]_ ;
  assign \new_[12784]_  = \new_[12783]_  & \new_[12778]_ ;
  assign \new_[12787]_  = A166 & A167;
  assign \new_[12791]_  = ~A265 & A200;
  assign \new_[12792]_  = A199 & \new_[12791]_ ;
  assign \new_[12793]_  = \new_[12792]_  & \new_[12787]_ ;
  assign \new_[12796]_  = A267 & A266;
  assign \new_[12800]_  = A301 & ~A300;
  assign \new_[12801]_  = A269 & \new_[12800]_ ;
  assign \new_[12802]_  = \new_[12801]_  & \new_[12796]_ ;
  assign \new_[12805]_  = A166 & A167;
  assign \new_[12809]_  = ~A265 & A200;
  assign \new_[12810]_  = A199 & \new_[12809]_ ;
  assign \new_[12811]_  = \new_[12810]_  & \new_[12805]_ ;
  assign \new_[12814]_  = A267 & A266;
  assign \new_[12818]_  = A302 & ~A300;
  assign \new_[12819]_  = A269 & \new_[12818]_ ;
  assign \new_[12820]_  = \new_[12819]_  & \new_[12814]_ ;
  assign \new_[12823]_  = A166 & A167;
  assign \new_[12827]_  = ~A265 & A200;
  assign \new_[12828]_  = A199 & \new_[12827]_ ;
  assign \new_[12829]_  = \new_[12828]_  & \new_[12823]_ ;
  assign \new_[12832]_  = A267 & A266;
  assign \new_[12836]_  = A299 & A298;
  assign \new_[12837]_  = A269 & \new_[12836]_ ;
  assign \new_[12838]_  = \new_[12837]_  & \new_[12832]_ ;
  assign \new_[12841]_  = A166 & A167;
  assign \new_[12845]_  = ~A265 & A200;
  assign \new_[12846]_  = A199 & \new_[12845]_ ;
  assign \new_[12847]_  = \new_[12846]_  & \new_[12841]_ ;
  assign \new_[12850]_  = A267 & A266;
  assign \new_[12854]_  = ~A299 & ~A298;
  assign \new_[12855]_  = A269 & \new_[12854]_ ;
  assign \new_[12856]_  = \new_[12855]_  & \new_[12850]_ ;
  assign \new_[12859]_  = A166 & A167;
  assign \new_[12863]_  = A265 & A200;
  assign \new_[12864]_  = A199 & \new_[12863]_ ;
  assign \new_[12865]_  = \new_[12864]_  & \new_[12859]_ ;
  assign \new_[12868]_  = A267 & ~A266;
  assign \new_[12872]_  = A301 & ~A300;
  assign \new_[12873]_  = A268 & \new_[12872]_ ;
  assign \new_[12874]_  = \new_[12873]_  & \new_[12868]_ ;
  assign \new_[12877]_  = A166 & A167;
  assign \new_[12881]_  = A265 & A200;
  assign \new_[12882]_  = A199 & \new_[12881]_ ;
  assign \new_[12883]_  = \new_[12882]_  & \new_[12877]_ ;
  assign \new_[12886]_  = A267 & ~A266;
  assign \new_[12890]_  = A302 & ~A300;
  assign \new_[12891]_  = A268 & \new_[12890]_ ;
  assign \new_[12892]_  = \new_[12891]_  & \new_[12886]_ ;
  assign \new_[12895]_  = A166 & A167;
  assign \new_[12899]_  = A265 & A200;
  assign \new_[12900]_  = A199 & \new_[12899]_ ;
  assign \new_[12901]_  = \new_[12900]_  & \new_[12895]_ ;
  assign \new_[12904]_  = A267 & ~A266;
  assign \new_[12908]_  = A299 & A298;
  assign \new_[12909]_  = A268 & \new_[12908]_ ;
  assign \new_[12910]_  = \new_[12909]_  & \new_[12904]_ ;
  assign \new_[12913]_  = A166 & A167;
  assign \new_[12917]_  = A265 & A200;
  assign \new_[12918]_  = A199 & \new_[12917]_ ;
  assign \new_[12919]_  = \new_[12918]_  & \new_[12913]_ ;
  assign \new_[12922]_  = A267 & ~A266;
  assign \new_[12926]_  = ~A299 & ~A298;
  assign \new_[12927]_  = A268 & \new_[12926]_ ;
  assign \new_[12928]_  = \new_[12927]_  & \new_[12922]_ ;
  assign \new_[12931]_  = A166 & A167;
  assign \new_[12935]_  = A265 & A200;
  assign \new_[12936]_  = A199 & \new_[12935]_ ;
  assign \new_[12937]_  = \new_[12936]_  & \new_[12931]_ ;
  assign \new_[12940]_  = A267 & ~A266;
  assign \new_[12944]_  = A301 & ~A300;
  assign \new_[12945]_  = A269 & \new_[12944]_ ;
  assign \new_[12946]_  = \new_[12945]_  & \new_[12940]_ ;
  assign \new_[12949]_  = A166 & A167;
  assign \new_[12953]_  = A265 & A200;
  assign \new_[12954]_  = A199 & \new_[12953]_ ;
  assign \new_[12955]_  = \new_[12954]_  & \new_[12949]_ ;
  assign \new_[12958]_  = A267 & ~A266;
  assign \new_[12962]_  = A302 & ~A300;
  assign \new_[12963]_  = A269 & \new_[12962]_ ;
  assign \new_[12964]_  = \new_[12963]_  & \new_[12958]_ ;
  assign \new_[12967]_  = A166 & A167;
  assign \new_[12971]_  = A265 & A200;
  assign \new_[12972]_  = A199 & \new_[12971]_ ;
  assign \new_[12973]_  = \new_[12972]_  & \new_[12967]_ ;
  assign \new_[12976]_  = A267 & ~A266;
  assign \new_[12980]_  = A299 & A298;
  assign \new_[12981]_  = A269 & \new_[12980]_ ;
  assign \new_[12982]_  = \new_[12981]_  & \new_[12976]_ ;
  assign \new_[12985]_  = A166 & A167;
  assign \new_[12989]_  = A265 & A200;
  assign \new_[12990]_  = A199 & \new_[12989]_ ;
  assign \new_[12991]_  = \new_[12990]_  & \new_[12985]_ ;
  assign \new_[12994]_  = A267 & ~A266;
  assign \new_[12998]_  = ~A299 & ~A298;
  assign \new_[12999]_  = A269 & \new_[12998]_ ;
  assign \new_[13000]_  = \new_[12999]_  & \new_[12994]_ ;
  assign \new_[13003]_  = A166 & A167;
  assign \new_[13007]_  = ~A265 & ~A200;
  assign \new_[13008]_  = ~A199 & \new_[13007]_ ;
  assign \new_[13009]_  = \new_[13008]_  & \new_[13003]_ ;
  assign \new_[13012]_  = A267 & A266;
  assign \new_[13016]_  = A301 & ~A300;
  assign \new_[13017]_  = A268 & \new_[13016]_ ;
  assign \new_[13018]_  = \new_[13017]_  & \new_[13012]_ ;
  assign \new_[13021]_  = A166 & A167;
  assign \new_[13025]_  = ~A265 & ~A200;
  assign \new_[13026]_  = ~A199 & \new_[13025]_ ;
  assign \new_[13027]_  = \new_[13026]_  & \new_[13021]_ ;
  assign \new_[13030]_  = A267 & A266;
  assign \new_[13034]_  = A302 & ~A300;
  assign \new_[13035]_  = A268 & \new_[13034]_ ;
  assign \new_[13036]_  = \new_[13035]_  & \new_[13030]_ ;
  assign \new_[13039]_  = A166 & A167;
  assign \new_[13043]_  = ~A265 & ~A200;
  assign \new_[13044]_  = ~A199 & \new_[13043]_ ;
  assign \new_[13045]_  = \new_[13044]_  & \new_[13039]_ ;
  assign \new_[13048]_  = A267 & A266;
  assign \new_[13052]_  = A299 & A298;
  assign \new_[13053]_  = A268 & \new_[13052]_ ;
  assign \new_[13054]_  = \new_[13053]_  & \new_[13048]_ ;
  assign \new_[13057]_  = A166 & A167;
  assign \new_[13061]_  = ~A265 & ~A200;
  assign \new_[13062]_  = ~A199 & \new_[13061]_ ;
  assign \new_[13063]_  = \new_[13062]_  & \new_[13057]_ ;
  assign \new_[13066]_  = A267 & A266;
  assign \new_[13070]_  = ~A299 & ~A298;
  assign \new_[13071]_  = A268 & \new_[13070]_ ;
  assign \new_[13072]_  = \new_[13071]_  & \new_[13066]_ ;
  assign \new_[13075]_  = A166 & A167;
  assign \new_[13079]_  = ~A265 & ~A200;
  assign \new_[13080]_  = ~A199 & \new_[13079]_ ;
  assign \new_[13081]_  = \new_[13080]_  & \new_[13075]_ ;
  assign \new_[13084]_  = A267 & A266;
  assign \new_[13088]_  = A301 & ~A300;
  assign \new_[13089]_  = A269 & \new_[13088]_ ;
  assign \new_[13090]_  = \new_[13089]_  & \new_[13084]_ ;
  assign \new_[13093]_  = A166 & A167;
  assign \new_[13097]_  = ~A265 & ~A200;
  assign \new_[13098]_  = ~A199 & \new_[13097]_ ;
  assign \new_[13099]_  = \new_[13098]_  & \new_[13093]_ ;
  assign \new_[13102]_  = A267 & A266;
  assign \new_[13106]_  = A302 & ~A300;
  assign \new_[13107]_  = A269 & \new_[13106]_ ;
  assign \new_[13108]_  = \new_[13107]_  & \new_[13102]_ ;
  assign \new_[13111]_  = A166 & A167;
  assign \new_[13115]_  = ~A265 & ~A200;
  assign \new_[13116]_  = ~A199 & \new_[13115]_ ;
  assign \new_[13117]_  = \new_[13116]_  & \new_[13111]_ ;
  assign \new_[13120]_  = A267 & A266;
  assign \new_[13124]_  = A299 & A298;
  assign \new_[13125]_  = A269 & \new_[13124]_ ;
  assign \new_[13126]_  = \new_[13125]_  & \new_[13120]_ ;
  assign \new_[13129]_  = A166 & A167;
  assign \new_[13133]_  = ~A265 & ~A200;
  assign \new_[13134]_  = ~A199 & \new_[13133]_ ;
  assign \new_[13135]_  = \new_[13134]_  & \new_[13129]_ ;
  assign \new_[13138]_  = A267 & A266;
  assign \new_[13142]_  = ~A299 & ~A298;
  assign \new_[13143]_  = A269 & \new_[13142]_ ;
  assign \new_[13144]_  = \new_[13143]_  & \new_[13138]_ ;
  assign \new_[13147]_  = A166 & A167;
  assign \new_[13151]_  = A265 & ~A200;
  assign \new_[13152]_  = ~A199 & \new_[13151]_ ;
  assign \new_[13153]_  = \new_[13152]_  & \new_[13147]_ ;
  assign \new_[13156]_  = A267 & ~A266;
  assign \new_[13160]_  = A301 & ~A300;
  assign \new_[13161]_  = A268 & \new_[13160]_ ;
  assign \new_[13162]_  = \new_[13161]_  & \new_[13156]_ ;
  assign \new_[13165]_  = A166 & A167;
  assign \new_[13169]_  = A265 & ~A200;
  assign \new_[13170]_  = ~A199 & \new_[13169]_ ;
  assign \new_[13171]_  = \new_[13170]_  & \new_[13165]_ ;
  assign \new_[13174]_  = A267 & ~A266;
  assign \new_[13178]_  = A302 & ~A300;
  assign \new_[13179]_  = A268 & \new_[13178]_ ;
  assign \new_[13180]_  = \new_[13179]_  & \new_[13174]_ ;
  assign \new_[13183]_  = A166 & A167;
  assign \new_[13187]_  = A265 & ~A200;
  assign \new_[13188]_  = ~A199 & \new_[13187]_ ;
  assign \new_[13189]_  = \new_[13188]_  & \new_[13183]_ ;
  assign \new_[13192]_  = A267 & ~A266;
  assign \new_[13196]_  = A299 & A298;
  assign \new_[13197]_  = A268 & \new_[13196]_ ;
  assign \new_[13198]_  = \new_[13197]_  & \new_[13192]_ ;
  assign \new_[13201]_  = A166 & A167;
  assign \new_[13205]_  = A265 & ~A200;
  assign \new_[13206]_  = ~A199 & \new_[13205]_ ;
  assign \new_[13207]_  = \new_[13206]_  & \new_[13201]_ ;
  assign \new_[13210]_  = A267 & ~A266;
  assign \new_[13214]_  = ~A299 & ~A298;
  assign \new_[13215]_  = A268 & \new_[13214]_ ;
  assign \new_[13216]_  = \new_[13215]_  & \new_[13210]_ ;
  assign \new_[13219]_  = A166 & A167;
  assign \new_[13223]_  = A265 & ~A200;
  assign \new_[13224]_  = ~A199 & \new_[13223]_ ;
  assign \new_[13225]_  = \new_[13224]_  & \new_[13219]_ ;
  assign \new_[13228]_  = A267 & ~A266;
  assign \new_[13232]_  = A301 & ~A300;
  assign \new_[13233]_  = A269 & \new_[13232]_ ;
  assign \new_[13234]_  = \new_[13233]_  & \new_[13228]_ ;
  assign \new_[13237]_  = A166 & A167;
  assign \new_[13241]_  = A265 & ~A200;
  assign \new_[13242]_  = ~A199 & \new_[13241]_ ;
  assign \new_[13243]_  = \new_[13242]_  & \new_[13237]_ ;
  assign \new_[13246]_  = A267 & ~A266;
  assign \new_[13250]_  = A302 & ~A300;
  assign \new_[13251]_  = A269 & \new_[13250]_ ;
  assign \new_[13252]_  = \new_[13251]_  & \new_[13246]_ ;
  assign \new_[13255]_  = A166 & A167;
  assign \new_[13259]_  = A265 & ~A200;
  assign \new_[13260]_  = ~A199 & \new_[13259]_ ;
  assign \new_[13261]_  = \new_[13260]_  & \new_[13255]_ ;
  assign \new_[13264]_  = A267 & ~A266;
  assign \new_[13268]_  = A299 & A298;
  assign \new_[13269]_  = A269 & \new_[13268]_ ;
  assign \new_[13270]_  = \new_[13269]_  & \new_[13264]_ ;
  assign \new_[13273]_  = A166 & A167;
  assign \new_[13277]_  = A265 & ~A200;
  assign \new_[13278]_  = ~A199 & \new_[13277]_ ;
  assign \new_[13279]_  = \new_[13278]_  & \new_[13273]_ ;
  assign \new_[13282]_  = A267 & ~A266;
  assign \new_[13286]_  = ~A299 & ~A298;
  assign \new_[13287]_  = A269 & \new_[13286]_ ;
  assign \new_[13288]_  = \new_[13287]_  & \new_[13282]_ ;
  assign \new_[13291]_  = ~A166 & ~A167;
  assign \new_[13295]_  = ~A265 & A202;
  assign \new_[13296]_  = ~A201 & \new_[13295]_ ;
  assign \new_[13297]_  = \new_[13296]_  & \new_[13291]_ ;
  assign \new_[13300]_  = A267 & A266;
  assign \new_[13304]_  = A301 & ~A300;
  assign \new_[13305]_  = A268 & \new_[13304]_ ;
  assign \new_[13306]_  = \new_[13305]_  & \new_[13300]_ ;
  assign \new_[13309]_  = ~A166 & ~A167;
  assign \new_[13313]_  = ~A265 & A202;
  assign \new_[13314]_  = ~A201 & \new_[13313]_ ;
  assign \new_[13315]_  = \new_[13314]_  & \new_[13309]_ ;
  assign \new_[13318]_  = A267 & A266;
  assign \new_[13322]_  = A302 & ~A300;
  assign \new_[13323]_  = A268 & \new_[13322]_ ;
  assign \new_[13324]_  = \new_[13323]_  & \new_[13318]_ ;
  assign \new_[13327]_  = ~A166 & ~A167;
  assign \new_[13331]_  = ~A265 & A202;
  assign \new_[13332]_  = ~A201 & \new_[13331]_ ;
  assign \new_[13333]_  = \new_[13332]_  & \new_[13327]_ ;
  assign \new_[13336]_  = A267 & A266;
  assign \new_[13340]_  = A299 & A298;
  assign \new_[13341]_  = A268 & \new_[13340]_ ;
  assign \new_[13342]_  = \new_[13341]_  & \new_[13336]_ ;
  assign \new_[13345]_  = ~A166 & ~A167;
  assign \new_[13349]_  = ~A265 & A202;
  assign \new_[13350]_  = ~A201 & \new_[13349]_ ;
  assign \new_[13351]_  = \new_[13350]_  & \new_[13345]_ ;
  assign \new_[13354]_  = A267 & A266;
  assign \new_[13358]_  = ~A299 & ~A298;
  assign \new_[13359]_  = A268 & \new_[13358]_ ;
  assign \new_[13360]_  = \new_[13359]_  & \new_[13354]_ ;
  assign \new_[13363]_  = ~A166 & ~A167;
  assign \new_[13367]_  = ~A265 & A202;
  assign \new_[13368]_  = ~A201 & \new_[13367]_ ;
  assign \new_[13369]_  = \new_[13368]_  & \new_[13363]_ ;
  assign \new_[13372]_  = A267 & A266;
  assign \new_[13376]_  = A301 & ~A300;
  assign \new_[13377]_  = A269 & \new_[13376]_ ;
  assign \new_[13378]_  = \new_[13377]_  & \new_[13372]_ ;
  assign \new_[13381]_  = ~A166 & ~A167;
  assign \new_[13385]_  = ~A265 & A202;
  assign \new_[13386]_  = ~A201 & \new_[13385]_ ;
  assign \new_[13387]_  = \new_[13386]_  & \new_[13381]_ ;
  assign \new_[13390]_  = A267 & A266;
  assign \new_[13394]_  = A302 & ~A300;
  assign \new_[13395]_  = A269 & \new_[13394]_ ;
  assign \new_[13396]_  = \new_[13395]_  & \new_[13390]_ ;
  assign \new_[13399]_  = ~A166 & ~A167;
  assign \new_[13403]_  = ~A265 & A202;
  assign \new_[13404]_  = ~A201 & \new_[13403]_ ;
  assign \new_[13405]_  = \new_[13404]_  & \new_[13399]_ ;
  assign \new_[13408]_  = A267 & A266;
  assign \new_[13412]_  = A299 & A298;
  assign \new_[13413]_  = A269 & \new_[13412]_ ;
  assign \new_[13414]_  = \new_[13413]_  & \new_[13408]_ ;
  assign \new_[13417]_  = ~A166 & ~A167;
  assign \new_[13421]_  = ~A265 & A202;
  assign \new_[13422]_  = ~A201 & \new_[13421]_ ;
  assign \new_[13423]_  = \new_[13422]_  & \new_[13417]_ ;
  assign \new_[13426]_  = A267 & A266;
  assign \new_[13430]_  = ~A299 & ~A298;
  assign \new_[13431]_  = A269 & \new_[13430]_ ;
  assign \new_[13432]_  = \new_[13431]_  & \new_[13426]_ ;
  assign \new_[13435]_  = ~A166 & ~A167;
  assign \new_[13439]_  = A265 & A202;
  assign \new_[13440]_  = ~A201 & \new_[13439]_ ;
  assign \new_[13441]_  = \new_[13440]_  & \new_[13435]_ ;
  assign \new_[13444]_  = A267 & ~A266;
  assign \new_[13448]_  = A301 & ~A300;
  assign \new_[13449]_  = A268 & \new_[13448]_ ;
  assign \new_[13450]_  = \new_[13449]_  & \new_[13444]_ ;
  assign \new_[13453]_  = ~A166 & ~A167;
  assign \new_[13457]_  = A265 & A202;
  assign \new_[13458]_  = ~A201 & \new_[13457]_ ;
  assign \new_[13459]_  = \new_[13458]_  & \new_[13453]_ ;
  assign \new_[13462]_  = A267 & ~A266;
  assign \new_[13466]_  = A302 & ~A300;
  assign \new_[13467]_  = A268 & \new_[13466]_ ;
  assign \new_[13468]_  = \new_[13467]_  & \new_[13462]_ ;
  assign \new_[13471]_  = ~A166 & ~A167;
  assign \new_[13475]_  = A265 & A202;
  assign \new_[13476]_  = ~A201 & \new_[13475]_ ;
  assign \new_[13477]_  = \new_[13476]_  & \new_[13471]_ ;
  assign \new_[13480]_  = A267 & ~A266;
  assign \new_[13484]_  = A299 & A298;
  assign \new_[13485]_  = A268 & \new_[13484]_ ;
  assign \new_[13486]_  = \new_[13485]_  & \new_[13480]_ ;
  assign \new_[13489]_  = ~A166 & ~A167;
  assign \new_[13493]_  = A265 & A202;
  assign \new_[13494]_  = ~A201 & \new_[13493]_ ;
  assign \new_[13495]_  = \new_[13494]_  & \new_[13489]_ ;
  assign \new_[13498]_  = A267 & ~A266;
  assign \new_[13502]_  = ~A299 & ~A298;
  assign \new_[13503]_  = A268 & \new_[13502]_ ;
  assign \new_[13504]_  = \new_[13503]_  & \new_[13498]_ ;
  assign \new_[13507]_  = ~A166 & ~A167;
  assign \new_[13511]_  = A265 & A202;
  assign \new_[13512]_  = ~A201 & \new_[13511]_ ;
  assign \new_[13513]_  = \new_[13512]_  & \new_[13507]_ ;
  assign \new_[13516]_  = A267 & ~A266;
  assign \new_[13520]_  = A301 & ~A300;
  assign \new_[13521]_  = A269 & \new_[13520]_ ;
  assign \new_[13522]_  = \new_[13521]_  & \new_[13516]_ ;
  assign \new_[13525]_  = ~A166 & ~A167;
  assign \new_[13529]_  = A265 & A202;
  assign \new_[13530]_  = ~A201 & \new_[13529]_ ;
  assign \new_[13531]_  = \new_[13530]_  & \new_[13525]_ ;
  assign \new_[13534]_  = A267 & ~A266;
  assign \new_[13538]_  = A302 & ~A300;
  assign \new_[13539]_  = A269 & \new_[13538]_ ;
  assign \new_[13540]_  = \new_[13539]_  & \new_[13534]_ ;
  assign \new_[13543]_  = ~A166 & ~A167;
  assign \new_[13547]_  = A265 & A202;
  assign \new_[13548]_  = ~A201 & \new_[13547]_ ;
  assign \new_[13549]_  = \new_[13548]_  & \new_[13543]_ ;
  assign \new_[13552]_  = A267 & ~A266;
  assign \new_[13556]_  = A299 & A298;
  assign \new_[13557]_  = A269 & \new_[13556]_ ;
  assign \new_[13558]_  = \new_[13557]_  & \new_[13552]_ ;
  assign \new_[13561]_  = ~A166 & ~A167;
  assign \new_[13565]_  = A265 & A202;
  assign \new_[13566]_  = ~A201 & \new_[13565]_ ;
  assign \new_[13567]_  = \new_[13566]_  & \new_[13561]_ ;
  assign \new_[13570]_  = A267 & ~A266;
  assign \new_[13574]_  = ~A299 & ~A298;
  assign \new_[13575]_  = A269 & \new_[13574]_ ;
  assign \new_[13576]_  = \new_[13575]_  & \new_[13570]_ ;
  assign \new_[13579]_  = ~A166 & ~A167;
  assign \new_[13583]_  = ~A265 & A203;
  assign \new_[13584]_  = ~A201 & \new_[13583]_ ;
  assign \new_[13585]_  = \new_[13584]_  & \new_[13579]_ ;
  assign \new_[13588]_  = A267 & A266;
  assign \new_[13592]_  = A301 & ~A300;
  assign \new_[13593]_  = A268 & \new_[13592]_ ;
  assign \new_[13594]_  = \new_[13593]_  & \new_[13588]_ ;
  assign \new_[13597]_  = ~A166 & ~A167;
  assign \new_[13601]_  = ~A265 & A203;
  assign \new_[13602]_  = ~A201 & \new_[13601]_ ;
  assign \new_[13603]_  = \new_[13602]_  & \new_[13597]_ ;
  assign \new_[13606]_  = A267 & A266;
  assign \new_[13610]_  = A302 & ~A300;
  assign \new_[13611]_  = A268 & \new_[13610]_ ;
  assign \new_[13612]_  = \new_[13611]_  & \new_[13606]_ ;
  assign \new_[13615]_  = ~A166 & ~A167;
  assign \new_[13619]_  = ~A265 & A203;
  assign \new_[13620]_  = ~A201 & \new_[13619]_ ;
  assign \new_[13621]_  = \new_[13620]_  & \new_[13615]_ ;
  assign \new_[13624]_  = A267 & A266;
  assign \new_[13628]_  = A299 & A298;
  assign \new_[13629]_  = A268 & \new_[13628]_ ;
  assign \new_[13630]_  = \new_[13629]_  & \new_[13624]_ ;
  assign \new_[13633]_  = ~A166 & ~A167;
  assign \new_[13637]_  = ~A265 & A203;
  assign \new_[13638]_  = ~A201 & \new_[13637]_ ;
  assign \new_[13639]_  = \new_[13638]_  & \new_[13633]_ ;
  assign \new_[13642]_  = A267 & A266;
  assign \new_[13646]_  = ~A299 & ~A298;
  assign \new_[13647]_  = A268 & \new_[13646]_ ;
  assign \new_[13648]_  = \new_[13647]_  & \new_[13642]_ ;
  assign \new_[13651]_  = ~A166 & ~A167;
  assign \new_[13655]_  = ~A265 & A203;
  assign \new_[13656]_  = ~A201 & \new_[13655]_ ;
  assign \new_[13657]_  = \new_[13656]_  & \new_[13651]_ ;
  assign \new_[13660]_  = A267 & A266;
  assign \new_[13664]_  = A301 & ~A300;
  assign \new_[13665]_  = A269 & \new_[13664]_ ;
  assign \new_[13666]_  = \new_[13665]_  & \new_[13660]_ ;
  assign \new_[13669]_  = ~A166 & ~A167;
  assign \new_[13673]_  = ~A265 & A203;
  assign \new_[13674]_  = ~A201 & \new_[13673]_ ;
  assign \new_[13675]_  = \new_[13674]_  & \new_[13669]_ ;
  assign \new_[13678]_  = A267 & A266;
  assign \new_[13682]_  = A302 & ~A300;
  assign \new_[13683]_  = A269 & \new_[13682]_ ;
  assign \new_[13684]_  = \new_[13683]_  & \new_[13678]_ ;
  assign \new_[13687]_  = ~A166 & ~A167;
  assign \new_[13691]_  = ~A265 & A203;
  assign \new_[13692]_  = ~A201 & \new_[13691]_ ;
  assign \new_[13693]_  = \new_[13692]_  & \new_[13687]_ ;
  assign \new_[13696]_  = A267 & A266;
  assign \new_[13700]_  = A299 & A298;
  assign \new_[13701]_  = A269 & \new_[13700]_ ;
  assign \new_[13702]_  = \new_[13701]_  & \new_[13696]_ ;
  assign \new_[13705]_  = ~A166 & ~A167;
  assign \new_[13709]_  = ~A265 & A203;
  assign \new_[13710]_  = ~A201 & \new_[13709]_ ;
  assign \new_[13711]_  = \new_[13710]_  & \new_[13705]_ ;
  assign \new_[13714]_  = A267 & A266;
  assign \new_[13718]_  = ~A299 & ~A298;
  assign \new_[13719]_  = A269 & \new_[13718]_ ;
  assign \new_[13720]_  = \new_[13719]_  & \new_[13714]_ ;
  assign \new_[13723]_  = ~A166 & ~A167;
  assign \new_[13727]_  = A265 & A203;
  assign \new_[13728]_  = ~A201 & \new_[13727]_ ;
  assign \new_[13729]_  = \new_[13728]_  & \new_[13723]_ ;
  assign \new_[13732]_  = A267 & ~A266;
  assign \new_[13736]_  = A301 & ~A300;
  assign \new_[13737]_  = A268 & \new_[13736]_ ;
  assign \new_[13738]_  = \new_[13737]_  & \new_[13732]_ ;
  assign \new_[13741]_  = ~A166 & ~A167;
  assign \new_[13745]_  = A265 & A203;
  assign \new_[13746]_  = ~A201 & \new_[13745]_ ;
  assign \new_[13747]_  = \new_[13746]_  & \new_[13741]_ ;
  assign \new_[13750]_  = A267 & ~A266;
  assign \new_[13754]_  = A302 & ~A300;
  assign \new_[13755]_  = A268 & \new_[13754]_ ;
  assign \new_[13756]_  = \new_[13755]_  & \new_[13750]_ ;
  assign \new_[13759]_  = ~A166 & ~A167;
  assign \new_[13763]_  = A265 & A203;
  assign \new_[13764]_  = ~A201 & \new_[13763]_ ;
  assign \new_[13765]_  = \new_[13764]_  & \new_[13759]_ ;
  assign \new_[13768]_  = A267 & ~A266;
  assign \new_[13772]_  = A299 & A298;
  assign \new_[13773]_  = A268 & \new_[13772]_ ;
  assign \new_[13774]_  = \new_[13773]_  & \new_[13768]_ ;
  assign \new_[13777]_  = ~A166 & ~A167;
  assign \new_[13781]_  = A265 & A203;
  assign \new_[13782]_  = ~A201 & \new_[13781]_ ;
  assign \new_[13783]_  = \new_[13782]_  & \new_[13777]_ ;
  assign \new_[13786]_  = A267 & ~A266;
  assign \new_[13790]_  = ~A299 & ~A298;
  assign \new_[13791]_  = A268 & \new_[13790]_ ;
  assign \new_[13792]_  = \new_[13791]_  & \new_[13786]_ ;
  assign \new_[13795]_  = ~A166 & ~A167;
  assign \new_[13799]_  = A265 & A203;
  assign \new_[13800]_  = ~A201 & \new_[13799]_ ;
  assign \new_[13801]_  = \new_[13800]_  & \new_[13795]_ ;
  assign \new_[13804]_  = A267 & ~A266;
  assign \new_[13808]_  = A301 & ~A300;
  assign \new_[13809]_  = A269 & \new_[13808]_ ;
  assign \new_[13810]_  = \new_[13809]_  & \new_[13804]_ ;
  assign \new_[13813]_  = ~A166 & ~A167;
  assign \new_[13817]_  = A265 & A203;
  assign \new_[13818]_  = ~A201 & \new_[13817]_ ;
  assign \new_[13819]_  = \new_[13818]_  & \new_[13813]_ ;
  assign \new_[13822]_  = A267 & ~A266;
  assign \new_[13826]_  = A302 & ~A300;
  assign \new_[13827]_  = A269 & \new_[13826]_ ;
  assign \new_[13828]_  = \new_[13827]_  & \new_[13822]_ ;
  assign \new_[13831]_  = ~A166 & ~A167;
  assign \new_[13835]_  = A265 & A203;
  assign \new_[13836]_  = ~A201 & \new_[13835]_ ;
  assign \new_[13837]_  = \new_[13836]_  & \new_[13831]_ ;
  assign \new_[13840]_  = A267 & ~A266;
  assign \new_[13844]_  = A299 & A298;
  assign \new_[13845]_  = A269 & \new_[13844]_ ;
  assign \new_[13846]_  = \new_[13845]_  & \new_[13840]_ ;
  assign \new_[13849]_  = ~A166 & ~A167;
  assign \new_[13853]_  = A265 & A203;
  assign \new_[13854]_  = ~A201 & \new_[13853]_ ;
  assign \new_[13855]_  = \new_[13854]_  & \new_[13849]_ ;
  assign \new_[13858]_  = A267 & ~A266;
  assign \new_[13862]_  = ~A299 & ~A298;
  assign \new_[13863]_  = A269 & \new_[13862]_ ;
  assign \new_[13864]_  = \new_[13863]_  & \new_[13858]_ ;
  assign \new_[13867]_  = ~A166 & ~A167;
  assign \new_[13871]_  = ~A265 & A200;
  assign \new_[13872]_  = A199 & \new_[13871]_ ;
  assign \new_[13873]_  = \new_[13872]_  & \new_[13867]_ ;
  assign \new_[13876]_  = A267 & A266;
  assign \new_[13880]_  = A301 & ~A300;
  assign \new_[13881]_  = A268 & \new_[13880]_ ;
  assign \new_[13882]_  = \new_[13881]_  & \new_[13876]_ ;
  assign \new_[13885]_  = ~A166 & ~A167;
  assign \new_[13889]_  = ~A265 & A200;
  assign \new_[13890]_  = A199 & \new_[13889]_ ;
  assign \new_[13891]_  = \new_[13890]_  & \new_[13885]_ ;
  assign \new_[13894]_  = A267 & A266;
  assign \new_[13898]_  = A302 & ~A300;
  assign \new_[13899]_  = A268 & \new_[13898]_ ;
  assign \new_[13900]_  = \new_[13899]_  & \new_[13894]_ ;
  assign \new_[13903]_  = ~A166 & ~A167;
  assign \new_[13907]_  = ~A265 & A200;
  assign \new_[13908]_  = A199 & \new_[13907]_ ;
  assign \new_[13909]_  = \new_[13908]_  & \new_[13903]_ ;
  assign \new_[13912]_  = A267 & A266;
  assign \new_[13916]_  = A299 & A298;
  assign \new_[13917]_  = A268 & \new_[13916]_ ;
  assign \new_[13918]_  = \new_[13917]_  & \new_[13912]_ ;
  assign \new_[13921]_  = ~A166 & ~A167;
  assign \new_[13925]_  = ~A265 & A200;
  assign \new_[13926]_  = A199 & \new_[13925]_ ;
  assign \new_[13927]_  = \new_[13926]_  & \new_[13921]_ ;
  assign \new_[13930]_  = A267 & A266;
  assign \new_[13934]_  = ~A299 & ~A298;
  assign \new_[13935]_  = A268 & \new_[13934]_ ;
  assign \new_[13936]_  = \new_[13935]_  & \new_[13930]_ ;
  assign \new_[13939]_  = ~A166 & ~A167;
  assign \new_[13943]_  = ~A265 & A200;
  assign \new_[13944]_  = A199 & \new_[13943]_ ;
  assign \new_[13945]_  = \new_[13944]_  & \new_[13939]_ ;
  assign \new_[13948]_  = A267 & A266;
  assign \new_[13952]_  = A301 & ~A300;
  assign \new_[13953]_  = A269 & \new_[13952]_ ;
  assign \new_[13954]_  = \new_[13953]_  & \new_[13948]_ ;
  assign \new_[13957]_  = ~A166 & ~A167;
  assign \new_[13961]_  = ~A265 & A200;
  assign \new_[13962]_  = A199 & \new_[13961]_ ;
  assign \new_[13963]_  = \new_[13962]_  & \new_[13957]_ ;
  assign \new_[13966]_  = A267 & A266;
  assign \new_[13970]_  = A302 & ~A300;
  assign \new_[13971]_  = A269 & \new_[13970]_ ;
  assign \new_[13972]_  = \new_[13971]_  & \new_[13966]_ ;
  assign \new_[13975]_  = ~A166 & ~A167;
  assign \new_[13979]_  = ~A265 & A200;
  assign \new_[13980]_  = A199 & \new_[13979]_ ;
  assign \new_[13981]_  = \new_[13980]_  & \new_[13975]_ ;
  assign \new_[13984]_  = A267 & A266;
  assign \new_[13988]_  = A299 & A298;
  assign \new_[13989]_  = A269 & \new_[13988]_ ;
  assign \new_[13990]_  = \new_[13989]_  & \new_[13984]_ ;
  assign \new_[13993]_  = ~A166 & ~A167;
  assign \new_[13997]_  = ~A265 & A200;
  assign \new_[13998]_  = A199 & \new_[13997]_ ;
  assign \new_[13999]_  = \new_[13998]_  & \new_[13993]_ ;
  assign \new_[14002]_  = A267 & A266;
  assign \new_[14006]_  = ~A299 & ~A298;
  assign \new_[14007]_  = A269 & \new_[14006]_ ;
  assign \new_[14008]_  = \new_[14007]_  & \new_[14002]_ ;
  assign \new_[14011]_  = ~A166 & ~A167;
  assign \new_[14015]_  = A265 & A200;
  assign \new_[14016]_  = A199 & \new_[14015]_ ;
  assign \new_[14017]_  = \new_[14016]_  & \new_[14011]_ ;
  assign \new_[14020]_  = A267 & ~A266;
  assign \new_[14024]_  = A301 & ~A300;
  assign \new_[14025]_  = A268 & \new_[14024]_ ;
  assign \new_[14026]_  = \new_[14025]_  & \new_[14020]_ ;
  assign \new_[14029]_  = ~A166 & ~A167;
  assign \new_[14033]_  = A265 & A200;
  assign \new_[14034]_  = A199 & \new_[14033]_ ;
  assign \new_[14035]_  = \new_[14034]_  & \new_[14029]_ ;
  assign \new_[14038]_  = A267 & ~A266;
  assign \new_[14042]_  = A302 & ~A300;
  assign \new_[14043]_  = A268 & \new_[14042]_ ;
  assign \new_[14044]_  = \new_[14043]_  & \new_[14038]_ ;
  assign \new_[14047]_  = ~A166 & ~A167;
  assign \new_[14051]_  = A265 & A200;
  assign \new_[14052]_  = A199 & \new_[14051]_ ;
  assign \new_[14053]_  = \new_[14052]_  & \new_[14047]_ ;
  assign \new_[14056]_  = A267 & ~A266;
  assign \new_[14060]_  = A299 & A298;
  assign \new_[14061]_  = A268 & \new_[14060]_ ;
  assign \new_[14062]_  = \new_[14061]_  & \new_[14056]_ ;
  assign \new_[14065]_  = ~A166 & ~A167;
  assign \new_[14069]_  = A265 & A200;
  assign \new_[14070]_  = A199 & \new_[14069]_ ;
  assign \new_[14071]_  = \new_[14070]_  & \new_[14065]_ ;
  assign \new_[14074]_  = A267 & ~A266;
  assign \new_[14078]_  = ~A299 & ~A298;
  assign \new_[14079]_  = A268 & \new_[14078]_ ;
  assign \new_[14080]_  = \new_[14079]_  & \new_[14074]_ ;
  assign \new_[14083]_  = ~A166 & ~A167;
  assign \new_[14087]_  = A265 & A200;
  assign \new_[14088]_  = A199 & \new_[14087]_ ;
  assign \new_[14089]_  = \new_[14088]_  & \new_[14083]_ ;
  assign \new_[14092]_  = A267 & ~A266;
  assign \new_[14096]_  = A301 & ~A300;
  assign \new_[14097]_  = A269 & \new_[14096]_ ;
  assign \new_[14098]_  = \new_[14097]_  & \new_[14092]_ ;
  assign \new_[14101]_  = ~A166 & ~A167;
  assign \new_[14105]_  = A265 & A200;
  assign \new_[14106]_  = A199 & \new_[14105]_ ;
  assign \new_[14107]_  = \new_[14106]_  & \new_[14101]_ ;
  assign \new_[14110]_  = A267 & ~A266;
  assign \new_[14114]_  = A302 & ~A300;
  assign \new_[14115]_  = A269 & \new_[14114]_ ;
  assign \new_[14116]_  = \new_[14115]_  & \new_[14110]_ ;
  assign \new_[14119]_  = ~A166 & ~A167;
  assign \new_[14123]_  = A265 & A200;
  assign \new_[14124]_  = A199 & \new_[14123]_ ;
  assign \new_[14125]_  = \new_[14124]_  & \new_[14119]_ ;
  assign \new_[14128]_  = A267 & ~A266;
  assign \new_[14132]_  = A299 & A298;
  assign \new_[14133]_  = A269 & \new_[14132]_ ;
  assign \new_[14134]_  = \new_[14133]_  & \new_[14128]_ ;
  assign \new_[14137]_  = ~A166 & ~A167;
  assign \new_[14141]_  = A265 & A200;
  assign \new_[14142]_  = A199 & \new_[14141]_ ;
  assign \new_[14143]_  = \new_[14142]_  & \new_[14137]_ ;
  assign \new_[14146]_  = A267 & ~A266;
  assign \new_[14150]_  = ~A299 & ~A298;
  assign \new_[14151]_  = A269 & \new_[14150]_ ;
  assign \new_[14152]_  = \new_[14151]_  & \new_[14146]_ ;
  assign \new_[14155]_  = ~A166 & ~A167;
  assign \new_[14159]_  = ~A265 & ~A200;
  assign \new_[14160]_  = ~A199 & \new_[14159]_ ;
  assign \new_[14161]_  = \new_[14160]_  & \new_[14155]_ ;
  assign \new_[14164]_  = A267 & A266;
  assign \new_[14168]_  = A301 & ~A300;
  assign \new_[14169]_  = A268 & \new_[14168]_ ;
  assign \new_[14170]_  = \new_[14169]_  & \new_[14164]_ ;
  assign \new_[14173]_  = ~A166 & ~A167;
  assign \new_[14177]_  = ~A265 & ~A200;
  assign \new_[14178]_  = ~A199 & \new_[14177]_ ;
  assign \new_[14179]_  = \new_[14178]_  & \new_[14173]_ ;
  assign \new_[14182]_  = A267 & A266;
  assign \new_[14186]_  = A302 & ~A300;
  assign \new_[14187]_  = A268 & \new_[14186]_ ;
  assign \new_[14188]_  = \new_[14187]_  & \new_[14182]_ ;
  assign \new_[14191]_  = ~A166 & ~A167;
  assign \new_[14195]_  = ~A265 & ~A200;
  assign \new_[14196]_  = ~A199 & \new_[14195]_ ;
  assign \new_[14197]_  = \new_[14196]_  & \new_[14191]_ ;
  assign \new_[14200]_  = A267 & A266;
  assign \new_[14204]_  = A299 & A298;
  assign \new_[14205]_  = A268 & \new_[14204]_ ;
  assign \new_[14206]_  = \new_[14205]_  & \new_[14200]_ ;
  assign \new_[14209]_  = ~A166 & ~A167;
  assign \new_[14213]_  = ~A265 & ~A200;
  assign \new_[14214]_  = ~A199 & \new_[14213]_ ;
  assign \new_[14215]_  = \new_[14214]_  & \new_[14209]_ ;
  assign \new_[14218]_  = A267 & A266;
  assign \new_[14222]_  = ~A299 & ~A298;
  assign \new_[14223]_  = A268 & \new_[14222]_ ;
  assign \new_[14224]_  = \new_[14223]_  & \new_[14218]_ ;
  assign \new_[14227]_  = ~A166 & ~A167;
  assign \new_[14231]_  = ~A265 & ~A200;
  assign \new_[14232]_  = ~A199 & \new_[14231]_ ;
  assign \new_[14233]_  = \new_[14232]_  & \new_[14227]_ ;
  assign \new_[14236]_  = A267 & A266;
  assign \new_[14240]_  = A301 & ~A300;
  assign \new_[14241]_  = A269 & \new_[14240]_ ;
  assign \new_[14242]_  = \new_[14241]_  & \new_[14236]_ ;
  assign \new_[14245]_  = ~A166 & ~A167;
  assign \new_[14249]_  = ~A265 & ~A200;
  assign \new_[14250]_  = ~A199 & \new_[14249]_ ;
  assign \new_[14251]_  = \new_[14250]_  & \new_[14245]_ ;
  assign \new_[14254]_  = A267 & A266;
  assign \new_[14258]_  = A302 & ~A300;
  assign \new_[14259]_  = A269 & \new_[14258]_ ;
  assign \new_[14260]_  = \new_[14259]_  & \new_[14254]_ ;
  assign \new_[14263]_  = ~A166 & ~A167;
  assign \new_[14267]_  = ~A265 & ~A200;
  assign \new_[14268]_  = ~A199 & \new_[14267]_ ;
  assign \new_[14269]_  = \new_[14268]_  & \new_[14263]_ ;
  assign \new_[14272]_  = A267 & A266;
  assign \new_[14276]_  = A299 & A298;
  assign \new_[14277]_  = A269 & \new_[14276]_ ;
  assign \new_[14278]_  = \new_[14277]_  & \new_[14272]_ ;
  assign \new_[14281]_  = ~A166 & ~A167;
  assign \new_[14285]_  = ~A265 & ~A200;
  assign \new_[14286]_  = ~A199 & \new_[14285]_ ;
  assign \new_[14287]_  = \new_[14286]_  & \new_[14281]_ ;
  assign \new_[14290]_  = A267 & A266;
  assign \new_[14294]_  = ~A299 & ~A298;
  assign \new_[14295]_  = A269 & \new_[14294]_ ;
  assign \new_[14296]_  = \new_[14295]_  & \new_[14290]_ ;
  assign \new_[14299]_  = ~A166 & ~A167;
  assign \new_[14303]_  = A265 & ~A200;
  assign \new_[14304]_  = ~A199 & \new_[14303]_ ;
  assign \new_[14305]_  = \new_[14304]_  & \new_[14299]_ ;
  assign \new_[14308]_  = A267 & ~A266;
  assign \new_[14312]_  = A301 & ~A300;
  assign \new_[14313]_  = A268 & \new_[14312]_ ;
  assign \new_[14314]_  = \new_[14313]_  & \new_[14308]_ ;
  assign \new_[14317]_  = ~A166 & ~A167;
  assign \new_[14321]_  = A265 & ~A200;
  assign \new_[14322]_  = ~A199 & \new_[14321]_ ;
  assign \new_[14323]_  = \new_[14322]_  & \new_[14317]_ ;
  assign \new_[14326]_  = A267 & ~A266;
  assign \new_[14330]_  = A302 & ~A300;
  assign \new_[14331]_  = A268 & \new_[14330]_ ;
  assign \new_[14332]_  = \new_[14331]_  & \new_[14326]_ ;
  assign \new_[14335]_  = ~A166 & ~A167;
  assign \new_[14339]_  = A265 & ~A200;
  assign \new_[14340]_  = ~A199 & \new_[14339]_ ;
  assign \new_[14341]_  = \new_[14340]_  & \new_[14335]_ ;
  assign \new_[14344]_  = A267 & ~A266;
  assign \new_[14348]_  = A299 & A298;
  assign \new_[14349]_  = A268 & \new_[14348]_ ;
  assign \new_[14350]_  = \new_[14349]_  & \new_[14344]_ ;
  assign \new_[14353]_  = ~A166 & ~A167;
  assign \new_[14357]_  = A265 & ~A200;
  assign \new_[14358]_  = ~A199 & \new_[14357]_ ;
  assign \new_[14359]_  = \new_[14358]_  & \new_[14353]_ ;
  assign \new_[14362]_  = A267 & ~A266;
  assign \new_[14366]_  = ~A299 & ~A298;
  assign \new_[14367]_  = A268 & \new_[14366]_ ;
  assign \new_[14368]_  = \new_[14367]_  & \new_[14362]_ ;
  assign \new_[14371]_  = ~A166 & ~A167;
  assign \new_[14375]_  = A265 & ~A200;
  assign \new_[14376]_  = ~A199 & \new_[14375]_ ;
  assign \new_[14377]_  = \new_[14376]_  & \new_[14371]_ ;
  assign \new_[14380]_  = A267 & ~A266;
  assign \new_[14384]_  = A301 & ~A300;
  assign \new_[14385]_  = A269 & \new_[14384]_ ;
  assign \new_[14386]_  = \new_[14385]_  & \new_[14380]_ ;
  assign \new_[14389]_  = ~A166 & ~A167;
  assign \new_[14393]_  = A265 & ~A200;
  assign \new_[14394]_  = ~A199 & \new_[14393]_ ;
  assign \new_[14395]_  = \new_[14394]_  & \new_[14389]_ ;
  assign \new_[14398]_  = A267 & ~A266;
  assign \new_[14402]_  = A302 & ~A300;
  assign \new_[14403]_  = A269 & \new_[14402]_ ;
  assign \new_[14404]_  = \new_[14403]_  & \new_[14398]_ ;
  assign \new_[14407]_  = ~A166 & ~A167;
  assign \new_[14411]_  = A265 & ~A200;
  assign \new_[14412]_  = ~A199 & \new_[14411]_ ;
  assign \new_[14413]_  = \new_[14412]_  & \new_[14407]_ ;
  assign \new_[14416]_  = A267 & ~A266;
  assign \new_[14420]_  = A299 & A298;
  assign \new_[14421]_  = A269 & \new_[14420]_ ;
  assign \new_[14422]_  = \new_[14421]_  & \new_[14416]_ ;
  assign \new_[14425]_  = ~A166 & ~A167;
  assign \new_[14429]_  = A265 & ~A200;
  assign \new_[14430]_  = ~A199 & \new_[14429]_ ;
  assign \new_[14431]_  = \new_[14430]_  & \new_[14425]_ ;
  assign \new_[14434]_  = A267 & ~A266;
  assign \new_[14438]_  = ~A299 & ~A298;
  assign \new_[14439]_  = A269 & \new_[14438]_ ;
  assign \new_[14440]_  = \new_[14439]_  & \new_[14434]_ ;
  assign \new_[14443]_  = ~A168 & ~A170;
  assign \new_[14447]_  = ~A265 & A202;
  assign \new_[14448]_  = ~A201 & \new_[14447]_ ;
  assign \new_[14449]_  = \new_[14448]_  & \new_[14443]_ ;
  assign \new_[14452]_  = A267 & A266;
  assign \new_[14456]_  = A301 & ~A300;
  assign \new_[14457]_  = A268 & \new_[14456]_ ;
  assign \new_[14458]_  = \new_[14457]_  & \new_[14452]_ ;
  assign \new_[14461]_  = ~A168 & ~A170;
  assign \new_[14465]_  = ~A265 & A202;
  assign \new_[14466]_  = ~A201 & \new_[14465]_ ;
  assign \new_[14467]_  = \new_[14466]_  & \new_[14461]_ ;
  assign \new_[14470]_  = A267 & A266;
  assign \new_[14474]_  = A302 & ~A300;
  assign \new_[14475]_  = A268 & \new_[14474]_ ;
  assign \new_[14476]_  = \new_[14475]_  & \new_[14470]_ ;
  assign \new_[14479]_  = ~A168 & ~A170;
  assign \new_[14483]_  = ~A265 & A202;
  assign \new_[14484]_  = ~A201 & \new_[14483]_ ;
  assign \new_[14485]_  = \new_[14484]_  & \new_[14479]_ ;
  assign \new_[14488]_  = A267 & A266;
  assign \new_[14492]_  = A299 & A298;
  assign \new_[14493]_  = A268 & \new_[14492]_ ;
  assign \new_[14494]_  = \new_[14493]_  & \new_[14488]_ ;
  assign \new_[14497]_  = ~A168 & ~A170;
  assign \new_[14501]_  = ~A265 & A202;
  assign \new_[14502]_  = ~A201 & \new_[14501]_ ;
  assign \new_[14503]_  = \new_[14502]_  & \new_[14497]_ ;
  assign \new_[14506]_  = A267 & A266;
  assign \new_[14510]_  = ~A299 & ~A298;
  assign \new_[14511]_  = A268 & \new_[14510]_ ;
  assign \new_[14512]_  = \new_[14511]_  & \new_[14506]_ ;
  assign \new_[14515]_  = ~A168 & ~A170;
  assign \new_[14519]_  = ~A265 & A202;
  assign \new_[14520]_  = ~A201 & \new_[14519]_ ;
  assign \new_[14521]_  = \new_[14520]_  & \new_[14515]_ ;
  assign \new_[14524]_  = A267 & A266;
  assign \new_[14528]_  = A301 & ~A300;
  assign \new_[14529]_  = A269 & \new_[14528]_ ;
  assign \new_[14530]_  = \new_[14529]_  & \new_[14524]_ ;
  assign \new_[14533]_  = ~A168 & ~A170;
  assign \new_[14537]_  = ~A265 & A202;
  assign \new_[14538]_  = ~A201 & \new_[14537]_ ;
  assign \new_[14539]_  = \new_[14538]_  & \new_[14533]_ ;
  assign \new_[14542]_  = A267 & A266;
  assign \new_[14546]_  = A302 & ~A300;
  assign \new_[14547]_  = A269 & \new_[14546]_ ;
  assign \new_[14548]_  = \new_[14547]_  & \new_[14542]_ ;
  assign \new_[14551]_  = ~A168 & ~A170;
  assign \new_[14555]_  = ~A265 & A202;
  assign \new_[14556]_  = ~A201 & \new_[14555]_ ;
  assign \new_[14557]_  = \new_[14556]_  & \new_[14551]_ ;
  assign \new_[14560]_  = A267 & A266;
  assign \new_[14564]_  = A299 & A298;
  assign \new_[14565]_  = A269 & \new_[14564]_ ;
  assign \new_[14566]_  = \new_[14565]_  & \new_[14560]_ ;
  assign \new_[14569]_  = ~A168 & ~A170;
  assign \new_[14573]_  = ~A265 & A202;
  assign \new_[14574]_  = ~A201 & \new_[14573]_ ;
  assign \new_[14575]_  = \new_[14574]_  & \new_[14569]_ ;
  assign \new_[14578]_  = A267 & A266;
  assign \new_[14582]_  = ~A299 & ~A298;
  assign \new_[14583]_  = A269 & \new_[14582]_ ;
  assign \new_[14584]_  = \new_[14583]_  & \new_[14578]_ ;
  assign \new_[14587]_  = ~A168 & ~A170;
  assign \new_[14591]_  = A265 & A202;
  assign \new_[14592]_  = ~A201 & \new_[14591]_ ;
  assign \new_[14593]_  = \new_[14592]_  & \new_[14587]_ ;
  assign \new_[14596]_  = A267 & ~A266;
  assign \new_[14600]_  = A301 & ~A300;
  assign \new_[14601]_  = A268 & \new_[14600]_ ;
  assign \new_[14602]_  = \new_[14601]_  & \new_[14596]_ ;
  assign \new_[14605]_  = ~A168 & ~A170;
  assign \new_[14609]_  = A265 & A202;
  assign \new_[14610]_  = ~A201 & \new_[14609]_ ;
  assign \new_[14611]_  = \new_[14610]_  & \new_[14605]_ ;
  assign \new_[14614]_  = A267 & ~A266;
  assign \new_[14618]_  = A302 & ~A300;
  assign \new_[14619]_  = A268 & \new_[14618]_ ;
  assign \new_[14620]_  = \new_[14619]_  & \new_[14614]_ ;
  assign \new_[14623]_  = ~A168 & ~A170;
  assign \new_[14627]_  = A265 & A202;
  assign \new_[14628]_  = ~A201 & \new_[14627]_ ;
  assign \new_[14629]_  = \new_[14628]_  & \new_[14623]_ ;
  assign \new_[14632]_  = A267 & ~A266;
  assign \new_[14636]_  = A299 & A298;
  assign \new_[14637]_  = A268 & \new_[14636]_ ;
  assign \new_[14638]_  = \new_[14637]_  & \new_[14632]_ ;
  assign \new_[14641]_  = ~A168 & ~A170;
  assign \new_[14645]_  = A265 & A202;
  assign \new_[14646]_  = ~A201 & \new_[14645]_ ;
  assign \new_[14647]_  = \new_[14646]_  & \new_[14641]_ ;
  assign \new_[14650]_  = A267 & ~A266;
  assign \new_[14654]_  = ~A299 & ~A298;
  assign \new_[14655]_  = A268 & \new_[14654]_ ;
  assign \new_[14656]_  = \new_[14655]_  & \new_[14650]_ ;
  assign \new_[14659]_  = ~A168 & ~A170;
  assign \new_[14663]_  = A265 & A202;
  assign \new_[14664]_  = ~A201 & \new_[14663]_ ;
  assign \new_[14665]_  = \new_[14664]_  & \new_[14659]_ ;
  assign \new_[14668]_  = A267 & ~A266;
  assign \new_[14672]_  = A301 & ~A300;
  assign \new_[14673]_  = A269 & \new_[14672]_ ;
  assign \new_[14674]_  = \new_[14673]_  & \new_[14668]_ ;
  assign \new_[14677]_  = ~A168 & ~A170;
  assign \new_[14681]_  = A265 & A202;
  assign \new_[14682]_  = ~A201 & \new_[14681]_ ;
  assign \new_[14683]_  = \new_[14682]_  & \new_[14677]_ ;
  assign \new_[14686]_  = A267 & ~A266;
  assign \new_[14690]_  = A302 & ~A300;
  assign \new_[14691]_  = A269 & \new_[14690]_ ;
  assign \new_[14692]_  = \new_[14691]_  & \new_[14686]_ ;
  assign \new_[14695]_  = ~A168 & ~A170;
  assign \new_[14699]_  = A265 & A202;
  assign \new_[14700]_  = ~A201 & \new_[14699]_ ;
  assign \new_[14701]_  = \new_[14700]_  & \new_[14695]_ ;
  assign \new_[14704]_  = A267 & ~A266;
  assign \new_[14708]_  = A299 & A298;
  assign \new_[14709]_  = A269 & \new_[14708]_ ;
  assign \new_[14710]_  = \new_[14709]_  & \new_[14704]_ ;
  assign \new_[14713]_  = ~A168 & ~A170;
  assign \new_[14717]_  = A265 & A202;
  assign \new_[14718]_  = ~A201 & \new_[14717]_ ;
  assign \new_[14719]_  = \new_[14718]_  & \new_[14713]_ ;
  assign \new_[14722]_  = A267 & ~A266;
  assign \new_[14726]_  = ~A299 & ~A298;
  assign \new_[14727]_  = A269 & \new_[14726]_ ;
  assign \new_[14728]_  = \new_[14727]_  & \new_[14722]_ ;
  assign \new_[14731]_  = ~A168 & ~A170;
  assign \new_[14735]_  = ~A265 & A203;
  assign \new_[14736]_  = ~A201 & \new_[14735]_ ;
  assign \new_[14737]_  = \new_[14736]_  & \new_[14731]_ ;
  assign \new_[14740]_  = A267 & A266;
  assign \new_[14744]_  = A301 & ~A300;
  assign \new_[14745]_  = A268 & \new_[14744]_ ;
  assign \new_[14746]_  = \new_[14745]_  & \new_[14740]_ ;
  assign \new_[14749]_  = ~A168 & ~A170;
  assign \new_[14753]_  = ~A265 & A203;
  assign \new_[14754]_  = ~A201 & \new_[14753]_ ;
  assign \new_[14755]_  = \new_[14754]_  & \new_[14749]_ ;
  assign \new_[14758]_  = A267 & A266;
  assign \new_[14762]_  = A302 & ~A300;
  assign \new_[14763]_  = A268 & \new_[14762]_ ;
  assign \new_[14764]_  = \new_[14763]_  & \new_[14758]_ ;
  assign \new_[14767]_  = ~A168 & ~A170;
  assign \new_[14771]_  = ~A265 & A203;
  assign \new_[14772]_  = ~A201 & \new_[14771]_ ;
  assign \new_[14773]_  = \new_[14772]_  & \new_[14767]_ ;
  assign \new_[14776]_  = A267 & A266;
  assign \new_[14780]_  = A299 & A298;
  assign \new_[14781]_  = A268 & \new_[14780]_ ;
  assign \new_[14782]_  = \new_[14781]_  & \new_[14776]_ ;
  assign \new_[14785]_  = ~A168 & ~A170;
  assign \new_[14789]_  = ~A265 & A203;
  assign \new_[14790]_  = ~A201 & \new_[14789]_ ;
  assign \new_[14791]_  = \new_[14790]_  & \new_[14785]_ ;
  assign \new_[14794]_  = A267 & A266;
  assign \new_[14798]_  = ~A299 & ~A298;
  assign \new_[14799]_  = A268 & \new_[14798]_ ;
  assign \new_[14800]_  = \new_[14799]_  & \new_[14794]_ ;
  assign \new_[14803]_  = ~A168 & ~A170;
  assign \new_[14807]_  = ~A265 & A203;
  assign \new_[14808]_  = ~A201 & \new_[14807]_ ;
  assign \new_[14809]_  = \new_[14808]_  & \new_[14803]_ ;
  assign \new_[14812]_  = A267 & A266;
  assign \new_[14816]_  = A301 & ~A300;
  assign \new_[14817]_  = A269 & \new_[14816]_ ;
  assign \new_[14818]_  = \new_[14817]_  & \new_[14812]_ ;
  assign \new_[14821]_  = ~A168 & ~A170;
  assign \new_[14825]_  = ~A265 & A203;
  assign \new_[14826]_  = ~A201 & \new_[14825]_ ;
  assign \new_[14827]_  = \new_[14826]_  & \new_[14821]_ ;
  assign \new_[14830]_  = A267 & A266;
  assign \new_[14834]_  = A302 & ~A300;
  assign \new_[14835]_  = A269 & \new_[14834]_ ;
  assign \new_[14836]_  = \new_[14835]_  & \new_[14830]_ ;
  assign \new_[14839]_  = ~A168 & ~A170;
  assign \new_[14843]_  = ~A265 & A203;
  assign \new_[14844]_  = ~A201 & \new_[14843]_ ;
  assign \new_[14845]_  = \new_[14844]_  & \new_[14839]_ ;
  assign \new_[14848]_  = A267 & A266;
  assign \new_[14852]_  = A299 & A298;
  assign \new_[14853]_  = A269 & \new_[14852]_ ;
  assign \new_[14854]_  = \new_[14853]_  & \new_[14848]_ ;
  assign \new_[14857]_  = ~A168 & ~A170;
  assign \new_[14861]_  = ~A265 & A203;
  assign \new_[14862]_  = ~A201 & \new_[14861]_ ;
  assign \new_[14863]_  = \new_[14862]_  & \new_[14857]_ ;
  assign \new_[14866]_  = A267 & A266;
  assign \new_[14870]_  = ~A299 & ~A298;
  assign \new_[14871]_  = A269 & \new_[14870]_ ;
  assign \new_[14872]_  = \new_[14871]_  & \new_[14866]_ ;
  assign \new_[14875]_  = ~A168 & ~A170;
  assign \new_[14879]_  = A265 & A203;
  assign \new_[14880]_  = ~A201 & \new_[14879]_ ;
  assign \new_[14881]_  = \new_[14880]_  & \new_[14875]_ ;
  assign \new_[14884]_  = A267 & ~A266;
  assign \new_[14888]_  = A301 & ~A300;
  assign \new_[14889]_  = A268 & \new_[14888]_ ;
  assign \new_[14890]_  = \new_[14889]_  & \new_[14884]_ ;
  assign \new_[14893]_  = ~A168 & ~A170;
  assign \new_[14897]_  = A265 & A203;
  assign \new_[14898]_  = ~A201 & \new_[14897]_ ;
  assign \new_[14899]_  = \new_[14898]_  & \new_[14893]_ ;
  assign \new_[14902]_  = A267 & ~A266;
  assign \new_[14906]_  = A302 & ~A300;
  assign \new_[14907]_  = A268 & \new_[14906]_ ;
  assign \new_[14908]_  = \new_[14907]_  & \new_[14902]_ ;
  assign \new_[14911]_  = ~A168 & ~A170;
  assign \new_[14915]_  = A265 & A203;
  assign \new_[14916]_  = ~A201 & \new_[14915]_ ;
  assign \new_[14917]_  = \new_[14916]_  & \new_[14911]_ ;
  assign \new_[14920]_  = A267 & ~A266;
  assign \new_[14924]_  = A299 & A298;
  assign \new_[14925]_  = A268 & \new_[14924]_ ;
  assign \new_[14926]_  = \new_[14925]_  & \new_[14920]_ ;
  assign \new_[14929]_  = ~A168 & ~A170;
  assign \new_[14933]_  = A265 & A203;
  assign \new_[14934]_  = ~A201 & \new_[14933]_ ;
  assign \new_[14935]_  = \new_[14934]_  & \new_[14929]_ ;
  assign \new_[14938]_  = A267 & ~A266;
  assign \new_[14942]_  = ~A299 & ~A298;
  assign \new_[14943]_  = A268 & \new_[14942]_ ;
  assign \new_[14944]_  = \new_[14943]_  & \new_[14938]_ ;
  assign \new_[14947]_  = ~A168 & ~A170;
  assign \new_[14951]_  = A265 & A203;
  assign \new_[14952]_  = ~A201 & \new_[14951]_ ;
  assign \new_[14953]_  = \new_[14952]_  & \new_[14947]_ ;
  assign \new_[14956]_  = A267 & ~A266;
  assign \new_[14960]_  = A301 & ~A300;
  assign \new_[14961]_  = A269 & \new_[14960]_ ;
  assign \new_[14962]_  = \new_[14961]_  & \new_[14956]_ ;
  assign \new_[14965]_  = ~A168 & ~A170;
  assign \new_[14969]_  = A265 & A203;
  assign \new_[14970]_  = ~A201 & \new_[14969]_ ;
  assign \new_[14971]_  = \new_[14970]_  & \new_[14965]_ ;
  assign \new_[14974]_  = A267 & ~A266;
  assign \new_[14978]_  = A302 & ~A300;
  assign \new_[14979]_  = A269 & \new_[14978]_ ;
  assign \new_[14980]_  = \new_[14979]_  & \new_[14974]_ ;
  assign \new_[14983]_  = ~A168 & ~A170;
  assign \new_[14987]_  = A265 & A203;
  assign \new_[14988]_  = ~A201 & \new_[14987]_ ;
  assign \new_[14989]_  = \new_[14988]_  & \new_[14983]_ ;
  assign \new_[14992]_  = A267 & ~A266;
  assign \new_[14996]_  = A299 & A298;
  assign \new_[14997]_  = A269 & \new_[14996]_ ;
  assign \new_[14998]_  = \new_[14997]_  & \new_[14992]_ ;
  assign \new_[15001]_  = ~A168 & ~A170;
  assign \new_[15005]_  = A265 & A203;
  assign \new_[15006]_  = ~A201 & \new_[15005]_ ;
  assign \new_[15007]_  = \new_[15006]_  & \new_[15001]_ ;
  assign \new_[15010]_  = A267 & ~A266;
  assign \new_[15014]_  = ~A299 & ~A298;
  assign \new_[15015]_  = A269 & \new_[15014]_ ;
  assign \new_[15016]_  = \new_[15015]_  & \new_[15010]_ ;
  assign \new_[15019]_  = ~A168 & ~A170;
  assign \new_[15023]_  = ~A265 & A200;
  assign \new_[15024]_  = A199 & \new_[15023]_ ;
  assign \new_[15025]_  = \new_[15024]_  & \new_[15019]_ ;
  assign \new_[15028]_  = A267 & A266;
  assign \new_[15032]_  = A301 & ~A300;
  assign \new_[15033]_  = A268 & \new_[15032]_ ;
  assign \new_[15034]_  = \new_[15033]_  & \new_[15028]_ ;
  assign \new_[15037]_  = ~A168 & ~A170;
  assign \new_[15041]_  = ~A265 & A200;
  assign \new_[15042]_  = A199 & \new_[15041]_ ;
  assign \new_[15043]_  = \new_[15042]_  & \new_[15037]_ ;
  assign \new_[15046]_  = A267 & A266;
  assign \new_[15050]_  = A302 & ~A300;
  assign \new_[15051]_  = A268 & \new_[15050]_ ;
  assign \new_[15052]_  = \new_[15051]_  & \new_[15046]_ ;
  assign \new_[15055]_  = ~A168 & ~A170;
  assign \new_[15059]_  = ~A265 & A200;
  assign \new_[15060]_  = A199 & \new_[15059]_ ;
  assign \new_[15061]_  = \new_[15060]_  & \new_[15055]_ ;
  assign \new_[15064]_  = A267 & A266;
  assign \new_[15068]_  = A299 & A298;
  assign \new_[15069]_  = A268 & \new_[15068]_ ;
  assign \new_[15070]_  = \new_[15069]_  & \new_[15064]_ ;
  assign \new_[15073]_  = ~A168 & ~A170;
  assign \new_[15077]_  = ~A265 & A200;
  assign \new_[15078]_  = A199 & \new_[15077]_ ;
  assign \new_[15079]_  = \new_[15078]_  & \new_[15073]_ ;
  assign \new_[15082]_  = A267 & A266;
  assign \new_[15086]_  = ~A299 & ~A298;
  assign \new_[15087]_  = A268 & \new_[15086]_ ;
  assign \new_[15088]_  = \new_[15087]_  & \new_[15082]_ ;
  assign \new_[15091]_  = ~A168 & ~A170;
  assign \new_[15095]_  = ~A265 & A200;
  assign \new_[15096]_  = A199 & \new_[15095]_ ;
  assign \new_[15097]_  = \new_[15096]_  & \new_[15091]_ ;
  assign \new_[15100]_  = A267 & A266;
  assign \new_[15104]_  = A301 & ~A300;
  assign \new_[15105]_  = A269 & \new_[15104]_ ;
  assign \new_[15106]_  = \new_[15105]_  & \new_[15100]_ ;
  assign \new_[15109]_  = ~A168 & ~A170;
  assign \new_[15113]_  = ~A265 & A200;
  assign \new_[15114]_  = A199 & \new_[15113]_ ;
  assign \new_[15115]_  = \new_[15114]_  & \new_[15109]_ ;
  assign \new_[15118]_  = A267 & A266;
  assign \new_[15122]_  = A302 & ~A300;
  assign \new_[15123]_  = A269 & \new_[15122]_ ;
  assign \new_[15124]_  = \new_[15123]_  & \new_[15118]_ ;
  assign \new_[15127]_  = ~A168 & ~A170;
  assign \new_[15131]_  = ~A265 & A200;
  assign \new_[15132]_  = A199 & \new_[15131]_ ;
  assign \new_[15133]_  = \new_[15132]_  & \new_[15127]_ ;
  assign \new_[15136]_  = A267 & A266;
  assign \new_[15140]_  = A299 & A298;
  assign \new_[15141]_  = A269 & \new_[15140]_ ;
  assign \new_[15142]_  = \new_[15141]_  & \new_[15136]_ ;
  assign \new_[15145]_  = ~A168 & ~A170;
  assign \new_[15149]_  = ~A265 & A200;
  assign \new_[15150]_  = A199 & \new_[15149]_ ;
  assign \new_[15151]_  = \new_[15150]_  & \new_[15145]_ ;
  assign \new_[15154]_  = A267 & A266;
  assign \new_[15158]_  = ~A299 & ~A298;
  assign \new_[15159]_  = A269 & \new_[15158]_ ;
  assign \new_[15160]_  = \new_[15159]_  & \new_[15154]_ ;
  assign \new_[15163]_  = ~A168 & ~A170;
  assign \new_[15167]_  = A265 & A200;
  assign \new_[15168]_  = A199 & \new_[15167]_ ;
  assign \new_[15169]_  = \new_[15168]_  & \new_[15163]_ ;
  assign \new_[15172]_  = A267 & ~A266;
  assign \new_[15176]_  = A301 & ~A300;
  assign \new_[15177]_  = A268 & \new_[15176]_ ;
  assign \new_[15178]_  = \new_[15177]_  & \new_[15172]_ ;
  assign \new_[15181]_  = ~A168 & ~A170;
  assign \new_[15185]_  = A265 & A200;
  assign \new_[15186]_  = A199 & \new_[15185]_ ;
  assign \new_[15187]_  = \new_[15186]_  & \new_[15181]_ ;
  assign \new_[15190]_  = A267 & ~A266;
  assign \new_[15194]_  = A302 & ~A300;
  assign \new_[15195]_  = A268 & \new_[15194]_ ;
  assign \new_[15196]_  = \new_[15195]_  & \new_[15190]_ ;
  assign \new_[15199]_  = ~A168 & ~A170;
  assign \new_[15203]_  = A265 & A200;
  assign \new_[15204]_  = A199 & \new_[15203]_ ;
  assign \new_[15205]_  = \new_[15204]_  & \new_[15199]_ ;
  assign \new_[15208]_  = A267 & ~A266;
  assign \new_[15212]_  = A299 & A298;
  assign \new_[15213]_  = A268 & \new_[15212]_ ;
  assign \new_[15214]_  = \new_[15213]_  & \new_[15208]_ ;
  assign \new_[15217]_  = ~A168 & ~A170;
  assign \new_[15221]_  = A265 & A200;
  assign \new_[15222]_  = A199 & \new_[15221]_ ;
  assign \new_[15223]_  = \new_[15222]_  & \new_[15217]_ ;
  assign \new_[15226]_  = A267 & ~A266;
  assign \new_[15230]_  = ~A299 & ~A298;
  assign \new_[15231]_  = A268 & \new_[15230]_ ;
  assign \new_[15232]_  = \new_[15231]_  & \new_[15226]_ ;
  assign \new_[15235]_  = ~A168 & ~A170;
  assign \new_[15239]_  = A265 & A200;
  assign \new_[15240]_  = A199 & \new_[15239]_ ;
  assign \new_[15241]_  = \new_[15240]_  & \new_[15235]_ ;
  assign \new_[15244]_  = A267 & ~A266;
  assign \new_[15248]_  = A301 & ~A300;
  assign \new_[15249]_  = A269 & \new_[15248]_ ;
  assign \new_[15250]_  = \new_[15249]_  & \new_[15244]_ ;
  assign \new_[15253]_  = ~A168 & ~A170;
  assign \new_[15257]_  = A265 & A200;
  assign \new_[15258]_  = A199 & \new_[15257]_ ;
  assign \new_[15259]_  = \new_[15258]_  & \new_[15253]_ ;
  assign \new_[15262]_  = A267 & ~A266;
  assign \new_[15266]_  = A302 & ~A300;
  assign \new_[15267]_  = A269 & \new_[15266]_ ;
  assign \new_[15268]_  = \new_[15267]_  & \new_[15262]_ ;
  assign \new_[15271]_  = ~A168 & ~A170;
  assign \new_[15275]_  = A265 & A200;
  assign \new_[15276]_  = A199 & \new_[15275]_ ;
  assign \new_[15277]_  = \new_[15276]_  & \new_[15271]_ ;
  assign \new_[15280]_  = A267 & ~A266;
  assign \new_[15284]_  = A299 & A298;
  assign \new_[15285]_  = A269 & \new_[15284]_ ;
  assign \new_[15286]_  = \new_[15285]_  & \new_[15280]_ ;
  assign \new_[15289]_  = ~A168 & ~A170;
  assign \new_[15293]_  = A265 & A200;
  assign \new_[15294]_  = A199 & \new_[15293]_ ;
  assign \new_[15295]_  = \new_[15294]_  & \new_[15289]_ ;
  assign \new_[15298]_  = A267 & ~A266;
  assign \new_[15302]_  = ~A299 & ~A298;
  assign \new_[15303]_  = A269 & \new_[15302]_ ;
  assign \new_[15304]_  = \new_[15303]_  & \new_[15298]_ ;
  assign \new_[15307]_  = ~A168 & ~A170;
  assign \new_[15311]_  = ~A265 & ~A200;
  assign \new_[15312]_  = ~A199 & \new_[15311]_ ;
  assign \new_[15313]_  = \new_[15312]_  & \new_[15307]_ ;
  assign \new_[15316]_  = A267 & A266;
  assign \new_[15320]_  = A301 & ~A300;
  assign \new_[15321]_  = A268 & \new_[15320]_ ;
  assign \new_[15322]_  = \new_[15321]_  & \new_[15316]_ ;
  assign \new_[15325]_  = ~A168 & ~A170;
  assign \new_[15329]_  = ~A265 & ~A200;
  assign \new_[15330]_  = ~A199 & \new_[15329]_ ;
  assign \new_[15331]_  = \new_[15330]_  & \new_[15325]_ ;
  assign \new_[15334]_  = A267 & A266;
  assign \new_[15338]_  = A302 & ~A300;
  assign \new_[15339]_  = A268 & \new_[15338]_ ;
  assign \new_[15340]_  = \new_[15339]_  & \new_[15334]_ ;
  assign \new_[15343]_  = ~A168 & ~A170;
  assign \new_[15347]_  = ~A265 & ~A200;
  assign \new_[15348]_  = ~A199 & \new_[15347]_ ;
  assign \new_[15349]_  = \new_[15348]_  & \new_[15343]_ ;
  assign \new_[15352]_  = A267 & A266;
  assign \new_[15356]_  = A299 & A298;
  assign \new_[15357]_  = A268 & \new_[15356]_ ;
  assign \new_[15358]_  = \new_[15357]_  & \new_[15352]_ ;
  assign \new_[15361]_  = ~A168 & ~A170;
  assign \new_[15365]_  = ~A265 & ~A200;
  assign \new_[15366]_  = ~A199 & \new_[15365]_ ;
  assign \new_[15367]_  = \new_[15366]_  & \new_[15361]_ ;
  assign \new_[15370]_  = A267 & A266;
  assign \new_[15374]_  = ~A299 & ~A298;
  assign \new_[15375]_  = A268 & \new_[15374]_ ;
  assign \new_[15376]_  = \new_[15375]_  & \new_[15370]_ ;
  assign \new_[15379]_  = ~A168 & ~A170;
  assign \new_[15383]_  = ~A265 & ~A200;
  assign \new_[15384]_  = ~A199 & \new_[15383]_ ;
  assign \new_[15385]_  = \new_[15384]_  & \new_[15379]_ ;
  assign \new_[15388]_  = A267 & A266;
  assign \new_[15392]_  = A301 & ~A300;
  assign \new_[15393]_  = A269 & \new_[15392]_ ;
  assign \new_[15394]_  = \new_[15393]_  & \new_[15388]_ ;
  assign \new_[15397]_  = ~A168 & ~A170;
  assign \new_[15401]_  = ~A265 & ~A200;
  assign \new_[15402]_  = ~A199 & \new_[15401]_ ;
  assign \new_[15403]_  = \new_[15402]_  & \new_[15397]_ ;
  assign \new_[15406]_  = A267 & A266;
  assign \new_[15410]_  = A302 & ~A300;
  assign \new_[15411]_  = A269 & \new_[15410]_ ;
  assign \new_[15412]_  = \new_[15411]_  & \new_[15406]_ ;
  assign \new_[15415]_  = ~A168 & ~A170;
  assign \new_[15419]_  = ~A265 & ~A200;
  assign \new_[15420]_  = ~A199 & \new_[15419]_ ;
  assign \new_[15421]_  = \new_[15420]_  & \new_[15415]_ ;
  assign \new_[15424]_  = A267 & A266;
  assign \new_[15428]_  = A299 & A298;
  assign \new_[15429]_  = A269 & \new_[15428]_ ;
  assign \new_[15430]_  = \new_[15429]_  & \new_[15424]_ ;
  assign \new_[15433]_  = ~A168 & ~A170;
  assign \new_[15437]_  = ~A265 & ~A200;
  assign \new_[15438]_  = ~A199 & \new_[15437]_ ;
  assign \new_[15439]_  = \new_[15438]_  & \new_[15433]_ ;
  assign \new_[15442]_  = A267 & A266;
  assign \new_[15446]_  = ~A299 & ~A298;
  assign \new_[15447]_  = A269 & \new_[15446]_ ;
  assign \new_[15448]_  = \new_[15447]_  & \new_[15442]_ ;
  assign \new_[15451]_  = ~A168 & ~A170;
  assign \new_[15455]_  = A265 & ~A200;
  assign \new_[15456]_  = ~A199 & \new_[15455]_ ;
  assign \new_[15457]_  = \new_[15456]_  & \new_[15451]_ ;
  assign \new_[15460]_  = A267 & ~A266;
  assign \new_[15464]_  = A301 & ~A300;
  assign \new_[15465]_  = A268 & \new_[15464]_ ;
  assign \new_[15466]_  = \new_[15465]_  & \new_[15460]_ ;
  assign \new_[15469]_  = ~A168 & ~A170;
  assign \new_[15473]_  = A265 & ~A200;
  assign \new_[15474]_  = ~A199 & \new_[15473]_ ;
  assign \new_[15475]_  = \new_[15474]_  & \new_[15469]_ ;
  assign \new_[15478]_  = A267 & ~A266;
  assign \new_[15482]_  = A302 & ~A300;
  assign \new_[15483]_  = A268 & \new_[15482]_ ;
  assign \new_[15484]_  = \new_[15483]_  & \new_[15478]_ ;
  assign \new_[15487]_  = ~A168 & ~A170;
  assign \new_[15491]_  = A265 & ~A200;
  assign \new_[15492]_  = ~A199 & \new_[15491]_ ;
  assign \new_[15493]_  = \new_[15492]_  & \new_[15487]_ ;
  assign \new_[15496]_  = A267 & ~A266;
  assign \new_[15500]_  = A299 & A298;
  assign \new_[15501]_  = A268 & \new_[15500]_ ;
  assign \new_[15502]_  = \new_[15501]_  & \new_[15496]_ ;
  assign \new_[15505]_  = ~A168 & ~A170;
  assign \new_[15509]_  = A265 & ~A200;
  assign \new_[15510]_  = ~A199 & \new_[15509]_ ;
  assign \new_[15511]_  = \new_[15510]_  & \new_[15505]_ ;
  assign \new_[15514]_  = A267 & ~A266;
  assign \new_[15518]_  = ~A299 & ~A298;
  assign \new_[15519]_  = A268 & \new_[15518]_ ;
  assign \new_[15520]_  = \new_[15519]_  & \new_[15514]_ ;
  assign \new_[15523]_  = ~A168 & ~A170;
  assign \new_[15527]_  = A265 & ~A200;
  assign \new_[15528]_  = ~A199 & \new_[15527]_ ;
  assign \new_[15529]_  = \new_[15528]_  & \new_[15523]_ ;
  assign \new_[15532]_  = A267 & ~A266;
  assign \new_[15536]_  = A301 & ~A300;
  assign \new_[15537]_  = A269 & \new_[15536]_ ;
  assign \new_[15538]_  = \new_[15537]_  & \new_[15532]_ ;
  assign \new_[15541]_  = ~A168 & ~A170;
  assign \new_[15545]_  = A265 & ~A200;
  assign \new_[15546]_  = ~A199 & \new_[15545]_ ;
  assign \new_[15547]_  = \new_[15546]_  & \new_[15541]_ ;
  assign \new_[15550]_  = A267 & ~A266;
  assign \new_[15554]_  = A302 & ~A300;
  assign \new_[15555]_  = A269 & \new_[15554]_ ;
  assign \new_[15556]_  = \new_[15555]_  & \new_[15550]_ ;
  assign \new_[15559]_  = ~A168 & ~A170;
  assign \new_[15563]_  = A265 & ~A200;
  assign \new_[15564]_  = ~A199 & \new_[15563]_ ;
  assign \new_[15565]_  = \new_[15564]_  & \new_[15559]_ ;
  assign \new_[15568]_  = A267 & ~A266;
  assign \new_[15572]_  = A299 & A298;
  assign \new_[15573]_  = A269 & \new_[15572]_ ;
  assign \new_[15574]_  = \new_[15573]_  & \new_[15568]_ ;
  assign \new_[15577]_  = ~A168 & ~A170;
  assign \new_[15581]_  = A265 & ~A200;
  assign \new_[15582]_  = ~A199 & \new_[15581]_ ;
  assign \new_[15583]_  = \new_[15582]_  & \new_[15577]_ ;
  assign \new_[15586]_  = A267 & ~A266;
  assign \new_[15590]_  = ~A299 & ~A298;
  assign \new_[15591]_  = A269 & \new_[15590]_ ;
  assign \new_[15592]_  = \new_[15591]_  & \new_[15586]_ ;
  assign \new_[15595]_  = ~A168 & A169;
  assign \new_[15599]_  = ~A265 & A202;
  assign \new_[15600]_  = ~A201 & \new_[15599]_ ;
  assign \new_[15601]_  = \new_[15600]_  & \new_[15595]_ ;
  assign \new_[15604]_  = A267 & A266;
  assign \new_[15608]_  = A301 & ~A300;
  assign \new_[15609]_  = A268 & \new_[15608]_ ;
  assign \new_[15610]_  = \new_[15609]_  & \new_[15604]_ ;
  assign \new_[15613]_  = ~A168 & A169;
  assign \new_[15617]_  = ~A265 & A202;
  assign \new_[15618]_  = ~A201 & \new_[15617]_ ;
  assign \new_[15619]_  = \new_[15618]_  & \new_[15613]_ ;
  assign \new_[15622]_  = A267 & A266;
  assign \new_[15626]_  = A302 & ~A300;
  assign \new_[15627]_  = A268 & \new_[15626]_ ;
  assign \new_[15628]_  = \new_[15627]_  & \new_[15622]_ ;
  assign \new_[15631]_  = ~A168 & A169;
  assign \new_[15635]_  = ~A265 & A202;
  assign \new_[15636]_  = ~A201 & \new_[15635]_ ;
  assign \new_[15637]_  = \new_[15636]_  & \new_[15631]_ ;
  assign \new_[15640]_  = A267 & A266;
  assign \new_[15644]_  = A299 & A298;
  assign \new_[15645]_  = A268 & \new_[15644]_ ;
  assign \new_[15646]_  = \new_[15645]_  & \new_[15640]_ ;
  assign \new_[15649]_  = ~A168 & A169;
  assign \new_[15653]_  = ~A265 & A202;
  assign \new_[15654]_  = ~A201 & \new_[15653]_ ;
  assign \new_[15655]_  = \new_[15654]_  & \new_[15649]_ ;
  assign \new_[15658]_  = A267 & A266;
  assign \new_[15662]_  = ~A299 & ~A298;
  assign \new_[15663]_  = A268 & \new_[15662]_ ;
  assign \new_[15664]_  = \new_[15663]_  & \new_[15658]_ ;
  assign \new_[15667]_  = ~A168 & A169;
  assign \new_[15671]_  = ~A265 & A202;
  assign \new_[15672]_  = ~A201 & \new_[15671]_ ;
  assign \new_[15673]_  = \new_[15672]_  & \new_[15667]_ ;
  assign \new_[15676]_  = A267 & A266;
  assign \new_[15680]_  = A301 & ~A300;
  assign \new_[15681]_  = A269 & \new_[15680]_ ;
  assign \new_[15682]_  = \new_[15681]_  & \new_[15676]_ ;
  assign \new_[15685]_  = ~A168 & A169;
  assign \new_[15689]_  = ~A265 & A202;
  assign \new_[15690]_  = ~A201 & \new_[15689]_ ;
  assign \new_[15691]_  = \new_[15690]_  & \new_[15685]_ ;
  assign \new_[15694]_  = A267 & A266;
  assign \new_[15698]_  = A302 & ~A300;
  assign \new_[15699]_  = A269 & \new_[15698]_ ;
  assign \new_[15700]_  = \new_[15699]_  & \new_[15694]_ ;
  assign \new_[15703]_  = ~A168 & A169;
  assign \new_[15707]_  = ~A265 & A202;
  assign \new_[15708]_  = ~A201 & \new_[15707]_ ;
  assign \new_[15709]_  = \new_[15708]_  & \new_[15703]_ ;
  assign \new_[15712]_  = A267 & A266;
  assign \new_[15716]_  = A299 & A298;
  assign \new_[15717]_  = A269 & \new_[15716]_ ;
  assign \new_[15718]_  = \new_[15717]_  & \new_[15712]_ ;
  assign \new_[15721]_  = ~A168 & A169;
  assign \new_[15725]_  = ~A265 & A202;
  assign \new_[15726]_  = ~A201 & \new_[15725]_ ;
  assign \new_[15727]_  = \new_[15726]_  & \new_[15721]_ ;
  assign \new_[15730]_  = A267 & A266;
  assign \new_[15734]_  = ~A299 & ~A298;
  assign \new_[15735]_  = A269 & \new_[15734]_ ;
  assign \new_[15736]_  = \new_[15735]_  & \new_[15730]_ ;
  assign \new_[15739]_  = ~A168 & A169;
  assign \new_[15743]_  = A265 & A202;
  assign \new_[15744]_  = ~A201 & \new_[15743]_ ;
  assign \new_[15745]_  = \new_[15744]_  & \new_[15739]_ ;
  assign \new_[15748]_  = A267 & ~A266;
  assign \new_[15752]_  = A301 & ~A300;
  assign \new_[15753]_  = A268 & \new_[15752]_ ;
  assign \new_[15754]_  = \new_[15753]_  & \new_[15748]_ ;
  assign \new_[15757]_  = ~A168 & A169;
  assign \new_[15761]_  = A265 & A202;
  assign \new_[15762]_  = ~A201 & \new_[15761]_ ;
  assign \new_[15763]_  = \new_[15762]_  & \new_[15757]_ ;
  assign \new_[15766]_  = A267 & ~A266;
  assign \new_[15770]_  = A302 & ~A300;
  assign \new_[15771]_  = A268 & \new_[15770]_ ;
  assign \new_[15772]_  = \new_[15771]_  & \new_[15766]_ ;
  assign \new_[15775]_  = ~A168 & A169;
  assign \new_[15779]_  = A265 & A202;
  assign \new_[15780]_  = ~A201 & \new_[15779]_ ;
  assign \new_[15781]_  = \new_[15780]_  & \new_[15775]_ ;
  assign \new_[15784]_  = A267 & ~A266;
  assign \new_[15788]_  = A299 & A298;
  assign \new_[15789]_  = A268 & \new_[15788]_ ;
  assign \new_[15790]_  = \new_[15789]_  & \new_[15784]_ ;
  assign \new_[15793]_  = ~A168 & A169;
  assign \new_[15797]_  = A265 & A202;
  assign \new_[15798]_  = ~A201 & \new_[15797]_ ;
  assign \new_[15799]_  = \new_[15798]_  & \new_[15793]_ ;
  assign \new_[15802]_  = A267 & ~A266;
  assign \new_[15806]_  = ~A299 & ~A298;
  assign \new_[15807]_  = A268 & \new_[15806]_ ;
  assign \new_[15808]_  = \new_[15807]_  & \new_[15802]_ ;
  assign \new_[15811]_  = ~A168 & A169;
  assign \new_[15815]_  = A265 & A202;
  assign \new_[15816]_  = ~A201 & \new_[15815]_ ;
  assign \new_[15817]_  = \new_[15816]_  & \new_[15811]_ ;
  assign \new_[15820]_  = A267 & ~A266;
  assign \new_[15824]_  = A301 & ~A300;
  assign \new_[15825]_  = A269 & \new_[15824]_ ;
  assign \new_[15826]_  = \new_[15825]_  & \new_[15820]_ ;
  assign \new_[15829]_  = ~A168 & A169;
  assign \new_[15833]_  = A265 & A202;
  assign \new_[15834]_  = ~A201 & \new_[15833]_ ;
  assign \new_[15835]_  = \new_[15834]_  & \new_[15829]_ ;
  assign \new_[15838]_  = A267 & ~A266;
  assign \new_[15842]_  = A302 & ~A300;
  assign \new_[15843]_  = A269 & \new_[15842]_ ;
  assign \new_[15844]_  = \new_[15843]_  & \new_[15838]_ ;
  assign \new_[15847]_  = ~A168 & A169;
  assign \new_[15851]_  = A265 & A202;
  assign \new_[15852]_  = ~A201 & \new_[15851]_ ;
  assign \new_[15853]_  = \new_[15852]_  & \new_[15847]_ ;
  assign \new_[15856]_  = A267 & ~A266;
  assign \new_[15860]_  = A299 & A298;
  assign \new_[15861]_  = A269 & \new_[15860]_ ;
  assign \new_[15862]_  = \new_[15861]_  & \new_[15856]_ ;
  assign \new_[15865]_  = ~A168 & A169;
  assign \new_[15869]_  = A265 & A202;
  assign \new_[15870]_  = ~A201 & \new_[15869]_ ;
  assign \new_[15871]_  = \new_[15870]_  & \new_[15865]_ ;
  assign \new_[15874]_  = A267 & ~A266;
  assign \new_[15878]_  = ~A299 & ~A298;
  assign \new_[15879]_  = A269 & \new_[15878]_ ;
  assign \new_[15880]_  = \new_[15879]_  & \new_[15874]_ ;
  assign \new_[15883]_  = ~A168 & A169;
  assign \new_[15887]_  = ~A265 & A203;
  assign \new_[15888]_  = ~A201 & \new_[15887]_ ;
  assign \new_[15889]_  = \new_[15888]_  & \new_[15883]_ ;
  assign \new_[15892]_  = A267 & A266;
  assign \new_[15896]_  = A301 & ~A300;
  assign \new_[15897]_  = A268 & \new_[15896]_ ;
  assign \new_[15898]_  = \new_[15897]_  & \new_[15892]_ ;
  assign \new_[15901]_  = ~A168 & A169;
  assign \new_[15905]_  = ~A265 & A203;
  assign \new_[15906]_  = ~A201 & \new_[15905]_ ;
  assign \new_[15907]_  = \new_[15906]_  & \new_[15901]_ ;
  assign \new_[15910]_  = A267 & A266;
  assign \new_[15914]_  = A302 & ~A300;
  assign \new_[15915]_  = A268 & \new_[15914]_ ;
  assign \new_[15916]_  = \new_[15915]_  & \new_[15910]_ ;
  assign \new_[15919]_  = ~A168 & A169;
  assign \new_[15923]_  = ~A265 & A203;
  assign \new_[15924]_  = ~A201 & \new_[15923]_ ;
  assign \new_[15925]_  = \new_[15924]_  & \new_[15919]_ ;
  assign \new_[15928]_  = A267 & A266;
  assign \new_[15932]_  = A299 & A298;
  assign \new_[15933]_  = A268 & \new_[15932]_ ;
  assign \new_[15934]_  = \new_[15933]_  & \new_[15928]_ ;
  assign \new_[15937]_  = ~A168 & A169;
  assign \new_[15941]_  = ~A265 & A203;
  assign \new_[15942]_  = ~A201 & \new_[15941]_ ;
  assign \new_[15943]_  = \new_[15942]_  & \new_[15937]_ ;
  assign \new_[15946]_  = A267 & A266;
  assign \new_[15950]_  = ~A299 & ~A298;
  assign \new_[15951]_  = A268 & \new_[15950]_ ;
  assign \new_[15952]_  = \new_[15951]_  & \new_[15946]_ ;
  assign \new_[15955]_  = ~A168 & A169;
  assign \new_[15959]_  = ~A265 & A203;
  assign \new_[15960]_  = ~A201 & \new_[15959]_ ;
  assign \new_[15961]_  = \new_[15960]_  & \new_[15955]_ ;
  assign \new_[15964]_  = A267 & A266;
  assign \new_[15968]_  = A301 & ~A300;
  assign \new_[15969]_  = A269 & \new_[15968]_ ;
  assign \new_[15970]_  = \new_[15969]_  & \new_[15964]_ ;
  assign \new_[15973]_  = ~A168 & A169;
  assign \new_[15977]_  = ~A265 & A203;
  assign \new_[15978]_  = ~A201 & \new_[15977]_ ;
  assign \new_[15979]_  = \new_[15978]_  & \new_[15973]_ ;
  assign \new_[15982]_  = A267 & A266;
  assign \new_[15986]_  = A302 & ~A300;
  assign \new_[15987]_  = A269 & \new_[15986]_ ;
  assign \new_[15988]_  = \new_[15987]_  & \new_[15982]_ ;
  assign \new_[15991]_  = ~A168 & A169;
  assign \new_[15995]_  = ~A265 & A203;
  assign \new_[15996]_  = ~A201 & \new_[15995]_ ;
  assign \new_[15997]_  = \new_[15996]_  & \new_[15991]_ ;
  assign \new_[16000]_  = A267 & A266;
  assign \new_[16004]_  = A299 & A298;
  assign \new_[16005]_  = A269 & \new_[16004]_ ;
  assign \new_[16006]_  = \new_[16005]_  & \new_[16000]_ ;
  assign \new_[16009]_  = ~A168 & A169;
  assign \new_[16013]_  = ~A265 & A203;
  assign \new_[16014]_  = ~A201 & \new_[16013]_ ;
  assign \new_[16015]_  = \new_[16014]_  & \new_[16009]_ ;
  assign \new_[16018]_  = A267 & A266;
  assign \new_[16022]_  = ~A299 & ~A298;
  assign \new_[16023]_  = A269 & \new_[16022]_ ;
  assign \new_[16024]_  = \new_[16023]_  & \new_[16018]_ ;
  assign \new_[16027]_  = ~A168 & A169;
  assign \new_[16031]_  = A265 & A203;
  assign \new_[16032]_  = ~A201 & \new_[16031]_ ;
  assign \new_[16033]_  = \new_[16032]_  & \new_[16027]_ ;
  assign \new_[16036]_  = A267 & ~A266;
  assign \new_[16040]_  = A301 & ~A300;
  assign \new_[16041]_  = A268 & \new_[16040]_ ;
  assign \new_[16042]_  = \new_[16041]_  & \new_[16036]_ ;
  assign \new_[16045]_  = ~A168 & A169;
  assign \new_[16049]_  = A265 & A203;
  assign \new_[16050]_  = ~A201 & \new_[16049]_ ;
  assign \new_[16051]_  = \new_[16050]_  & \new_[16045]_ ;
  assign \new_[16054]_  = A267 & ~A266;
  assign \new_[16058]_  = A302 & ~A300;
  assign \new_[16059]_  = A268 & \new_[16058]_ ;
  assign \new_[16060]_  = \new_[16059]_  & \new_[16054]_ ;
  assign \new_[16063]_  = ~A168 & A169;
  assign \new_[16067]_  = A265 & A203;
  assign \new_[16068]_  = ~A201 & \new_[16067]_ ;
  assign \new_[16069]_  = \new_[16068]_  & \new_[16063]_ ;
  assign \new_[16072]_  = A267 & ~A266;
  assign \new_[16076]_  = A299 & A298;
  assign \new_[16077]_  = A268 & \new_[16076]_ ;
  assign \new_[16078]_  = \new_[16077]_  & \new_[16072]_ ;
  assign \new_[16081]_  = ~A168 & A169;
  assign \new_[16085]_  = A265 & A203;
  assign \new_[16086]_  = ~A201 & \new_[16085]_ ;
  assign \new_[16087]_  = \new_[16086]_  & \new_[16081]_ ;
  assign \new_[16090]_  = A267 & ~A266;
  assign \new_[16094]_  = ~A299 & ~A298;
  assign \new_[16095]_  = A268 & \new_[16094]_ ;
  assign \new_[16096]_  = \new_[16095]_  & \new_[16090]_ ;
  assign \new_[16099]_  = ~A168 & A169;
  assign \new_[16103]_  = A265 & A203;
  assign \new_[16104]_  = ~A201 & \new_[16103]_ ;
  assign \new_[16105]_  = \new_[16104]_  & \new_[16099]_ ;
  assign \new_[16108]_  = A267 & ~A266;
  assign \new_[16112]_  = A301 & ~A300;
  assign \new_[16113]_  = A269 & \new_[16112]_ ;
  assign \new_[16114]_  = \new_[16113]_  & \new_[16108]_ ;
  assign \new_[16117]_  = ~A168 & A169;
  assign \new_[16121]_  = A265 & A203;
  assign \new_[16122]_  = ~A201 & \new_[16121]_ ;
  assign \new_[16123]_  = \new_[16122]_  & \new_[16117]_ ;
  assign \new_[16126]_  = A267 & ~A266;
  assign \new_[16130]_  = A302 & ~A300;
  assign \new_[16131]_  = A269 & \new_[16130]_ ;
  assign \new_[16132]_  = \new_[16131]_  & \new_[16126]_ ;
  assign \new_[16135]_  = ~A168 & A169;
  assign \new_[16139]_  = A265 & A203;
  assign \new_[16140]_  = ~A201 & \new_[16139]_ ;
  assign \new_[16141]_  = \new_[16140]_  & \new_[16135]_ ;
  assign \new_[16144]_  = A267 & ~A266;
  assign \new_[16148]_  = A299 & A298;
  assign \new_[16149]_  = A269 & \new_[16148]_ ;
  assign \new_[16150]_  = \new_[16149]_  & \new_[16144]_ ;
  assign \new_[16153]_  = ~A168 & A169;
  assign \new_[16157]_  = A265 & A203;
  assign \new_[16158]_  = ~A201 & \new_[16157]_ ;
  assign \new_[16159]_  = \new_[16158]_  & \new_[16153]_ ;
  assign \new_[16162]_  = A267 & ~A266;
  assign \new_[16166]_  = ~A299 & ~A298;
  assign \new_[16167]_  = A269 & \new_[16166]_ ;
  assign \new_[16168]_  = \new_[16167]_  & \new_[16162]_ ;
  assign \new_[16171]_  = ~A168 & A169;
  assign \new_[16175]_  = ~A265 & A200;
  assign \new_[16176]_  = A199 & \new_[16175]_ ;
  assign \new_[16177]_  = \new_[16176]_  & \new_[16171]_ ;
  assign \new_[16180]_  = A267 & A266;
  assign \new_[16184]_  = A301 & ~A300;
  assign \new_[16185]_  = A268 & \new_[16184]_ ;
  assign \new_[16186]_  = \new_[16185]_  & \new_[16180]_ ;
  assign \new_[16189]_  = ~A168 & A169;
  assign \new_[16193]_  = ~A265 & A200;
  assign \new_[16194]_  = A199 & \new_[16193]_ ;
  assign \new_[16195]_  = \new_[16194]_  & \new_[16189]_ ;
  assign \new_[16198]_  = A267 & A266;
  assign \new_[16202]_  = A302 & ~A300;
  assign \new_[16203]_  = A268 & \new_[16202]_ ;
  assign \new_[16204]_  = \new_[16203]_  & \new_[16198]_ ;
  assign \new_[16207]_  = ~A168 & A169;
  assign \new_[16211]_  = ~A265 & A200;
  assign \new_[16212]_  = A199 & \new_[16211]_ ;
  assign \new_[16213]_  = \new_[16212]_  & \new_[16207]_ ;
  assign \new_[16216]_  = A267 & A266;
  assign \new_[16220]_  = A299 & A298;
  assign \new_[16221]_  = A268 & \new_[16220]_ ;
  assign \new_[16222]_  = \new_[16221]_  & \new_[16216]_ ;
  assign \new_[16225]_  = ~A168 & A169;
  assign \new_[16229]_  = ~A265 & A200;
  assign \new_[16230]_  = A199 & \new_[16229]_ ;
  assign \new_[16231]_  = \new_[16230]_  & \new_[16225]_ ;
  assign \new_[16234]_  = A267 & A266;
  assign \new_[16238]_  = ~A299 & ~A298;
  assign \new_[16239]_  = A268 & \new_[16238]_ ;
  assign \new_[16240]_  = \new_[16239]_  & \new_[16234]_ ;
  assign \new_[16243]_  = ~A168 & A169;
  assign \new_[16247]_  = ~A265 & A200;
  assign \new_[16248]_  = A199 & \new_[16247]_ ;
  assign \new_[16249]_  = \new_[16248]_  & \new_[16243]_ ;
  assign \new_[16252]_  = A267 & A266;
  assign \new_[16256]_  = A301 & ~A300;
  assign \new_[16257]_  = A269 & \new_[16256]_ ;
  assign \new_[16258]_  = \new_[16257]_  & \new_[16252]_ ;
  assign \new_[16261]_  = ~A168 & A169;
  assign \new_[16265]_  = ~A265 & A200;
  assign \new_[16266]_  = A199 & \new_[16265]_ ;
  assign \new_[16267]_  = \new_[16266]_  & \new_[16261]_ ;
  assign \new_[16270]_  = A267 & A266;
  assign \new_[16274]_  = A302 & ~A300;
  assign \new_[16275]_  = A269 & \new_[16274]_ ;
  assign \new_[16276]_  = \new_[16275]_  & \new_[16270]_ ;
  assign \new_[16279]_  = ~A168 & A169;
  assign \new_[16283]_  = ~A265 & A200;
  assign \new_[16284]_  = A199 & \new_[16283]_ ;
  assign \new_[16285]_  = \new_[16284]_  & \new_[16279]_ ;
  assign \new_[16288]_  = A267 & A266;
  assign \new_[16292]_  = A299 & A298;
  assign \new_[16293]_  = A269 & \new_[16292]_ ;
  assign \new_[16294]_  = \new_[16293]_  & \new_[16288]_ ;
  assign \new_[16297]_  = ~A168 & A169;
  assign \new_[16301]_  = ~A265 & A200;
  assign \new_[16302]_  = A199 & \new_[16301]_ ;
  assign \new_[16303]_  = \new_[16302]_  & \new_[16297]_ ;
  assign \new_[16306]_  = A267 & A266;
  assign \new_[16310]_  = ~A299 & ~A298;
  assign \new_[16311]_  = A269 & \new_[16310]_ ;
  assign \new_[16312]_  = \new_[16311]_  & \new_[16306]_ ;
  assign \new_[16315]_  = ~A168 & A169;
  assign \new_[16319]_  = A265 & A200;
  assign \new_[16320]_  = A199 & \new_[16319]_ ;
  assign \new_[16321]_  = \new_[16320]_  & \new_[16315]_ ;
  assign \new_[16324]_  = A267 & ~A266;
  assign \new_[16328]_  = A301 & ~A300;
  assign \new_[16329]_  = A268 & \new_[16328]_ ;
  assign \new_[16330]_  = \new_[16329]_  & \new_[16324]_ ;
  assign \new_[16333]_  = ~A168 & A169;
  assign \new_[16337]_  = A265 & A200;
  assign \new_[16338]_  = A199 & \new_[16337]_ ;
  assign \new_[16339]_  = \new_[16338]_  & \new_[16333]_ ;
  assign \new_[16342]_  = A267 & ~A266;
  assign \new_[16346]_  = A302 & ~A300;
  assign \new_[16347]_  = A268 & \new_[16346]_ ;
  assign \new_[16348]_  = \new_[16347]_  & \new_[16342]_ ;
  assign \new_[16351]_  = ~A168 & A169;
  assign \new_[16355]_  = A265 & A200;
  assign \new_[16356]_  = A199 & \new_[16355]_ ;
  assign \new_[16357]_  = \new_[16356]_  & \new_[16351]_ ;
  assign \new_[16360]_  = A267 & ~A266;
  assign \new_[16364]_  = A299 & A298;
  assign \new_[16365]_  = A268 & \new_[16364]_ ;
  assign \new_[16366]_  = \new_[16365]_  & \new_[16360]_ ;
  assign \new_[16369]_  = ~A168 & A169;
  assign \new_[16373]_  = A265 & A200;
  assign \new_[16374]_  = A199 & \new_[16373]_ ;
  assign \new_[16375]_  = \new_[16374]_  & \new_[16369]_ ;
  assign \new_[16378]_  = A267 & ~A266;
  assign \new_[16382]_  = ~A299 & ~A298;
  assign \new_[16383]_  = A268 & \new_[16382]_ ;
  assign \new_[16384]_  = \new_[16383]_  & \new_[16378]_ ;
  assign \new_[16387]_  = ~A168 & A169;
  assign \new_[16391]_  = A265 & A200;
  assign \new_[16392]_  = A199 & \new_[16391]_ ;
  assign \new_[16393]_  = \new_[16392]_  & \new_[16387]_ ;
  assign \new_[16396]_  = A267 & ~A266;
  assign \new_[16400]_  = A301 & ~A300;
  assign \new_[16401]_  = A269 & \new_[16400]_ ;
  assign \new_[16402]_  = \new_[16401]_  & \new_[16396]_ ;
  assign \new_[16405]_  = ~A168 & A169;
  assign \new_[16409]_  = A265 & A200;
  assign \new_[16410]_  = A199 & \new_[16409]_ ;
  assign \new_[16411]_  = \new_[16410]_  & \new_[16405]_ ;
  assign \new_[16414]_  = A267 & ~A266;
  assign \new_[16418]_  = A302 & ~A300;
  assign \new_[16419]_  = A269 & \new_[16418]_ ;
  assign \new_[16420]_  = \new_[16419]_  & \new_[16414]_ ;
  assign \new_[16423]_  = ~A168 & A169;
  assign \new_[16427]_  = A265 & A200;
  assign \new_[16428]_  = A199 & \new_[16427]_ ;
  assign \new_[16429]_  = \new_[16428]_  & \new_[16423]_ ;
  assign \new_[16432]_  = A267 & ~A266;
  assign \new_[16436]_  = A299 & A298;
  assign \new_[16437]_  = A269 & \new_[16436]_ ;
  assign \new_[16438]_  = \new_[16437]_  & \new_[16432]_ ;
  assign \new_[16441]_  = ~A168 & A169;
  assign \new_[16445]_  = A265 & A200;
  assign \new_[16446]_  = A199 & \new_[16445]_ ;
  assign \new_[16447]_  = \new_[16446]_  & \new_[16441]_ ;
  assign \new_[16450]_  = A267 & ~A266;
  assign \new_[16454]_  = ~A299 & ~A298;
  assign \new_[16455]_  = A269 & \new_[16454]_ ;
  assign \new_[16456]_  = \new_[16455]_  & \new_[16450]_ ;
  assign \new_[16459]_  = ~A168 & A169;
  assign \new_[16463]_  = ~A265 & ~A200;
  assign \new_[16464]_  = ~A199 & \new_[16463]_ ;
  assign \new_[16465]_  = \new_[16464]_  & \new_[16459]_ ;
  assign \new_[16468]_  = A267 & A266;
  assign \new_[16472]_  = A301 & ~A300;
  assign \new_[16473]_  = A268 & \new_[16472]_ ;
  assign \new_[16474]_  = \new_[16473]_  & \new_[16468]_ ;
  assign \new_[16477]_  = ~A168 & A169;
  assign \new_[16481]_  = ~A265 & ~A200;
  assign \new_[16482]_  = ~A199 & \new_[16481]_ ;
  assign \new_[16483]_  = \new_[16482]_  & \new_[16477]_ ;
  assign \new_[16486]_  = A267 & A266;
  assign \new_[16490]_  = A302 & ~A300;
  assign \new_[16491]_  = A268 & \new_[16490]_ ;
  assign \new_[16492]_  = \new_[16491]_  & \new_[16486]_ ;
  assign \new_[16495]_  = ~A168 & A169;
  assign \new_[16499]_  = ~A265 & ~A200;
  assign \new_[16500]_  = ~A199 & \new_[16499]_ ;
  assign \new_[16501]_  = \new_[16500]_  & \new_[16495]_ ;
  assign \new_[16504]_  = A267 & A266;
  assign \new_[16508]_  = A299 & A298;
  assign \new_[16509]_  = A268 & \new_[16508]_ ;
  assign \new_[16510]_  = \new_[16509]_  & \new_[16504]_ ;
  assign \new_[16513]_  = ~A168 & A169;
  assign \new_[16517]_  = ~A265 & ~A200;
  assign \new_[16518]_  = ~A199 & \new_[16517]_ ;
  assign \new_[16519]_  = \new_[16518]_  & \new_[16513]_ ;
  assign \new_[16522]_  = A267 & A266;
  assign \new_[16526]_  = ~A299 & ~A298;
  assign \new_[16527]_  = A268 & \new_[16526]_ ;
  assign \new_[16528]_  = \new_[16527]_  & \new_[16522]_ ;
  assign \new_[16531]_  = ~A168 & A169;
  assign \new_[16535]_  = ~A265 & ~A200;
  assign \new_[16536]_  = ~A199 & \new_[16535]_ ;
  assign \new_[16537]_  = \new_[16536]_  & \new_[16531]_ ;
  assign \new_[16540]_  = A267 & A266;
  assign \new_[16544]_  = A301 & ~A300;
  assign \new_[16545]_  = A269 & \new_[16544]_ ;
  assign \new_[16546]_  = \new_[16545]_  & \new_[16540]_ ;
  assign \new_[16549]_  = ~A168 & A169;
  assign \new_[16553]_  = ~A265 & ~A200;
  assign \new_[16554]_  = ~A199 & \new_[16553]_ ;
  assign \new_[16555]_  = \new_[16554]_  & \new_[16549]_ ;
  assign \new_[16558]_  = A267 & A266;
  assign \new_[16562]_  = A302 & ~A300;
  assign \new_[16563]_  = A269 & \new_[16562]_ ;
  assign \new_[16564]_  = \new_[16563]_  & \new_[16558]_ ;
  assign \new_[16567]_  = ~A168 & A169;
  assign \new_[16571]_  = ~A265 & ~A200;
  assign \new_[16572]_  = ~A199 & \new_[16571]_ ;
  assign \new_[16573]_  = \new_[16572]_  & \new_[16567]_ ;
  assign \new_[16576]_  = A267 & A266;
  assign \new_[16580]_  = A299 & A298;
  assign \new_[16581]_  = A269 & \new_[16580]_ ;
  assign \new_[16582]_  = \new_[16581]_  & \new_[16576]_ ;
  assign \new_[16585]_  = ~A168 & A169;
  assign \new_[16589]_  = ~A265 & ~A200;
  assign \new_[16590]_  = ~A199 & \new_[16589]_ ;
  assign \new_[16591]_  = \new_[16590]_  & \new_[16585]_ ;
  assign \new_[16594]_  = A267 & A266;
  assign \new_[16598]_  = ~A299 & ~A298;
  assign \new_[16599]_  = A269 & \new_[16598]_ ;
  assign \new_[16600]_  = \new_[16599]_  & \new_[16594]_ ;
  assign \new_[16603]_  = ~A168 & A169;
  assign \new_[16607]_  = A265 & ~A200;
  assign \new_[16608]_  = ~A199 & \new_[16607]_ ;
  assign \new_[16609]_  = \new_[16608]_  & \new_[16603]_ ;
  assign \new_[16612]_  = A267 & ~A266;
  assign \new_[16616]_  = A301 & ~A300;
  assign \new_[16617]_  = A268 & \new_[16616]_ ;
  assign \new_[16618]_  = \new_[16617]_  & \new_[16612]_ ;
  assign \new_[16621]_  = ~A168 & A169;
  assign \new_[16625]_  = A265 & ~A200;
  assign \new_[16626]_  = ~A199 & \new_[16625]_ ;
  assign \new_[16627]_  = \new_[16626]_  & \new_[16621]_ ;
  assign \new_[16630]_  = A267 & ~A266;
  assign \new_[16634]_  = A302 & ~A300;
  assign \new_[16635]_  = A268 & \new_[16634]_ ;
  assign \new_[16636]_  = \new_[16635]_  & \new_[16630]_ ;
  assign \new_[16639]_  = ~A168 & A169;
  assign \new_[16643]_  = A265 & ~A200;
  assign \new_[16644]_  = ~A199 & \new_[16643]_ ;
  assign \new_[16645]_  = \new_[16644]_  & \new_[16639]_ ;
  assign \new_[16648]_  = A267 & ~A266;
  assign \new_[16652]_  = A299 & A298;
  assign \new_[16653]_  = A268 & \new_[16652]_ ;
  assign \new_[16654]_  = \new_[16653]_  & \new_[16648]_ ;
  assign \new_[16657]_  = ~A168 & A169;
  assign \new_[16661]_  = A265 & ~A200;
  assign \new_[16662]_  = ~A199 & \new_[16661]_ ;
  assign \new_[16663]_  = \new_[16662]_  & \new_[16657]_ ;
  assign \new_[16666]_  = A267 & ~A266;
  assign \new_[16670]_  = ~A299 & ~A298;
  assign \new_[16671]_  = A268 & \new_[16670]_ ;
  assign \new_[16672]_  = \new_[16671]_  & \new_[16666]_ ;
  assign \new_[16675]_  = ~A168 & A169;
  assign \new_[16679]_  = A265 & ~A200;
  assign \new_[16680]_  = ~A199 & \new_[16679]_ ;
  assign \new_[16681]_  = \new_[16680]_  & \new_[16675]_ ;
  assign \new_[16684]_  = A267 & ~A266;
  assign \new_[16688]_  = A301 & ~A300;
  assign \new_[16689]_  = A269 & \new_[16688]_ ;
  assign \new_[16690]_  = \new_[16689]_  & \new_[16684]_ ;
  assign \new_[16693]_  = ~A168 & A169;
  assign \new_[16697]_  = A265 & ~A200;
  assign \new_[16698]_  = ~A199 & \new_[16697]_ ;
  assign \new_[16699]_  = \new_[16698]_  & \new_[16693]_ ;
  assign \new_[16702]_  = A267 & ~A266;
  assign \new_[16706]_  = A302 & ~A300;
  assign \new_[16707]_  = A269 & \new_[16706]_ ;
  assign \new_[16708]_  = \new_[16707]_  & \new_[16702]_ ;
  assign \new_[16711]_  = ~A168 & A169;
  assign \new_[16715]_  = A265 & ~A200;
  assign \new_[16716]_  = ~A199 & \new_[16715]_ ;
  assign \new_[16717]_  = \new_[16716]_  & \new_[16711]_ ;
  assign \new_[16720]_  = A267 & ~A266;
  assign \new_[16724]_  = A299 & A298;
  assign \new_[16725]_  = A269 & \new_[16724]_ ;
  assign \new_[16726]_  = \new_[16725]_  & \new_[16720]_ ;
  assign \new_[16729]_  = ~A168 & A169;
  assign \new_[16733]_  = A265 & ~A200;
  assign \new_[16734]_  = ~A199 & \new_[16733]_ ;
  assign \new_[16735]_  = \new_[16734]_  & \new_[16729]_ ;
  assign \new_[16738]_  = A267 & ~A266;
  assign \new_[16742]_  = ~A299 & ~A298;
  assign \new_[16743]_  = A269 & \new_[16742]_ ;
  assign \new_[16744]_  = \new_[16743]_  & \new_[16738]_ ;
  assign \new_[16747]_  = ~A169 & A170;
  assign \new_[16751]_  = ~A166 & A167;
  assign \new_[16752]_  = ~A168 & \new_[16751]_ ;
  assign \new_[16753]_  = \new_[16752]_  & \new_[16747]_ ;
  assign \new_[16756]_  = A233 & ~A232;
  assign \new_[16760]_  = ~A236 & ~A235;
  assign \new_[16761]_  = ~A234 & \new_[16760]_ ;
  assign \new_[16762]_  = \new_[16761]_  & \new_[16756]_ ;
  assign \new_[16765]_  = ~A169 & A170;
  assign \new_[16769]_  = ~A166 & A167;
  assign \new_[16770]_  = ~A168 & \new_[16769]_ ;
  assign \new_[16771]_  = \new_[16770]_  & \new_[16765]_ ;
  assign \new_[16774]_  = ~A233 & A232;
  assign \new_[16778]_  = ~A236 & ~A235;
  assign \new_[16779]_  = ~A234 & \new_[16778]_ ;
  assign \new_[16780]_  = \new_[16779]_  & \new_[16774]_ ;
  assign \new_[16783]_  = ~A169 & A170;
  assign \new_[16787]_  = A166 & ~A167;
  assign \new_[16788]_  = ~A168 & \new_[16787]_ ;
  assign \new_[16789]_  = \new_[16788]_  & \new_[16783]_ ;
  assign \new_[16792]_  = A233 & ~A232;
  assign \new_[16796]_  = ~A236 & ~A235;
  assign \new_[16797]_  = ~A234 & \new_[16796]_ ;
  assign \new_[16798]_  = \new_[16797]_  & \new_[16792]_ ;
  assign \new_[16801]_  = ~A169 & A170;
  assign \new_[16805]_  = A166 & ~A167;
  assign \new_[16806]_  = ~A168 & \new_[16805]_ ;
  assign \new_[16807]_  = \new_[16806]_  & \new_[16801]_ ;
  assign \new_[16810]_  = ~A233 & A232;
  assign \new_[16814]_  = ~A236 & ~A235;
  assign \new_[16815]_  = ~A234 & \new_[16814]_ ;
  assign \new_[16816]_  = \new_[16815]_  & \new_[16810]_ ;
  assign \new_[16819]_  = A166 & A167;
  assign \new_[16823]_  = ~A203 & ~A202;
  assign \new_[16824]_  = A201 & \new_[16823]_ ;
  assign \new_[16825]_  = \new_[16824]_  & \new_[16819]_ ;
  assign \new_[16829]_  = A267 & A266;
  assign \new_[16830]_  = ~A265 & \new_[16829]_ ;
  assign \new_[16834]_  = A301 & ~A300;
  assign \new_[16835]_  = A268 & \new_[16834]_ ;
  assign \new_[16836]_  = \new_[16835]_  & \new_[16830]_ ;
  assign \new_[16839]_  = A166 & A167;
  assign \new_[16843]_  = ~A203 & ~A202;
  assign \new_[16844]_  = A201 & \new_[16843]_ ;
  assign \new_[16845]_  = \new_[16844]_  & \new_[16839]_ ;
  assign \new_[16849]_  = A267 & A266;
  assign \new_[16850]_  = ~A265 & \new_[16849]_ ;
  assign \new_[16854]_  = A302 & ~A300;
  assign \new_[16855]_  = A268 & \new_[16854]_ ;
  assign \new_[16856]_  = \new_[16855]_  & \new_[16850]_ ;
  assign \new_[16859]_  = A166 & A167;
  assign \new_[16863]_  = ~A203 & ~A202;
  assign \new_[16864]_  = A201 & \new_[16863]_ ;
  assign \new_[16865]_  = \new_[16864]_  & \new_[16859]_ ;
  assign \new_[16869]_  = A267 & A266;
  assign \new_[16870]_  = ~A265 & \new_[16869]_ ;
  assign \new_[16874]_  = A299 & A298;
  assign \new_[16875]_  = A268 & \new_[16874]_ ;
  assign \new_[16876]_  = \new_[16875]_  & \new_[16870]_ ;
  assign \new_[16879]_  = A166 & A167;
  assign \new_[16883]_  = ~A203 & ~A202;
  assign \new_[16884]_  = A201 & \new_[16883]_ ;
  assign \new_[16885]_  = \new_[16884]_  & \new_[16879]_ ;
  assign \new_[16889]_  = A267 & A266;
  assign \new_[16890]_  = ~A265 & \new_[16889]_ ;
  assign \new_[16894]_  = ~A299 & ~A298;
  assign \new_[16895]_  = A268 & \new_[16894]_ ;
  assign \new_[16896]_  = \new_[16895]_  & \new_[16890]_ ;
  assign \new_[16899]_  = A166 & A167;
  assign \new_[16903]_  = ~A203 & ~A202;
  assign \new_[16904]_  = A201 & \new_[16903]_ ;
  assign \new_[16905]_  = \new_[16904]_  & \new_[16899]_ ;
  assign \new_[16909]_  = A267 & A266;
  assign \new_[16910]_  = ~A265 & \new_[16909]_ ;
  assign \new_[16914]_  = A301 & ~A300;
  assign \new_[16915]_  = A269 & \new_[16914]_ ;
  assign \new_[16916]_  = \new_[16915]_  & \new_[16910]_ ;
  assign \new_[16919]_  = A166 & A167;
  assign \new_[16923]_  = ~A203 & ~A202;
  assign \new_[16924]_  = A201 & \new_[16923]_ ;
  assign \new_[16925]_  = \new_[16924]_  & \new_[16919]_ ;
  assign \new_[16929]_  = A267 & A266;
  assign \new_[16930]_  = ~A265 & \new_[16929]_ ;
  assign \new_[16934]_  = A302 & ~A300;
  assign \new_[16935]_  = A269 & \new_[16934]_ ;
  assign \new_[16936]_  = \new_[16935]_  & \new_[16930]_ ;
  assign \new_[16939]_  = A166 & A167;
  assign \new_[16943]_  = ~A203 & ~A202;
  assign \new_[16944]_  = A201 & \new_[16943]_ ;
  assign \new_[16945]_  = \new_[16944]_  & \new_[16939]_ ;
  assign \new_[16949]_  = A267 & A266;
  assign \new_[16950]_  = ~A265 & \new_[16949]_ ;
  assign \new_[16954]_  = A299 & A298;
  assign \new_[16955]_  = A269 & \new_[16954]_ ;
  assign \new_[16956]_  = \new_[16955]_  & \new_[16950]_ ;
  assign \new_[16959]_  = A166 & A167;
  assign \new_[16963]_  = ~A203 & ~A202;
  assign \new_[16964]_  = A201 & \new_[16963]_ ;
  assign \new_[16965]_  = \new_[16964]_  & \new_[16959]_ ;
  assign \new_[16969]_  = A267 & A266;
  assign \new_[16970]_  = ~A265 & \new_[16969]_ ;
  assign \new_[16974]_  = ~A299 & ~A298;
  assign \new_[16975]_  = A269 & \new_[16974]_ ;
  assign \new_[16976]_  = \new_[16975]_  & \new_[16970]_ ;
  assign \new_[16979]_  = A166 & A167;
  assign \new_[16983]_  = ~A203 & ~A202;
  assign \new_[16984]_  = A201 & \new_[16983]_ ;
  assign \new_[16985]_  = \new_[16984]_  & \new_[16979]_ ;
  assign \new_[16989]_  = A267 & ~A266;
  assign \new_[16990]_  = A265 & \new_[16989]_ ;
  assign \new_[16994]_  = A301 & ~A300;
  assign \new_[16995]_  = A268 & \new_[16994]_ ;
  assign \new_[16996]_  = \new_[16995]_  & \new_[16990]_ ;
  assign \new_[16999]_  = A166 & A167;
  assign \new_[17003]_  = ~A203 & ~A202;
  assign \new_[17004]_  = A201 & \new_[17003]_ ;
  assign \new_[17005]_  = \new_[17004]_  & \new_[16999]_ ;
  assign \new_[17009]_  = A267 & ~A266;
  assign \new_[17010]_  = A265 & \new_[17009]_ ;
  assign \new_[17014]_  = A302 & ~A300;
  assign \new_[17015]_  = A268 & \new_[17014]_ ;
  assign \new_[17016]_  = \new_[17015]_  & \new_[17010]_ ;
  assign \new_[17019]_  = A166 & A167;
  assign \new_[17023]_  = ~A203 & ~A202;
  assign \new_[17024]_  = A201 & \new_[17023]_ ;
  assign \new_[17025]_  = \new_[17024]_  & \new_[17019]_ ;
  assign \new_[17029]_  = A267 & ~A266;
  assign \new_[17030]_  = A265 & \new_[17029]_ ;
  assign \new_[17034]_  = A299 & A298;
  assign \new_[17035]_  = A268 & \new_[17034]_ ;
  assign \new_[17036]_  = \new_[17035]_  & \new_[17030]_ ;
  assign \new_[17039]_  = A166 & A167;
  assign \new_[17043]_  = ~A203 & ~A202;
  assign \new_[17044]_  = A201 & \new_[17043]_ ;
  assign \new_[17045]_  = \new_[17044]_  & \new_[17039]_ ;
  assign \new_[17049]_  = A267 & ~A266;
  assign \new_[17050]_  = A265 & \new_[17049]_ ;
  assign \new_[17054]_  = ~A299 & ~A298;
  assign \new_[17055]_  = A268 & \new_[17054]_ ;
  assign \new_[17056]_  = \new_[17055]_  & \new_[17050]_ ;
  assign \new_[17059]_  = A166 & A167;
  assign \new_[17063]_  = ~A203 & ~A202;
  assign \new_[17064]_  = A201 & \new_[17063]_ ;
  assign \new_[17065]_  = \new_[17064]_  & \new_[17059]_ ;
  assign \new_[17069]_  = A267 & ~A266;
  assign \new_[17070]_  = A265 & \new_[17069]_ ;
  assign \new_[17074]_  = A301 & ~A300;
  assign \new_[17075]_  = A269 & \new_[17074]_ ;
  assign \new_[17076]_  = \new_[17075]_  & \new_[17070]_ ;
  assign \new_[17079]_  = A166 & A167;
  assign \new_[17083]_  = ~A203 & ~A202;
  assign \new_[17084]_  = A201 & \new_[17083]_ ;
  assign \new_[17085]_  = \new_[17084]_  & \new_[17079]_ ;
  assign \new_[17089]_  = A267 & ~A266;
  assign \new_[17090]_  = A265 & \new_[17089]_ ;
  assign \new_[17094]_  = A302 & ~A300;
  assign \new_[17095]_  = A269 & \new_[17094]_ ;
  assign \new_[17096]_  = \new_[17095]_  & \new_[17090]_ ;
  assign \new_[17099]_  = A166 & A167;
  assign \new_[17103]_  = ~A203 & ~A202;
  assign \new_[17104]_  = A201 & \new_[17103]_ ;
  assign \new_[17105]_  = \new_[17104]_  & \new_[17099]_ ;
  assign \new_[17109]_  = A267 & ~A266;
  assign \new_[17110]_  = A265 & \new_[17109]_ ;
  assign \new_[17114]_  = A299 & A298;
  assign \new_[17115]_  = A269 & \new_[17114]_ ;
  assign \new_[17116]_  = \new_[17115]_  & \new_[17110]_ ;
  assign \new_[17119]_  = A166 & A167;
  assign \new_[17123]_  = ~A203 & ~A202;
  assign \new_[17124]_  = A201 & \new_[17123]_ ;
  assign \new_[17125]_  = \new_[17124]_  & \new_[17119]_ ;
  assign \new_[17129]_  = A267 & ~A266;
  assign \new_[17130]_  = A265 & \new_[17129]_ ;
  assign \new_[17134]_  = ~A299 & ~A298;
  assign \new_[17135]_  = A269 & \new_[17134]_ ;
  assign \new_[17136]_  = \new_[17135]_  & \new_[17130]_ ;
  assign \new_[17139]_  = A166 & A167;
  assign \new_[17143]_  = ~A265 & A202;
  assign \new_[17144]_  = ~A201 & \new_[17143]_ ;
  assign \new_[17145]_  = \new_[17144]_  & \new_[17139]_ ;
  assign \new_[17149]_  = A268 & A267;
  assign \new_[17150]_  = A266 & \new_[17149]_ ;
  assign \new_[17154]_  = ~A302 & ~A301;
  assign \new_[17155]_  = A300 & \new_[17154]_ ;
  assign \new_[17156]_  = \new_[17155]_  & \new_[17150]_ ;
  assign \new_[17159]_  = A166 & A167;
  assign \new_[17163]_  = ~A265 & A202;
  assign \new_[17164]_  = ~A201 & \new_[17163]_ ;
  assign \new_[17165]_  = \new_[17164]_  & \new_[17159]_ ;
  assign \new_[17169]_  = A269 & A267;
  assign \new_[17170]_  = A266 & \new_[17169]_ ;
  assign \new_[17174]_  = ~A302 & ~A301;
  assign \new_[17175]_  = A300 & \new_[17174]_ ;
  assign \new_[17176]_  = \new_[17175]_  & \new_[17170]_ ;
  assign \new_[17179]_  = A166 & A167;
  assign \new_[17183]_  = ~A265 & A202;
  assign \new_[17184]_  = ~A201 & \new_[17183]_ ;
  assign \new_[17185]_  = \new_[17184]_  & \new_[17179]_ ;
  assign \new_[17189]_  = ~A268 & ~A267;
  assign \new_[17190]_  = A266 & \new_[17189]_ ;
  assign \new_[17194]_  = A301 & ~A300;
  assign \new_[17195]_  = ~A269 & \new_[17194]_ ;
  assign \new_[17196]_  = \new_[17195]_  & \new_[17190]_ ;
  assign \new_[17199]_  = A166 & A167;
  assign \new_[17203]_  = ~A265 & A202;
  assign \new_[17204]_  = ~A201 & \new_[17203]_ ;
  assign \new_[17205]_  = \new_[17204]_  & \new_[17199]_ ;
  assign \new_[17209]_  = ~A268 & ~A267;
  assign \new_[17210]_  = A266 & \new_[17209]_ ;
  assign \new_[17214]_  = A302 & ~A300;
  assign \new_[17215]_  = ~A269 & \new_[17214]_ ;
  assign \new_[17216]_  = \new_[17215]_  & \new_[17210]_ ;
  assign \new_[17219]_  = A166 & A167;
  assign \new_[17223]_  = ~A265 & A202;
  assign \new_[17224]_  = ~A201 & \new_[17223]_ ;
  assign \new_[17225]_  = \new_[17224]_  & \new_[17219]_ ;
  assign \new_[17229]_  = ~A268 & ~A267;
  assign \new_[17230]_  = A266 & \new_[17229]_ ;
  assign \new_[17234]_  = A299 & A298;
  assign \new_[17235]_  = ~A269 & \new_[17234]_ ;
  assign \new_[17236]_  = \new_[17235]_  & \new_[17230]_ ;
  assign \new_[17239]_  = A166 & A167;
  assign \new_[17243]_  = ~A265 & A202;
  assign \new_[17244]_  = ~A201 & \new_[17243]_ ;
  assign \new_[17245]_  = \new_[17244]_  & \new_[17239]_ ;
  assign \new_[17249]_  = ~A268 & ~A267;
  assign \new_[17250]_  = A266 & \new_[17249]_ ;
  assign \new_[17254]_  = ~A299 & ~A298;
  assign \new_[17255]_  = ~A269 & \new_[17254]_ ;
  assign \new_[17256]_  = \new_[17255]_  & \new_[17250]_ ;
  assign \new_[17259]_  = A166 & A167;
  assign \new_[17263]_  = A265 & A202;
  assign \new_[17264]_  = ~A201 & \new_[17263]_ ;
  assign \new_[17265]_  = \new_[17264]_  & \new_[17259]_ ;
  assign \new_[17269]_  = A268 & A267;
  assign \new_[17270]_  = ~A266 & \new_[17269]_ ;
  assign \new_[17274]_  = ~A302 & ~A301;
  assign \new_[17275]_  = A300 & \new_[17274]_ ;
  assign \new_[17276]_  = \new_[17275]_  & \new_[17270]_ ;
  assign \new_[17279]_  = A166 & A167;
  assign \new_[17283]_  = A265 & A202;
  assign \new_[17284]_  = ~A201 & \new_[17283]_ ;
  assign \new_[17285]_  = \new_[17284]_  & \new_[17279]_ ;
  assign \new_[17289]_  = A269 & A267;
  assign \new_[17290]_  = ~A266 & \new_[17289]_ ;
  assign \new_[17294]_  = ~A302 & ~A301;
  assign \new_[17295]_  = A300 & \new_[17294]_ ;
  assign \new_[17296]_  = \new_[17295]_  & \new_[17290]_ ;
  assign \new_[17299]_  = A166 & A167;
  assign \new_[17303]_  = A265 & A202;
  assign \new_[17304]_  = ~A201 & \new_[17303]_ ;
  assign \new_[17305]_  = \new_[17304]_  & \new_[17299]_ ;
  assign \new_[17309]_  = ~A268 & ~A267;
  assign \new_[17310]_  = ~A266 & \new_[17309]_ ;
  assign \new_[17314]_  = A301 & ~A300;
  assign \new_[17315]_  = ~A269 & \new_[17314]_ ;
  assign \new_[17316]_  = \new_[17315]_  & \new_[17310]_ ;
  assign \new_[17319]_  = A166 & A167;
  assign \new_[17323]_  = A265 & A202;
  assign \new_[17324]_  = ~A201 & \new_[17323]_ ;
  assign \new_[17325]_  = \new_[17324]_  & \new_[17319]_ ;
  assign \new_[17329]_  = ~A268 & ~A267;
  assign \new_[17330]_  = ~A266 & \new_[17329]_ ;
  assign \new_[17334]_  = A302 & ~A300;
  assign \new_[17335]_  = ~A269 & \new_[17334]_ ;
  assign \new_[17336]_  = \new_[17335]_  & \new_[17330]_ ;
  assign \new_[17339]_  = A166 & A167;
  assign \new_[17343]_  = A265 & A202;
  assign \new_[17344]_  = ~A201 & \new_[17343]_ ;
  assign \new_[17345]_  = \new_[17344]_  & \new_[17339]_ ;
  assign \new_[17349]_  = ~A268 & ~A267;
  assign \new_[17350]_  = ~A266 & \new_[17349]_ ;
  assign \new_[17354]_  = A299 & A298;
  assign \new_[17355]_  = ~A269 & \new_[17354]_ ;
  assign \new_[17356]_  = \new_[17355]_  & \new_[17350]_ ;
  assign \new_[17359]_  = A166 & A167;
  assign \new_[17363]_  = A265 & A202;
  assign \new_[17364]_  = ~A201 & \new_[17363]_ ;
  assign \new_[17365]_  = \new_[17364]_  & \new_[17359]_ ;
  assign \new_[17369]_  = ~A268 & ~A267;
  assign \new_[17370]_  = ~A266 & \new_[17369]_ ;
  assign \new_[17374]_  = ~A299 & ~A298;
  assign \new_[17375]_  = ~A269 & \new_[17374]_ ;
  assign \new_[17376]_  = \new_[17375]_  & \new_[17370]_ ;
  assign \new_[17379]_  = A166 & A167;
  assign \new_[17383]_  = ~A265 & A203;
  assign \new_[17384]_  = ~A201 & \new_[17383]_ ;
  assign \new_[17385]_  = \new_[17384]_  & \new_[17379]_ ;
  assign \new_[17389]_  = A268 & A267;
  assign \new_[17390]_  = A266 & \new_[17389]_ ;
  assign \new_[17394]_  = ~A302 & ~A301;
  assign \new_[17395]_  = A300 & \new_[17394]_ ;
  assign \new_[17396]_  = \new_[17395]_  & \new_[17390]_ ;
  assign \new_[17399]_  = A166 & A167;
  assign \new_[17403]_  = ~A265 & A203;
  assign \new_[17404]_  = ~A201 & \new_[17403]_ ;
  assign \new_[17405]_  = \new_[17404]_  & \new_[17399]_ ;
  assign \new_[17409]_  = A269 & A267;
  assign \new_[17410]_  = A266 & \new_[17409]_ ;
  assign \new_[17414]_  = ~A302 & ~A301;
  assign \new_[17415]_  = A300 & \new_[17414]_ ;
  assign \new_[17416]_  = \new_[17415]_  & \new_[17410]_ ;
  assign \new_[17419]_  = A166 & A167;
  assign \new_[17423]_  = ~A265 & A203;
  assign \new_[17424]_  = ~A201 & \new_[17423]_ ;
  assign \new_[17425]_  = \new_[17424]_  & \new_[17419]_ ;
  assign \new_[17429]_  = ~A268 & ~A267;
  assign \new_[17430]_  = A266 & \new_[17429]_ ;
  assign \new_[17434]_  = A301 & ~A300;
  assign \new_[17435]_  = ~A269 & \new_[17434]_ ;
  assign \new_[17436]_  = \new_[17435]_  & \new_[17430]_ ;
  assign \new_[17439]_  = A166 & A167;
  assign \new_[17443]_  = ~A265 & A203;
  assign \new_[17444]_  = ~A201 & \new_[17443]_ ;
  assign \new_[17445]_  = \new_[17444]_  & \new_[17439]_ ;
  assign \new_[17449]_  = ~A268 & ~A267;
  assign \new_[17450]_  = A266 & \new_[17449]_ ;
  assign \new_[17454]_  = A302 & ~A300;
  assign \new_[17455]_  = ~A269 & \new_[17454]_ ;
  assign \new_[17456]_  = \new_[17455]_  & \new_[17450]_ ;
  assign \new_[17459]_  = A166 & A167;
  assign \new_[17463]_  = ~A265 & A203;
  assign \new_[17464]_  = ~A201 & \new_[17463]_ ;
  assign \new_[17465]_  = \new_[17464]_  & \new_[17459]_ ;
  assign \new_[17469]_  = ~A268 & ~A267;
  assign \new_[17470]_  = A266 & \new_[17469]_ ;
  assign \new_[17474]_  = A299 & A298;
  assign \new_[17475]_  = ~A269 & \new_[17474]_ ;
  assign \new_[17476]_  = \new_[17475]_  & \new_[17470]_ ;
  assign \new_[17479]_  = A166 & A167;
  assign \new_[17483]_  = ~A265 & A203;
  assign \new_[17484]_  = ~A201 & \new_[17483]_ ;
  assign \new_[17485]_  = \new_[17484]_  & \new_[17479]_ ;
  assign \new_[17489]_  = ~A268 & ~A267;
  assign \new_[17490]_  = A266 & \new_[17489]_ ;
  assign \new_[17494]_  = ~A299 & ~A298;
  assign \new_[17495]_  = ~A269 & \new_[17494]_ ;
  assign \new_[17496]_  = \new_[17495]_  & \new_[17490]_ ;
  assign \new_[17499]_  = A166 & A167;
  assign \new_[17503]_  = A265 & A203;
  assign \new_[17504]_  = ~A201 & \new_[17503]_ ;
  assign \new_[17505]_  = \new_[17504]_  & \new_[17499]_ ;
  assign \new_[17509]_  = A268 & A267;
  assign \new_[17510]_  = ~A266 & \new_[17509]_ ;
  assign \new_[17514]_  = ~A302 & ~A301;
  assign \new_[17515]_  = A300 & \new_[17514]_ ;
  assign \new_[17516]_  = \new_[17515]_  & \new_[17510]_ ;
  assign \new_[17519]_  = A166 & A167;
  assign \new_[17523]_  = A265 & A203;
  assign \new_[17524]_  = ~A201 & \new_[17523]_ ;
  assign \new_[17525]_  = \new_[17524]_  & \new_[17519]_ ;
  assign \new_[17529]_  = A269 & A267;
  assign \new_[17530]_  = ~A266 & \new_[17529]_ ;
  assign \new_[17534]_  = ~A302 & ~A301;
  assign \new_[17535]_  = A300 & \new_[17534]_ ;
  assign \new_[17536]_  = \new_[17535]_  & \new_[17530]_ ;
  assign \new_[17539]_  = A166 & A167;
  assign \new_[17543]_  = A265 & A203;
  assign \new_[17544]_  = ~A201 & \new_[17543]_ ;
  assign \new_[17545]_  = \new_[17544]_  & \new_[17539]_ ;
  assign \new_[17549]_  = ~A268 & ~A267;
  assign \new_[17550]_  = ~A266 & \new_[17549]_ ;
  assign \new_[17554]_  = A301 & ~A300;
  assign \new_[17555]_  = ~A269 & \new_[17554]_ ;
  assign \new_[17556]_  = \new_[17555]_  & \new_[17550]_ ;
  assign \new_[17559]_  = A166 & A167;
  assign \new_[17563]_  = A265 & A203;
  assign \new_[17564]_  = ~A201 & \new_[17563]_ ;
  assign \new_[17565]_  = \new_[17564]_  & \new_[17559]_ ;
  assign \new_[17569]_  = ~A268 & ~A267;
  assign \new_[17570]_  = ~A266 & \new_[17569]_ ;
  assign \new_[17574]_  = A302 & ~A300;
  assign \new_[17575]_  = ~A269 & \new_[17574]_ ;
  assign \new_[17576]_  = \new_[17575]_  & \new_[17570]_ ;
  assign \new_[17579]_  = A166 & A167;
  assign \new_[17583]_  = A265 & A203;
  assign \new_[17584]_  = ~A201 & \new_[17583]_ ;
  assign \new_[17585]_  = \new_[17584]_  & \new_[17579]_ ;
  assign \new_[17589]_  = ~A268 & ~A267;
  assign \new_[17590]_  = ~A266 & \new_[17589]_ ;
  assign \new_[17594]_  = A299 & A298;
  assign \new_[17595]_  = ~A269 & \new_[17594]_ ;
  assign \new_[17596]_  = \new_[17595]_  & \new_[17590]_ ;
  assign \new_[17599]_  = A166 & A167;
  assign \new_[17603]_  = A265 & A203;
  assign \new_[17604]_  = ~A201 & \new_[17603]_ ;
  assign \new_[17605]_  = \new_[17604]_  & \new_[17599]_ ;
  assign \new_[17609]_  = ~A268 & ~A267;
  assign \new_[17610]_  = ~A266 & \new_[17609]_ ;
  assign \new_[17614]_  = ~A299 & ~A298;
  assign \new_[17615]_  = ~A269 & \new_[17614]_ ;
  assign \new_[17616]_  = \new_[17615]_  & \new_[17610]_ ;
  assign \new_[17619]_  = A166 & A167;
  assign \new_[17623]_  = ~A265 & A200;
  assign \new_[17624]_  = A199 & \new_[17623]_ ;
  assign \new_[17625]_  = \new_[17624]_  & \new_[17619]_ ;
  assign \new_[17629]_  = A268 & A267;
  assign \new_[17630]_  = A266 & \new_[17629]_ ;
  assign \new_[17634]_  = ~A302 & ~A301;
  assign \new_[17635]_  = A300 & \new_[17634]_ ;
  assign \new_[17636]_  = \new_[17635]_  & \new_[17630]_ ;
  assign \new_[17639]_  = A166 & A167;
  assign \new_[17643]_  = ~A265 & A200;
  assign \new_[17644]_  = A199 & \new_[17643]_ ;
  assign \new_[17645]_  = \new_[17644]_  & \new_[17639]_ ;
  assign \new_[17649]_  = A269 & A267;
  assign \new_[17650]_  = A266 & \new_[17649]_ ;
  assign \new_[17654]_  = ~A302 & ~A301;
  assign \new_[17655]_  = A300 & \new_[17654]_ ;
  assign \new_[17656]_  = \new_[17655]_  & \new_[17650]_ ;
  assign \new_[17659]_  = A166 & A167;
  assign \new_[17663]_  = ~A265 & A200;
  assign \new_[17664]_  = A199 & \new_[17663]_ ;
  assign \new_[17665]_  = \new_[17664]_  & \new_[17659]_ ;
  assign \new_[17669]_  = ~A268 & ~A267;
  assign \new_[17670]_  = A266 & \new_[17669]_ ;
  assign \new_[17674]_  = A301 & ~A300;
  assign \new_[17675]_  = ~A269 & \new_[17674]_ ;
  assign \new_[17676]_  = \new_[17675]_  & \new_[17670]_ ;
  assign \new_[17679]_  = A166 & A167;
  assign \new_[17683]_  = ~A265 & A200;
  assign \new_[17684]_  = A199 & \new_[17683]_ ;
  assign \new_[17685]_  = \new_[17684]_  & \new_[17679]_ ;
  assign \new_[17689]_  = ~A268 & ~A267;
  assign \new_[17690]_  = A266 & \new_[17689]_ ;
  assign \new_[17694]_  = A302 & ~A300;
  assign \new_[17695]_  = ~A269 & \new_[17694]_ ;
  assign \new_[17696]_  = \new_[17695]_  & \new_[17690]_ ;
  assign \new_[17699]_  = A166 & A167;
  assign \new_[17703]_  = ~A265 & A200;
  assign \new_[17704]_  = A199 & \new_[17703]_ ;
  assign \new_[17705]_  = \new_[17704]_  & \new_[17699]_ ;
  assign \new_[17709]_  = ~A268 & ~A267;
  assign \new_[17710]_  = A266 & \new_[17709]_ ;
  assign \new_[17714]_  = A299 & A298;
  assign \new_[17715]_  = ~A269 & \new_[17714]_ ;
  assign \new_[17716]_  = \new_[17715]_  & \new_[17710]_ ;
  assign \new_[17719]_  = A166 & A167;
  assign \new_[17723]_  = ~A265 & A200;
  assign \new_[17724]_  = A199 & \new_[17723]_ ;
  assign \new_[17725]_  = \new_[17724]_  & \new_[17719]_ ;
  assign \new_[17729]_  = ~A268 & ~A267;
  assign \new_[17730]_  = A266 & \new_[17729]_ ;
  assign \new_[17734]_  = ~A299 & ~A298;
  assign \new_[17735]_  = ~A269 & \new_[17734]_ ;
  assign \new_[17736]_  = \new_[17735]_  & \new_[17730]_ ;
  assign \new_[17739]_  = A166 & A167;
  assign \new_[17743]_  = A265 & A200;
  assign \new_[17744]_  = A199 & \new_[17743]_ ;
  assign \new_[17745]_  = \new_[17744]_  & \new_[17739]_ ;
  assign \new_[17749]_  = A268 & A267;
  assign \new_[17750]_  = ~A266 & \new_[17749]_ ;
  assign \new_[17754]_  = ~A302 & ~A301;
  assign \new_[17755]_  = A300 & \new_[17754]_ ;
  assign \new_[17756]_  = \new_[17755]_  & \new_[17750]_ ;
  assign \new_[17759]_  = A166 & A167;
  assign \new_[17763]_  = A265 & A200;
  assign \new_[17764]_  = A199 & \new_[17763]_ ;
  assign \new_[17765]_  = \new_[17764]_  & \new_[17759]_ ;
  assign \new_[17769]_  = A269 & A267;
  assign \new_[17770]_  = ~A266 & \new_[17769]_ ;
  assign \new_[17774]_  = ~A302 & ~A301;
  assign \new_[17775]_  = A300 & \new_[17774]_ ;
  assign \new_[17776]_  = \new_[17775]_  & \new_[17770]_ ;
  assign \new_[17779]_  = A166 & A167;
  assign \new_[17783]_  = A265 & A200;
  assign \new_[17784]_  = A199 & \new_[17783]_ ;
  assign \new_[17785]_  = \new_[17784]_  & \new_[17779]_ ;
  assign \new_[17789]_  = ~A268 & ~A267;
  assign \new_[17790]_  = ~A266 & \new_[17789]_ ;
  assign \new_[17794]_  = A301 & ~A300;
  assign \new_[17795]_  = ~A269 & \new_[17794]_ ;
  assign \new_[17796]_  = \new_[17795]_  & \new_[17790]_ ;
  assign \new_[17799]_  = A166 & A167;
  assign \new_[17803]_  = A265 & A200;
  assign \new_[17804]_  = A199 & \new_[17803]_ ;
  assign \new_[17805]_  = \new_[17804]_  & \new_[17799]_ ;
  assign \new_[17809]_  = ~A268 & ~A267;
  assign \new_[17810]_  = ~A266 & \new_[17809]_ ;
  assign \new_[17814]_  = A302 & ~A300;
  assign \new_[17815]_  = ~A269 & \new_[17814]_ ;
  assign \new_[17816]_  = \new_[17815]_  & \new_[17810]_ ;
  assign \new_[17819]_  = A166 & A167;
  assign \new_[17823]_  = A265 & A200;
  assign \new_[17824]_  = A199 & \new_[17823]_ ;
  assign \new_[17825]_  = \new_[17824]_  & \new_[17819]_ ;
  assign \new_[17829]_  = ~A268 & ~A267;
  assign \new_[17830]_  = ~A266 & \new_[17829]_ ;
  assign \new_[17834]_  = A299 & A298;
  assign \new_[17835]_  = ~A269 & \new_[17834]_ ;
  assign \new_[17836]_  = \new_[17835]_  & \new_[17830]_ ;
  assign \new_[17839]_  = A166 & A167;
  assign \new_[17843]_  = A265 & A200;
  assign \new_[17844]_  = A199 & \new_[17843]_ ;
  assign \new_[17845]_  = \new_[17844]_  & \new_[17839]_ ;
  assign \new_[17849]_  = ~A268 & ~A267;
  assign \new_[17850]_  = ~A266 & \new_[17849]_ ;
  assign \new_[17854]_  = ~A299 & ~A298;
  assign \new_[17855]_  = ~A269 & \new_[17854]_ ;
  assign \new_[17856]_  = \new_[17855]_  & \new_[17850]_ ;
  assign \new_[17859]_  = A166 & A167;
  assign \new_[17863]_  = ~A265 & ~A200;
  assign \new_[17864]_  = ~A199 & \new_[17863]_ ;
  assign \new_[17865]_  = \new_[17864]_  & \new_[17859]_ ;
  assign \new_[17869]_  = A268 & A267;
  assign \new_[17870]_  = A266 & \new_[17869]_ ;
  assign \new_[17874]_  = ~A302 & ~A301;
  assign \new_[17875]_  = A300 & \new_[17874]_ ;
  assign \new_[17876]_  = \new_[17875]_  & \new_[17870]_ ;
  assign \new_[17879]_  = A166 & A167;
  assign \new_[17883]_  = ~A265 & ~A200;
  assign \new_[17884]_  = ~A199 & \new_[17883]_ ;
  assign \new_[17885]_  = \new_[17884]_  & \new_[17879]_ ;
  assign \new_[17889]_  = A269 & A267;
  assign \new_[17890]_  = A266 & \new_[17889]_ ;
  assign \new_[17894]_  = ~A302 & ~A301;
  assign \new_[17895]_  = A300 & \new_[17894]_ ;
  assign \new_[17896]_  = \new_[17895]_  & \new_[17890]_ ;
  assign \new_[17899]_  = A166 & A167;
  assign \new_[17903]_  = ~A265 & ~A200;
  assign \new_[17904]_  = ~A199 & \new_[17903]_ ;
  assign \new_[17905]_  = \new_[17904]_  & \new_[17899]_ ;
  assign \new_[17909]_  = ~A268 & ~A267;
  assign \new_[17910]_  = A266 & \new_[17909]_ ;
  assign \new_[17914]_  = A301 & ~A300;
  assign \new_[17915]_  = ~A269 & \new_[17914]_ ;
  assign \new_[17916]_  = \new_[17915]_  & \new_[17910]_ ;
  assign \new_[17919]_  = A166 & A167;
  assign \new_[17923]_  = ~A265 & ~A200;
  assign \new_[17924]_  = ~A199 & \new_[17923]_ ;
  assign \new_[17925]_  = \new_[17924]_  & \new_[17919]_ ;
  assign \new_[17929]_  = ~A268 & ~A267;
  assign \new_[17930]_  = A266 & \new_[17929]_ ;
  assign \new_[17934]_  = A302 & ~A300;
  assign \new_[17935]_  = ~A269 & \new_[17934]_ ;
  assign \new_[17936]_  = \new_[17935]_  & \new_[17930]_ ;
  assign \new_[17939]_  = A166 & A167;
  assign \new_[17943]_  = ~A265 & ~A200;
  assign \new_[17944]_  = ~A199 & \new_[17943]_ ;
  assign \new_[17945]_  = \new_[17944]_  & \new_[17939]_ ;
  assign \new_[17949]_  = ~A268 & ~A267;
  assign \new_[17950]_  = A266 & \new_[17949]_ ;
  assign \new_[17954]_  = A299 & A298;
  assign \new_[17955]_  = ~A269 & \new_[17954]_ ;
  assign \new_[17956]_  = \new_[17955]_  & \new_[17950]_ ;
  assign \new_[17959]_  = A166 & A167;
  assign \new_[17963]_  = ~A265 & ~A200;
  assign \new_[17964]_  = ~A199 & \new_[17963]_ ;
  assign \new_[17965]_  = \new_[17964]_  & \new_[17959]_ ;
  assign \new_[17969]_  = ~A268 & ~A267;
  assign \new_[17970]_  = A266 & \new_[17969]_ ;
  assign \new_[17974]_  = ~A299 & ~A298;
  assign \new_[17975]_  = ~A269 & \new_[17974]_ ;
  assign \new_[17976]_  = \new_[17975]_  & \new_[17970]_ ;
  assign \new_[17979]_  = A166 & A167;
  assign \new_[17983]_  = A265 & ~A200;
  assign \new_[17984]_  = ~A199 & \new_[17983]_ ;
  assign \new_[17985]_  = \new_[17984]_  & \new_[17979]_ ;
  assign \new_[17989]_  = A268 & A267;
  assign \new_[17990]_  = ~A266 & \new_[17989]_ ;
  assign \new_[17994]_  = ~A302 & ~A301;
  assign \new_[17995]_  = A300 & \new_[17994]_ ;
  assign \new_[17996]_  = \new_[17995]_  & \new_[17990]_ ;
  assign \new_[17999]_  = A166 & A167;
  assign \new_[18003]_  = A265 & ~A200;
  assign \new_[18004]_  = ~A199 & \new_[18003]_ ;
  assign \new_[18005]_  = \new_[18004]_  & \new_[17999]_ ;
  assign \new_[18009]_  = A269 & A267;
  assign \new_[18010]_  = ~A266 & \new_[18009]_ ;
  assign \new_[18014]_  = ~A302 & ~A301;
  assign \new_[18015]_  = A300 & \new_[18014]_ ;
  assign \new_[18016]_  = \new_[18015]_  & \new_[18010]_ ;
  assign \new_[18019]_  = A166 & A167;
  assign \new_[18023]_  = A265 & ~A200;
  assign \new_[18024]_  = ~A199 & \new_[18023]_ ;
  assign \new_[18025]_  = \new_[18024]_  & \new_[18019]_ ;
  assign \new_[18029]_  = ~A268 & ~A267;
  assign \new_[18030]_  = ~A266 & \new_[18029]_ ;
  assign \new_[18034]_  = A301 & ~A300;
  assign \new_[18035]_  = ~A269 & \new_[18034]_ ;
  assign \new_[18036]_  = \new_[18035]_  & \new_[18030]_ ;
  assign \new_[18039]_  = A166 & A167;
  assign \new_[18043]_  = A265 & ~A200;
  assign \new_[18044]_  = ~A199 & \new_[18043]_ ;
  assign \new_[18045]_  = \new_[18044]_  & \new_[18039]_ ;
  assign \new_[18049]_  = ~A268 & ~A267;
  assign \new_[18050]_  = ~A266 & \new_[18049]_ ;
  assign \new_[18054]_  = A302 & ~A300;
  assign \new_[18055]_  = ~A269 & \new_[18054]_ ;
  assign \new_[18056]_  = \new_[18055]_  & \new_[18050]_ ;
  assign \new_[18059]_  = A166 & A167;
  assign \new_[18063]_  = A265 & ~A200;
  assign \new_[18064]_  = ~A199 & \new_[18063]_ ;
  assign \new_[18065]_  = \new_[18064]_  & \new_[18059]_ ;
  assign \new_[18069]_  = ~A268 & ~A267;
  assign \new_[18070]_  = ~A266 & \new_[18069]_ ;
  assign \new_[18074]_  = A299 & A298;
  assign \new_[18075]_  = ~A269 & \new_[18074]_ ;
  assign \new_[18076]_  = \new_[18075]_  & \new_[18070]_ ;
  assign \new_[18079]_  = A166 & A167;
  assign \new_[18083]_  = A265 & ~A200;
  assign \new_[18084]_  = ~A199 & \new_[18083]_ ;
  assign \new_[18085]_  = \new_[18084]_  & \new_[18079]_ ;
  assign \new_[18089]_  = ~A268 & ~A267;
  assign \new_[18090]_  = ~A266 & \new_[18089]_ ;
  assign \new_[18094]_  = ~A299 & ~A298;
  assign \new_[18095]_  = ~A269 & \new_[18094]_ ;
  assign \new_[18096]_  = \new_[18095]_  & \new_[18090]_ ;
  assign \new_[18099]_  = ~A166 & ~A167;
  assign \new_[18103]_  = ~A203 & ~A202;
  assign \new_[18104]_  = A201 & \new_[18103]_ ;
  assign \new_[18105]_  = \new_[18104]_  & \new_[18099]_ ;
  assign \new_[18109]_  = A267 & A266;
  assign \new_[18110]_  = ~A265 & \new_[18109]_ ;
  assign \new_[18114]_  = A301 & ~A300;
  assign \new_[18115]_  = A268 & \new_[18114]_ ;
  assign \new_[18116]_  = \new_[18115]_  & \new_[18110]_ ;
  assign \new_[18119]_  = ~A166 & ~A167;
  assign \new_[18123]_  = ~A203 & ~A202;
  assign \new_[18124]_  = A201 & \new_[18123]_ ;
  assign \new_[18125]_  = \new_[18124]_  & \new_[18119]_ ;
  assign \new_[18129]_  = A267 & A266;
  assign \new_[18130]_  = ~A265 & \new_[18129]_ ;
  assign \new_[18134]_  = A302 & ~A300;
  assign \new_[18135]_  = A268 & \new_[18134]_ ;
  assign \new_[18136]_  = \new_[18135]_  & \new_[18130]_ ;
  assign \new_[18139]_  = ~A166 & ~A167;
  assign \new_[18143]_  = ~A203 & ~A202;
  assign \new_[18144]_  = A201 & \new_[18143]_ ;
  assign \new_[18145]_  = \new_[18144]_  & \new_[18139]_ ;
  assign \new_[18149]_  = A267 & A266;
  assign \new_[18150]_  = ~A265 & \new_[18149]_ ;
  assign \new_[18154]_  = A299 & A298;
  assign \new_[18155]_  = A268 & \new_[18154]_ ;
  assign \new_[18156]_  = \new_[18155]_  & \new_[18150]_ ;
  assign \new_[18159]_  = ~A166 & ~A167;
  assign \new_[18163]_  = ~A203 & ~A202;
  assign \new_[18164]_  = A201 & \new_[18163]_ ;
  assign \new_[18165]_  = \new_[18164]_  & \new_[18159]_ ;
  assign \new_[18169]_  = A267 & A266;
  assign \new_[18170]_  = ~A265 & \new_[18169]_ ;
  assign \new_[18174]_  = ~A299 & ~A298;
  assign \new_[18175]_  = A268 & \new_[18174]_ ;
  assign \new_[18176]_  = \new_[18175]_  & \new_[18170]_ ;
  assign \new_[18179]_  = ~A166 & ~A167;
  assign \new_[18183]_  = ~A203 & ~A202;
  assign \new_[18184]_  = A201 & \new_[18183]_ ;
  assign \new_[18185]_  = \new_[18184]_  & \new_[18179]_ ;
  assign \new_[18189]_  = A267 & A266;
  assign \new_[18190]_  = ~A265 & \new_[18189]_ ;
  assign \new_[18194]_  = A301 & ~A300;
  assign \new_[18195]_  = A269 & \new_[18194]_ ;
  assign \new_[18196]_  = \new_[18195]_  & \new_[18190]_ ;
  assign \new_[18199]_  = ~A166 & ~A167;
  assign \new_[18203]_  = ~A203 & ~A202;
  assign \new_[18204]_  = A201 & \new_[18203]_ ;
  assign \new_[18205]_  = \new_[18204]_  & \new_[18199]_ ;
  assign \new_[18209]_  = A267 & A266;
  assign \new_[18210]_  = ~A265 & \new_[18209]_ ;
  assign \new_[18214]_  = A302 & ~A300;
  assign \new_[18215]_  = A269 & \new_[18214]_ ;
  assign \new_[18216]_  = \new_[18215]_  & \new_[18210]_ ;
  assign \new_[18219]_  = ~A166 & ~A167;
  assign \new_[18223]_  = ~A203 & ~A202;
  assign \new_[18224]_  = A201 & \new_[18223]_ ;
  assign \new_[18225]_  = \new_[18224]_  & \new_[18219]_ ;
  assign \new_[18229]_  = A267 & A266;
  assign \new_[18230]_  = ~A265 & \new_[18229]_ ;
  assign \new_[18234]_  = A299 & A298;
  assign \new_[18235]_  = A269 & \new_[18234]_ ;
  assign \new_[18236]_  = \new_[18235]_  & \new_[18230]_ ;
  assign \new_[18239]_  = ~A166 & ~A167;
  assign \new_[18243]_  = ~A203 & ~A202;
  assign \new_[18244]_  = A201 & \new_[18243]_ ;
  assign \new_[18245]_  = \new_[18244]_  & \new_[18239]_ ;
  assign \new_[18249]_  = A267 & A266;
  assign \new_[18250]_  = ~A265 & \new_[18249]_ ;
  assign \new_[18254]_  = ~A299 & ~A298;
  assign \new_[18255]_  = A269 & \new_[18254]_ ;
  assign \new_[18256]_  = \new_[18255]_  & \new_[18250]_ ;
  assign \new_[18259]_  = ~A166 & ~A167;
  assign \new_[18263]_  = ~A203 & ~A202;
  assign \new_[18264]_  = A201 & \new_[18263]_ ;
  assign \new_[18265]_  = \new_[18264]_  & \new_[18259]_ ;
  assign \new_[18269]_  = A267 & ~A266;
  assign \new_[18270]_  = A265 & \new_[18269]_ ;
  assign \new_[18274]_  = A301 & ~A300;
  assign \new_[18275]_  = A268 & \new_[18274]_ ;
  assign \new_[18276]_  = \new_[18275]_  & \new_[18270]_ ;
  assign \new_[18279]_  = ~A166 & ~A167;
  assign \new_[18283]_  = ~A203 & ~A202;
  assign \new_[18284]_  = A201 & \new_[18283]_ ;
  assign \new_[18285]_  = \new_[18284]_  & \new_[18279]_ ;
  assign \new_[18289]_  = A267 & ~A266;
  assign \new_[18290]_  = A265 & \new_[18289]_ ;
  assign \new_[18294]_  = A302 & ~A300;
  assign \new_[18295]_  = A268 & \new_[18294]_ ;
  assign \new_[18296]_  = \new_[18295]_  & \new_[18290]_ ;
  assign \new_[18299]_  = ~A166 & ~A167;
  assign \new_[18303]_  = ~A203 & ~A202;
  assign \new_[18304]_  = A201 & \new_[18303]_ ;
  assign \new_[18305]_  = \new_[18304]_  & \new_[18299]_ ;
  assign \new_[18309]_  = A267 & ~A266;
  assign \new_[18310]_  = A265 & \new_[18309]_ ;
  assign \new_[18314]_  = A299 & A298;
  assign \new_[18315]_  = A268 & \new_[18314]_ ;
  assign \new_[18316]_  = \new_[18315]_  & \new_[18310]_ ;
  assign \new_[18319]_  = ~A166 & ~A167;
  assign \new_[18323]_  = ~A203 & ~A202;
  assign \new_[18324]_  = A201 & \new_[18323]_ ;
  assign \new_[18325]_  = \new_[18324]_  & \new_[18319]_ ;
  assign \new_[18329]_  = A267 & ~A266;
  assign \new_[18330]_  = A265 & \new_[18329]_ ;
  assign \new_[18334]_  = ~A299 & ~A298;
  assign \new_[18335]_  = A268 & \new_[18334]_ ;
  assign \new_[18336]_  = \new_[18335]_  & \new_[18330]_ ;
  assign \new_[18339]_  = ~A166 & ~A167;
  assign \new_[18343]_  = ~A203 & ~A202;
  assign \new_[18344]_  = A201 & \new_[18343]_ ;
  assign \new_[18345]_  = \new_[18344]_  & \new_[18339]_ ;
  assign \new_[18349]_  = A267 & ~A266;
  assign \new_[18350]_  = A265 & \new_[18349]_ ;
  assign \new_[18354]_  = A301 & ~A300;
  assign \new_[18355]_  = A269 & \new_[18354]_ ;
  assign \new_[18356]_  = \new_[18355]_  & \new_[18350]_ ;
  assign \new_[18359]_  = ~A166 & ~A167;
  assign \new_[18363]_  = ~A203 & ~A202;
  assign \new_[18364]_  = A201 & \new_[18363]_ ;
  assign \new_[18365]_  = \new_[18364]_  & \new_[18359]_ ;
  assign \new_[18369]_  = A267 & ~A266;
  assign \new_[18370]_  = A265 & \new_[18369]_ ;
  assign \new_[18374]_  = A302 & ~A300;
  assign \new_[18375]_  = A269 & \new_[18374]_ ;
  assign \new_[18376]_  = \new_[18375]_  & \new_[18370]_ ;
  assign \new_[18379]_  = ~A166 & ~A167;
  assign \new_[18383]_  = ~A203 & ~A202;
  assign \new_[18384]_  = A201 & \new_[18383]_ ;
  assign \new_[18385]_  = \new_[18384]_  & \new_[18379]_ ;
  assign \new_[18389]_  = A267 & ~A266;
  assign \new_[18390]_  = A265 & \new_[18389]_ ;
  assign \new_[18394]_  = A299 & A298;
  assign \new_[18395]_  = A269 & \new_[18394]_ ;
  assign \new_[18396]_  = \new_[18395]_  & \new_[18390]_ ;
  assign \new_[18399]_  = ~A166 & ~A167;
  assign \new_[18403]_  = ~A203 & ~A202;
  assign \new_[18404]_  = A201 & \new_[18403]_ ;
  assign \new_[18405]_  = \new_[18404]_  & \new_[18399]_ ;
  assign \new_[18409]_  = A267 & ~A266;
  assign \new_[18410]_  = A265 & \new_[18409]_ ;
  assign \new_[18414]_  = ~A299 & ~A298;
  assign \new_[18415]_  = A269 & \new_[18414]_ ;
  assign \new_[18416]_  = \new_[18415]_  & \new_[18410]_ ;
  assign \new_[18419]_  = ~A166 & ~A167;
  assign \new_[18423]_  = ~A265 & A202;
  assign \new_[18424]_  = ~A201 & \new_[18423]_ ;
  assign \new_[18425]_  = \new_[18424]_  & \new_[18419]_ ;
  assign \new_[18429]_  = A268 & A267;
  assign \new_[18430]_  = A266 & \new_[18429]_ ;
  assign \new_[18434]_  = ~A302 & ~A301;
  assign \new_[18435]_  = A300 & \new_[18434]_ ;
  assign \new_[18436]_  = \new_[18435]_  & \new_[18430]_ ;
  assign \new_[18439]_  = ~A166 & ~A167;
  assign \new_[18443]_  = ~A265 & A202;
  assign \new_[18444]_  = ~A201 & \new_[18443]_ ;
  assign \new_[18445]_  = \new_[18444]_  & \new_[18439]_ ;
  assign \new_[18449]_  = A269 & A267;
  assign \new_[18450]_  = A266 & \new_[18449]_ ;
  assign \new_[18454]_  = ~A302 & ~A301;
  assign \new_[18455]_  = A300 & \new_[18454]_ ;
  assign \new_[18456]_  = \new_[18455]_  & \new_[18450]_ ;
  assign \new_[18459]_  = ~A166 & ~A167;
  assign \new_[18463]_  = ~A265 & A202;
  assign \new_[18464]_  = ~A201 & \new_[18463]_ ;
  assign \new_[18465]_  = \new_[18464]_  & \new_[18459]_ ;
  assign \new_[18469]_  = ~A268 & ~A267;
  assign \new_[18470]_  = A266 & \new_[18469]_ ;
  assign \new_[18474]_  = A301 & ~A300;
  assign \new_[18475]_  = ~A269 & \new_[18474]_ ;
  assign \new_[18476]_  = \new_[18475]_  & \new_[18470]_ ;
  assign \new_[18479]_  = ~A166 & ~A167;
  assign \new_[18483]_  = ~A265 & A202;
  assign \new_[18484]_  = ~A201 & \new_[18483]_ ;
  assign \new_[18485]_  = \new_[18484]_  & \new_[18479]_ ;
  assign \new_[18489]_  = ~A268 & ~A267;
  assign \new_[18490]_  = A266 & \new_[18489]_ ;
  assign \new_[18494]_  = A302 & ~A300;
  assign \new_[18495]_  = ~A269 & \new_[18494]_ ;
  assign \new_[18496]_  = \new_[18495]_  & \new_[18490]_ ;
  assign \new_[18499]_  = ~A166 & ~A167;
  assign \new_[18503]_  = ~A265 & A202;
  assign \new_[18504]_  = ~A201 & \new_[18503]_ ;
  assign \new_[18505]_  = \new_[18504]_  & \new_[18499]_ ;
  assign \new_[18509]_  = ~A268 & ~A267;
  assign \new_[18510]_  = A266 & \new_[18509]_ ;
  assign \new_[18514]_  = A299 & A298;
  assign \new_[18515]_  = ~A269 & \new_[18514]_ ;
  assign \new_[18516]_  = \new_[18515]_  & \new_[18510]_ ;
  assign \new_[18519]_  = ~A166 & ~A167;
  assign \new_[18523]_  = ~A265 & A202;
  assign \new_[18524]_  = ~A201 & \new_[18523]_ ;
  assign \new_[18525]_  = \new_[18524]_  & \new_[18519]_ ;
  assign \new_[18529]_  = ~A268 & ~A267;
  assign \new_[18530]_  = A266 & \new_[18529]_ ;
  assign \new_[18534]_  = ~A299 & ~A298;
  assign \new_[18535]_  = ~A269 & \new_[18534]_ ;
  assign \new_[18536]_  = \new_[18535]_  & \new_[18530]_ ;
  assign \new_[18539]_  = ~A166 & ~A167;
  assign \new_[18543]_  = A265 & A202;
  assign \new_[18544]_  = ~A201 & \new_[18543]_ ;
  assign \new_[18545]_  = \new_[18544]_  & \new_[18539]_ ;
  assign \new_[18549]_  = A268 & A267;
  assign \new_[18550]_  = ~A266 & \new_[18549]_ ;
  assign \new_[18554]_  = ~A302 & ~A301;
  assign \new_[18555]_  = A300 & \new_[18554]_ ;
  assign \new_[18556]_  = \new_[18555]_  & \new_[18550]_ ;
  assign \new_[18559]_  = ~A166 & ~A167;
  assign \new_[18563]_  = A265 & A202;
  assign \new_[18564]_  = ~A201 & \new_[18563]_ ;
  assign \new_[18565]_  = \new_[18564]_  & \new_[18559]_ ;
  assign \new_[18569]_  = A269 & A267;
  assign \new_[18570]_  = ~A266 & \new_[18569]_ ;
  assign \new_[18574]_  = ~A302 & ~A301;
  assign \new_[18575]_  = A300 & \new_[18574]_ ;
  assign \new_[18576]_  = \new_[18575]_  & \new_[18570]_ ;
  assign \new_[18579]_  = ~A166 & ~A167;
  assign \new_[18583]_  = A265 & A202;
  assign \new_[18584]_  = ~A201 & \new_[18583]_ ;
  assign \new_[18585]_  = \new_[18584]_  & \new_[18579]_ ;
  assign \new_[18589]_  = ~A268 & ~A267;
  assign \new_[18590]_  = ~A266 & \new_[18589]_ ;
  assign \new_[18594]_  = A301 & ~A300;
  assign \new_[18595]_  = ~A269 & \new_[18594]_ ;
  assign \new_[18596]_  = \new_[18595]_  & \new_[18590]_ ;
  assign \new_[18599]_  = ~A166 & ~A167;
  assign \new_[18603]_  = A265 & A202;
  assign \new_[18604]_  = ~A201 & \new_[18603]_ ;
  assign \new_[18605]_  = \new_[18604]_  & \new_[18599]_ ;
  assign \new_[18609]_  = ~A268 & ~A267;
  assign \new_[18610]_  = ~A266 & \new_[18609]_ ;
  assign \new_[18614]_  = A302 & ~A300;
  assign \new_[18615]_  = ~A269 & \new_[18614]_ ;
  assign \new_[18616]_  = \new_[18615]_  & \new_[18610]_ ;
  assign \new_[18619]_  = ~A166 & ~A167;
  assign \new_[18623]_  = A265 & A202;
  assign \new_[18624]_  = ~A201 & \new_[18623]_ ;
  assign \new_[18625]_  = \new_[18624]_  & \new_[18619]_ ;
  assign \new_[18629]_  = ~A268 & ~A267;
  assign \new_[18630]_  = ~A266 & \new_[18629]_ ;
  assign \new_[18634]_  = A299 & A298;
  assign \new_[18635]_  = ~A269 & \new_[18634]_ ;
  assign \new_[18636]_  = \new_[18635]_  & \new_[18630]_ ;
  assign \new_[18639]_  = ~A166 & ~A167;
  assign \new_[18643]_  = A265 & A202;
  assign \new_[18644]_  = ~A201 & \new_[18643]_ ;
  assign \new_[18645]_  = \new_[18644]_  & \new_[18639]_ ;
  assign \new_[18649]_  = ~A268 & ~A267;
  assign \new_[18650]_  = ~A266 & \new_[18649]_ ;
  assign \new_[18654]_  = ~A299 & ~A298;
  assign \new_[18655]_  = ~A269 & \new_[18654]_ ;
  assign \new_[18656]_  = \new_[18655]_  & \new_[18650]_ ;
  assign \new_[18659]_  = ~A166 & ~A167;
  assign \new_[18663]_  = ~A265 & A203;
  assign \new_[18664]_  = ~A201 & \new_[18663]_ ;
  assign \new_[18665]_  = \new_[18664]_  & \new_[18659]_ ;
  assign \new_[18669]_  = A268 & A267;
  assign \new_[18670]_  = A266 & \new_[18669]_ ;
  assign \new_[18674]_  = ~A302 & ~A301;
  assign \new_[18675]_  = A300 & \new_[18674]_ ;
  assign \new_[18676]_  = \new_[18675]_  & \new_[18670]_ ;
  assign \new_[18679]_  = ~A166 & ~A167;
  assign \new_[18683]_  = ~A265 & A203;
  assign \new_[18684]_  = ~A201 & \new_[18683]_ ;
  assign \new_[18685]_  = \new_[18684]_  & \new_[18679]_ ;
  assign \new_[18689]_  = A269 & A267;
  assign \new_[18690]_  = A266 & \new_[18689]_ ;
  assign \new_[18694]_  = ~A302 & ~A301;
  assign \new_[18695]_  = A300 & \new_[18694]_ ;
  assign \new_[18696]_  = \new_[18695]_  & \new_[18690]_ ;
  assign \new_[18699]_  = ~A166 & ~A167;
  assign \new_[18703]_  = ~A265 & A203;
  assign \new_[18704]_  = ~A201 & \new_[18703]_ ;
  assign \new_[18705]_  = \new_[18704]_  & \new_[18699]_ ;
  assign \new_[18709]_  = ~A268 & ~A267;
  assign \new_[18710]_  = A266 & \new_[18709]_ ;
  assign \new_[18714]_  = A301 & ~A300;
  assign \new_[18715]_  = ~A269 & \new_[18714]_ ;
  assign \new_[18716]_  = \new_[18715]_  & \new_[18710]_ ;
  assign \new_[18719]_  = ~A166 & ~A167;
  assign \new_[18723]_  = ~A265 & A203;
  assign \new_[18724]_  = ~A201 & \new_[18723]_ ;
  assign \new_[18725]_  = \new_[18724]_  & \new_[18719]_ ;
  assign \new_[18729]_  = ~A268 & ~A267;
  assign \new_[18730]_  = A266 & \new_[18729]_ ;
  assign \new_[18734]_  = A302 & ~A300;
  assign \new_[18735]_  = ~A269 & \new_[18734]_ ;
  assign \new_[18736]_  = \new_[18735]_  & \new_[18730]_ ;
  assign \new_[18739]_  = ~A166 & ~A167;
  assign \new_[18743]_  = ~A265 & A203;
  assign \new_[18744]_  = ~A201 & \new_[18743]_ ;
  assign \new_[18745]_  = \new_[18744]_  & \new_[18739]_ ;
  assign \new_[18749]_  = ~A268 & ~A267;
  assign \new_[18750]_  = A266 & \new_[18749]_ ;
  assign \new_[18754]_  = A299 & A298;
  assign \new_[18755]_  = ~A269 & \new_[18754]_ ;
  assign \new_[18756]_  = \new_[18755]_  & \new_[18750]_ ;
  assign \new_[18759]_  = ~A166 & ~A167;
  assign \new_[18763]_  = ~A265 & A203;
  assign \new_[18764]_  = ~A201 & \new_[18763]_ ;
  assign \new_[18765]_  = \new_[18764]_  & \new_[18759]_ ;
  assign \new_[18769]_  = ~A268 & ~A267;
  assign \new_[18770]_  = A266 & \new_[18769]_ ;
  assign \new_[18774]_  = ~A299 & ~A298;
  assign \new_[18775]_  = ~A269 & \new_[18774]_ ;
  assign \new_[18776]_  = \new_[18775]_  & \new_[18770]_ ;
  assign \new_[18779]_  = ~A166 & ~A167;
  assign \new_[18783]_  = A265 & A203;
  assign \new_[18784]_  = ~A201 & \new_[18783]_ ;
  assign \new_[18785]_  = \new_[18784]_  & \new_[18779]_ ;
  assign \new_[18789]_  = A268 & A267;
  assign \new_[18790]_  = ~A266 & \new_[18789]_ ;
  assign \new_[18794]_  = ~A302 & ~A301;
  assign \new_[18795]_  = A300 & \new_[18794]_ ;
  assign \new_[18796]_  = \new_[18795]_  & \new_[18790]_ ;
  assign \new_[18799]_  = ~A166 & ~A167;
  assign \new_[18803]_  = A265 & A203;
  assign \new_[18804]_  = ~A201 & \new_[18803]_ ;
  assign \new_[18805]_  = \new_[18804]_  & \new_[18799]_ ;
  assign \new_[18809]_  = A269 & A267;
  assign \new_[18810]_  = ~A266 & \new_[18809]_ ;
  assign \new_[18814]_  = ~A302 & ~A301;
  assign \new_[18815]_  = A300 & \new_[18814]_ ;
  assign \new_[18816]_  = \new_[18815]_  & \new_[18810]_ ;
  assign \new_[18819]_  = ~A166 & ~A167;
  assign \new_[18823]_  = A265 & A203;
  assign \new_[18824]_  = ~A201 & \new_[18823]_ ;
  assign \new_[18825]_  = \new_[18824]_  & \new_[18819]_ ;
  assign \new_[18829]_  = ~A268 & ~A267;
  assign \new_[18830]_  = ~A266 & \new_[18829]_ ;
  assign \new_[18834]_  = A301 & ~A300;
  assign \new_[18835]_  = ~A269 & \new_[18834]_ ;
  assign \new_[18836]_  = \new_[18835]_  & \new_[18830]_ ;
  assign \new_[18839]_  = ~A166 & ~A167;
  assign \new_[18843]_  = A265 & A203;
  assign \new_[18844]_  = ~A201 & \new_[18843]_ ;
  assign \new_[18845]_  = \new_[18844]_  & \new_[18839]_ ;
  assign \new_[18849]_  = ~A268 & ~A267;
  assign \new_[18850]_  = ~A266 & \new_[18849]_ ;
  assign \new_[18854]_  = A302 & ~A300;
  assign \new_[18855]_  = ~A269 & \new_[18854]_ ;
  assign \new_[18856]_  = \new_[18855]_  & \new_[18850]_ ;
  assign \new_[18859]_  = ~A166 & ~A167;
  assign \new_[18863]_  = A265 & A203;
  assign \new_[18864]_  = ~A201 & \new_[18863]_ ;
  assign \new_[18865]_  = \new_[18864]_  & \new_[18859]_ ;
  assign \new_[18869]_  = ~A268 & ~A267;
  assign \new_[18870]_  = ~A266 & \new_[18869]_ ;
  assign \new_[18874]_  = A299 & A298;
  assign \new_[18875]_  = ~A269 & \new_[18874]_ ;
  assign \new_[18876]_  = \new_[18875]_  & \new_[18870]_ ;
  assign \new_[18879]_  = ~A166 & ~A167;
  assign \new_[18883]_  = A265 & A203;
  assign \new_[18884]_  = ~A201 & \new_[18883]_ ;
  assign \new_[18885]_  = \new_[18884]_  & \new_[18879]_ ;
  assign \new_[18889]_  = ~A268 & ~A267;
  assign \new_[18890]_  = ~A266 & \new_[18889]_ ;
  assign \new_[18894]_  = ~A299 & ~A298;
  assign \new_[18895]_  = ~A269 & \new_[18894]_ ;
  assign \new_[18896]_  = \new_[18895]_  & \new_[18890]_ ;
  assign \new_[18899]_  = ~A166 & ~A167;
  assign \new_[18903]_  = ~A265 & A200;
  assign \new_[18904]_  = A199 & \new_[18903]_ ;
  assign \new_[18905]_  = \new_[18904]_  & \new_[18899]_ ;
  assign \new_[18909]_  = A268 & A267;
  assign \new_[18910]_  = A266 & \new_[18909]_ ;
  assign \new_[18914]_  = ~A302 & ~A301;
  assign \new_[18915]_  = A300 & \new_[18914]_ ;
  assign \new_[18916]_  = \new_[18915]_  & \new_[18910]_ ;
  assign \new_[18919]_  = ~A166 & ~A167;
  assign \new_[18923]_  = ~A265 & A200;
  assign \new_[18924]_  = A199 & \new_[18923]_ ;
  assign \new_[18925]_  = \new_[18924]_  & \new_[18919]_ ;
  assign \new_[18929]_  = A269 & A267;
  assign \new_[18930]_  = A266 & \new_[18929]_ ;
  assign \new_[18934]_  = ~A302 & ~A301;
  assign \new_[18935]_  = A300 & \new_[18934]_ ;
  assign \new_[18936]_  = \new_[18935]_  & \new_[18930]_ ;
  assign \new_[18939]_  = ~A166 & ~A167;
  assign \new_[18943]_  = ~A265 & A200;
  assign \new_[18944]_  = A199 & \new_[18943]_ ;
  assign \new_[18945]_  = \new_[18944]_  & \new_[18939]_ ;
  assign \new_[18949]_  = ~A268 & ~A267;
  assign \new_[18950]_  = A266 & \new_[18949]_ ;
  assign \new_[18954]_  = A301 & ~A300;
  assign \new_[18955]_  = ~A269 & \new_[18954]_ ;
  assign \new_[18956]_  = \new_[18955]_  & \new_[18950]_ ;
  assign \new_[18959]_  = ~A166 & ~A167;
  assign \new_[18963]_  = ~A265 & A200;
  assign \new_[18964]_  = A199 & \new_[18963]_ ;
  assign \new_[18965]_  = \new_[18964]_  & \new_[18959]_ ;
  assign \new_[18969]_  = ~A268 & ~A267;
  assign \new_[18970]_  = A266 & \new_[18969]_ ;
  assign \new_[18974]_  = A302 & ~A300;
  assign \new_[18975]_  = ~A269 & \new_[18974]_ ;
  assign \new_[18976]_  = \new_[18975]_  & \new_[18970]_ ;
  assign \new_[18979]_  = ~A166 & ~A167;
  assign \new_[18983]_  = ~A265 & A200;
  assign \new_[18984]_  = A199 & \new_[18983]_ ;
  assign \new_[18985]_  = \new_[18984]_  & \new_[18979]_ ;
  assign \new_[18989]_  = ~A268 & ~A267;
  assign \new_[18990]_  = A266 & \new_[18989]_ ;
  assign \new_[18994]_  = A299 & A298;
  assign \new_[18995]_  = ~A269 & \new_[18994]_ ;
  assign \new_[18996]_  = \new_[18995]_  & \new_[18990]_ ;
  assign \new_[18999]_  = ~A166 & ~A167;
  assign \new_[19003]_  = ~A265 & A200;
  assign \new_[19004]_  = A199 & \new_[19003]_ ;
  assign \new_[19005]_  = \new_[19004]_  & \new_[18999]_ ;
  assign \new_[19009]_  = ~A268 & ~A267;
  assign \new_[19010]_  = A266 & \new_[19009]_ ;
  assign \new_[19014]_  = ~A299 & ~A298;
  assign \new_[19015]_  = ~A269 & \new_[19014]_ ;
  assign \new_[19016]_  = \new_[19015]_  & \new_[19010]_ ;
  assign \new_[19019]_  = ~A166 & ~A167;
  assign \new_[19023]_  = A265 & A200;
  assign \new_[19024]_  = A199 & \new_[19023]_ ;
  assign \new_[19025]_  = \new_[19024]_  & \new_[19019]_ ;
  assign \new_[19029]_  = A268 & A267;
  assign \new_[19030]_  = ~A266 & \new_[19029]_ ;
  assign \new_[19034]_  = ~A302 & ~A301;
  assign \new_[19035]_  = A300 & \new_[19034]_ ;
  assign \new_[19036]_  = \new_[19035]_  & \new_[19030]_ ;
  assign \new_[19039]_  = ~A166 & ~A167;
  assign \new_[19043]_  = A265 & A200;
  assign \new_[19044]_  = A199 & \new_[19043]_ ;
  assign \new_[19045]_  = \new_[19044]_  & \new_[19039]_ ;
  assign \new_[19049]_  = A269 & A267;
  assign \new_[19050]_  = ~A266 & \new_[19049]_ ;
  assign \new_[19054]_  = ~A302 & ~A301;
  assign \new_[19055]_  = A300 & \new_[19054]_ ;
  assign \new_[19056]_  = \new_[19055]_  & \new_[19050]_ ;
  assign \new_[19059]_  = ~A166 & ~A167;
  assign \new_[19063]_  = A265 & A200;
  assign \new_[19064]_  = A199 & \new_[19063]_ ;
  assign \new_[19065]_  = \new_[19064]_  & \new_[19059]_ ;
  assign \new_[19069]_  = ~A268 & ~A267;
  assign \new_[19070]_  = ~A266 & \new_[19069]_ ;
  assign \new_[19074]_  = A301 & ~A300;
  assign \new_[19075]_  = ~A269 & \new_[19074]_ ;
  assign \new_[19076]_  = \new_[19075]_  & \new_[19070]_ ;
  assign \new_[19079]_  = ~A166 & ~A167;
  assign \new_[19083]_  = A265 & A200;
  assign \new_[19084]_  = A199 & \new_[19083]_ ;
  assign \new_[19085]_  = \new_[19084]_  & \new_[19079]_ ;
  assign \new_[19089]_  = ~A268 & ~A267;
  assign \new_[19090]_  = ~A266 & \new_[19089]_ ;
  assign \new_[19094]_  = A302 & ~A300;
  assign \new_[19095]_  = ~A269 & \new_[19094]_ ;
  assign \new_[19096]_  = \new_[19095]_  & \new_[19090]_ ;
  assign \new_[19099]_  = ~A166 & ~A167;
  assign \new_[19103]_  = A265 & A200;
  assign \new_[19104]_  = A199 & \new_[19103]_ ;
  assign \new_[19105]_  = \new_[19104]_  & \new_[19099]_ ;
  assign \new_[19109]_  = ~A268 & ~A267;
  assign \new_[19110]_  = ~A266 & \new_[19109]_ ;
  assign \new_[19114]_  = A299 & A298;
  assign \new_[19115]_  = ~A269 & \new_[19114]_ ;
  assign \new_[19116]_  = \new_[19115]_  & \new_[19110]_ ;
  assign \new_[19119]_  = ~A166 & ~A167;
  assign \new_[19123]_  = A265 & A200;
  assign \new_[19124]_  = A199 & \new_[19123]_ ;
  assign \new_[19125]_  = \new_[19124]_  & \new_[19119]_ ;
  assign \new_[19129]_  = ~A268 & ~A267;
  assign \new_[19130]_  = ~A266 & \new_[19129]_ ;
  assign \new_[19134]_  = ~A299 & ~A298;
  assign \new_[19135]_  = ~A269 & \new_[19134]_ ;
  assign \new_[19136]_  = \new_[19135]_  & \new_[19130]_ ;
  assign \new_[19139]_  = ~A166 & ~A167;
  assign \new_[19143]_  = ~A265 & ~A200;
  assign \new_[19144]_  = ~A199 & \new_[19143]_ ;
  assign \new_[19145]_  = \new_[19144]_  & \new_[19139]_ ;
  assign \new_[19149]_  = A268 & A267;
  assign \new_[19150]_  = A266 & \new_[19149]_ ;
  assign \new_[19154]_  = ~A302 & ~A301;
  assign \new_[19155]_  = A300 & \new_[19154]_ ;
  assign \new_[19156]_  = \new_[19155]_  & \new_[19150]_ ;
  assign \new_[19159]_  = ~A166 & ~A167;
  assign \new_[19163]_  = ~A265 & ~A200;
  assign \new_[19164]_  = ~A199 & \new_[19163]_ ;
  assign \new_[19165]_  = \new_[19164]_  & \new_[19159]_ ;
  assign \new_[19169]_  = A269 & A267;
  assign \new_[19170]_  = A266 & \new_[19169]_ ;
  assign \new_[19174]_  = ~A302 & ~A301;
  assign \new_[19175]_  = A300 & \new_[19174]_ ;
  assign \new_[19176]_  = \new_[19175]_  & \new_[19170]_ ;
  assign \new_[19179]_  = ~A166 & ~A167;
  assign \new_[19183]_  = ~A265 & ~A200;
  assign \new_[19184]_  = ~A199 & \new_[19183]_ ;
  assign \new_[19185]_  = \new_[19184]_  & \new_[19179]_ ;
  assign \new_[19189]_  = ~A268 & ~A267;
  assign \new_[19190]_  = A266 & \new_[19189]_ ;
  assign \new_[19194]_  = A301 & ~A300;
  assign \new_[19195]_  = ~A269 & \new_[19194]_ ;
  assign \new_[19196]_  = \new_[19195]_  & \new_[19190]_ ;
  assign \new_[19199]_  = ~A166 & ~A167;
  assign \new_[19203]_  = ~A265 & ~A200;
  assign \new_[19204]_  = ~A199 & \new_[19203]_ ;
  assign \new_[19205]_  = \new_[19204]_  & \new_[19199]_ ;
  assign \new_[19209]_  = ~A268 & ~A267;
  assign \new_[19210]_  = A266 & \new_[19209]_ ;
  assign \new_[19214]_  = A302 & ~A300;
  assign \new_[19215]_  = ~A269 & \new_[19214]_ ;
  assign \new_[19216]_  = \new_[19215]_  & \new_[19210]_ ;
  assign \new_[19219]_  = ~A166 & ~A167;
  assign \new_[19223]_  = ~A265 & ~A200;
  assign \new_[19224]_  = ~A199 & \new_[19223]_ ;
  assign \new_[19225]_  = \new_[19224]_  & \new_[19219]_ ;
  assign \new_[19229]_  = ~A268 & ~A267;
  assign \new_[19230]_  = A266 & \new_[19229]_ ;
  assign \new_[19234]_  = A299 & A298;
  assign \new_[19235]_  = ~A269 & \new_[19234]_ ;
  assign \new_[19236]_  = \new_[19235]_  & \new_[19230]_ ;
  assign \new_[19239]_  = ~A166 & ~A167;
  assign \new_[19243]_  = ~A265 & ~A200;
  assign \new_[19244]_  = ~A199 & \new_[19243]_ ;
  assign \new_[19245]_  = \new_[19244]_  & \new_[19239]_ ;
  assign \new_[19249]_  = ~A268 & ~A267;
  assign \new_[19250]_  = A266 & \new_[19249]_ ;
  assign \new_[19254]_  = ~A299 & ~A298;
  assign \new_[19255]_  = ~A269 & \new_[19254]_ ;
  assign \new_[19256]_  = \new_[19255]_  & \new_[19250]_ ;
  assign \new_[19259]_  = ~A166 & ~A167;
  assign \new_[19263]_  = A265 & ~A200;
  assign \new_[19264]_  = ~A199 & \new_[19263]_ ;
  assign \new_[19265]_  = \new_[19264]_  & \new_[19259]_ ;
  assign \new_[19269]_  = A268 & A267;
  assign \new_[19270]_  = ~A266 & \new_[19269]_ ;
  assign \new_[19274]_  = ~A302 & ~A301;
  assign \new_[19275]_  = A300 & \new_[19274]_ ;
  assign \new_[19276]_  = \new_[19275]_  & \new_[19270]_ ;
  assign \new_[19279]_  = ~A166 & ~A167;
  assign \new_[19283]_  = A265 & ~A200;
  assign \new_[19284]_  = ~A199 & \new_[19283]_ ;
  assign \new_[19285]_  = \new_[19284]_  & \new_[19279]_ ;
  assign \new_[19289]_  = A269 & A267;
  assign \new_[19290]_  = ~A266 & \new_[19289]_ ;
  assign \new_[19294]_  = ~A302 & ~A301;
  assign \new_[19295]_  = A300 & \new_[19294]_ ;
  assign \new_[19296]_  = \new_[19295]_  & \new_[19290]_ ;
  assign \new_[19299]_  = ~A166 & ~A167;
  assign \new_[19303]_  = A265 & ~A200;
  assign \new_[19304]_  = ~A199 & \new_[19303]_ ;
  assign \new_[19305]_  = \new_[19304]_  & \new_[19299]_ ;
  assign \new_[19309]_  = ~A268 & ~A267;
  assign \new_[19310]_  = ~A266 & \new_[19309]_ ;
  assign \new_[19314]_  = A301 & ~A300;
  assign \new_[19315]_  = ~A269 & \new_[19314]_ ;
  assign \new_[19316]_  = \new_[19315]_  & \new_[19310]_ ;
  assign \new_[19319]_  = ~A166 & ~A167;
  assign \new_[19323]_  = A265 & ~A200;
  assign \new_[19324]_  = ~A199 & \new_[19323]_ ;
  assign \new_[19325]_  = \new_[19324]_  & \new_[19319]_ ;
  assign \new_[19329]_  = ~A268 & ~A267;
  assign \new_[19330]_  = ~A266 & \new_[19329]_ ;
  assign \new_[19334]_  = A302 & ~A300;
  assign \new_[19335]_  = ~A269 & \new_[19334]_ ;
  assign \new_[19336]_  = \new_[19335]_  & \new_[19330]_ ;
  assign \new_[19339]_  = ~A166 & ~A167;
  assign \new_[19343]_  = A265 & ~A200;
  assign \new_[19344]_  = ~A199 & \new_[19343]_ ;
  assign \new_[19345]_  = \new_[19344]_  & \new_[19339]_ ;
  assign \new_[19349]_  = ~A268 & ~A267;
  assign \new_[19350]_  = ~A266 & \new_[19349]_ ;
  assign \new_[19354]_  = A299 & A298;
  assign \new_[19355]_  = ~A269 & \new_[19354]_ ;
  assign \new_[19356]_  = \new_[19355]_  & \new_[19350]_ ;
  assign \new_[19359]_  = ~A166 & ~A167;
  assign \new_[19363]_  = A265 & ~A200;
  assign \new_[19364]_  = ~A199 & \new_[19363]_ ;
  assign \new_[19365]_  = \new_[19364]_  & \new_[19359]_ ;
  assign \new_[19369]_  = ~A268 & ~A267;
  assign \new_[19370]_  = ~A266 & \new_[19369]_ ;
  assign \new_[19374]_  = ~A299 & ~A298;
  assign \new_[19375]_  = ~A269 & \new_[19374]_ ;
  assign \new_[19376]_  = \new_[19375]_  & \new_[19370]_ ;
  assign \new_[19379]_  = ~A168 & ~A170;
  assign \new_[19383]_  = ~A203 & ~A202;
  assign \new_[19384]_  = A201 & \new_[19383]_ ;
  assign \new_[19385]_  = \new_[19384]_  & \new_[19379]_ ;
  assign \new_[19389]_  = A267 & A266;
  assign \new_[19390]_  = ~A265 & \new_[19389]_ ;
  assign \new_[19394]_  = A301 & ~A300;
  assign \new_[19395]_  = A268 & \new_[19394]_ ;
  assign \new_[19396]_  = \new_[19395]_  & \new_[19390]_ ;
  assign \new_[19399]_  = ~A168 & ~A170;
  assign \new_[19403]_  = ~A203 & ~A202;
  assign \new_[19404]_  = A201 & \new_[19403]_ ;
  assign \new_[19405]_  = \new_[19404]_  & \new_[19399]_ ;
  assign \new_[19409]_  = A267 & A266;
  assign \new_[19410]_  = ~A265 & \new_[19409]_ ;
  assign \new_[19414]_  = A302 & ~A300;
  assign \new_[19415]_  = A268 & \new_[19414]_ ;
  assign \new_[19416]_  = \new_[19415]_  & \new_[19410]_ ;
  assign \new_[19419]_  = ~A168 & ~A170;
  assign \new_[19423]_  = ~A203 & ~A202;
  assign \new_[19424]_  = A201 & \new_[19423]_ ;
  assign \new_[19425]_  = \new_[19424]_  & \new_[19419]_ ;
  assign \new_[19429]_  = A267 & A266;
  assign \new_[19430]_  = ~A265 & \new_[19429]_ ;
  assign \new_[19434]_  = A299 & A298;
  assign \new_[19435]_  = A268 & \new_[19434]_ ;
  assign \new_[19436]_  = \new_[19435]_  & \new_[19430]_ ;
  assign \new_[19439]_  = ~A168 & ~A170;
  assign \new_[19443]_  = ~A203 & ~A202;
  assign \new_[19444]_  = A201 & \new_[19443]_ ;
  assign \new_[19445]_  = \new_[19444]_  & \new_[19439]_ ;
  assign \new_[19449]_  = A267 & A266;
  assign \new_[19450]_  = ~A265 & \new_[19449]_ ;
  assign \new_[19454]_  = ~A299 & ~A298;
  assign \new_[19455]_  = A268 & \new_[19454]_ ;
  assign \new_[19456]_  = \new_[19455]_  & \new_[19450]_ ;
  assign \new_[19459]_  = ~A168 & ~A170;
  assign \new_[19463]_  = ~A203 & ~A202;
  assign \new_[19464]_  = A201 & \new_[19463]_ ;
  assign \new_[19465]_  = \new_[19464]_  & \new_[19459]_ ;
  assign \new_[19469]_  = A267 & A266;
  assign \new_[19470]_  = ~A265 & \new_[19469]_ ;
  assign \new_[19474]_  = A301 & ~A300;
  assign \new_[19475]_  = A269 & \new_[19474]_ ;
  assign \new_[19476]_  = \new_[19475]_  & \new_[19470]_ ;
  assign \new_[19479]_  = ~A168 & ~A170;
  assign \new_[19483]_  = ~A203 & ~A202;
  assign \new_[19484]_  = A201 & \new_[19483]_ ;
  assign \new_[19485]_  = \new_[19484]_  & \new_[19479]_ ;
  assign \new_[19489]_  = A267 & A266;
  assign \new_[19490]_  = ~A265 & \new_[19489]_ ;
  assign \new_[19494]_  = A302 & ~A300;
  assign \new_[19495]_  = A269 & \new_[19494]_ ;
  assign \new_[19496]_  = \new_[19495]_  & \new_[19490]_ ;
  assign \new_[19499]_  = ~A168 & ~A170;
  assign \new_[19503]_  = ~A203 & ~A202;
  assign \new_[19504]_  = A201 & \new_[19503]_ ;
  assign \new_[19505]_  = \new_[19504]_  & \new_[19499]_ ;
  assign \new_[19509]_  = A267 & A266;
  assign \new_[19510]_  = ~A265 & \new_[19509]_ ;
  assign \new_[19514]_  = A299 & A298;
  assign \new_[19515]_  = A269 & \new_[19514]_ ;
  assign \new_[19516]_  = \new_[19515]_  & \new_[19510]_ ;
  assign \new_[19519]_  = ~A168 & ~A170;
  assign \new_[19523]_  = ~A203 & ~A202;
  assign \new_[19524]_  = A201 & \new_[19523]_ ;
  assign \new_[19525]_  = \new_[19524]_  & \new_[19519]_ ;
  assign \new_[19529]_  = A267 & A266;
  assign \new_[19530]_  = ~A265 & \new_[19529]_ ;
  assign \new_[19534]_  = ~A299 & ~A298;
  assign \new_[19535]_  = A269 & \new_[19534]_ ;
  assign \new_[19536]_  = \new_[19535]_  & \new_[19530]_ ;
  assign \new_[19539]_  = ~A168 & ~A170;
  assign \new_[19543]_  = ~A203 & ~A202;
  assign \new_[19544]_  = A201 & \new_[19543]_ ;
  assign \new_[19545]_  = \new_[19544]_  & \new_[19539]_ ;
  assign \new_[19549]_  = A267 & ~A266;
  assign \new_[19550]_  = A265 & \new_[19549]_ ;
  assign \new_[19554]_  = A301 & ~A300;
  assign \new_[19555]_  = A268 & \new_[19554]_ ;
  assign \new_[19556]_  = \new_[19555]_  & \new_[19550]_ ;
  assign \new_[19559]_  = ~A168 & ~A170;
  assign \new_[19563]_  = ~A203 & ~A202;
  assign \new_[19564]_  = A201 & \new_[19563]_ ;
  assign \new_[19565]_  = \new_[19564]_  & \new_[19559]_ ;
  assign \new_[19569]_  = A267 & ~A266;
  assign \new_[19570]_  = A265 & \new_[19569]_ ;
  assign \new_[19574]_  = A302 & ~A300;
  assign \new_[19575]_  = A268 & \new_[19574]_ ;
  assign \new_[19576]_  = \new_[19575]_  & \new_[19570]_ ;
  assign \new_[19579]_  = ~A168 & ~A170;
  assign \new_[19583]_  = ~A203 & ~A202;
  assign \new_[19584]_  = A201 & \new_[19583]_ ;
  assign \new_[19585]_  = \new_[19584]_  & \new_[19579]_ ;
  assign \new_[19589]_  = A267 & ~A266;
  assign \new_[19590]_  = A265 & \new_[19589]_ ;
  assign \new_[19594]_  = A299 & A298;
  assign \new_[19595]_  = A268 & \new_[19594]_ ;
  assign \new_[19596]_  = \new_[19595]_  & \new_[19590]_ ;
  assign \new_[19599]_  = ~A168 & ~A170;
  assign \new_[19603]_  = ~A203 & ~A202;
  assign \new_[19604]_  = A201 & \new_[19603]_ ;
  assign \new_[19605]_  = \new_[19604]_  & \new_[19599]_ ;
  assign \new_[19609]_  = A267 & ~A266;
  assign \new_[19610]_  = A265 & \new_[19609]_ ;
  assign \new_[19614]_  = ~A299 & ~A298;
  assign \new_[19615]_  = A268 & \new_[19614]_ ;
  assign \new_[19616]_  = \new_[19615]_  & \new_[19610]_ ;
  assign \new_[19619]_  = ~A168 & ~A170;
  assign \new_[19623]_  = ~A203 & ~A202;
  assign \new_[19624]_  = A201 & \new_[19623]_ ;
  assign \new_[19625]_  = \new_[19624]_  & \new_[19619]_ ;
  assign \new_[19629]_  = A267 & ~A266;
  assign \new_[19630]_  = A265 & \new_[19629]_ ;
  assign \new_[19634]_  = A301 & ~A300;
  assign \new_[19635]_  = A269 & \new_[19634]_ ;
  assign \new_[19636]_  = \new_[19635]_  & \new_[19630]_ ;
  assign \new_[19639]_  = ~A168 & ~A170;
  assign \new_[19643]_  = ~A203 & ~A202;
  assign \new_[19644]_  = A201 & \new_[19643]_ ;
  assign \new_[19645]_  = \new_[19644]_  & \new_[19639]_ ;
  assign \new_[19649]_  = A267 & ~A266;
  assign \new_[19650]_  = A265 & \new_[19649]_ ;
  assign \new_[19654]_  = A302 & ~A300;
  assign \new_[19655]_  = A269 & \new_[19654]_ ;
  assign \new_[19656]_  = \new_[19655]_  & \new_[19650]_ ;
  assign \new_[19659]_  = ~A168 & ~A170;
  assign \new_[19663]_  = ~A203 & ~A202;
  assign \new_[19664]_  = A201 & \new_[19663]_ ;
  assign \new_[19665]_  = \new_[19664]_  & \new_[19659]_ ;
  assign \new_[19669]_  = A267 & ~A266;
  assign \new_[19670]_  = A265 & \new_[19669]_ ;
  assign \new_[19674]_  = A299 & A298;
  assign \new_[19675]_  = A269 & \new_[19674]_ ;
  assign \new_[19676]_  = \new_[19675]_  & \new_[19670]_ ;
  assign \new_[19679]_  = ~A168 & ~A170;
  assign \new_[19683]_  = ~A203 & ~A202;
  assign \new_[19684]_  = A201 & \new_[19683]_ ;
  assign \new_[19685]_  = \new_[19684]_  & \new_[19679]_ ;
  assign \new_[19689]_  = A267 & ~A266;
  assign \new_[19690]_  = A265 & \new_[19689]_ ;
  assign \new_[19694]_  = ~A299 & ~A298;
  assign \new_[19695]_  = A269 & \new_[19694]_ ;
  assign \new_[19696]_  = \new_[19695]_  & \new_[19690]_ ;
  assign \new_[19699]_  = ~A168 & ~A170;
  assign \new_[19703]_  = ~A265 & A202;
  assign \new_[19704]_  = ~A201 & \new_[19703]_ ;
  assign \new_[19705]_  = \new_[19704]_  & \new_[19699]_ ;
  assign \new_[19709]_  = A268 & A267;
  assign \new_[19710]_  = A266 & \new_[19709]_ ;
  assign \new_[19714]_  = ~A302 & ~A301;
  assign \new_[19715]_  = A300 & \new_[19714]_ ;
  assign \new_[19716]_  = \new_[19715]_  & \new_[19710]_ ;
  assign \new_[19719]_  = ~A168 & ~A170;
  assign \new_[19723]_  = ~A265 & A202;
  assign \new_[19724]_  = ~A201 & \new_[19723]_ ;
  assign \new_[19725]_  = \new_[19724]_  & \new_[19719]_ ;
  assign \new_[19729]_  = A269 & A267;
  assign \new_[19730]_  = A266 & \new_[19729]_ ;
  assign \new_[19734]_  = ~A302 & ~A301;
  assign \new_[19735]_  = A300 & \new_[19734]_ ;
  assign \new_[19736]_  = \new_[19735]_  & \new_[19730]_ ;
  assign \new_[19739]_  = ~A168 & ~A170;
  assign \new_[19743]_  = ~A265 & A202;
  assign \new_[19744]_  = ~A201 & \new_[19743]_ ;
  assign \new_[19745]_  = \new_[19744]_  & \new_[19739]_ ;
  assign \new_[19749]_  = ~A268 & ~A267;
  assign \new_[19750]_  = A266 & \new_[19749]_ ;
  assign \new_[19754]_  = A301 & ~A300;
  assign \new_[19755]_  = ~A269 & \new_[19754]_ ;
  assign \new_[19756]_  = \new_[19755]_  & \new_[19750]_ ;
  assign \new_[19759]_  = ~A168 & ~A170;
  assign \new_[19763]_  = ~A265 & A202;
  assign \new_[19764]_  = ~A201 & \new_[19763]_ ;
  assign \new_[19765]_  = \new_[19764]_  & \new_[19759]_ ;
  assign \new_[19769]_  = ~A268 & ~A267;
  assign \new_[19770]_  = A266 & \new_[19769]_ ;
  assign \new_[19774]_  = A302 & ~A300;
  assign \new_[19775]_  = ~A269 & \new_[19774]_ ;
  assign \new_[19776]_  = \new_[19775]_  & \new_[19770]_ ;
  assign \new_[19779]_  = ~A168 & ~A170;
  assign \new_[19783]_  = ~A265 & A202;
  assign \new_[19784]_  = ~A201 & \new_[19783]_ ;
  assign \new_[19785]_  = \new_[19784]_  & \new_[19779]_ ;
  assign \new_[19789]_  = ~A268 & ~A267;
  assign \new_[19790]_  = A266 & \new_[19789]_ ;
  assign \new_[19794]_  = A299 & A298;
  assign \new_[19795]_  = ~A269 & \new_[19794]_ ;
  assign \new_[19796]_  = \new_[19795]_  & \new_[19790]_ ;
  assign \new_[19799]_  = ~A168 & ~A170;
  assign \new_[19803]_  = ~A265 & A202;
  assign \new_[19804]_  = ~A201 & \new_[19803]_ ;
  assign \new_[19805]_  = \new_[19804]_  & \new_[19799]_ ;
  assign \new_[19809]_  = ~A268 & ~A267;
  assign \new_[19810]_  = A266 & \new_[19809]_ ;
  assign \new_[19814]_  = ~A299 & ~A298;
  assign \new_[19815]_  = ~A269 & \new_[19814]_ ;
  assign \new_[19816]_  = \new_[19815]_  & \new_[19810]_ ;
  assign \new_[19819]_  = ~A168 & ~A170;
  assign \new_[19823]_  = A265 & A202;
  assign \new_[19824]_  = ~A201 & \new_[19823]_ ;
  assign \new_[19825]_  = \new_[19824]_  & \new_[19819]_ ;
  assign \new_[19829]_  = A268 & A267;
  assign \new_[19830]_  = ~A266 & \new_[19829]_ ;
  assign \new_[19834]_  = ~A302 & ~A301;
  assign \new_[19835]_  = A300 & \new_[19834]_ ;
  assign \new_[19836]_  = \new_[19835]_  & \new_[19830]_ ;
  assign \new_[19839]_  = ~A168 & ~A170;
  assign \new_[19843]_  = A265 & A202;
  assign \new_[19844]_  = ~A201 & \new_[19843]_ ;
  assign \new_[19845]_  = \new_[19844]_  & \new_[19839]_ ;
  assign \new_[19849]_  = A269 & A267;
  assign \new_[19850]_  = ~A266 & \new_[19849]_ ;
  assign \new_[19854]_  = ~A302 & ~A301;
  assign \new_[19855]_  = A300 & \new_[19854]_ ;
  assign \new_[19856]_  = \new_[19855]_  & \new_[19850]_ ;
  assign \new_[19859]_  = ~A168 & ~A170;
  assign \new_[19863]_  = A265 & A202;
  assign \new_[19864]_  = ~A201 & \new_[19863]_ ;
  assign \new_[19865]_  = \new_[19864]_  & \new_[19859]_ ;
  assign \new_[19869]_  = ~A268 & ~A267;
  assign \new_[19870]_  = ~A266 & \new_[19869]_ ;
  assign \new_[19874]_  = A301 & ~A300;
  assign \new_[19875]_  = ~A269 & \new_[19874]_ ;
  assign \new_[19876]_  = \new_[19875]_  & \new_[19870]_ ;
  assign \new_[19879]_  = ~A168 & ~A170;
  assign \new_[19883]_  = A265 & A202;
  assign \new_[19884]_  = ~A201 & \new_[19883]_ ;
  assign \new_[19885]_  = \new_[19884]_  & \new_[19879]_ ;
  assign \new_[19889]_  = ~A268 & ~A267;
  assign \new_[19890]_  = ~A266 & \new_[19889]_ ;
  assign \new_[19894]_  = A302 & ~A300;
  assign \new_[19895]_  = ~A269 & \new_[19894]_ ;
  assign \new_[19896]_  = \new_[19895]_  & \new_[19890]_ ;
  assign \new_[19899]_  = ~A168 & ~A170;
  assign \new_[19903]_  = A265 & A202;
  assign \new_[19904]_  = ~A201 & \new_[19903]_ ;
  assign \new_[19905]_  = \new_[19904]_  & \new_[19899]_ ;
  assign \new_[19909]_  = ~A268 & ~A267;
  assign \new_[19910]_  = ~A266 & \new_[19909]_ ;
  assign \new_[19914]_  = A299 & A298;
  assign \new_[19915]_  = ~A269 & \new_[19914]_ ;
  assign \new_[19916]_  = \new_[19915]_  & \new_[19910]_ ;
  assign \new_[19919]_  = ~A168 & ~A170;
  assign \new_[19923]_  = A265 & A202;
  assign \new_[19924]_  = ~A201 & \new_[19923]_ ;
  assign \new_[19925]_  = \new_[19924]_  & \new_[19919]_ ;
  assign \new_[19929]_  = ~A268 & ~A267;
  assign \new_[19930]_  = ~A266 & \new_[19929]_ ;
  assign \new_[19934]_  = ~A299 & ~A298;
  assign \new_[19935]_  = ~A269 & \new_[19934]_ ;
  assign \new_[19936]_  = \new_[19935]_  & \new_[19930]_ ;
  assign \new_[19939]_  = ~A168 & ~A170;
  assign \new_[19943]_  = ~A265 & A203;
  assign \new_[19944]_  = ~A201 & \new_[19943]_ ;
  assign \new_[19945]_  = \new_[19944]_  & \new_[19939]_ ;
  assign \new_[19949]_  = A268 & A267;
  assign \new_[19950]_  = A266 & \new_[19949]_ ;
  assign \new_[19954]_  = ~A302 & ~A301;
  assign \new_[19955]_  = A300 & \new_[19954]_ ;
  assign \new_[19956]_  = \new_[19955]_  & \new_[19950]_ ;
  assign \new_[19959]_  = ~A168 & ~A170;
  assign \new_[19963]_  = ~A265 & A203;
  assign \new_[19964]_  = ~A201 & \new_[19963]_ ;
  assign \new_[19965]_  = \new_[19964]_  & \new_[19959]_ ;
  assign \new_[19969]_  = A269 & A267;
  assign \new_[19970]_  = A266 & \new_[19969]_ ;
  assign \new_[19974]_  = ~A302 & ~A301;
  assign \new_[19975]_  = A300 & \new_[19974]_ ;
  assign \new_[19976]_  = \new_[19975]_  & \new_[19970]_ ;
  assign \new_[19979]_  = ~A168 & ~A170;
  assign \new_[19983]_  = ~A265 & A203;
  assign \new_[19984]_  = ~A201 & \new_[19983]_ ;
  assign \new_[19985]_  = \new_[19984]_  & \new_[19979]_ ;
  assign \new_[19989]_  = ~A268 & ~A267;
  assign \new_[19990]_  = A266 & \new_[19989]_ ;
  assign \new_[19994]_  = A301 & ~A300;
  assign \new_[19995]_  = ~A269 & \new_[19994]_ ;
  assign \new_[19996]_  = \new_[19995]_  & \new_[19990]_ ;
  assign \new_[19999]_  = ~A168 & ~A170;
  assign \new_[20003]_  = ~A265 & A203;
  assign \new_[20004]_  = ~A201 & \new_[20003]_ ;
  assign \new_[20005]_  = \new_[20004]_  & \new_[19999]_ ;
  assign \new_[20009]_  = ~A268 & ~A267;
  assign \new_[20010]_  = A266 & \new_[20009]_ ;
  assign \new_[20014]_  = A302 & ~A300;
  assign \new_[20015]_  = ~A269 & \new_[20014]_ ;
  assign \new_[20016]_  = \new_[20015]_  & \new_[20010]_ ;
  assign \new_[20019]_  = ~A168 & ~A170;
  assign \new_[20023]_  = ~A265 & A203;
  assign \new_[20024]_  = ~A201 & \new_[20023]_ ;
  assign \new_[20025]_  = \new_[20024]_  & \new_[20019]_ ;
  assign \new_[20029]_  = ~A268 & ~A267;
  assign \new_[20030]_  = A266 & \new_[20029]_ ;
  assign \new_[20034]_  = A299 & A298;
  assign \new_[20035]_  = ~A269 & \new_[20034]_ ;
  assign \new_[20036]_  = \new_[20035]_  & \new_[20030]_ ;
  assign \new_[20039]_  = ~A168 & ~A170;
  assign \new_[20043]_  = ~A265 & A203;
  assign \new_[20044]_  = ~A201 & \new_[20043]_ ;
  assign \new_[20045]_  = \new_[20044]_  & \new_[20039]_ ;
  assign \new_[20049]_  = ~A268 & ~A267;
  assign \new_[20050]_  = A266 & \new_[20049]_ ;
  assign \new_[20054]_  = ~A299 & ~A298;
  assign \new_[20055]_  = ~A269 & \new_[20054]_ ;
  assign \new_[20056]_  = \new_[20055]_  & \new_[20050]_ ;
  assign \new_[20059]_  = ~A168 & ~A170;
  assign \new_[20063]_  = A265 & A203;
  assign \new_[20064]_  = ~A201 & \new_[20063]_ ;
  assign \new_[20065]_  = \new_[20064]_  & \new_[20059]_ ;
  assign \new_[20069]_  = A268 & A267;
  assign \new_[20070]_  = ~A266 & \new_[20069]_ ;
  assign \new_[20074]_  = ~A302 & ~A301;
  assign \new_[20075]_  = A300 & \new_[20074]_ ;
  assign \new_[20076]_  = \new_[20075]_  & \new_[20070]_ ;
  assign \new_[20079]_  = ~A168 & ~A170;
  assign \new_[20083]_  = A265 & A203;
  assign \new_[20084]_  = ~A201 & \new_[20083]_ ;
  assign \new_[20085]_  = \new_[20084]_  & \new_[20079]_ ;
  assign \new_[20089]_  = A269 & A267;
  assign \new_[20090]_  = ~A266 & \new_[20089]_ ;
  assign \new_[20094]_  = ~A302 & ~A301;
  assign \new_[20095]_  = A300 & \new_[20094]_ ;
  assign \new_[20096]_  = \new_[20095]_  & \new_[20090]_ ;
  assign \new_[20099]_  = ~A168 & ~A170;
  assign \new_[20103]_  = A265 & A203;
  assign \new_[20104]_  = ~A201 & \new_[20103]_ ;
  assign \new_[20105]_  = \new_[20104]_  & \new_[20099]_ ;
  assign \new_[20109]_  = ~A268 & ~A267;
  assign \new_[20110]_  = ~A266 & \new_[20109]_ ;
  assign \new_[20114]_  = A301 & ~A300;
  assign \new_[20115]_  = ~A269 & \new_[20114]_ ;
  assign \new_[20116]_  = \new_[20115]_  & \new_[20110]_ ;
  assign \new_[20119]_  = ~A168 & ~A170;
  assign \new_[20123]_  = A265 & A203;
  assign \new_[20124]_  = ~A201 & \new_[20123]_ ;
  assign \new_[20125]_  = \new_[20124]_  & \new_[20119]_ ;
  assign \new_[20129]_  = ~A268 & ~A267;
  assign \new_[20130]_  = ~A266 & \new_[20129]_ ;
  assign \new_[20134]_  = A302 & ~A300;
  assign \new_[20135]_  = ~A269 & \new_[20134]_ ;
  assign \new_[20136]_  = \new_[20135]_  & \new_[20130]_ ;
  assign \new_[20139]_  = ~A168 & ~A170;
  assign \new_[20143]_  = A265 & A203;
  assign \new_[20144]_  = ~A201 & \new_[20143]_ ;
  assign \new_[20145]_  = \new_[20144]_  & \new_[20139]_ ;
  assign \new_[20149]_  = ~A268 & ~A267;
  assign \new_[20150]_  = ~A266 & \new_[20149]_ ;
  assign \new_[20154]_  = A299 & A298;
  assign \new_[20155]_  = ~A269 & \new_[20154]_ ;
  assign \new_[20156]_  = \new_[20155]_  & \new_[20150]_ ;
  assign \new_[20159]_  = ~A168 & ~A170;
  assign \new_[20163]_  = A265 & A203;
  assign \new_[20164]_  = ~A201 & \new_[20163]_ ;
  assign \new_[20165]_  = \new_[20164]_  & \new_[20159]_ ;
  assign \new_[20169]_  = ~A268 & ~A267;
  assign \new_[20170]_  = ~A266 & \new_[20169]_ ;
  assign \new_[20174]_  = ~A299 & ~A298;
  assign \new_[20175]_  = ~A269 & \new_[20174]_ ;
  assign \new_[20176]_  = \new_[20175]_  & \new_[20170]_ ;
  assign \new_[20179]_  = ~A168 & ~A170;
  assign \new_[20183]_  = ~A265 & A200;
  assign \new_[20184]_  = A199 & \new_[20183]_ ;
  assign \new_[20185]_  = \new_[20184]_  & \new_[20179]_ ;
  assign \new_[20189]_  = A268 & A267;
  assign \new_[20190]_  = A266 & \new_[20189]_ ;
  assign \new_[20194]_  = ~A302 & ~A301;
  assign \new_[20195]_  = A300 & \new_[20194]_ ;
  assign \new_[20196]_  = \new_[20195]_  & \new_[20190]_ ;
  assign \new_[20199]_  = ~A168 & ~A170;
  assign \new_[20203]_  = ~A265 & A200;
  assign \new_[20204]_  = A199 & \new_[20203]_ ;
  assign \new_[20205]_  = \new_[20204]_  & \new_[20199]_ ;
  assign \new_[20209]_  = A269 & A267;
  assign \new_[20210]_  = A266 & \new_[20209]_ ;
  assign \new_[20214]_  = ~A302 & ~A301;
  assign \new_[20215]_  = A300 & \new_[20214]_ ;
  assign \new_[20216]_  = \new_[20215]_  & \new_[20210]_ ;
  assign \new_[20219]_  = ~A168 & ~A170;
  assign \new_[20223]_  = ~A265 & A200;
  assign \new_[20224]_  = A199 & \new_[20223]_ ;
  assign \new_[20225]_  = \new_[20224]_  & \new_[20219]_ ;
  assign \new_[20229]_  = ~A268 & ~A267;
  assign \new_[20230]_  = A266 & \new_[20229]_ ;
  assign \new_[20234]_  = A301 & ~A300;
  assign \new_[20235]_  = ~A269 & \new_[20234]_ ;
  assign \new_[20236]_  = \new_[20235]_  & \new_[20230]_ ;
  assign \new_[20239]_  = ~A168 & ~A170;
  assign \new_[20243]_  = ~A265 & A200;
  assign \new_[20244]_  = A199 & \new_[20243]_ ;
  assign \new_[20245]_  = \new_[20244]_  & \new_[20239]_ ;
  assign \new_[20249]_  = ~A268 & ~A267;
  assign \new_[20250]_  = A266 & \new_[20249]_ ;
  assign \new_[20254]_  = A302 & ~A300;
  assign \new_[20255]_  = ~A269 & \new_[20254]_ ;
  assign \new_[20256]_  = \new_[20255]_  & \new_[20250]_ ;
  assign \new_[20259]_  = ~A168 & ~A170;
  assign \new_[20263]_  = ~A265 & A200;
  assign \new_[20264]_  = A199 & \new_[20263]_ ;
  assign \new_[20265]_  = \new_[20264]_  & \new_[20259]_ ;
  assign \new_[20269]_  = ~A268 & ~A267;
  assign \new_[20270]_  = A266 & \new_[20269]_ ;
  assign \new_[20274]_  = A299 & A298;
  assign \new_[20275]_  = ~A269 & \new_[20274]_ ;
  assign \new_[20276]_  = \new_[20275]_  & \new_[20270]_ ;
  assign \new_[20279]_  = ~A168 & ~A170;
  assign \new_[20283]_  = ~A265 & A200;
  assign \new_[20284]_  = A199 & \new_[20283]_ ;
  assign \new_[20285]_  = \new_[20284]_  & \new_[20279]_ ;
  assign \new_[20289]_  = ~A268 & ~A267;
  assign \new_[20290]_  = A266 & \new_[20289]_ ;
  assign \new_[20294]_  = ~A299 & ~A298;
  assign \new_[20295]_  = ~A269 & \new_[20294]_ ;
  assign \new_[20296]_  = \new_[20295]_  & \new_[20290]_ ;
  assign \new_[20299]_  = ~A168 & ~A170;
  assign \new_[20303]_  = A265 & A200;
  assign \new_[20304]_  = A199 & \new_[20303]_ ;
  assign \new_[20305]_  = \new_[20304]_  & \new_[20299]_ ;
  assign \new_[20309]_  = A268 & A267;
  assign \new_[20310]_  = ~A266 & \new_[20309]_ ;
  assign \new_[20314]_  = ~A302 & ~A301;
  assign \new_[20315]_  = A300 & \new_[20314]_ ;
  assign \new_[20316]_  = \new_[20315]_  & \new_[20310]_ ;
  assign \new_[20319]_  = ~A168 & ~A170;
  assign \new_[20323]_  = A265 & A200;
  assign \new_[20324]_  = A199 & \new_[20323]_ ;
  assign \new_[20325]_  = \new_[20324]_  & \new_[20319]_ ;
  assign \new_[20329]_  = A269 & A267;
  assign \new_[20330]_  = ~A266 & \new_[20329]_ ;
  assign \new_[20334]_  = ~A302 & ~A301;
  assign \new_[20335]_  = A300 & \new_[20334]_ ;
  assign \new_[20336]_  = \new_[20335]_  & \new_[20330]_ ;
  assign \new_[20339]_  = ~A168 & ~A170;
  assign \new_[20343]_  = A265 & A200;
  assign \new_[20344]_  = A199 & \new_[20343]_ ;
  assign \new_[20345]_  = \new_[20344]_  & \new_[20339]_ ;
  assign \new_[20349]_  = ~A268 & ~A267;
  assign \new_[20350]_  = ~A266 & \new_[20349]_ ;
  assign \new_[20354]_  = A301 & ~A300;
  assign \new_[20355]_  = ~A269 & \new_[20354]_ ;
  assign \new_[20356]_  = \new_[20355]_  & \new_[20350]_ ;
  assign \new_[20359]_  = ~A168 & ~A170;
  assign \new_[20363]_  = A265 & A200;
  assign \new_[20364]_  = A199 & \new_[20363]_ ;
  assign \new_[20365]_  = \new_[20364]_  & \new_[20359]_ ;
  assign \new_[20369]_  = ~A268 & ~A267;
  assign \new_[20370]_  = ~A266 & \new_[20369]_ ;
  assign \new_[20374]_  = A302 & ~A300;
  assign \new_[20375]_  = ~A269 & \new_[20374]_ ;
  assign \new_[20376]_  = \new_[20375]_  & \new_[20370]_ ;
  assign \new_[20379]_  = ~A168 & ~A170;
  assign \new_[20383]_  = A265 & A200;
  assign \new_[20384]_  = A199 & \new_[20383]_ ;
  assign \new_[20385]_  = \new_[20384]_  & \new_[20379]_ ;
  assign \new_[20389]_  = ~A268 & ~A267;
  assign \new_[20390]_  = ~A266 & \new_[20389]_ ;
  assign \new_[20394]_  = A299 & A298;
  assign \new_[20395]_  = ~A269 & \new_[20394]_ ;
  assign \new_[20396]_  = \new_[20395]_  & \new_[20390]_ ;
  assign \new_[20399]_  = ~A168 & ~A170;
  assign \new_[20403]_  = A265 & A200;
  assign \new_[20404]_  = A199 & \new_[20403]_ ;
  assign \new_[20405]_  = \new_[20404]_  & \new_[20399]_ ;
  assign \new_[20409]_  = ~A268 & ~A267;
  assign \new_[20410]_  = ~A266 & \new_[20409]_ ;
  assign \new_[20414]_  = ~A299 & ~A298;
  assign \new_[20415]_  = ~A269 & \new_[20414]_ ;
  assign \new_[20416]_  = \new_[20415]_  & \new_[20410]_ ;
  assign \new_[20419]_  = ~A168 & ~A170;
  assign \new_[20423]_  = ~A265 & ~A200;
  assign \new_[20424]_  = ~A199 & \new_[20423]_ ;
  assign \new_[20425]_  = \new_[20424]_  & \new_[20419]_ ;
  assign \new_[20429]_  = A268 & A267;
  assign \new_[20430]_  = A266 & \new_[20429]_ ;
  assign \new_[20434]_  = ~A302 & ~A301;
  assign \new_[20435]_  = A300 & \new_[20434]_ ;
  assign \new_[20436]_  = \new_[20435]_  & \new_[20430]_ ;
  assign \new_[20439]_  = ~A168 & ~A170;
  assign \new_[20443]_  = ~A265 & ~A200;
  assign \new_[20444]_  = ~A199 & \new_[20443]_ ;
  assign \new_[20445]_  = \new_[20444]_  & \new_[20439]_ ;
  assign \new_[20449]_  = A269 & A267;
  assign \new_[20450]_  = A266 & \new_[20449]_ ;
  assign \new_[20454]_  = ~A302 & ~A301;
  assign \new_[20455]_  = A300 & \new_[20454]_ ;
  assign \new_[20456]_  = \new_[20455]_  & \new_[20450]_ ;
  assign \new_[20459]_  = ~A168 & ~A170;
  assign \new_[20463]_  = ~A265 & ~A200;
  assign \new_[20464]_  = ~A199 & \new_[20463]_ ;
  assign \new_[20465]_  = \new_[20464]_  & \new_[20459]_ ;
  assign \new_[20469]_  = ~A268 & ~A267;
  assign \new_[20470]_  = A266 & \new_[20469]_ ;
  assign \new_[20474]_  = A301 & ~A300;
  assign \new_[20475]_  = ~A269 & \new_[20474]_ ;
  assign \new_[20476]_  = \new_[20475]_  & \new_[20470]_ ;
  assign \new_[20479]_  = ~A168 & ~A170;
  assign \new_[20483]_  = ~A265 & ~A200;
  assign \new_[20484]_  = ~A199 & \new_[20483]_ ;
  assign \new_[20485]_  = \new_[20484]_  & \new_[20479]_ ;
  assign \new_[20489]_  = ~A268 & ~A267;
  assign \new_[20490]_  = A266 & \new_[20489]_ ;
  assign \new_[20494]_  = A302 & ~A300;
  assign \new_[20495]_  = ~A269 & \new_[20494]_ ;
  assign \new_[20496]_  = \new_[20495]_  & \new_[20490]_ ;
  assign \new_[20499]_  = ~A168 & ~A170;
  assign \new_[20503]_  = ~A265 & ~A200;
  assign \new_[20504]_  = ~A199 & \new_[20503]_ ;
  assign \new_[20505]_  = \new_[20504]_  & \new_[20499]_ ;
  assign \new_[20509]_  = ~A268 & ~A267;
  assign \new_[20510]_  = A266 & \new_[20509]_ ;
  assign \new_[20514]_  = A299 & A298;
  assign \new_[20515]_  = ~A269 & \new_[20514]_ ;
  assign \new_[20516]_  = \new_[20515]_  & \new_[20510]_ ;
  assign \new_[20519]_  = ~A168 & ~A170;
  assign \new_[20523]_  = ~A265 & ~A200;
  assign \new_[20524]_  = ~A199 & \new_[20523]_ ;
  assign \new_[20525]_  = \new_[20524]_  & \new_[20519]_ ;
  assign \new_[20529]_  = ~A268 & ~A267;
  assign \new_[20530]_  = A266 & \new_[20529]_ ;
  assign \new_[20534]_  = ~A299 & ~A298;
  assign \new_[20535]_  = ~A269 & \new_[20534]_ ;
  assign \new_[20536]_  = \new_[20535]_  & \new_[20530]_ ;
  assign \new_[20539]_  = ~A168 & ~A170;
  assign \new_[20543]_  = A265 & ~A200;
  assign \new_[20544]_  = ~A199 & \new_[20543]_ ;
  assign \new_[20545]_  = \new_[20544]_  & \new_[20539]_ ;
  assign \new_[20549]_  = A268 & A267;
  assign \new_[20550]_  = ~A266 & \new_[20549]_ ;
  assign \new_[20554]_  = ~A302 & ~A301;
  assign \new_[20555]_  = A300 & \new_[20554]_ ;
  assign \new_[20556]_  = \new_[20555]_  & \new_[20550]_ ;
  assign \new_[20559]_  = ~A168 & ~A170;
  assign \new_[20563]_  = A265 & ~A200;
  assign \new_[20564]_  = ~A199 & \new_[20563]_ ;
  assign \new_[20565]_  = \new_[20564]_  & \new_[20559]_ ;
  assign \new_[20569]_  = A269 & A267;
  assign \new_[20570]_  = ~A266 & \new_[20569]_ ;
  assign \new_[20574]_  = ~A302 & ~A301;
  assign \new_[20575]_  = A300 & \new_[20574]_ ;
  assign \new_[20576]_  = \new_[20575]_  & \new_[20570]_ ;
  assign \new_[20579]_  = ~A168 & ~A170;
  assign \new_[20583]_  = A265 & ~A200;
  assign \new_[20584]_  = ~A199 & \new_[20583]_ ;
  assign \new_[20585]_  = \new_[20584]_  & \new_[20579]_ ;
  assign \new_[20589]_  = ~A268 & ~A267;
  assign \new_[20590]_  = ~A266 & \new_[20589]_ ;
  assign \new_[20594]_  = A301 & ~A300;
  assign \new_[20595]_  = ~A269 & \new_[20594]_ ;
  assign \new_[20596]_  = \new_[20595]_  & \new_[20590]_ ;
  assign \new_[20599]_  = ~A168 & ~A170;
  assign \new_[20603]_  = A265 & ~A200;
  assign \new_[20604]_  = ~A199 & \new_[20603]_ ;
  assign \new_[20605]_  = \new_[20604]_  & \new_[20599]_ ;
  assign \new_[20609]_  = ~A268 & ~A267;
  assign \new_[20610]_  = ~A266 & \new_[20609]_ ;
  assign \new_[20614]_  = A302 & ~A300;
  assign \new_[20615]_  = ~A269 & \new_[20614]_ ;
  assign \new_[20616]_  = \new_[20615]_  & \new_[20610]_ ;
  assign \new_[20619]_  = ~A168 & ~A170;
  assign \new_[20623]_  = A265 & ~A200;
  assign \new_[20624]_  = ~A199 & \new_[20623]_ ;
  assign \new_[20625]_  = \new_[20624]_  & \new_[20619]_ ;
  assign \new_[20629]_  = ~A268 & ~A267;
  assign \new_[20630]_  = ~A266 & \new_[20629]_ ;
  assign \new_[20634]_  = A299 & A298;
  assign \new_[20635]_  = ~A269 & \new_[20634]_ ;
  assign \new_[20636]_  = \new_[20635]_  & \new_[20630]_ ;
  assign \new_[20639]_  = ~A168 & ~A170;
  assign \new_[20643]_  = A265 & ~A200;
  assign \new_[20644]_  = ~A199 & \new_[20643]_ ;
  assign \new_[20645]_  = \new_[20644]_  & \new_[20639]_ ;
  assign \new_[20649]_  = ~A268 & ~A267;
  assign \new_[20650]_  = ~A266 & \new_[20649]_ ;
  assign \new_[20654]_  = ~A299 & ~A298;
  assign \new_[20655]_  = ~A269 & \new_[20654]_ ;
  assign \new_[20656]_  = \new_[20655]_  & \new_[20650]_ ;
  assign \new_[20659]_  = ~A168 & A169;
  assign \new_[20663]_  = ~A203 & ~A202;
  assign \new_[20664]_  = A201 & \new_[20663]_ ;
  assign \new_[20665]_  = \new_[20664]_  & \new_[20659]_ ;
  assign \new_[20669]_  = A267 & A266;
  assign \new_[20670]_  = ~A265 & \new_[20669]_ ;
  assign \new_[20674]_  = A301 & ~A300;
  assign \new_[20675]_  = A268 & \new_[20674]_ ;
  assign \new_[20676]_  = \new_[20675]_  & \new_[20670]_ ;
  assign \new_[20679]_  = ~A168 & A169;
  assign \new_[20683]_  = ~A203 & ~A202;
  assign \new_[20684]_  = A201 & \new_[20683]_ ;
  assign \new_[20685]_  = \new_[20684]_  & \new_[20679]_ ;
  assign \new_[20689]_  = A267 & A266;
  assign \new_[20690]_  = ~A265 & \new_[20689]_ ;
  assign \new_[20694]_  = A302 & ~A300;
  assign \new_[20695]_  = A268 & \new_[20694]_ ;
  assign \new_[20696]_  = \new_[20695]_  & \new_[20690]_ ;
  assign \new_[20699]_  = ~A168 & A169;
  assign \new_[20703]_  = ~A203 & ~A202;
  assign \new_[20704]_  = A201 & \new_[20703]_ ;
  assign \new_[20705]_  = \new_[20704]_  & \new_[20699]_ ;
  assign \new_[20709]_  = A267 & A266;
  assign \new_[20710]_  = ~A265 & \new_[20709]_ ;
  assign \new_[20714]_  = A299 & A298;
  assign \new_[20715]_  = A268 & \new_[20714]_ ;
  assign \new_[20716]_  = \new_[20715]_  & \new_[20710]_ ;
  assign \new_[20719]_  = ~A168 & A169;
  assign \new_[20723]_  = ~A203 & ~A202;
  assign \new_[20724]_  = A201 & \new_[20723]_ ;
  assign \new_[20725]_  = \new_[20724]_  & \new_[20719]_ ;
  assign \new_[20729]_  = A267 & A266;
  assign \new_[20730]_  = ~A265 & \new_[20729]_ ;
  assign \new_[20734]_  = ~A299 & ~A298;
  assign \new_[20735]_  = A268 & \new_[20734]_ ;
  assign \new_[20736]_  = \new_[20735]_  & \new_[20730]_ ;
  assign \new_[20739]_  = ~A168 & A169;
  assign \new_[20743]_  = ~A203 & ~A202;
  assign \new_[20744]_  = A201 & \new_[20743]_ ;
  assign \new_[20745]_  = \new_[20744]_  & \new_[20739]_ ;
  assign \new_[20749]_  = A267 & A266;
  assign \new_[20750]_  = ~A265 & \new_[20749]_ ;
  assign \new_[20754]_  = A301 & ~A300;
  assign \new_[20755]_  = A269 & \new_[20754]_ ;
  assign \new_[20756]_  = \new_[20755]_  & \new_[20750]_ ;
  assign \new_[20759]_  = ~A168 & A169;
  assign \new_[20763]_  = ~A203 & ~A202;
  assign \new_[20764]_  = A201 & \new_[20763]_ ;
  assign \new_[20765]_  = \new_[20764]_  & \new_[20759]_ ;
  assign \new_[20769]_  = A267 & A266;
  assign \new_[20770]_  = ~A265 & \new_[20769]_ ;
  assign \new_[20774]_  = A302 & ~A300;
  assign \new_[20775]_  = A269 & \new_[20774]_ ;
  assign \new_[20776]_  = \new_[20775]_  & \new_[20770]_ ;
  assign \new_[20779]_  = ~A168 & A169;
  assign \new_[20783]_  = ~A203 & ~A202;
  assign \new_[20784]_  = A201 & \new_[20783]_ ;
  assign \new_[20785]_  = \new_[20784]_  & \new_[20779]_ ;
  assign \new_[20789]_  = A267 & A266;
  assign \new_[20790]_  = ~A265 & \new_[20789]_ ;
  assign \new_[20794]_  = A299 & A298;
  assign \new_[20795]_  = A269 & \new_[20794]_ ;
  assign \new_[20796]_  = \new_[20795]_  & \new_[20790]_ ;
  assign \new_[20799]_  = ~A168 & A169;
  assign \new_[20803]_  = ~A203 & ~A202;
  assign \new_[20804]_  = A201 & \new_[20803]_ ;
  assign \new_[20805]_  = \new_[20804]_  & \new_[20799]_ ;
  assign \new_[20809]_  = A267 & A266;
  assign \new_[20810]_  = ~A265 & \new_[20809]_ ;
  assign \new_[20814]_  = ~A299 & ~A298;
  assign \new_[20815]_  = A269 & \new_[20814]_ ;
  assign \new_[20816]_  = \new_[20815]_  & \new_[20810]_ ;
  assign \new_[20819]_  = ~A168 & A169;
  assign \new_[20823]_  = ~A203 & ~A202;
  assign \new_[20824]_  = A201 & \new_[20823]_ ;
  assign \new_[20825]_  = \new_[20824]_  & \new_[20819]_ ;
  assign \new_[20829]_  = A267 & ~A266;
  assign \new_[20830]_  = A265 & \new_[20829]_ ;
  assign \new_[20834]_  = A301 & ~A300;
  assign \new_[20835]_  = A268 & \new_[20834]_ ;
  assign \new_[20836]_  = \new_[20835]_  & \new_[20830]_ ;
  assign \new_[20839]_  = ~A168 & A169;
  assign \new_[20843]_  = ~A203 & ~A202;
  assign \new_[20844]_  = A201 & \new_[20843]_ ;
  assign \new_[20845]_  = \new_[20844]_  & \new_[20839]_ ;
  assign \new_[20849]_  = A267 & ~A266;
  assign \new_[20850]_  = A265 & \new_[20849]_ ;
  assign \new_[20854]_  = A302 & ~A300;
  assign \new_[20855]_  = A268 & \new_[20854]_ ;
  assign \new_[20856]_  = \new_[20855]_  & \new_[20850]_ ;
  assign \new_[20859]_  = ~A168 & A169;
  assign \new_[20863]_  = ~A203 & ~A202;
  assign \new_[20864]_  = A201 & \new_[20863]_ ;
  assign \new_[20865]_  = \new_[20864]_  & \new_[20859]_ ;
  assign \new_[20869]_  = A267 & ~A266;
  assign \new_[20870]_  = A265 & \new_[20869]_ ;
  assign \new_[20874]_  = A299 & A298;
  assign \new_[20875]_  = A268 & \new_[20874]_ ;
  assign \new_[20876]_  = \new_[20875]_  & \new_[20870]_ ;
  assign \new_[20879]_  = ~A168 & A169;
  assign \new_[20883]_  = ~A203 & ~A202;
  assign \new_[20884]_  = A201 & \new_[20883]_ ;
  assign \new_[20885]_  = \new_[20884]_  & \new_[20879]_ ;
  assign \new_[20889]_  = A267 & ~A266;
  assign \new_[20890]_  = A265 & \new_[20889]_ ;
  assign \new_[20894]_  = ~A299 & ~A298;
  assign \new_[20895]_  = A268 & \new_[20894]_ ;
  assign \new_[20896]_  = \new_[20895]_  & \new_[20890]_ ;
  assign \new_[20899]_  = ~A168 & A169;
  assign \new_[20903]_  = ~A203 & ~A202;
  assign \new_[20904]_  = A201 & \new_[20903]_ ;
  assign \new_[20905]_  = \new_[20904]_  & \new_[20899]_ ;
  assign \new_[20909]_  = A267 & ~A266;
  assign \new_[20910]_  = A265 & \new_[20909]_ ;
  assign \new_[20914]_  = A301 & ~A300;
  assign \new_[20915]_  = A269 & \new_[20914]_ ;
  assign \new_[20916]_  = \new_[20915]_  & \new_[20910]_ ;
  assign \new_[20919]_  = ~A168 & A169;
  assign \new_[20923]_  = ~A203 & ~A202;
  assign \new_[20924]_  = A201 & \new_[20923]_ ;
  assign \new_[20925]_  = \new_[20924]_  & \new_[20919]_ ;
  assign \new_[20929]_  = A267 & ~A266;
  assign \new_[20930]_  = A265 & \new_[20929]_ ;
  assign \new_[20934]_  = A302 & ~A300;
  assign \new_[20935]_  = A269 & \new_[20934]_ ;
  assign \new_[20936]_  = \new_[20935]_  & \new_[20930]_ ;
  assign \new_[20939]_  = ~A168 & A169;
  assign \new_[20943]_  = ~A203 & ~A202;
  assign \new_[20944]_  = A201 & \new_[20943]_ ;
  assign \new_[20945]_  = \new_[20944]_  & \new_[20939]_ ;
  assign \new_[20949]_  = A267 & ~A266;
  assign \new_[20950]_  = A265 & \new_[20949]_ ;
  assign \new_[20954]_  = A299 & A298;
  assign \new_[20955]_  = A269 & \new_[20954]_ ;
  assign \new_[20956]_  = \new_[20955]_  & \new_[20950]_ ;
  assign \new_[20959]_  = ~A168 & A169;
  assign \new_[20963]_  = ~A203 & ~A202;
  assign \new_[20964]_  = A201 & \new_[20963]_ ;
  assign \new_[20965]_  = \new_[20964]_  & \new_[20959]_ ;
  assign \new_[20969]_  = A267 & ~A266;
  assign \new_[20970]_  = A265 & \new_[20969]_ ;
  assign \new_[20974]_  = ~A299 & ~A298;
  assign \new_[20975]_  = A269 & \new_[20974]_ ;
  assign \new_[20976]_  = \new_[20975]_  & \new_[20970]_ ;
  assign \new_[20979]_  = ~A168 & A169;
  assign \new_[20983]_  = ~A265 & A202;
  assign \new_[20984]_  = ~A201 & \new_[20983]_ ;
  assign \new_[20985]_  = \new_[20984]_  & \new_[20979]_ ;
  assign \new_[20989]_  = A268 & A267;
  assign \new_[20990]_  = A266 & \new_[20989]_ ;
  assign \new_[20994]_  = ~A302 & ~A301;
  assign \new_[20995]_  = A300 & \new_[20994]_ ;
  assign \new_[20996]_  = \new_[20995]_  & \new_[20990]_ ;
  assign \new_[20999]_  = ~A168 & A169;
  assign \new_[21003]_  = ~A265 & A202;
  assign \new_[21004]_  = ~A201 & \new_[21003]_ ;
  assign \new_[21005]_  = \new_[21004]_  & \new_[20999]_ ;
  assign \new_[21009]_  = A269 & A267;
  assign \new_[21010]_  = A266 & \new_[21009]_ ;
  assign \new_[21014]_  = ~A302 & ~A301;
  assign \new_[21015]_  = A300 & \new_[21014]_ ;
  assign \new_[21016]_  = \new_[21015]_  & \new_[21010]_ ;
  assign \new_[21019]_  = ~A168 & A169;
  assign \new_[21023]_  = ~A265 & A202;
  assign \new_[21024]_  = ~A201 & \new_[21023]_ ;
  assign \new_[21025]_  = \new_[21024]_  & \new_[21019]_ ;
  assign \new_[21029]_  = ~A268 & ~A267;
  assign \new_[21030]_  = A266 & \new_[21029]_ ;
  assign \new_[21034]_  = A301 & ~A300;
  assign \new_[21035]_  = ~A269 & \new_[21034]_ ;
  assign \new_[21036]_  = \new_[21035]_  & \new_[21030]_ ;
  assign \new_[21039]_  = ~A168 & A169;
  assign \new_[21043]_  = ~A265 & A202;
  assign \new_[21044]_  = ~A201 & \new_[21043]_ ;
  assign \new_[21045]_  = \new_[21044]_  & \new_[21039]_ ;
  assign \new_[21049]_  = ~A268 & ~A267;
  assign \new_[21050]_  = A266 & \new_[21049]_ ;
  assign \new_[21054]_  = A302 & ~A300;
  assign \new_[21055]_  = ~A269 & \new_[21054]_ ;
  assign \new_[21056]_  = \new_[21055]_  & \new_[21050]_ ;
  assign \new_[21059]_  = ~A168 & A169;
  assign \new_[21063]_  = ~A265 & A202;
  assign \new_[21064]_  = ~A201 & \new_[21063]_ ;
  assign \new_[21065]_  = \new_[21064]_  & \new_[21059]_ ;
  assign \new_[21069]_  = ~A268 & ~A267;
  assign \new_[21070]_  = A266 & \new_[21069]_ ;
  assign \new_[21074]_  = A299 & A298;
  assign \new_[21075]_  = ~A269 & \new_[21074]_ ;
  assign \new_[21076]_  = \new_[21075]_  & \new_[21070]_ ;
  assign \new_[21079]_  = ~A168 & A169;
  assign \new_[21083]_  = ~A265 & A202;
  assign \new_[21084]_  = ~A201 & \new_[21083]_ ;
  assign \new_[21085]_  = \new_[21084]_  & \new_[21079]_ ;
  assign \new_[21089]_  = ~A268 & ~A267;
  assign \new_[21090]_  = A266 & \new_[21089]_ ;
  assign \new_[21094]_  = ~A299 & ~A298;
  assign \new_[21095]_  = ~A269 & \new_[21094]_ ;
  assign \new_[21096]_  = \new_[21095]_  & \new_[21090]_ ;
  assign \new_[21099]_  = ~A168 & A169;
  assign \new_[21103]_  = A265 & A202;
  assign \new_[21104]_  = ~A201 & \new_[21103]_ ;
  assign \new_[21105]_  = \new_[21104]_  & \new_[21099]_ ;
  assign \new_[21109]_  = A268 & A267;
  assign \new_[21110]_  = ~A266 & \new_[21109]_ ;
  assign \new_[21114]_  = ~A302 & ~A301;
  assign \new_[21115]_  = A300 & \new_[21114]_ ;
  assign \new_[21116]_  = \new_[21115]_  & \new_[21110]_ ;
  assign \new_[21119]_  = ~A168 & A169;
  assign \new_[21123]_  = A265 & A202;
  assign \new_[21124]_  = ~A201 & \new_[21123]_ ;
  assign \new_[21125]_  = \new_[21124]_  & \new_[21119]_ ;
  assign \new_[21129]_  = A269 & A267;
  assign \new_[21130]_  = ~A266 & \new_[21129]_ ;
  assign \new_[21134]_  = ~A302 & ~A301;
  assign \new_[21135]_  = A300 & \new_[21134]_ ;
  assign \new_[21136]_  = \new_[21135]_  & \new_[21130]_ ;
  assign \new_[21139]_  = ~A168 & A169;
  assign \new_[21143]_  = A265 & A202;
  assign \new_[21144]_  = ~A201 & \new_[21143]_ ;
  assign \new_[21145]_  = \new_[21144]_  & \new_[21139]_ ;
  assign \new_[21149]_  = ~A268 & ~A267;
  assign \new_[21150]_  = ~A266 & \new_[21149]_ ;
  assign \new_[21154]_  = A301 & ~A300;
  assign \new_[21155]_  = ~A269 & \new_[21154]_ ;
  assign \new_[21156]_  = \new_[21155]_  & \new_[21150]_ ;
  assign \new_[21159]_  = ~A168 & A169;
  assign \new_[21163]_  = A265 & A202;
  assign \new_[21164]_  = ~A201 & \new_[21163]_ ;
  assign \new_[21165]_  = \new_[21164]_  & \new_[21159]_ ;
  assign \new_[21169]_  = ~A268 & ~A267;
  assign \new_[21170]_  = ~A266 & \new_[21169]_ ;
  assign \new_[21174]_  = A302 & ~A300;
  assign \new_[21175]_  = ~A269 & \new_[21174]_ ;
  assign \new_[21176]_  = \new_[21175]_  & \new_[21170]_ ;
  assign \new_[21179]_  = ~A168 & A169;
  assign \new_[21183]_  = A265 & A202;
  assign \new_[21184]_  = ~A201 & \new_[21183]_ ;
  assign \new_[21185]_  = \new_[21184]_  & \new_[21179]_ ;
  assign \new_[21189]_  = ~A268 & ~A267;
  assign \new_[21190]_  = ~A266 & \new_[21189]_ ;
  assign \new_[21194]_  = A299 & A298;
  assign \new_[21195]_  = ~A269 & \new_[21194]_ ;
  assign \new_[21196]_  = \new_[21195]_  & \new_[21190]_ ;
  assign \new_[21199]_  = ~A168 & A169;
  assign \new_[21203]_  = A265 & A202;
  assign \new_[21204]_  = ~A201 & \new_[21203]_ ;
  assign \new_[21205]_  = \new_[21204]_  & \new_[21199]_ ;
  assign \new_[21209]_  = ~A268 & ~A267;
  assign \new_[21210]_  = ~A266 & \new_[21209]_ ;
  assign \new_[21214]_  = ~A299 & ~A298;
  assign \new_[21215]_  = ~A269 & \new_[21214]_ ;
  assign \new_[21216]_  = \new_[21215]_  & \new_[21210]_ ;
  assign \new_[21219]_  = ~A168 & A169;
  assign \new_[21223]_  = ~A265 & A203;
  assign \new_[21224]_  = ~A201 & \new_[21223]_ ;
  assign \new_[21225]_  = \new_[21224]_  & \new_[21219]_ ;
  assign \new_[21229]_  = A268 & A267;
  assign \new_[21230]_  = A266 & \new_[21229]_ ;
  assign \new_[21234]_  = ~A302 & ~A301;
  assign \new_[21235]_  = A300 & \new_[21234]_ ;
  assign \new_[21236]_  = \new_[21235]_  & \new_[21230]_ ;
  assign \new_[21239]_  = ~A168 & A169;
  assign \new_[21243]_  = ~A265 & A203;
  assign \new_[21244]_  = ~A201 & \new_[21243]_ ;
  assign \new_[21245]_  = \new_[21244]_  & \new_[21239]_ ;
  assign \new_[21249]_  = A269 & A267;
  assign \new_[21250]_  = A266 & \new_[21249]_ ;
  assign \new_[21254]_  = ~A302 & ~A301;
  assign \new_[21255]_  = A300 & \new_[21254]_ ;
  assign \new_[21256]_  = \new_[21255]_  & \new_[21250]_ ;
  assign \new_[21259]_  = ~A168 & A169;
  assign \new_[21263]_  = ~A265 & A203;
  assign \new_[21264]_  = ~A201 & \new_[21263]_ ;
  assign \new_[21265]_  = \new_[21264]_  & \new_[21259]_ ;
  assign \new_[21269]_  = ~A268 & ~A267;
  assign \new_[21270]_  = A266 & \new_[21269]_ ;
  assign \new_[21274]_  = A301 & ~A300;
  assign \new_[21275]_  = ~A269 & \new_[21274]_ ;
  assign \new_[21276]_  = \new_[21275]_  & \new_[21270]_ ;
  assign \new_[21279]_  = ~A168 & A169;
  assign \new_[21283]_  = ~A265 & A203;
  assign \new_[21284]_  = ~A201 & \new_[21283]_ ;
  assign \new_[21285]_  = \new_[21284]_  & \new_[21279]_ ;
  assign \new_[21289]_  = ~A268 & ~A267;
  assign \new_[21290]_  = A266 & \new_[21289]_ ;
  assign \new_[21294]_  = A302 & ~A300;
  assign \new_[21295]_  = ~A269 & \new_[21294]_ ;
  assign \new_[21296]_  = \new_[21295]_  & \new_[21290]_ ;
  assign \new_[21299]_  = ~A168 & A169;
  assign \new_[21303]_  = ~A265 & A203;
  assign \new_[21304]_  = ~A201 & \new_[21303]_ ;
  assign \new_[21305]_  = \new_[21304]_  & \new_[21299]_ ;
  assign \new_[21309]_  = ~A268 & ~A267;
  assign \new_[21310]_  = A266 & \new_[21309]_ ;
  assign \new_[21314]_  = A299 & A298;
  assign \new_[21315]_  = ~A269 & \new_[21314]_ ;
  assign \new_[21316]_  = \new_[21315]_  & \new_[21310]_ ;
  assign \new_[21319]_  = ~A168 & A169;
  assign \new_[21323]_  = ~A265 & A203;
  assign \new_[21324]_  = ~A201 & \new_[21323]_ ;
  assign \new_[21325]_  = \new_[21324]_  & \new_[21319]_ ;
  assign \new_[21329]_  = ~A268 & ~A267;
  assign \new_[21330]_  = A266 & \new_[21329]_ ;
  assign \new_[21334]_  = ~A299 & ~A298;
  assign \new_[21335]_  = ~A269 & \new_[21334]_ ;
  assign \new_[21336]_  = \new_[21335]_  & \new_[21330]_ ;
  assign \new_[21339]_  = ~A168 & A169;
  assign \new_[21343]_  = A265 & A203;
  assign \new_[21344]_  = ~A201 & \new_[21343]_ ;
  assign \new_[21345]_  = \new_[21344]_  & \new_[21339]_ ;
  assign \new_[21349]_  = A268 & A267;
  assign \new_[21350]_  = ~A266 & \new_[21349]_ ;
  assign \new_[21354]_  = ~A302 & ~A301;
  assign \new_[21355]_  = A300 & \new_[21354]_ ;
  assign \new_[21356]_  = \new_[21355]_  & \new_[21350]_ ;
  assign \new_[21359]_  = ~A168 & A169;
  assign \new_[21363]_  = A265 & A203;
  assign \new_[21364]_  = ~A201 & \new_[21363]_ ;
  assign \new_[21365]_  = \new_[21364]_  & \new_[21359]_ ;
  assign \new_[21369]_  = A269 & A267;
  assign \new_[21370]_  = ~A266 & \new_[21369]_ ;
  assign \new_[21374]_  = ~A302 & ~A301;
  assign \new_[21375]_  = A300 & \new_[21374]_ ;
  assign \new_[21376]_  = \new_[21375]_  & \new_[21370]_ ;
  assign \new_[21379]_  = ~A168 & A169;
  assign \new_[21383]_  = A265 & A203;
  assign \new_[21384]_  = ~A201 & \new_[21383]_ ;
  assign \new_[21385]_  = \new_[21384]_  & \new_[21379]_ ;
  assign \new_[21389]_  = ~A268 & ~A267;
  assign \new_[21390]_  = ~A266 & \new_[21389]_ ;
  assign \new_[21394]_  = A301 & ~A300;
  assign \new_[21395]_  = ~A269 & \new_[21394]_ ;
  assign \new_[21396]_  = \new_[21395]_  & \new_[21390]_ ;
  assign \new_[21399]_  = ~A168 & A169;
  assign \new_[21403]_  = A265 & A203;
  assign \new_[21404]_  = ~A201 & \new_[21403]_ ;
  assign \new_[21405]_  = \new_[21404]_  & \new_[21399]_ ;
  assign \new_[21409]_  = ~A268 & ~A267;
  assign \new_[21410]_  = ~A266 & \new_[21409]_ ;
  assign \new_[21414]_  = A302 & ~A300;
  assign \new_[21415]_  = ~A269 & \new_[21414]_ ;
  assign \new_[21416]_  = \new_[21415]_  & \new_[21410]_ ;
  assign \new_[21419]_  = ~A168 & A169;
  assign \new_[21423]_  = A265 & A203;
  assign \new_[21424]_  = ~A201 & \new_[21423]_ ;
  assign \new_[21425]_  = \new_[21424]_  & \new_[21419]_ ;
  assign \new_[21429]_  = ~A268 & ~A267;
  assign \new_[21430]_  = ~A266 & \new_[21429]_ ;
  assign \new_[21434]_  = A299 & A298;
  assign \new_[21435]_  = ~A269 & \new_[21434]_ ;
  assign \new_[21436]_  = \new_[21435]_  & \new_[21430]_ ;
  assign \new_[21439]_  = ~A168 & A169;
  assign \new_[21443]_  = A265 & A203;
  assign \new_[21444]_  = ~A201 & \new_[21443]_ ;
  assign \new_[21445]_  = \new_[21444]_  & \new_[21439]_ ;
  assign \new_[21449]_  = ~A268 & ~A267;
  assign \new_[21450]_  = ~A266 & \new_[21449]_ ;
  assign \new_[21454]_  = ~A299 & ~A298;
  assign \new_[21455]_  = ~A269 & \new_[21454]_ ;
  assign \new_[21456]_  = \new_[21455]_  & \new_[21450]_ ;
  assign \new_[21459]_  = ~A168 & A169;
  assign \new_[21463]_  = ~A265 & A200;
  assign \new_[21464]_  = A199 & \new_[21463]_ ;
  assign \new_[21465]_  = \new_[21464]_  & \new_[21459]_ ;
  assign \new_[21469]_  = A268 & A267;
  assign \new_[21470]_  = A266 & \new_[21469]_ ;
  assign \new_[21474]_  = ~A302 & ~A301;
  assign \new_[21475]_  = A300 & \new_[21474]_ ;
  assign \new_[21476]_  = \new_[21475]_  & \new_[21470]_ ;
  assign \new_[21479]_  = ~A168 & A169;
  assign \new_[21483]_  = ~A265 & A200;
  assign \new_[21484]_  = A199 & \new_[21483]_ ;
  assign \new_[21485]_  = \new_[21484]_  & \new_[21479]_ ;
  assign \new_[21489]_  = A269 & A267;
  assign \new_[21490]_  = A266 & \new_[21489]_ ;
  assign \new_[21494]_  = ~A302 & ~A301;
  assign \new_[21495]_  = A300 & \new_[21494]_ ;
  assign \new_[21496]_  = \new_[21495]_  & \new_[21490]_ ;
  assign \new_[21499]_  = ~A168 & A169;
  assign \new_[21503]_  = ~A265 & A200;
  assign \new_[21504]_  = A199 & \new_[21503]_ ;
  assign \new_[21505]_  = \new_[21504]_  & \new_[21499]_ ;
  assign \new_[21509]_  = ~A268 & ~A267;
  assign \new_[21510]_  = A266 & \new_[21509]_ ;
  assign \new_[21514]_  = A301 & ~A300;
  assign \new_[21515]_  = ~A269 & \new_[21514]_ ;
  assign \new_[21516]_  = \new_[21515]_  & \new_[21510]_ ;
  assign \new_[21519]_  = ~A168 & A169;
  assign \new_[21523]_  = ~A265 & A200;
  assign \new_[21524]_  = A199 & \new_[21523]_ ;
  assign \new_[21525]_  = \new_[21524]_  & \new_[21519]_ ;
  assign \new_[21529]_  = ~A268 & ~A267;
  assign \new_[21530]_  = A266 & \new_[21529]_ ;
  assign \new_[21534]_  = A302 & ~A300;
  assign \new_[21535]_  = ~A269 & \new_[21534]_ ;
  assign \new_[21536]_  = \new_[21535]_  & \new_[21530]_ ;
  assign \new_[21539]_  = ~A168 & A169;
  assign \new_[21543]_  = ~A265 & A200;
  assign \new_[21544]_  = A199 & \new_[21543]_ ;
  assign \new_[21545]_  = \new_[21544]_  & \new_[21539]_ ;
  assign \new_[21549]_  = ~A268 & ~A267;
  assign \new_[21550]_  = A266 & \new_[21549]_ ;
  assign \new_[21554]_  = A299 & A298;
  assign \new_[21555]_  = ~A269 & \new_[21554]_ ;
  assign \new_[21556]_  = \new_[21555]_  & \new_[21550]_ ;
  assign \new_[21559]_  = ~A168 & A169;
  assign \new_[21563]_  = ~A265 & A200;
  assign \new_[21564]_  = A199 & \new_[21563]_ ;
  assign \new_[21565]_  = \new_[21564]_  & \new_[21559]_ ;
  assign \new_[21569]_  = ~A268 & ~A267;
  assign \new_[21570]_  = A266 & \new_[21569]_ ;
  assign \new_[21574]_  = ~A299 & ~A298;
  assign \new_[21575]_  = ~A269 & \new_[21574]_ ;
  assign \new_[21576]_  = \new_[21575]_  & \new_[21570]_ ;
  assign \new_[21579]_  = ~A168 & A169;
  assign \new_[21583]_  = A265 & A200;
  assign \new_[21584]_  = A199 & \new_[21583]_ ;
  assign \new_[21585]_  = \new_[21584]_  & \new_[21579]_ ;
  assign \new_[21589]_  = A268 & A267;
  assign \new_[21590]_  = ~A266 & \new_[21589]_ ;
  assign \new_[21594]_  = ~A302 & ~A301;
  assign \new_[21595]_  = A300 & \new_[21594]_ ;
  assign \new_[21596]_  = \new_[21595]_  & \new_[21590]_ ;
  assign \new_[21599]_  = ~A168 & A169;
  assign \new_[21603]_  = A265 & A200;
  assign \new_[21604]_  = A199 & \new_[21603]_ ;
  assign \new_[21605]_  = \new_[21604]_  & \new_[21599]_ ;
  assign \new_[21609]_  = A269 & A267;
  assign \new_[21610]_  = ~A266 & \new_[21609]_ ;
  assign \new_[21614]_  = ~A302 & ~A301;
  assign \new_[21615]_  = A300 & \new_[21614]_ ;
  assign \new_[21616]_  = \new_[21615]_  & \new_[21610]_ ;
  assign \new_[21619]_  = ~A168 & A169;
  assign \new_[21623]_  = A265 & A200;
  assign \new_[21624]_  = A199 & \new_[21623]_ ;
  assign \new_[21625]_  = \new_[21624]_  & \new_[21619]_ ;
  assign \new_[21629]_  = ~A268 & ~A267;
  assign \new_[21630]_  = ~A266 & \new_[21629]_ ;
  assign \new_[21634]_  = A301 & ~A300;
  assign \new_[21635]_  = ~A269 & \new_[21634]_ ;
  assign \new_[21636]_  = \new_[21635]_  & \new_[21630]_ ;
  assign \new_[21639]_  = ~A168 & A169;
  assign \new_[21643]_  = A265 & A200;
  assign \new_[21644]_  = A199 & \new_[21643]_ ;
  assign \new_[21645]_  = \new_[21644]_  & \new_[21639]_ ;
  assign \new_[21649]_  = ~A268 & ~A267;
  assign \new_[21650]_  = ~A266 & \new_[21649]_ ;
  assign \new_[21654]_  = A302 & ~A300;
  assign \new_[21655]_  = ~A269 & \new_[21654]_ ;
  assign \new_[21656]_  = \new_[21655]_  & \new_[21650]_ ;
  assign \new_[21659]_  = ~A168 & A169;
  assign \new_[21663]_  = A265 & A200;
  assign \new_[21664]_  = A199 & \new_[21663]_ ;
  assign \new_[21665]_  = \new_[21664]_  & \new_[21659]_ ;
  assign \new_[21669]_  = ~A268 & ~A267;
  assign \new_[21670]_  = ~A266 & \new_[21669]_ ;
  assign \new_[21674]_  = A299 & A298;
  assign \new_[21675]_  = ~A269 & \new_[21674]_ ;
  assign \new_[21676]_  = \new_[21675]_  & \new_[21670]_ ;
  assign \new_[21679]_  = ~A168 & A169;
  assign \new_[21683]_  = A265 & A200;
  assign \new_[21684]_  = A199 & \new_[21683]_ ;
  assign \new_[21685]_  = \new_[21684]_  & \new_[21679]_ ;
  assign \new_[21689]_  = ~A268 & ~A267;
  assign \new_[21690]_  = ~A266 & \new_[21689]_ ;
  assign \new_[21694]_  = ~A299 & ~A298;
  assign \new_[21695]_  = ~A269 & \new_[21694]_ ;
  assign \new_[21696]_  = \new_[21695]_  & \new_[21690]_ ;
  assign \new_[21699]_  = ~A168 & A169;
  assign \new_[21703]_  = ~A265 & ~A200;
  assign \new_[21704]_  = ~A199 & \new_[21703]_ ;
  assign \new_[21705]_  = \new_[21704]_  & \new_[21699]_ ;
  assign \new_[21709]_  = A268 & A267;
  assign \new_[21710]_  = A266 & \new_[21709]_ ;
  assign \new_[21714]_  = ~A302 & ~A301;
  assign \new_[21715]_  = A300 & \new_[21714]_ ;
  assign \new_[21716]_  = \new_[21715]_  & \new_[21710]_ ;
  assign \new_[21719]_  = ~A168 & A169;
  assign \new_[21723]_  = ~A265 & ~A200;
  assign \new_[21724]_  = ~A199 & \new_[21723]_ ;
  assign \new_[21725]_  = \new_[21724]_  & \new_[21719]_ ;
  assign \new_[21729]_  = A269 & A267;
  assign \new_[21730]_  = A266 & \new_[21729]_ ;
  assign \new_[21734]_  = ~A302 & ~A301;
  assign \new_[21735]_  = A300 & \new_[21734]_ ;
  assign \new_[21736]_  = \new_[21735]_  & \new_[21730]_ ;
  assign \new_[21739]_  = ~A168 & A169;
  assign \new_[21743]_  = ~A265 & ~A200;
  assign \new_[21744]_  = ~A199 & \new_[21743]_ ;
  assign \new_[21745]_  = \new_[21744]_  & \new_[21739]_ ;
  assign \new_[21749]_  = ~A268 & ~A267;
  assign \new_[21750]_  = A266 & \new_[21749]_ ;
  assign \new_[21754]_  = A301 & ~A300;
  assign \new_[21755]_  = ~A269 & \new_[21754]_ ;
  assign \new_[21756]_  = \new_[21755]_  & \new_[21750]_ ;
  assign \new_[21759]_  = ~A168 & A169;
  assign \new_[21763]_  = ~A265 & ~A200;
  assign \new_[21764]_  = ~A199 & \new_[21763]_ ;
  assign \new_[21765]_  = \new_[21764]_  & \new_[21759]_ ;
  assign \new_[21769]_  = ~A268 & ~A267;
  assign \new_[21770]_  = A266 & \new_[21769]_ ;
  assign \new_[21774]_  = A302 & ~A300;
  assign \new_[21775]_  = ~A269 & \new_[21774]_ ;
  assign \new_[21776]_  = \new_[21775]_  & \new_[21770]_ ;
  assign \new_[21779]_  = ~A168 & A169;
  assign \new_[21783]_  = ~A265 & ~A200;
  assign \new_[21784]_  = ~A199 & \new_[21783]_ ;
  assign \new_[21785]_  = \new_[21784]_  & \new_[21779]_ ;
  assign \new_[21789]_  = ~A268 & ~A267;
  assign \new_[21790]_  = A266 & \new_[21789]_ ;
  assign \new_[21794]_  = A299 & A298;
  assign \new_[21795]_  = ~A269 & \new_[21794]_ ;
  assign \new_[21796]_  = \new_[21795]_  & \new_[21790]_ ;
  assign \new_[21799]_  = ~A168 & A169;
  assign \new_[21803]_  = ~A265 & ~A200;
  assign \new_[21804]_  = ~A199 & \new_[21803]_ ;
  assign \new_[21805]_  = \new_[21804]_  & \new_[21799]_ ;
  assign \new_[21809]_  = ~A268 & ~A267;
  assign \new_[21810]_  = A266 & \new_[21809]_ ;
  assign \new_[21814]_  = ~A299 & ~A298;
  assign \new_[21815]_  = ~A269 & \new_[21814]_ ;
  assign \new_[21816]_  = \new_[21815]_  & \new_[21810]_ ;
  assign \new_[21819]_  = ~A168 & A169;
  assign \new_[21823]_  = A265 & ~A200;
  assign \new_[21824]_  = ~A199 & \new_[21823]_ ;
  assign \new_[21825]_  = \new_[21824]_  & \new_[21819]_ ;
  assign \new_[21829]_  = A268 & A267;
  assign \new_[21830]_  = ~A266 & \new_[21829]_ ;
  assign \new_[21834]_  = ~A302 & ~A301;
  assign \new_[21835]_  = A300 & \new_[21834]_ ;
  assign \new_[21836]_  = \new_[21835]_  & \new_[21830]_ ;
  assign \new_[21839]_  = ~A168 & A169;
  assign \new_[21843]_  = A265 & ~A200;
  assign \new_[21844]_  = ~A199 & \new_[21843]_ ;
  assign \new_[21845]_  = \new_[21844]_  & \new_[21839]_ ;
  assign \new_[21849]_  = A269 & A267;
  assign \new_[21850]_  = ~A266 & \new_[21849]_ ;
  assign \new_[21854]_  = ~A302 & ~A301;
  assign \new_[21855]_  = A300 & \new_[21854]_ ;
  assign \new_[21856]_  = \new_[21855]_  & \new_[21850]_ ;
  assign \new_[21859]_  = ~A168 & A169;
  assign \new_[21863]_  = A265 & ~A200;
  assign \new_[21864]_  = ~A199 & \new_[21863]_ ;
  assign \new_[21865]_  = \new_[21864]_  & \new_[21859]_ ;
  assign \new_[21869]_  = ~A268 & ~A267;
  assign \new_[21870]_  = ~A266 & \new_[21869]_ ;
  assign \new_[21874]_  = A301 & ~A300;
  assign \new_[21875]_  = ~A269 & \new_[21874]_ ;
  assign \new_[21876]_  = \new_[21875]_  & \new_[21870]_ ;
  assign \new_[21879]_  = ~A168 & A169;
  assign \new_[21883]_  = A265 & ~A200;
  assign \new_[21884]_  = ~A199 & \new_[21883]_ ;
  assign \new_[21885]_  = \new_[21884]_  & \new_[21879]_ ;
  assign \new_[21889]_  = ~A268 & ~A267;
  assign \new_[21890]_  = ~A266 & \new_[21889]_ ;
  assign \new_[21894]_  = A302 & ~A300;
  assign \new_[21895]_  = ~A269 & \new_[21894]_ ;
  assign \new_[21896]_  = \new_[21895]_  & \new_[21890]_ ;
  assign \new_[21899]_  = ~A168 & A169;
  assign \new_[21903]_  = A265 & ~A200;
  assign \new_[21904]_  = ~A199 & \new_[21903]_ ;
  assign \new_[21905]_  = \new_[21904]_  & \new_[21899]_ ;
  assign \new_[21909]_  = ~A268 & ~A267;
  assign \new_[21910]_  = ~A266 & \new_[21909]_ ;
  assign \new_[21914]_  = A299 & A298;
  assign \new_[21915]_  = ~A269 & \new_[21914]_ ;
  assign \new_[21916]_  = \new_[21915]_  & \new_[21910]_ ;
  assign \new_[21919]_  = ~A168 & A169;
  assign \new_[21923]_  = A265 & ~A200;
  assign \new_[21924]_  = ~A199 & \new_[21923]_ ;
  assign \new_[21925]_  = \new_[21924]_  & \new_[21919]_ ;
  assign \new_[21929]_  = ~A268 & ~A267;
  assign \new_[21930]_  = ~A266 & \new_[21929]_ ;
  assign \new_[21934]_  = ~A299 & ~A298;
  assign \new_[21935]_  = ~A269 & \new_[21934]_ ;
  assign \new_[21936]_  = \new_[21935]_  & \new_[21930]_ ;
  assign \new_[21939]_  = ~A169 & A170;
  assign \new_[21943]_  = A202 & ~A201;
  assign \new_[21944]_  = A168 & \new_[21943]_ ;
  assign \new_[21945]_  = \new_[21944]_  & \new_[21939]_ ;
  assign \new_[21949]_  = A267 & A266;
  assign \new_[21950]_  = ~A265 & \new_[21949]_ ;
  assign \new_[21954]_  = A301 & ~A300;
  assign \new_[21955]_  = A268 & \new_[21954]_ ;
  assign \new_[21956]_  = \new_[21955]_  & \new_[21950]_ ;
  assign \new_[21959]_  = ~A169 & A170;
  assign \new_[21963]_  = A202 & ~A201;
  assign \new_[21964]_  = A168 & \new_[21963]_ ;
  assign \new_[21965]_  = \new_[21964]_  & \new_[21959]_ ;
  assign \new_[21969]_  = A267 & A266;
  assign \new_[21970]_  = ~A265 & \new_[21969]_ ;
  assign \new_[21974]_  = A302 & ~A300;
  assign \new_[21975]_  = A268 & \new_[21974]_ ;
  assign \new_[21976]_  = \new_[21975]_  & \new_[21970]_ ;
  assign \new_[21979]_  = ~A169 & A170;
  assign \new_[21983]_  = A202 & ~A201;
  assign \new_[21984]_  = A168 & \new_[21983]_ ;
  assign \new_[21985]_  = \new_[21984]_  & \new_[21979]_ ;
  assign \new_[21989]_  = A267 & A266;
  assign \new_[21990]_  = ~A265 & \new_[21989]_ ;
  assign \new_[21994]_  = A299 & A298;
  assign \new_[21995]_  = A268 & \new_[21994]_ ;
  assign \new_[21996]_  = \new_[21995]_  & \new_[21990]_ ;
  assign \new_[21999]_  = ~A169 & A170;
  assign \new_[22003]_  = A202 & ~A201;
  assign \new_[22004]_  = A168 & \new_[22003]_ ;
  assign \new_[22005]_  = \new_[22004]_  & \new_[21999]_ ;
  assign \new_[22009]_  = A267 & A266;
  assign \new_[22010]_  = ~A265 & \new_[22009]_ ;
  assign \new_[22014]_  = ~A299 & ~A298;
  assign \new_[22015]_  = A268 & \new_[22014]_ ;
  assign \new_[22016]_  = \new_[22015]_  & \new_[22010]_ ;
  assign \new_[22019]_  = ~A169 & A170;
  assign \new_[22023]_  = A202 & ~A201;
  assign \new_[22024]_  = A168 & \new_[22023]_ ;
  assign \new_[22025]_  = \new_[22024]_  & \new_[22019]_ ;
  assign \new_[22029]_  = A267 & A266;
  assign \new_[22030]_  = ~A265 & \new_[22029]_ ;
  assign \new_[22034]_  = A301 & ~A300;
  assign \new_[22035]_  = A269 & \new_[22034]_ ;
  assign \new_[22036]_  = \new_[22035]_  & \new_[22030]_ ;
  assign \new_[22039]_  = ~A169 & A170;
  assign \new_[22043]_  = A202 & ~A201;
  assign \new_[22044]_  = A168 & \new_[22043]_ ;
  assign \new_[22045]_  = \new_[22044]_  & \new_[22039]_ ;
  assign \new_[22049]_  = A267 & A266;
  assign \new_[22050]_  = ~A265 & \new_[22049]_ ;
  assign \new_[22054]_  = A302 & ~A300;
  assign \new_[22055]_  = A269 & \new_[22054]_ ;
  assign \new_[22056]_  = \new_[22055]_  & \new_[22050]_ ;
  assign \new_[22059]_  = ~A169 & A170;
  assign \new_[22063]_  = A202 & ~A201;
  assign \new_[22064]_  = A168 & \new_[22063]_ ;
  assign \new_[22065]_  = \new_[22064]_  & \new_[22059]_ ;
  assign \new_[22069]_  = A267 & A266;
  assign \new_[22070]_  = ~A265 & \new_[22069]_ ;
  assign \new_[22074]_  = A299 & A298;
  assign \new_[22075]_  = A269 & \new_[22074]_ ;
  assign \new_[22076]_  = \new_[22075]_  & \new_[22070]_ ;
  assign \new_[22079]_  = ~A169 & A170;
  assign \new_[22083]_  = A202 & ~A201;
  assign \new_[22084]_  = A168 & \new_[22083]_ ;
  assign \new_[22085]_  = \new_[22084]_  & \new_[22079]_ ;
  assign \new_[22089]_  = A267 & A266;
  assign \new_[22090]_  = ~A265 & \new_[22089]_ ;
  assign \new_[22094]_  = ~A299 & ~A298;
  assign \new_[22095]_  = A269 & \new_[22094]_ ;
  assign \new_[22096]_  = \new_[22095]_  & \new_[22090]_ ;
  assign \new_[22099]_  = ~A169 & A170;
  assign \new_[22103]_  = A202 & ~A201;
  assign \new_[22104]_  = A168 & \new_[22103]_ ;
  assign \new_[22105]_  = \new_[22104]_  & \new_[22099]_ ;
  assign \new_[22109]_  = A267 & ~A266;
  assign \new_[22110]_  = A265 & \new_[22109]_ ;
  assign \new_[22114]_  = A301 & ~A300;
  assign \new_[22115]_  = A268 & \new_[22114]_ ;
  assign \new_[22116]_  = \new_[22115]_  & \new_[22110]_ ;
  assign \new_[22119]_  = ~A169 & A170;
  assign \new_[22123]_  = A202 & ~A201;
  assign \new_[22124]_  = A168 & \new_[22123]_ ;
  assign \new_[22125]_  = \new_[22124]_  & \new_[22119]_ ;
  assign \new_[22129]_  = A267 & ~A266;
  assign \new_[22130]_  = A265 & \new_[22129]_ ;
  assign \new_[22134]_  = A302 & ~A300;
  assign \new_[22135]_  = A268 & \new_[22134]_ ;
  assign \new_[22136]_  = \new_[22135]_  & \new_[22130]_ ;
  assign \new_[22139]_  = ~A169 & A170;
  assign \new_[22143]_  = A202 & ~A201;
  assign \new_[22144]_  = A168 & \new_[22143]_ ;
  assign \new_[22145]_  = \new_[22144]_  & \new_[22139]_ ;
  assign \new_[22149]_  = A267 & ~A266;
  assign \new_[22150]_  = A265 & \new_[22149]_ ;
  assign \new_[22154]_  = A299 & A298;
  assign \new_[22155]_  = A268 & \new_[22154]_ ;
  assign \new_[22156]_  = \new_[22155]_  & \new_[22150]_ ;
  assign \new_[22159]_  = ~A169 & A170;
  assign \new_[22163]_  = A202 & ~A201;
  assign \new_[22164]_  = A168 & \new_[22163]_ ;
  assign \new_[22165]_  = \new_[22164]_  & \new_[22159]_ ;
  assign \new_[22169]_  = A267 & ~A266;
  assign \new_[22170]_  = A265 & \new_[22169]_ ;
  assign \new_[22174]_  = ~A299 & ~A298;
  assign \new_[22175]_  = A268 & \new_[22174]_ ;
  assign \new_[22176]_  = \new_[22175]_  & \new_[22170]_ ;
  assign \new_[22179]_  = ~A169 & A170;
  assign \new_[22183]_  = A202 & ~A201;
  assign \new_[22184]_  = A168 & \new_[22183]_ ;
  assign \new_[22185]_  = \new_[22184]_  & \new_[22179]_ ;
  assign \new_[22189]_  = A267 & ~A266;
  assign \new_[22190]_  = A265 & \new_[22189]_ ;
  assign \new_[22194]_  = A301 & ~A300;
  assign \new_[22195]_  = A269 & \new_[22194]_ ;
  assign \new_[22196]_  = \new_[22195]_  & \new_[22190]_ ;
  assign \new_[22199]_  = ~A169 & A170;
  assign \new_[22203]_  = A202 & ~A201;
  assign \new_[22204]_  = A168 & \new_[22203]_ ;
  assign \new_[22205]_  = \new_[22204]_  & \new_[22199]_ ;
  assign \new_[22209]_  = A267 & ~A266;
  assign \new_[22210]_  = A265 & \new_[22209]_ ;
  assign \new_[22214]_  = A302 & ~A300;
  assign \new_[22215]_  = A269 & \new_[22214]_ ;
  assign \new_[22216]_  = \new_[22215]_  & \new_[22210]_ ;
  assign \new_[22219]_  = ~A169 & A170;
  assign \new_[22223]_  = A202 & ~A201;
  assign \new_[22224]_  = A168 & \new_[22223]_ ;
  assign \new_[22225]_  = \new_[22224]_  & \new_[22219]_ ;
  assign \new_[22229]_  = A267 & ~A266;
  assign \new_[22230]_  = A265 & \new_[22229]_ ;
  assign \new_[22234]_  = A299 & A298;
  assign \new_[22235]_  = A269 & \new_[22234]_ ;
  assign \new_[22236]_  = \new_[22235]_  & \new_[22230]_ ;
  assign \new_[22239]_  = ~A169 & A170;
  assign \new_[22243]_  = A202 & ~A201;
  assign \new_[22244]_  = A168 & \new_[22243]_ ;
  assign \new_[22245]_  = \new_[22244]_  & \new_[22239]_ ;
  assign \new_[22249]_  = A267 & ~A266;
  assign \new_[22250]_  = A265 & \new_[22249]_ ;
  assign \new_[22254]_  = ~A299 & ~A298;
  assign \new_[22255]_  = A269 & \new_[22254]_ ;
  assign \new_[22256]_  = \new_[22255]_  & \new_[22250]_ ;
  assign \new_[22259]_  = ~A169 & A170;
  assign \new_[22263]_  = A203 & ~A201;
  assign \new_[22264]_  = A168 & \new_[22263]_ ;
  assign \new_[22265]_  = \new_[22264]_  & \new_[22259]_ ;
  assign \new_[22269]_  = A267 & A266;
  assign \new_[22270]_  = ~A265 & \new_[22269]_ ;
  assign \new_[22274]_  = A301 & ~A300;
  assign \new_[22275]_  = A268 & \new_[22274]_ ;
  assign \new_[22276]_  = \new_[22275]_  & \new_[22270]_ ;
  assign \new_[22279]_  = ~A169 & A170;
  assign \new_[22283]_  = A203 & ~A201;
  assign \new_[22284]_  = A168 & \new_[22283]_ ;
  assign \new_[22285]_  = \new_[22284]_  & \new_[22279]_ ;
  assign \new_[22289]_  = A267 & A266;
  assign \new_[22290]_  = ~A265 & \new_[22289]_ ;
  assign \new_[22294]_  = A302 & ~A300;
  assign \new_[22295]_  = A268 & \new_[22294]_ ;
  assign \new_[22296]_  = \new_[22295]_  & \new_[22290]_ ;
  assign \new_[22299]_  = ~A169 & A170;
  assign \new_[22303]_  = A203 & ~A201;
  assign \new_[22304]_  = A168 & \new_[22303]_ ;
  assign \new_[22305]_  = \new_[22304]_  & \new_[22299]_ ;
  assign \new_[22309]_  = A267 & A266;
  assign \new_[22310]_  = ~A265 & \new_[22309]_ ;
  assign \new_[22314]_  = A299 & A298;
  assign \new_[22315]_  = A268 & \new_[22314]_ ;
  assign \new_[22316]_  = \new_[22315]_  & \new_[22310]_ ;
  assign \new_[22319]_  = ~A169 & A170;
  assign \new_[22323]_  = A203 & ~A201;
  assign \new_[22324]_  = A168 & \new_[22323]_ ;
  assign \new_[22325]_  = \new_[22324]_  & \new_[22319]_ ;
  assign \new_[22329]_  = A267 & A266;
  assign \new_[22330]_  = ~A265 & \new_[22329]_ ;
  assign \new_[22334]_  = ~A299 & ~A298;
  assign \new_[22335]_  = A268 & \new_[22334]_ ;
  assign \new_[22336]_  = \new_[22335]_  & \new_[22330]_ ;
  assign \new_[22339]_  = ~A169 & A170;
  assign \new_[22343]_  = A203 & ~A201;
  assign \new_[22344]_  = A168 & \new_[22343]_ ;
  assign \new_[22345]_  = \new_[22344]_  & \new_[22339]_ ;
  assign \new_[22349]_  = A267 & A266;
  assign \new_[22350]_  = ~A265 & \new_[22349]_ ;
  assign \new_[22354]_  = A301 & ~A300;
  assign \new_[22355]_  = A269 & \new_[22354]_ ;
  assign \new_[22356]_  = \new_[22355]_  & \new_[22350]_ ;
  assign \new_[22359]_  = ~A169 & A170;
  assign \new_[22363]_  = A203 & ~A201;
  assign \new_[22364]_  = A168 & \new_[22363]_ ;
  assign \new_[22365]_  = \new_[22364]_  & \new_[22359]_ ;
  assign \new_[22369]_  = A267 & A266;
  assign \new_[22370]_  = ~A265 & \new_[22369]_ ;
  assign \new_[22374]_  = A302 & ~A300;
  assign \new_[22375]_  = A269 & \new_[22374]_ ;
  assign \new_[22376]_  = \new_[22375]_  & \new_[22370]_ ;
  assign \new_[22379]_  = ~A169 & A170;
  assign \new_[22383]_  = A203 & ~A201;
  assign \new_[22384]_  = A168 & \new_[22383]_ ;
  assign \new_[22385]_  = \new_[22384]_  & \new_[22379]_ ;
  assign \new_[22389]_  = A267 & A266;
  assign \new_[22390]_  = ~A265 & \new_[22389]_ ;
  assign \new_[22394]_  = A299 & A298;
  assign \new_[22395]_  = A269 & \new_[22394]_ ;
  assign \new_[22396]_  = \new_[22395]_  & \new_[22390]_ ;
  assign \new_[22399]_  = ~A169 & A170;
  assign \new_[22403]_  = A203 & ~A201;
  assign \new_[22404]_  = A168 & \new_[22403]_ ;
  assign \new_[22405]_  = \new_[22404]_  & \new_[22399]_ ;
  assign \new_[22409]_  = A267 & A266;
  assign \new_[22410]_  = ~A265 & \new_[22409]_ ;
  assign \new_[22414]_  = ~A299 & ~A298;
  assign \new_[22415]_  = A269 & \new_[22414]_ ;
  assign \new_[22416]_  = \new_[22415]_  & \new_[22410]_ ;
  assign \new_[22419]_  = ~A169 & A170;
  assign \new_[22423]_  = A203 & ~A201;
  assign \new_[22424]_  = A168 & \new_[22423]_ ;
  assign \new_[22425]_  = \new_[22424]_  & \new_[22419]_ ;
  assign \new_[22429]_  = A267 & ~A266;
  assign \new_[22430]_  = A265 & \new_[22429]_ ;
  assign \new_[22434]_  = A301 & ~A300;
  assign \new_[22435]_  = A268 & \new_[22434]_ ;
  assign \new_[22436]_  = \new_[22435]_  & \new_[22430]_ ;
  assign \new_[22439]_  = ~A169 & A170;
  assign \new_[22443]_  = A203 & ~A201;
  assign \new_[22444]_  = A168 & \new_[22443]_ ;
  assign \new_[22445]_  = \new_[22444]_  & \new_[22439]_ ;
  assign \new_[22449]_  = A267 & ~A266;
  assign \new_[22450]_  = A265 & \new_[22449]_ ;
  assign \new_[22454]_  = A302 & ~A300;
  assign \new_[22455]_  = A268 & \new_[22454]_ ;
  assign \new_[22456]_  = \new_[22455]_  & \new_[22450]_ ;
  assign \new_[22459]_  = ~A169 & A170;
  assign \new_[22463]_  = A203 & ~A201;
  assign \new_[22464]_  = A168 & \new_[22463]_ ;
  assign \new_[22465]_  = \new_[22464]_  & \new_[22459]_ ;
  assign \new_[22469]_  = A267 & ~A266;
  assign \new_[22470]_  = A265 & \new_[22469]_ ;
  assign \new_[22474]_  = A299 & A298;
  assign \new_[22475]_  = A268 & \new_[22474]_ ;
  assign \new_[22476]_  = \new_[22475]_  & \new_[22470]_ ;
  assign \new_[22479]_  = ~A169 & A170;
  assign \new_[22483]_  = A203 & ~A201;
  assign \new_[22484]_  = A168 & \new_[22483]_ ;
  assign \new_[22485]_  = \new_[22484]_  & \new_[22479]_ ;
  assign \new_[22489]_  = A267 & ~A266;
  assign \new_[22490]_  = A265 & \new_[22489]_ ;
  assign \new_[22494]_  = ~A299 & ~A298;
  assign \new_[22495]_  = A268 & \new_[22494]_ ;
  assign \new_[22496]_  = \new_[22495]_  & \new_[22490]_ ;
  assign \new_[22499]_  = ~A169 & A170;
  assign \new_[22503]_  = A203 & ~A201;
  assign \new_[22504]_  = A168 & \new_[22503]_ ;
  assign \new_[22505]_  = \new_[22504]_  & \new_[22499]_ ;
  assign \new_[22509]_  = A267 & ~A266;
  assign \new_[22510]_  = A265 & \new_[22509]_ ;
  assign \new_[22514]_  = A301 & ~A300;
  assign \new_[22515]_  = A269 & \new_[22514]_ ;
  assign \new_[22516]_  = \new_[22515]_  & \new_[22510]_ ;
  assign \new_[22519]_  = ~A169 & A170;
  assign \new_[22523]_  = A203 & ~A201;
  assign \new_[22524]_  = A168 & \new_[22523]_ ;
  assign \new_[22525]_  = \new_[22524]_  & \new_[22519]_ ;
  assign \new_[22529]_  = A267 & ~A266;
  assign \new_[22530]_  = A265 & \new_[22529]_ ;
  assign \new_[22534]_  = A302 & ~A300;
  assign \new_[22535]_  = A269 & \new_[22534]_ ;
  assign \new_[22536]_  = \new_[22535]_  & \new_[22530]_ ;
  assign \new_[22539]_  = ~A169 & A170;
  assign \new_[22543]_  = A203 & ~A201;
  assign \new_[22544]_  = A168 & \new_[22543]_ ;
  assign \new_[22545]_  = \new_[22544]_  & \new_[22539]_ ;
  assign \new_[22549]_  = A267 & ~A266;
  assign \new_[22550]_  = A265 & \new_[22549]_ ;
  assign \new_[22554]_  = A299 & A298;
  assign \new_[22555]_  = A269 & \new_[22554]_ ;
  assign \new_[22556]_  = \new_[22555]_  & \new_[22550]_ ;
  assign \new_[22559]_  = ~A169 & A170;
  assign \new_[22563]_  = A203 & ~A201;
  assign \new_[22564]_  = A168 & \new_[22563]_ ;
  assign \new_[22565]_  = \new_[22564]_  & \new_[22559]_ ;
  assign \new_[22569]_  = A267 & ~A266;
  assign \new_[22570]_  = A265 & \new_[22569]_ ;
  assign \new_[22574]_  = ~A299 & ~A298;
  assign \new_[22575]_  = A269 & \new_[22574]_ ;
  assign \new_[22576]_  = \new_[22575]_  & \new_[22570]_ ;
  assign \new_[22579]_  = ~A169 & A170;
  assign \new_[22583]_  = A200 & A199;
  assign \new_[22584]_  = A168 & \new_[22583]_ ;
  assign \new_[22585]_  = \new_[22584]_  & \new_[22579]_ ;
  assign \new_[22589]_  = A267 & A266;
  assign \new_[22590]_  = ~A265 & \new_[22589]_ ;
  assign \new_[22594]_  = A301 & ~A300;
  assign \new_[22595]_  = A268 & \new_[22594]_ ;
  assign \new_[22596]_  = \new_[22595]_  & \new_[22590]_ ;
  assign \new_[22599]_  = ~A169 & A170;
  assign \new_[22603]_  = A200 & A199;
  assign \new_[22604]_  = A168 & \new_[22603]_ ;
  assign \new_[22605]_  = \new_[22604]_  & \new_[22599]_ ;
  assign \new_[22609]_  = A267 & A266;
  assign \new_[22610]_  = ~A265 & \new_[22609]_ ;
  assign \new_[22614]_  = A302 & ~A300;
  assign \new_[22615]_  = A268 & \new_[22614]_ ;
  assign \new_[22616]_  = \new_[22615]_  & \new_[22610]_ ;
  assign \new_[22619]_  = ~A169 & A170;
  assign \new_[22623]_  = A200 & A199;
  assign \new_[22624]_  = A168 & \new_[22623]_ ;
  assign \new_[22625]_  = \new_[22624]_  & \new_[22619]_ ;
  assign \new_[22629]_  = A267 & A266;
  assign \new_[22630]_  = ~A265 & \new_[22629]_ ;
  assign \new_[22634]_  = A299 & A298;
  assign \new_[22635]_  = A268 & \new_[22634]_ ;
  assign \new_[22636]_  = \new_[22635]_  & \new_[22630]_ ;
  assign \new_[22639]_  = ~A169 & A170;
  assign \new_[22643]_  = A200 & A199;
  assign \new_[22644]_  = A168 & \new_[22643]_ ;
  assign \new_[22645]_  = \new_[22644]_  & \new_[22639]_ ;
  assign \new_[22649]_  = A267 & A266;
  assign \new_[22650]_  = ~A265 & \new_[22649]_ ;
  assign \new_[22654]_  = ~A299 & ~A298;
  assign \new_[22655]_  = A268 & \new_[22654]_ ;
  assign \new_[22656]_  = \new_[22655]_  & \new_[22650]_ ;
  assign \new_[22659]_  = ~A169 & A170;
  assign \new_[22663]_  = A200 & A199;
  assign \new_[22664]_  = A168 & \new_[22663]_ ;
  assign \new_[22665]_  = \new_[22664]_  & \new_[22659]_ ;
  assign \new_[22669]_  = A267 & A266;
  assign \new_[22670]_  = ~A265 & \new_[22669]_ ;
  assign \new_[22674]_  = A301 & ~A300;
  assign \new_[22675]_  = A269 & \new_[22674]_ ;
  assign \new_[22676]_  = \new_[22675]_  & \new_[22670]_ ;
  assign \new_[22679]_  = ~A169 & A170;
  assign \new_[22683]_  = A200 & A199;
  assign \new_[22684]_  = A168 & \new_[22683]_ ;
  assign \new_[22685]_  = \new_[22684]_  & \new_[22679]_ ;
  assign \new_[22689]_  = A267 & A266;
  assign \new_[22690]_  = ~A265 & \new_[22689]_ ;
  assign \new_[22694]_  = A302 & ~A300;
  assign \new_[22695]_  = A269 & \new_[22694]_ ;
  assign \new_[22696]_  = \new_[22695]_  & \new_[22690]_ ;
  assign \new_[22699]_  = ~A169 & A170;
  assign \new_[22703]_  = A200 & A199;
  assign \new_[22704]_  = A168 & \new_[22703]_ ;
  assign \new_[22705]_  = \new_[22704]_  & \new_[22699]_ ;
  assign \new_[22709]_  = A267 & A266;
  assign \new_[22710]_  = ~A265 & \new_[22709]_ ;
  assign \new_[22714]_  = A299 & A298;
  assign \new_[22715]_  = A269 & \new_[22714]_ ;
  assign \new_[22716]_  = \new_[22715]_  & \new_[22710]_ ;
  assign \new_[22719]_  = ~A169 & A170;
  assign \new_[22723]_  = A200 & A199;
  assign \new_[22724]_  = A168 & \new_[22723]_ ;
  assign \new_[22725]_  = \new_[22724]_  & \new_[22719]_ ;
  assign \new_[22729]_  = A267 & A266;
  assign \new_[22730]_  = ~A265 & \new_[22729]_ ;
  assign \new_[22734]_  = ~A299 & ~A298;
  assign \new_[22735]_  = A269 & \new_[22734]_ ;
  assign \new_[22736]_  = \new_[22735]_  & \new_[22730]_ ;
  assign \new_[22739]_  = ~A169 & A170;
  assign \new_[22743]_  = A200 & A199;
  assign \new_[22744]_  = A168 & \new_[22743]_ ;
  assign \new_[22745]_  = \new_[22744]_  & \new_[22739]_ ;
  assign \new_[22749]_  = A267 & ~A266;
  assign \new_[22750]_  = A265 & \new_[22749]_ ;
  assign \new_[22754]_  = A301 & ~A300;
  assign \new_[22755]_  = A268 & \new_[22754]_ ;
  assign \new_[22756]_  = \new_[22755]_  & \new_[22750]_ ;
  assign \new_[22759]_  = ~A169 & A170;
  assign \new_[22763]_  = A200 & A199;
  assign \new_[22764]_  = A168 & \new_[22763]_ ;
  assign \new_[22765]_  = \new_[22764]_  & \new_[22759]_ ;
  assign \new_[22769]_  = A267 & ~A266;
  assign \new_[22770]_  = A265 & \new_[22769]_ ;
  assign \new_[22774]_  = A302 & ~A300;
  assign \new_[22775]_  = A268 & \new_[22774]_ ;
  assign \new_[22776]_  = \new_[22775]_  & \new_[22770]_ ;
  assign \new_[22779]_  = ~A169 & A170;
  assign \new_[22783]_  = A200 & A199;
  assign \new_[22784]_  = A168 & \new_[22783]_ ;
  assign \new_[22785]_  = \new_[22784]_  & \new_[22779]_ ;
  assign \new_[22789]_  = A267 & ~A266;
  assign \new_[22790]_  = A265 & \new_[22789]_ ;
  assign \new_[22794]_  = A299 & A298;
  assign \new_[22795]_  = A268 & \new_[22794]_ ;
  assign \new_[22796]_  = \new_[22795]_  & \new_[22790]_ ;
  assign \new_[22799]_  = ~A169 & A170;
  assign \new_[22803]_  = A200 & A199;
  assign \new_[22804]_  = A168 & \new_[22803]_ ;
  assign \new_[22805]_  = \new_[22804]_  & \new_[22799]_ ;
  assign \new_[22809]_  = A267 & ~A266;
  assign \new_[22810]_  = A265 & \new_[22809]_ ;
  assign \new_[22814]_  = ~A299 & ~A298;
  assign \new_[22815]_  = A268 & \new_[22814]_ ;
  assign \new_[22816]_  = \new_[22815]_  & \new_[22810]_ ;
  assign \new_[22819]_  = ~A169 & A170;
  assign \new_[22823]_  = A200 & A199;
  assign \new_[22824]_  = A168 & \new_[22823]_ ;
  assign \new_[22825]_  = \new_[22824]_  & \new_[22819]_ ;
  assign \new_[22829]_  = A267 & ~A266;
  assign \new_[22830]_  = A265 & \new_[22829]_ ;
  assign \new_[22834]_  = A301 & ~A300;
  assign \new_[22835]_  = A269 & \new_[22834]_ ;
  assign \new_[22836]_  = \new_[22835]_  & \new_[22830]_ ;
  assign \new_[22839]_  = ~A169 & A170;
  assign \new_[22843]_  = A200 & A199;
  assign \new_[22844]_  = A168 & \new_[22843]_ ;
  assign \new_[22845]_  = \new_[22844]_  & \new_[22839]_ ;
  assign \new_[22849]_  = A267 & ~A266;
  assign \new_[22850]_  = A265 & \new_[22849]_ ;
  assign \new_[22854]_  = A302 & ~A300;
  assign \new_[22855]_  = A269 & \new_[22854]_ ;
  assign \new_[22856]_  = \new_[22855]_  & \new_[22850]_ ;
  assign \new_[22859]_  = ~A169 & A170;
  assign \new_[22863]_  = A200 & A199;
  assign \new_[22864]_  = A168 & \new_[22863]_ ;
  assign \new_[22865]_  = \new_[22864]_  & \new_[22859]_ ;
  assign \new_[22869]_  = A267 & ~A266;
  assign \new_[22870]_  = A265 & \new_[22869]_ ;
  assign \new_[22874]_  = A299 & A298;
  assign \new_[22875]_  = A269 & \new_[22874]_ ;
  assign \new_[22876]_  = \new_[22875]_  & \new_[22870]_ ;
  assign \new_[22879]_  = ~A169 & A170;
  assign \new_[22883]_  = A200 & A199;
  assign \new_[22884]_  = A168 & \new_[22883]_ ;
  assign \new_[22885]_  = \new_[22884]_  & \new_[22879]_ ;
  assign \new_[22889]_  = A267 & ~A266;
  assign \new_[22890]_  = A265 & \new_[22889]_ ;
  assign \new_[22894]_  = ~A299 & ~A298;
  assign \new_[22895]_  = A269 & \new_[22894]_ ;
  assign \new_[22896]_  = \new_[22895]_  & \new_[22890]_ ;
  assign \new_[22899]_  = ~A169 & A170;
  assign \new_[22903]_  = ~A200 & ~A199;
  assign \new_[22904]_  = A168 & \new_[22903]_ ;
  assign \new_[22905]_  = \new_[22904]_  & \new_[22899]_ ;
  assign \new_[22909]_  = A267 & A266;
  assign \new_[22910]_  = ~A265 & \new_[22909]_ ;
  assign \new_[22914]_  = A301 & ~A300;
  assign \new_[22915]_  = A268 & \new_[22914]_ ;
  assign \new_[22916]_  = \new_[22915]_  & \new_[22910]_ ;
  assign \new_[22919]_  = ~A169 & A170;
  assign \new_[22923]_  = ~A200 & ~A199;
  assign \new_[22924]_  = A168 & \new_[22923]_ ;
  assign \new_[22925]_  = \new_[22924]_  & \new_[22919]_ ;
  assign \new_[22929]_  = A267 & A266;
  assign \new_[22930]_  = ~A265 & \new_[22929]_ ;
  assign \new_[22934]_  = A302 & ~A300;
  assign \new_[22935]_  = A268 & \new_[22934]_ ;
  assign \new_[22936]_  = \new_[22935]_  & \new_[22930]_ ;
  assign \new_[22939]_  = ~A169 & A170;
  assign \new_[22943]_  = ~A200 & ~A199;
  assign \new_[22944]_  = A168 & \new_[22943]_ ;
  assign \new_[22945]_  = \new_[22944]_  & \new_[22939]_ ;
  assign \new_[22949]_  = A267 & A266;
  assign \new_[22950]_  = ~A265 & \new_[22949]_ ;
  assign \new_[22954]_  = A299 & A298;
  assign \new_[22955]_  = A268 & \new_[22954]_ ;
  assign \new_[22956]_  = \new_[22955]_  & \new_[22950]_ ;
  assign \new_[22959]_  = ~A169 & A170;
  assign \new_[22963]_  = ~A200 & ~A199;
  assign \new_[22964]_  = A168 & \new_[22963]_ ;
  assign \new_[22965]_  = \new_[22964]_  & \new_[22959]_ ;
  assign \new_[22969]_  = A267 & A266;
  assign \new_[22970]_  = ~A265 & \new_[22969]_ ;
  assign \new_[22974]_  = ~A299 & ~A298;
  assign \new_[22975]_  = A268 & \new_[22974]_ ;
  assign \new_[22976]_  = \new_[22975]_  & \new_[22970]_ ;
  assign \new_[22979]_  = ~A169 & A170;
  assign \new_[22983]_  = ~A200 & ~A199;
  assign \new_[22984]_  = A168 & \new_[22983]_ ;
  assign \new_[22985]_  = \new_[22984]_  & \new_[22979]_ ;
  assign \new_[22989]_  = A267 & A266;
  assign \new_[22990]_  = ~A265 & \new_[22989]_ ;
  assign \new_[22994]_  = A301 & ~A300;
  assign \new_[22995]_  = A269 & \new_[22994]_ ;
  assign \new_[22996]_  = \new_[22995]_  & \new_[22990]_ ;
  assign \new_[22999]_  = ~A169 & A170;
  assign \new_[23003]_  = ~A200 & ~A199;
  assign \new_[23004]_  = A168 & \new_[23003]_ ;
  assign \new_[23005]_  = \new_[23004]_  & \new_[22999]_ ;
  assign \new_[23009]_  = A267 & A266;
  assign \new_[23010]_  = ~A265 & \new_[23009]_ ;
  assign \new_[23014]_  = A302 & ~A300;
  assign \new_[23015]_  = A269 & \new_[23014]_ ;
  assign \new_[23016]_  = \new_[23015]_  & \new_[23010]_ ;
  assign \new_[23019]_  = ~A169 & A170;
  assign \new_[23023]_  = ~A200 & ~A199;
  assign \new_[23024]_  = A168 & \new_[23023]_ ;
  assign \new_[23025]_  = \new_[23024]_  & \new_[23019]_ ;
  assign \new_[23029]_  = A267 & A266;
  assign \new_[23030]_  = ~A265 & \new_[23029]_ ;
  assign \new_[23034]_  = A299 & A298;
  assign \new_[23035]_  = A269 & \new_[23034]_ ;
  assign \new_[23036]_  = \new_[23035]_  & \new_[23030]_ ;
  assign \new_[23039]_  = ~A169 & A170;
  assign \new_[23043]_  = ~A200 & ~A199;
  assign \new_[23044]_  = A168 & \new_[23043]_ ;
  assign \new_[23045]_  = \new_[23044]_  & \new_[23039]_ ;
  assign \new_[23049]_  = A267 & A266;
  assign \new_[23050]_  = ~A265 & \new_[23049]_ ;
  assign \new_[23054]_  = ~A299 & ~A298;
  assign \new_[23055]_  = A269 & \new_[23054]_ ;
  assign \new_[23056]_  = \new_[23055]_  & \new_[23050]_ ;
  assign \new_[23059]_  = ~A169 & A170;
  assign \new_[23063]_  = ~A200 & ~A199;
  assign \new_[23064]_  = A168 & \new_[23063]_ ;
  assign \new_[23065]_  = \new_[23064]_  & \new_[23059]_ ;
  assign \new_[23069]_  = A267 & ~A266;
  assign \new_[23070]_  = A265 & \new_[23069]_ ;
  assign \new_[23074]_  = A301 & ~A300;
  assign \new_[23075]_  = A268 & \new_[23074]_ ;
  assign \new_[23076]_  = \new_[23075]_  & \new_[23070]_ ;
  assign \new_[23079]_  = ~A169 & A170;
  assign \new_[23083]_  = ~A200 & ~A199;
  assign \new_[23084]_  = A168 & \new_[23083]_ ;
  assign \new_[23085]_  = \new_[23084]_  & \new_[23079]_ ;
  assign \new_[23089]_  = A267 & ~A266;
  assign \new_[23090]_  = A265 & \new_[23089]_ ;
  assign \new_[23094]_  = A302 & ~A300;
  assign \new_[23095]_  = A268 & \new_[23094]_ ;
  assign \new_[23096]_  = \new_[23095]_  & \new_[23090]_ ;
  assign \new_[23099]_  = ~A169 & A170;
  assign \new_[23103]_  = ~A200 & ~A199;
  assign \new_[23104]_  = A168 & \new_[23103]_ ;
  assign \new_[23105]_  = \new_[23104]_  & \new_[23099]_ ;
  assign \new_[23109]_  = A267 & ~A266;
  assign \new_[23110]_  = A265 & \new_[23109]_ ;
  assign \new_[23114]_  = A299 & A298;
  assign \new_[23115]_  = A268 & \new_[23114]_ ;
  assign \new_[23116]_  = \new_[23115]_  & \new_[23110]_ ;
  assign \new_[23119]_  = ~A169 & A170;
  assign \new_[23123]_  = ~A200 & ~A199;
  assign \new_[23124]_  = A168 & \new_[23123]_ ;
  assign \new_[23125]_  = \new_[23124]_  & \new_[23119]_ ;
  assign \new_[23129]_  = A267 & ~A266;
  assign \new_[23130]_  = A265 & \new_[23129]_ ;
  assign \new_[23134]_  = ~A299 & ~A298;
  assign \new_[23135]_  = A268 & \new_[23134]_ ;
  assign \new_[23136]_  = \new_[23135]_  & \new_[23130]_ ;
  assign \new_[23139]_  = ~A169 & A170;
  assign \new_[23143]_  = ~A200 & ~A199;
  assign \new_[23144]_  = A168 & \new_[23143]_ ;
  assign \new_[23145]_  = \new_[23144]_  & \new_[23139]_ ;
  assign \new_[23149]_  = A267 & ~A266;
  assign \new_[23150]_  = A265 & \new_[23149]_ ;
  assign \new_[23154]_  = A301 & ~A300;
  assign \new_[23155]_  = A269 & \new_[23154]_ ;
  assign \new_[23156]_  = \new_[23155]_  & \new_[23150]_ ;
  assign \new_[23159]_  = ~A169 & A170;
  assign \new_[23163]_  = ~A200 & ~A199;
  assign \new_[23164]_  = A168 & \new_[23163]_ ;
  assign \new_[23165]_  = \new_[23164]_  & \new_[23159]_ ;
  assign \new_[23169]_  = A267 & ~A266;
  assign \new_[23170]_  = A265 & \new_[23169]_ ;
  assign \new_[23174]_  = A302 & ~A300;
  assign \new_[23175]_  = A269 & \new_[23174]_ ;
  assign \new_[23176]_  = \new_[23175]_  & \new_[23170]_ ;
  assign \new_[23179]_  = ~A169 & A170;
  assign \new_[23183]_  = ~A200 & ~A199;
  assign \new_[23184]_  = A168 & \new_[23183]_ ;
  assign \new_[23185]_  = \new_[23184]_  & \new_[23179]_ ;
  assign \new_[23189]_  = A267 & ~A266;
  assign \new_[23190]_  = A265 & \new_[23189]_ ;
  assign \new_[23194]_  = A299 & A298;
  assign \new_[23195]_  = A269 & \new_[23194]_ ;
  assign \new_[23196]_  = \new_[23195]_  & \new_[23190]_ ;
  assign \new_[23199]_  = ~A169 & A170;
  assign \new_[23203]_  = ~A200 & ~A199;
  assign \new_[23204]_  = A168 & \new_[23203]_ ;
  assign \new_[23205]_  = \new_[23204]_  & \new_[23199]_ ;
  assign \new_[23209]_  = A267 & ~A266;
  assign \new_[23210]_  = A265 & \new_[23209]_ ;
  assign \new_[23214]_  = ~A299 & ~A298;
  assign \new_[23215]_  = A269 & \new_[23214]_ ;
  assign \new_[23216]_  = \new_[23215]_  & \new_[23210]_ ;
  assign \new_[23220]_  = A201 & A166;
  assign \new_[23221]_  = A167 & \new_[23220]_ ;
  assign \new_[23225]_  = ~A265 & ~A203;
  assign \new_[23226]_  = ~A202 & \new_[23225]_ ;
  assign \new_[23227]_  = \new_[23226]_  & \new_[23221]_ ;
  assign \new_[23231]_  = A268 & A267;
  assign \new_[23232]_  = A266 & \new_[23231]_ ;
  assign \new_[23236]_  = ~A302 & ~A301;
  assign \new_[23237]_  = A300 & \new_[23236]_ ;
  assign \new_[23238]_  = \new_[23237]_  & \new_[23232]_ ;
  assign \new_[23242]_  = A201 & A166;
  assign \new_[23243]_  = A167 & \new_[23242]_ ;
  assign \new_[23247]_  = ~A265 & ~A203;
  assign \new_[23248]_  = ~A202 & \new_[23247]_ ;
  assign \new_[23249]_  = \new_[23248]_  & \new_[23243]_ ;
  assign \new_[23253]_  = A269 & A267;
  assign \new_[23254]_  = A266 & \new_[23253]_ ;
  assign \new_[23258]_  = ~A302 & ~A301;
  assign \new_[23259]_  = A300 & \new_[23258]_ ;
  assign \new_[23260]_  = \new_[23259]_  & \new_[23254]_ ;
  assign \new_[23264]_  = A201 & A166;
  assign \new_[23265]_  = A167 & \new_[23264]_ ;
  assign \new_[23269]_  = ~A265 & ~A203;
  assign \new_[23270]_  = ~A202 & \new_[23269]_ ;
  assign \new_[23271]_  = \new_[23270]_  & \new_[23265]_ ;
  assign \new_[23275]_  = ~A268 & ~A267;
  assign \new_[23276]_  = A266 & \new_[23275]_ ;
  assign \new_[23280]_  = A301 & ~A300;
  assign \new_[23281]_  = ~A269 & \new_[23280]_ ;
  assign \new_[23282]_  = \new_[23281]_  & \new_[23276]_ ;
  assign \new_[23286]_  = A201 & A166;
  assign \new_[23287]_  = A167 & \new_[23286]_ ;
  assign \new_[23291]_  = ~A265 & ~A203;
  assign \new_[23292]_  = ~A202 & \new_[23291]_ ;
  assign \new_[23293]_  = \new_[23292]_  & \new_[23287]_ ;
  assign \new_[23297]_  = ~A268 & ~A267;
  assign \new_[23298]_  = A266 & \new_[23297]_ ;
  assign \new_[23302]_  = A302 & ~A300;
  assign \new_[23303]_  = ~A269 & \new_[23302]_ ;
  assign \new_[23304]_  = \new_[23303]_  & \new_[23298]_ ;
  assign \new_[23308]_  = A201 & A166;
  assign \new_[23309]_  = A167 & \new_[23308]_ ;
  assign \new_[23313]_  = ~A265 & ~A203;
  assign \new_[23314]_  = ~A202 & \new_[23313]_ ;
  assign \new_[23315]_  = \new_[23314]_  & \new_[23309]_ ;
  assign \new_[23319]_  = ~A268 & ~A267;
  assign \new_[23320]_  = A266 & \new_[23319]_ ;
  assign \new_[23324]_  = A299 & A298;
  assign \new_[23325]_  = ~A269 & \new_[23324]_ ;
  assign \new_[23326]_  = \new_[23325]_  & \new_[23320]_ ;
  assign \new_[23330]_  = A201 & A166;
  assign \new_[23331]_  = A167 & \new_[23330]_ ;
  assign \new_[23335]_  = ~A265 & ~A203;
  assign \new_[23336]_  = ~A202 & \new_[23335]_ ;
  assign \new_[23337]_  = \new_[23336]_  & \new_[23331]_ ;
  assign \new_[23341]_  = ~A268 & ~A267;
  assign \new_[23342]_  = A266 & \new_[23341]_ ;
  assign \new_[23346]_  = ~A299 & ~A298;
  assign \new_[23347]_  = ~A269 & \new_[23346]_ ;
  assign \new_[23348]_  = \new_[23347]_  & \new_[23342]_ ;
  assign \new_[23352]_  = A201 & A166;
  assign \new_[23353]_  = A167 & \new_[23352]_ ;
  assign \new_[23357]_  = A265 & ~A203;
  assign \new_[23358]_  = ~A202 & \new_[23357]_ ;
  assign \new_[23359]_  = \new_[23358]_  & \new_[23353]_ ;
  assign \new_[23363]_  = A268 & A267;
  assign \new_[23364]_  = ~A266 & \new_[23363]_ ;
  assign \new_[23368]_  = ~A302 & ~A301;
  assign \new_[23369]_  = A300 & \new_[23368]_ ;
  assign \new_[23370]_  = \new_[23369]_  & \new_[23364]_ ;
  assign \new_[23374]_  = A201 & A166;
  assign \new_[23375]_  = A167 & \new_[23374]_ ;
  assign \new_[23379]_  = A265 & ~A203;
  assign \new_[23380]_  = ~A202 & \new_[23379]_ ;
  assign \new_[23381]_  = \new_[23380]_  & \new_[23375]_ ;
  assign \new_[23385]_  = A269 & A267;
  assign \new_[23386]_  = ~A266 & \new_[23385]_ ;
  assign \new_[23390]_  = ~A302 & ~A301;
  assign \new_[23391]_  = A300 & \new_[23390]_ ;
  assign \new_[23392]_  = \new_[23391]_  & \new_[23386]_ ;
  assign \new_[23396]_  = A201 & A166;
  assign \new_[23397]_  = A167 & \new_[23396]_ ;
  assign \new_[23401]_  = A265 & ~A203;
  assign \new_[23402]_  = ~A202 & \new_[23401]_ ;
  assign \new_[23403]_  = \new_[23402]_  & \new_[23397]_ ;
  assign \new_[23407]_  = ~A268 & ~A267;
  assign \new_[23408]_  = ~A266 & \new_[23407]_ ;
  assign \new_[23412]_  = A301 & ~A300;
  assign \new_[23413]_  = ~A269 & \new_[23412]_ ;
  assign \new_[23414]_  = \new_[23413]_  & \new_[23408]_ ;
  assign \new_[23418]_  = A201 & A166;
  assign \new_[23419]_  = A167 & \new_[23418]_ ;
  assign \new_[23423]_  = A265 & ~A203;
  assign \new_[23424]_  = ~A202 & \new_[23423]_ ;
  assign \new_[23425]_  = \new_[23424]_  & \new_[23419]_ ;
  assign \new_[23429]_  = ~A268 & ~A267;
  assign \new_[23430]_  = ~A266 & \new_[23429]_ ;
  assign \new_[23434]_  = A302 & ~A300;
  assign \new_[23435]_  = ~A269 & \new_[23434]_ ;
  assign \new_[23436]_  = \new_[23435]_  & \new_[23430]_ ;
  assign \new_[23440]_  = A201 & A166;
  assign \new_[23441]_  = A167 & \new_[23440]_ ;
  assign \new_[23445]_  = A265 & ~A203;
  assign \new_[23446]_  = ~A202 & \new_[23445]_ ;
  assign \new_[23447]_  = \new_[23446]_  & \new_[23441]_ ;
  assign \new_[23451]_  = ~A268 & ~A267;
  assign \new_[23452]_  = ~A266 & \new_[23451]_ ;
  assign \new_[23456]_  = A299 & A298;
  assign \new_[23457]_  = ~A269 & \new_[23456]_ ;
  assign \new_[23458]_  = \new_[23457]_  & \new_[23452]_ ;
  assign \new_[23462]_  = A201 & A166;
  assign \new_[23463]_  = A167 & \new_[23462]_ ;
  assign \new_[23467]_  = A265 & ~A203;
  assign \new_[23468]_  = ~A202 & \new_[23467]_ ;
  assign \new_[23469]_  = \new_[23468]_  & \new_[23463]_ ;
  assign \new_[23473]_  = ~A268 & ~A267;
  assign \new_[23474]_  = ~A266 & \new_[23473]_ ;
  assign \new_[23478]_  = ~A299 & ~A298;
  assign \new_[23479]_  = ~A269 & \new_[23478]_ ;
  assign \new_[23480]_  = \new_[23479]_  & \new_[23474]_ ;
  assign \new_[23484]_  = ~A201 & A166;
  assign \new_[23485]_  = A167 & \new_[23484]_ ;
  assign \new_[23489]_  = A266 & ~A265;
  assign \new_[23490]_  = A202 & \new_[23489]_ ;
  assign \new_[23491]_  = \new_[23490]_  & \new_[23485]_ ;
  assign \new_[23495]_  = ~A269 & ~A268;
  assign \new_[23496]_  = ~A267 & \new_[23495]_ ;
  assign \new_[23500]_  = ~A302 & ~A301;
  assign \new_[23501]_  = A300 & \new_[23500]_ ;
  assign \new_[23502]_  = \new_[23501]_  & \new_[23496]_ ;
  assign \new_[23506]_  = ~A201 & A166;
  assign \new_[23507]_  = A167 & \new_[23506]_ ;
  assign \new_[23511]_  = ~A266 & A265;
  assign \new_[23512]_  = A202 & \new_[23511]_ ;
  assign \new_[23513]_  = \new_[23512]_  & \new_[23507]_ ;
  assign \new_[23517]_  = ~A269 & ~A268;
  assign \new_[23518]_  = ~A267 & \new_[23517]_ ;
  assign \new_[23522]_  = ~A302 & ~A301;
  assign \new_[23523]_  = A300 & \new_[23522]_ ;
  assign \new_[23524]_  = \new_[23523]_  & \new_[23518]_ ;
  assign \new_[23528]_  = ~A201 & A166;
  assign \new_[23529]_  = A167 & \new_[23528]_ ;
  assign \new_[23533]_  = A266 & ~A265;
  assign \new_[23534]_  = A203 & \new_[23533]_ ;
  assign \new_[23535]_  = \new_[23534]_  & \new_[23529]_ ;
  assign \new_[23539]_  = ~A269 & ~A268;
  assign \new_[23540]_  = ~A267 & \new_[23539]_ ;
  assign \new_[23544]_  = ~A302 & ~A301;
  assign \new_[23545]_  = A300 & \new_[23544]_ ;
  assign \new_[23546]_  = \new_[23545]_  & \new_[23540]_ ;
  assign \new_[23550]_  = ~A201 & A166;
  assign \new_[23551]_  = A167 & \new_[23550]_ ;
  assign \new_[23555]_  = ~A266 & A265;
  assign \new_[23556]_  = A203 & \new_[23555]_ ;
  assign \new_[23557]_  = \new_[23556]_  & \new_[23551]_ ;
  assign \new_[23561]_  = ~A269 & ~A268;
  assign \new_[23562]_  = ~A267 & \new_[23561]_ ;
  assign \new_[23566]_  = ~A302 & ~A301;
  assign \new_[23567]_  = A300 & \new_[23566]_ ;
  assign \new_[23568]_  = \new_[23567]_  & \new_[23562]_ ;
  assign \new_[23572]_  = A199 & A166;
  assign \new_[23573]_  = A167 & \new_[23572]_ ;
  assign \new_[23577]_  = A266 & ~A265;
  assign \new_[23578]_  = A200 & \new_[23577]_ ;
  assign \new_[23579]_  = \new_[23578]_  & \new_[23573]_ ;
  assign \new_[23583]_  = ~A269 & ~A268;
  assign \new_[23584]_  = ~A267 & \new_[23583]_ ;
  assign \new_[23588]_  = ~A302 & ~A301;
  assign \new_[23589]_  = A300 & \new_[23588]_ ;
  assign \new_[23590]_  = \new_[23589]_  & \new_[23584]_ ;
  assign \new_[23594]_  = A199 & A166;
  assign \new_[23595]_  = A167 & \new_[23594]_ ;
  assign \new_[23599]_  = ~A266 & A265;
  assign \new_[23600]_  = A200 & \new_[23599]_ ;
  assign \new_[23601]_  = \new_[23600]_  & \new_[23595]_ ;
  assign \new_[23605]_  = ~A269 & ~A268;
  assign \new_[23606]_  = ~A267 & \new_[23605]_ ;
  assign \new_[23610]_  = ~A302 & ~A301;
  assign \new_[23611]_  = A300 & \new_[23610]_ ;
  assign \new_[23612]_  = \new_[23611]_  & \new_[23606]_ ;
  assign \new_[23616]_  = ~A199 & A166;
  assign \new_[23617]_  = A167 & \new_[23616]_ ;
  assign \new_[23621]_  = A202 & A201;
  assign \new_[23622]_  = A200 & \new_[23621]_ ;
  assign \new_[23623]_  = \new_[23622]_  & \new_[23617]_ ;
  assign \new_[23627]_  = A298 & A268;
  assign \new_[23628]_  = ~A267 & \new_[23627]_ ;
  assign \new_[23632]_  = A301 & A300;
  assign \new_[23633]_  = ~A299 & \new_[23632]_ ;
  assign \new_[23634]_  = \new_[23633]_  & \new_[23628]_ ;
  assign \new_[23638]_  = ~A199 & A166;
  assign \new_[23639]_  = A167 & \new_[23638]_ ;
  assign \new_[23643]_  = A202 & A201;
  assign \new_[23644]_  = A200 & \new_[23643]_ ;
  assign \new_[23645]_  = \new_[23644]_  & \new_[23639]_ ;
  assign \new_[23649]_  = A298 & A268;
  assign \new_[23650]_  = ~A267 & \new_[23649]_ ;
  assign \new_[23654]_  = A302 & A300;
  assign \new_[23655]_  = ~A299 & \new_[23654]_ ;
  assign \new_[23656]_  = \new_[23655]_  & \new_[23650]_ ;
  assign \new_[23660]_  = ~A199 & A166;
  assign \new_[23661]_  = A167 & \new_[23660]_ ;
  assign \new_[23665]_  = A202 & A201;
  assign \new_[23666]_  = A200 & \new_[23665]_ ;
  assign \new_[23667]_  = \new_[23666]_  & \new_[23661]_ ;
  assign \new_[23671]_  = ~A298 & A268;
  assign \new_[23672]_  = ~A267 & \new_[23671]_ ;
  assign \new_[23676]_  = A301 & A300;
  assign \new_[23677]_  = A299 & \new_[23676]_ ;
  assign \new_[23678]_  = \new_[23677]_  & \new_[23672]_ ;
  assign \new_[23682]_  = ~A199 & A166;
  assign \new_[23683]_  = A167 & \new_[23682]_ ;
  assign \new_[23687]_  = A202 & A201;
  assign \new_[23688]_  = A200 & \new_[23687]_ ;
  assign \new_[23689]_  = \new_[23688]_  & \new_[23683]_ ;
  assign \new_[23693]_  = ~A298 & A268;
  assign \new_[23694]_  = ~A267 & \new_[23693]_ ;
  assign \new_[23698]_  = A302 & A300;
  assign \new_[23699]_  = A299 & \new_[23698]_ ;
  assign \new_[23700]_  = \new_[23699]_  & \new_[23694]_ ;
  assign \new_[23704]_  = ~A199 & A166;
  assign \new_[23705]_  = A167 & \new_[23704]_ ;
  assign \new_[23709]_  = A202 & A201;
  assign \new_[23710]_  = A200 & \new_[23709]_ ;
  assign \new_[23711]_  = \new_[23710]_  & \new_[23705]_ ;
  assign \new_[23715]_  = A298 & A269;
  assign \new_[23716]_  = ~A267 & \new_[23715]_ ;
  assign \new_[23720]_  = A301 & A300;
  assign \new_[23721]_  = ~A299 & \new_[23720]_ ;
  assign \new_[23722]_  = \new_[23721]_  & \new_[23716]_ ;
  assign \new_[23726]_  = ~A199 & A166;
  assign \new_[23727]_  = A167 & \new_[23726]_ ;
  assign \new_[23731]_  = A202 & A201;
  assign \new_[23732]_  = A200 & \new_[23731]_ ;
  assign \new_[23733]_  = \new_[23732]_  & \new_[23727]_ ;
  assign \new_[23737]_  = A298 & A269;
  assign \new_[23738]_  = ~A267 & \new_[23737]_ ;
  assign \new_[23742]_  = A302 & A300;
  assign \new_[23743]_  = ~A299 & \new_[23742]_ ;
  assign \new_[23744]_  = \new_[23743]_  & \new_[23738]_ ;
  assign \new_[23748]_  = ~A199 & A166;
  assign \new_[23749]_  = A167 & \new_[23748]_ ;
  assign \new_[23753]_  = A202 & A201;
  assign \new_[23754]_  = A200 & \new_[23753]_ ;
  assign \new_[23755]_  = \new_[23754]_  & \new_[23749]_ ;
  assign \new_[23759]_  = ~A298 & A269;
  assign \new_[23760]_  = ~A267 & \new_[23759]_ ;
  assign \new_[23764]_  = A301 & A300;
  assign \new_[23765]_  = A299 & \new_[23764]_ ;
  assign \new_[23766]_  = \new_[23765]_  & \new_[23760]_ ;
  assign \new_[23770]_  = ~A199 & A166;
  assign \new_[23771]_  = A167 & \new_[23770]_ ;
  assign \new_[23775]_  = A202 & A201;
  assign \new_[23776]_  = A200 & \new_[23775]_ ;
  assign \new_[23777]_  = \new_[23776]_  & \new_[23771]_ ;
  assign \new_[23781]_  = ~A298 & A269;
  assign \new_[23782]_  = ~A267 & \new_[23781]_ ;
  assign \new_[23786]_  = A302 & A300;
  assign \new_[23787]_  = A299 & \new_[23786]_ ;
  assign \new_[23788]_  = \new_[23787]_  & \new_[23782]_ ;
  assign \new_[23792]_  = ~A199 & A166;
  assign \new_[23793]_  = A167 & \new_[23792]_ ;
  assign \new_[23797]_  = A202 & A201;
  assign \new_[23798]_  = A200 & \new_[23797]_ ;
  assign \new_[23799]_  = \new_[23798]_  & \new_[23793]_ ;
  assign \new_[23803]_  = A298 & A266;
  assign \new_[23804]_  = A265 & \new_[23803]_ ;
  assign \new_[23808]_  = A301 & A300;
  assign \new_[23809]_  = ~A299 & \new_[23808]_ ;
  assign \new_[23810]_  = \new_[23809]_  & \new_[23804]_ ;
  assign \new_[23814]_  = ~A199 & A166;
  assign \new_[23815]_  = A167 & \new_[23814]_ ;
  assign \new_[23819]_  = A202 & A201;
  assign \new_[23820]_  = A200 & \new_[23819]_ ;
  assign \new_[23821]_  = \new_[23820]_  & \new_[23815]_ ;
  assign \new_[23825]_  = A298 & A266;
  assign \new_[23826]_  = A265 & \new_[23825]_ ;
  assign \new_[23830]_  = A302 & A300;
  assign \new_[23831]_  = ~A299 & \new_[23830]_ ;
  assign \new_[23832]_  = \new_[23831]_  & \new_[23826]_ ;
  assign \new_[23836]_  = ~A199 & A166;
  assign \new_[23837]_  = A167 & \new_[23836]_ ;
  assign \new_[23841]_  = A202 & A201;
  assign \new_[23842]_  = A200 & \new_[23841]_ ;
  assign \new_[23843]_  = \new_[23842]_  & \new_[23837]_ ;
  assign \new_[23847]_  = ~A298 & A266;
  assign \new_[23848]_  = A265 & \new_[23847]_ ;
  assign \new_[23852]_  = A301 & A300;
  assign \new_[23853]_  = A299 & \new_[23852]_ ;
  assign \new_[23854]_  = \new_[23853]_  & \new_[23848]_ ;
  assign \new_[23858]_  = ~A199 & A166;
  assign \new_[23859]_  = A167 & \new_[23858]_ ;
  assign \new_[23863]_  = A202 & A201;
  assign \new_[23864]_  = A200 & \new_[23863]_ ;
  assign \new_[23865]_  = \new_[23864]_  & \new_[23859]_ ;
  assign \new_[23869]_  = ~A298 & A266;
  assign \new_[23870]_  = A265 & \new_[23869]_ ;
  assign \new_[23874]_  = A302 & A300;
  assign \new_[23875]_  = A299 & \new_[23874]_ ;
  assign \new_[23876]_  = \new_[23875]_  & \new_[23870]_ ;
  assign \new_[23880]_  = ~A199 & A166;
  assign \new_[23881]_  = A167 & \new_[23880]_ ;
  assign \new_[23885]_  = A202 & A201;
  assign \new_[23886]_  = A200 & \new_[23885]_ ;
  assign \new_[23887]_  = \new_[23886]_  & \new_[23881]_ ;
  assign \new_[23891]_  = A298 & ~A266;
  assign \new_[23892]_  = ~A265 & \new_[23891]_ ;
  assign \new_[23896]_  = A301 & A300;
  assign \new_[23897]_  = ~A299 & \new_[23896]_ ;
  assign \new_[23898]_  = \new_[23897]_  & \new_[23892]_ ;
  assign \new_[23902]_  = ~A199 & A166;
  assign \new_[23903]_  = A167 & \new_[23902]_ ;
  assign \new_[23907]_  = A202 & A201;
  assign \new_[23908]_  = A200 & \new_[23907]_ ;
  assign \new_[23909]_  = \new_[23908]_  & \new_[23903]_ ;
  assign \new_[23913]_  = A298 & ~A266;
  assign \new_[23914]_  = ~A265 & \new_[23913]_ ;
  assign \new_[23918]_  = A302 & A300;
  assign \new_[23919]_  = ~A299 & \new_[23918]_ ;
  assign \new_[23920]_  = \new_[23919]_  & \new_[23914]_ ;
  assign \new_[23924]_  = ~A199 & A166;
  assign \new_[23925]_  = A167 & \new_[23924]_ ;
  assign \new_[23929]_  = A202 & A201;
  assign \new_[23930]_  = A200 & \new_[23929]_ ;
  assign \new_[23931]_  = \new_[23930]_  & \new_[23925]_ ;
  assign \new_[23935]_  = ~A298 & ~A266;
  assign \new_[23936]_  = ~A265 & \new_[23935]_ ;
  assign \new_[23940]_  = A301 & A300;
  assign \new_[23941]_  = A299 & \new_[23940]_ ;
  assign \new_[23942]_  = \new_[23941]_  & \new_[23936]_ ;
  assign \new_[23946]_  = ~A199 & A166;
  assign \new_[23947]_  = A167 & \new_[23946]_ ;
  assign \new_[23951]_  = A202 & A201;
  assign \new_[23952]_  = A200 & \new_[23951]_ ;
  assign \new_[23953]_  = \new_[23952]_  & \new_[23947]_ ;
  assign \new_[23957]_  = ~A298 & ~A266;
  assign \new_[23958]_  = ~A265 & \new_[23957]_ ;
  assign \new_[23962]_  = A302 & A300;
  assign \new_[23963]_  = A299 & \new_[23962]_ ;
  assign \new_[23964]_  = \new_[23963]_  & \new_[23958]_ ;
  assign \new_[23968]_  = ~A199 & A166;
  assign \new_[23969]_  = A167 & \new_[23968]_ ;
  assign \new_[23973]_  = A203 & A201;
  assign \new_[23974]_  = A200 & \new_[23973]_ ;
  assign \new_[23975]_  = \new_[23974]_  & \new_[23969]_ ;
  assign \new_[23979]_  = A298 & A268;
  assign \new_[23980]_  = ~A267 & \new_[23979]_ ;
  assign \new_[23984]_  = A301 & A300;
  assign \new_[23985]_  = ~A299 & \new_[23984]_ ;
  assign \new_[23986]_  = \new_[23985]_  & \new_[23980]_ ;
  assign \new_[23990]_  = ~A199 & A166;
  assign \new_[23991]_  = A167 & \new_[23990]_ ;
  assign \new_[23995]_  = A203 & A201;
  assign \new_[23996]_  = A200 & \new_[23995]_ ;
  assign \new_[23997]_  = \new_[23996]_  & \new_[23991]_ ;
  assign \new_[24001]_  = A298 & A268;
  assign \new_[24002]_  = ~A267 & \new_[24001]_ ;
  assign \new_[24006]_  = A302 & A300;
  assign \new_[24007]_  = ~A299 & \new_[24006]_ ;
  assign \new_[24008]_  = \new_[24007]_  & \new_[24002]_ ;
  assign \new_[24012]_  = ~A199 & A166;
  assign \new_[24013]_  = A167 & \new_[24012]_ ;
  assign \new_[24017]_  = A203 & A201;
  assign \new_[24018]_  = A200 & \new_[24017]_ ;
  assign \new_[24019]_  = \new_[24018]_  & \new_[24013]_ ;
  assign \new_[24023]_  = ~A298 & A268;
  assign \new_[24024]_  = ~A267 & \new_[24023]_ ;
  assign \new_[24028]_  = A301 & A300;
  assign \new_[24029]_  = A299 & \new_[24028]_ ;
  assign \new_[24030]_  = \new_[24029]_  & \new_[24024]_ ;
  assign \new_[24034]_  = ~A199 & A166;
  assign \new_[24035]_  = A167 & \new_[24034]_ ;
  assign \new_[24039]_  = A203 & A201;
  assign \new_[24040]_  = A200 & \new_[24039]_ ;
  assign \new_[24041]_  = \new_[24040]_  & \new_[24035]_ ;
  assign \new_[24045]_  = ~A298 & A268;
  assign \new_[24046]_  = ~A267 & \new_[24045]_ ;
  assign \new_[24050]_  = A302 & A300;
  assign \new_[24051]_  = A299 & \new_[24050]_ ;
  assign \new_[24052]_  = \new_[24051]_  & \new_[24046]_ ;
  assign \new_[24056]_  = ~A199 & A166;
  assign \new_[24057]_  = A167 & \new_[24056]_ ;
  assign \new_[24061]_  = A203 & A201;
  assign \new_[24062]_  = A200 & \new_[24061]_ ;
  assign \new_[24063]_  = \new_[24062]_  & \new_[24057]_ ;
  assign \new_[24067]_  = A298 & A269;
  assign \new_[24068]_  = ~A267 & \new_[24067]_ ;
  assign \new_[24072]_  = A301 & A300;
  assign \new_[24073]_  = ~A299 & \new_[24072]_ ;
  assign \new_[24074]_  = \new_[24073]_  & \new_[24068]_ ;
  assign \new_[24078]_  = ~A199 & A166;
  assign \new_[24079]_  = A167 & \new_[24078]_ ;
  assign \new_[24083]_  = A203 & A201;
  assign \new_[24084]_  = A200 & \new_[24083]_ ;
  assign \new_[24085]_  = \new_[24084]_  & \new_[24079]_ ;
  assign \new_[24089]_  = A298 & A269;
  assign \new_[24090]_  = ~A267 & \new_[24089]_ ;
  assign \new_[24094]_  = A302 & A300;
  assign \new_[24095]_  = ~A299 & \new_[24094]_ ;
  assign \new_[24096]_  = \new_[24095]_  & \new_[24090]_ ;
  assign \new_[24100]_  = ~A199 & A166;
  assign \new_[24101]_  = A167 & \new_[24100]_ ;
  assign \new_[24105]_  = A203 & A201;
  assign \new_[24106]_  = A200 & \new_[24105]_ ;
  assign \new_[24107]_  = \new_[24106]_  & \new_[24101]_ ;
  assign \new_[24111]_  = ~A298 & A269;
  assign \new_[24112]_  = ~A267 & \new_[24111]_ ;
  assign \new_[24116]_  = A301 & A300;
  assign \new_[24117]_  = A299 & \new_[24116]_ ;
  assign \new_[24118]_  = \new_[24117]_  & \new_[24112]_ ;
  assign \new_[24122]_  = ~A199 & A166;
  assign \new_[24123]_  = A167 & \new_[24122]_ ;
  assign \new_[24127]_  = A203 & A201;
  assign \new_[24128]_  = A200 & \new_[24127]_ ;
  assign \new_[24129]_  = \new_[24128]_  & \new_[24123]_ ;
  assign \new_[24133]_  = ~A298 & A269;
  assign \new_[24134]_  = ~A267 & \new_[24133]_ ;
  assign \new_[24138]_  = A302 & A300;
  assign \new_[24139]_  = A299 & \new_[24138]_ ;
  assign \new_[24140]_  = \new_[24139]_  & \new_[24134]_ ;
  assign \new_[24144]_  = ~A199 & A166;
  assign \new_[24145]_  = A167 & \new_[24144]_ ;
  assign \new_[24149]_  = A203 & A201;
  assign \new_[24150]_  = A200 & \new_[24149]_ ;
  assign \new_[24151]_  = \new_[24150]_  & \new_[24145]_ ;
  assign \new_[24155]_  = A298 & A266;
  assign \new_[24156]_  = A265 & \new_[24155]_ ;
  assign \new_[24160]_  = A301 & A300;
  assign \new_[24161]_  = ~A299 & \new_[24160]_ ;
  assign \new_[24162]_  = \new_[24161]_  & \new_[24156]_ ;
  assign \new_[24166]_  = ~A199 & A166;
  assign \new_[24167]_  = A167 & \new_[24166]_ ;
  assign \new_[24171]_  = A203 & A201;
  assign \new_[24172]_  = A200 & \new_[24171]_ ;
  assign \new_[24173]_  = \new_[24172]_  & \new_[24167]_ ;
  assign \new_[24177]_  = A298 & A266;
  assign \new_[24178]_  = A265 & \new_[24177]_ ;
  assign \new_[24182]_  = A302 & A300;
  assign \new_[24183]_  = ~A299 & \new_[24182]_ ;
  assign \new_[24184]_  = \new_[24183]_  & \new_[24178]_ ;
  assign \new_[24188]_  = ~A199 & A166;
  assign \new_[24189]_  = A167 & \new_[24188]_ ;
  assign \new_[24193]_  = A203 & A201;
  assign \new_[24194]_  = A200 & \new_[24193]_ ;
  assign \new_[24195]_  = \new_[24194]_  & \new_[24189]_ ;
  assign \new_[24199]_  = ~A298 & A266;
  assign \new_[24200]_  = A265 & \new_[24199]_ ;
  assign \new_[24204]_  = A301 & A300;
  assign \new_[24205]_  = A299 & \new_[24204]_ ;
  assign \new_[24206]_  = \new_[24205]_  & \new_[24200]_ ;
  assign \new_[24210]_  = ~A199 & A166;
  assign \new_[24211]_  = A167 & \new_[24210]_ ;
  assign \new_[24215]_  = A203 & A201;
  assign \new_[24216]_  = A200 & \new_[24215]_ ;
  assign \new_[24217]_  = \new_[24216]_  & \new_[24211]_ ;
  assign \new_[24221]_  = ~A298 & A266;
  assign \new_[24222]_  = A265 & \new_[24221]_ ;
  assign \new_[24226]_  = A302 & A300;
  assign \new_[24227]_  = A299 & \new_[24226]_ ;
  assign \new_[24228]_  = \new_[24227]_  & \new_[24222]_ ;
  assign \new_[24232]_  = ~A199 & A166;
  assign \new_[24233]_  = A167 & \new_[24232]_ ;
  assign \new_[24237]_  = A203 & A201;
  assign \new_[24238]_  = A200 & \new_[24237]_ ;
  assign \new_[24239]_  = \new_[24238]_  & \new_[24233]_ ;
  assign \new_[24243]_  = A298 & ~A266;
  assign \new_[24244]_  = ~A265 & \new_[24243]_ ;
  assign \new_[24248]_  = A301 & A300;
  assign \new_[24249]_  = ~A299 & \new_[24248]_ ;
  assign \new_[24250]_  = \new_[24249]_  & \new_[24244]_ ;
  assign \new_[24254]_  = ~A199 & A166;
  assign \new_[24255]_  = A167 & \new_[24254]_ ;
  assign \new_[24259]_  = A203 & A201;
  assign \new_[24260]_  = A200 & \new_[24259]_ ;
  assign \new_[24261]_  = \new_[24260]_  & \new_[24255]_ ;
  assign \new_[24265]_  = A298 & ~A266;
  assign \new_[24266]_  = ~A265 & \new_[24265]_ ;
  assign \new_[24270]_  = A302 & A300;
  assign \new_[24271]_  = ~A299 & \new_[24270]_ ;
  assign \new_[24272]_  = \new_[24271]_  & \new_[24266]_ ;
  assign \new_[24276]_  = ~A199 & A166;
  assign \new_[24277]_  = A167 & \new_[24276]_ ;
  assign \new_[24281]_  = A203 & A201;
  assign \new_[24282]_  = A200 & \new_[24281]_ ;
  assign \new_[24283]_  = \new_[24282]_  & \new_[24277]_ ;
  assign \new_[24287]_  = ~A298 & ~A266;
  assign \new_[24288]_  = ~A265 & \new_[24287]_ ;
  assign \new_[24292]_  = A301 & A300;
  assign \new_[24293]_  = A299 & \new_[24292]_ ;
  assign \new_[24294]_  = \new_[24293]_  & \new_[24288]_ ;
  assign \new_[24298]_  = ~A199 & A166;
  assign \new_[24299]_  = A167 & \new_[24298]_ ;
  assign \new_[24303]_  = A203 & A201;
  assign \new_[24304]_  = A200 & \new_[24303]_ ;
  assign \new_[24305]_  = \new_[24304]_  & \new_[24299]_ ;
  assign \new_[24309]_  = ~A298 & ~A266;
  assign \new_[24310]_  = ~A265 & \new_[24309]_ ;
  assign \new_[24314]_  = A302 & A300;
  assign \new_[24315]_  = A299 & \new_[24314]_ ;
  assign \new_[24316]_  = \new_[24315]_  & \new_[24310]_ ;
  assign \new_[24320]_  = A199 & A166;
  assign \new_[24321]_  = A167 & \new_[24320]_ ;
  assign \new_[24325]_  = A202 & A201;
  assign \new_[24326]_  = ~A200 & \new_[24325]_ ;
  assign \new_[24327]_  = \new_[24326]_  & \new_[24321]_ ;
  assign \new_[24331]_  = A298 & A268;
  assign \new_[24332]_  = ~A267 & \new_[24331]_ ;
  assign \new_[24336]_  = A301 & A300;
  assign \new_[24337]_  = ~A299 & \new_[24336]_ ;
  assign \new_[24338]_  = \new_[24337]_  & \new_[24332]_ ;
  assign \new_[24342]_  = A199 & A166;
  assign \new_[24343]_  = A167 & \new_[24342]_ ;
  assign \new_[24347]_  = A202 & A201;
  assign \new_[24348]_  = ~A200 & \new_[24347]_ ;
  assign \new_[24349]_  = \new_[24348]_  & \new_[24343]_ ;
  assign \new_[24353]_  = A298 & A268;
  assign \new_[24354]_  = ~A267 & \new_[24353]_ ;
  assign \new_[24358]_  = A302 & A300;
  assign \new_[24359]_  = ~A299 & \new_[24358]_ ;
  assign \new_[24360]_  = \new_[24359]_  & \new_[24354]_ ;
  assign \new_[24364]_  = A199 & A166;
  assign \new_[24365]_  = A167 & \new_[24364]_ ;
  assign \new_[24369]_  = A202 & A201;
  assign \new_[24370]_  = ~A200 & \new_[24369]_ ;
  assign \new_[24371]_  = \new_[24370]_  & \new_[24365]_ ;
  assign \new_[24375]_  = ~A298 & A268;
  assign \new_[24376]_  = ~A267 & \new_[24375]_ ;
  assign \new_[24380]_  = A301 & A300;
  assign \new_[24381]_  = A299 & \new_[24380]_ ;
  assign \new_[24382]_  = \new_[24381]_  & \new_[24376]_ ;
  assign \new_[24386]_  = A199 & A166;
  assign \new_[24387]_  = A167 & \new_[24386]_ ;
  assign \new_[24391]_  = A202 & A201;
  assign \new_[24392]_  = ~A200 & \new_[24391]_ ;
  assign \new_[24393]_  = \new_[24392]_  & \new_[24387]_ ;
  assign \new_[24397]_  = ~A298 & A268;
  assign \new_[24398]_  = ~A267 & \new_[24397]_ ;
  assign \new_[24402]_  = A302 & A300;
  assign \new_[24403]_  = A299 & \new_[24402]_ ;
  assign \new_[24404]_  = \new_[24403]_  & \new_[24398]_ ;
  assign \new_[24408]_  = A199 & A166;
  assign \new_[24409]_  = A167 & \new_[24408]_ ;
  assign \new_[24413]_  = A202 & A201;
  assign \new_[24414]_  = ~A200 & \new_[24413]_ ;
  assign \new_[24415]_  = \new_[24414]_  & \new_[24409]_ ;
  assign \new_[24419]_  = A298 & A269;
  assign \new_[24420]_  = ~A267 & \new_[24419]_ ;
  assign \new_[24424]_  = A301 & A300;
  assign \new_[24425]_  = ~A299 & \new_[24424]_ ;
  assign \new_[24426]_  = \new_[24425]_  & \new_[24420]_ ;
  assign \new_[24430]_  = A199 & A166;
  assign \new_[24431]_  = A167 & \new_[24430]_ ;
  assign \new_[24435]_  = A202 & A201;
  assign \new_[24436]_  = ~A200 & \new_[24435]_ ;
  assign \new_[24437]_  = \new_[24436]_  & \new_[24431]_ ;
  assign \new_[24441]_  = A298 & A269;
  assign \new_[24442]_  = ~A267 & \new_[24441]_ ;
  assign \new_[24446]_  = A302 & A300;
  assign \new_[24447]_  = ~A299 & \new_[24446]_ ;
  assign \new_[24448]_  = \new_[24447]_  & \new_[24442]_ ;
  assign \new_[24452]_  = A199 & A166;
  assign \new_[24453]_  = A167 & \new_[24452]_ ;
  assign \new_[24457]_  = A202 & A201;
  assign \new_[24458]_  = ~A200 & \new_[24457]_ ;
  assign \new_[24459]_  = \new_[24458]_  & \new_[24453]_ ;
  assign \new_[24463]_  = ~A298 & A269;
  assign \new_[24464]_  = ~A267 & \new_[24463]_ ;
  assign \new_[24468]_  = A301 & A300;
  assign \new_[24469]_  = A299 & \new_[24468]_ ;
  assign \new_[24470]_  = \new_[24469]_  & \new_[24464]_ ;
  assign \new_[24474]_  = A199 & A166;
  assign \new_[24475]_  = A167 & \new_[24474]_ ;
  assign \new_[24479]_  = A202 & A201;
  assign \new_[24480]_  = ~A200 & \new_[24479]_ ;
  assign \new_[24481]_  = \new_[24480]_  & \new_[24475]_ ;
  assign \new_[24485]_  = ~A298 & A269;
  assign \new_[24486]_  = ~A267 & \new_[24485]_ ;
  assign \new_[24490]_  = A302 & A300;
  assign \new_[24491]_  = A299 & \new_[24490]_ ;
  assign \new_[24492]_  = \new_[24491]_  & \new_[24486]_ ;
  assign \new_[24496]_  = A199 & A166;
  assign \new_[24497]_  = A167 & \new_[24496]_ ;
  assign \new_[24501]_  = A202 & A201;
  assign \new_[24502]_  = ~A200 & \new_[24501]_ ;
  assign \new_[24503]_  = \new_[24502]_  & \new_[24497]_ ;
  assign \new_[24507]_  = A298 & A266;
  assign \new_[24508]_  = A265 & \new_[24507]_ ;
  assign \new_[24512]_  = A301 & A300;
  assign \new_[24513]_  = ~A299 & \new_[24512]_ ;
  assign \new_[24514]_  = \new_[24513]_  & \new_[24508]_ ;
  assign \new_[24518]_  = A199 & A166;
  assign \new_[24519]_  = A167 & \new_[24518]_ ;
  assign \new_[24523]_  = A202 & A201;
  assign \new_[24524]_  = ~A200 & \new_[24523]_ ;
  assign \new_[24525]_  = \new_[24524]_  & \new_[24519]_ ;
  assign \new_[24529]_  = A298 & A266;
  assign \new_[24530]_  = A265 & \new_[24529]_ ;
  assign \new_[24534]_  = A302 & A300;
  assign \new_[24535]_  = ~A299 & \new_[24534]_ ;
  assign \new_[24536]_  = \new_[24535]_  & \new_[24530]_ ;
  assign \new_[24540]_  = A199 & A166;
  assign \new_[24541]_  = A167 & \new_[24540]_ ;
  assign \new_[24545]_  = A202 & A201;
  assign \new_[24546]_  = ~A200 & \new_[24545]_ ;
  assign \new_[24547]_  = \new_[24546]_  & \new_[24541]_ ;
  assign \new_[24551]_  = ~A298 & A266;
  assign \new_[24552]_  = A265 & \new_[24551]_ ;
  assign \new_[24556]_  = A301 & A300;
  assign \new_[24557]_  = A299 & \new_[24556]_ ;
  assign \new_[24558]_  = \new_[24557]_  & \new_[24552]_ ;
  assign \new_[24562]_  = A199 & A166;
  assign \new_[24563]_  = A167 & \new_[24562]_ ;
  assign \new_[24567]_  = A202 & A201;
  assign \new_[24568]_  = ~A200 & \new_[24567]_ ;
  assign \new_[24569]_  = \new_[24568]_  & \new_[24563]_ ;
  assign \new_[24573]_  = ~A298 & A266;
  assign \new_[24574]_  = A265 & \new_[24573]_ ;
  assign \new_[24578]_  = A302 & A300;
  assign \new_[24579]_  = A299 & \new_[24578]_ ;
  assign \new_[24580]_  = \new_[24579]_  & \new_[24574]_ ;
  assign \new_[24584]_  = A199 & A166;
  assign \new_[24585]_  = A167 & \new_[24584]_ ;
  assign \new_[24589]_  = A202 & A201;
  assign \new_[24590]_  = ~A200 & \new_[24589]_ ;
  assign \new_[24591]_  = \new_[24590]_  & \new_[24585]_ ;
  assign \new_[24595]_  = A298 & ~A266;
  assign \new_[24596]_  = ~A265 & \new_[24595]_ ;
  assign \new_[24600]_  = A301 & A300;
  assign \new_[24601]_  = ~A299 & \new_[24600]_ ;
  assign \new_[24602]_  = \new_[24601]_  & \new_[24596]_ ;
  assign \new_[24606]_  = A199 & A166;
  assign \new_[24607]_  = A167 & \new_[24606]_ ;
  assign \new_[24611]_  = A202 & A201;
  assign \new_[24612]_  = ~A200 & \new_[24611]_ ;
  assign \new_[24613]_  = \new_[24612]_  & \new_[24607]_ ;
  assign \new_[24617]_  = A298 & ~A266;
  assign \new_[24618]_  = ~A265 & \new_[24617]_ ;
  assign \new_[24622]_  = A302 & A300;
  assign \new_[24623]_  = ~A299 & \new_[24622]_ ;
  assign \new_[24624]_  = \new_[24623]_  & \new_[24618]_ ;
  assign \new_[24628]_  = A199 & A166;
  assign \new_[24629]_  = A167 & \new_[24628]_ ;
  assign \new_[24633]_  = A202 & A201;
  assign \new_[24634]_  = ~A200 & \new_[24633]_ ;
  assign \new_[24635]_  = \new_[24634]_  & \new_[24629]_ ;
  assign \new_[24639]_  = ~A298 & ~A266;
  assign \new_[24640]_  = ~A265 & \new_[24639]_ ;
  assign \new_[24644]_  = A301 & A300;
  assign \new_[24645]_  = A299 & \new_[24644]_ ;
  assign \new_[24646]_  = \new_[24645]_  & \new_[24640]_ ;
  assign \new_[24650]_  = A199 & A166;
  assign \new_[24651]_  = A167 & \new_[24650]_ ;
  assign \new_[24655]_  = A202 & A201;
  assign \new_[24656]_  = ~A200 & \new_[24655]_ ;
  assign \new_[24657]_  = \new_[24656]_  & \new_[24651]_ ;
  assign \new_[24661]_  = ~A298 & ~A266;
  assign \new_[24662]_  = ~A265 & \new_[24661]_ ;
  assign \new_[24666]_  = A302 & A300;
  assign \new_[24667]_  = A299 & \new_[24666]_ ;
  assign \new_[24668]_  = \new_[24667]_  & \new_[24662]_ ;
  assign \new_[24672]_  = A199 & A166;
  assign \new_[24673]_  = A167 & \new_[24672]_ ;
  assign \new_[24677]_  = A203 & A201;
  assign \new_[24678]_  = ~A200 & \new_[24677]_ ;
  assign \new_[24679]_  = \new_[24678]_  & \new_[24673]_ ;
  assign \new_[24683]_  = A298 & A268;
  assign \new_[24684]_  = ~A267 & \new_[24683]_ ;
  assign \new_[24688]_  = A301 & A300;
  assign \new_[24689]_  = ~A299 & \new_[24688]_ ;
  assign \new_[24690]_  = \new_[24689]_  & \new_[24684]_ ;
  assign \new_[24694]_  = A199 & A166;
  assign \new_[24695]_  = A167 & \new_[24694]_ ;
  assign \new_[24699]_  = A203 & A201;
  assign \new_[24700]_  = ~A200 & \new_[24699]_ ;
  assign \new_[24701]_  = \new_[24700]_  & \new_[24695]_ ;
  assign \new_[24705]_  = A298 & A268;
  assign \new_[24706]_  = ~A267 & \new_[24705]_ ;
  assign \new_[24710]_  = A302 & A300;
  assign \new_[24711]_  = ~A299 & \new_[24710]_ ;
  assign \new_[24712]_  = \new_[24711]_  & \new_[24706]_ ;
  assign \new_[24716]_  = A199 & A166;
  assign \new_[24717]_  = A167 & \new_[24716]_ ;
  assign \new_[24721]_  = A203 & A201;
  assign \new_[24722]_  = ~A200 & \new_[24721]_ ;
  assign \new_[24723]_  = \new_[24722]_  & \new_[24717]_ ;
  assign \new_[24727]_  = ~A298 & A268;
  assign \new_[24728]_  = ~A267 & \new_[24727]_ ;
  assign \new_[24732]_  = A301 & A300;
  assign \new_[24733]_  = A299 & \new_[24732]_ ;
  assign \new_[24734]_  = \new_[24733]_  & \new_[24728]_ ;
  assign \new_[24738]_  = A199 & A166;
  assign \new_[24739]_  = A167 & \new_[24738]_ ;
  assign \new_[24743]_  = A203 & A201;
  assign \new_[24744]_  = ~A200 & \new_[24743]_ ;
  assign \new_[24745]_  = \new_[24744]_  & \new_[24739]_ ;
  assign \new_[24749]_  = ~A298 & A268;
  assign \new_[24750]_  = ~A267 & \new_[24749]_ ;
  assign \new_[24754]_  = A302 & A300;
  assign \new_[24755]_  = A299 & \new_[24754]_ ;
  assign \new_[24756]_  = \new_[24755]_  & \new_[24750]_ ;
  assign \new_[24760]_  = A199 & A166;
  assign \new_[24761]_  = A167 & \new_[24760]_ ;
  assign \new_[24765]_  = A203 & A201;
  assign \new_[24766]_  = ~A200 & \new_[24765]_ ;
  assign \new_[24767]_  = \new_[24766]_  & \new_[24761]_ ;
  assign \new_[24771]_  = A298 & A269;
  assign \new_[24772]_  = ~A267 & \new_[24771]_ ;
  assign \new_[24776]_  = A301 & A300;
  assign \new_[24777]_  = ~A299 & \new_[24776]_ ;
  assign \new_[24778]_  = \new_[24777]_  & \new_[24772]_ ;
  assign \new_[24782]_  = A199 & A166;
  assign \new_[24783]_  = A167 & \new_[24782]_ ;
  assign \new_[24787]_  = A203 & A201;
  assign \new_[24788]_  = ~A200 & \new_[24787]_ ;
  assign \new_[24789]_  = \new_[24788]_  & \new_[24783]_ ;
  assign \new_[24793]_  = A298 & A269;
  assign \new_[24794]_  = ~A267 & \new_[24793]_ ;
  assign \new_[24798]_  = A302 & A300;
  assign \new_[24799]_  = ~A299 & \new_[24798]_ ;
  assign \new_[24800]_  = \new_[24799]_  & \new_[24794]_ ;
  assign \new_[24804]_  = A199 & A166;
  assign \new_[24805]_  = A167 & \new_[24804]_ ;
  assign \new_[24809]_  = A203 & A201;
  assign \new_[24810]_  = ~A200 & \new_[24809]_ ;
  assign \new_[24811]_  = \new_[24810]_  & \new_[24805]_ ;
  assign \new_[24815]_  = ~A298 & A269;
  assign \new_[24816]_  = ~A267 & \new_[24815]_ ;
  assign \new_[24820]_  = A301 & A300;
  assign \new_[24821]_  = A299 & \new_[24820]_ ;
  assign \new_[24822]_  = \new_[24821]_  & \new_[24816]_ ;
  assign \new_[24826]_  = A199 & A166;
  assign \new_[24827]_  = A167 & \new_[24826]_ ;
  assign \new_[24831]_  = A203 & A201;
  assign \new_[24832]_  = ~A200 & \new_[24831]_ ;
  assign \new_[24833]_  = \new_[24832]_  & \new_[24827]_ ;
  assign \new_[24837]_  = ~A298 & A269;
  assign \new_[24838]_  = ~A267 & \new_[24837]_ ;
  assign \new_[24842]_  = A302 & A300;
  assign \new_[24843]_  = A299 & \new_[24842]_ ;
  assign \new_[24844]_  = \new_[24843]_  & \new_[24838]_ ;
  assign \new_[24848]_  = A199 & A166;
  assign \new_[24849]_  = A167 & \new_[24848]_ ;
  assign \new_[24853]_  = A203 & A201;
  assign \new_[24854]_  = ~A200 & \new_[24853]_ ;
  assign \new_[24855]_  = \new_[24854]_  & \new_[24849]_ ;
  assign \new_[24859]_  = A298 & A266;
  assign \new_[24860]_  = A265 & \new_[24859]_ ;
  assign \new_[24864]_  = A301 & A300;
  assign \new_[24865]_  = ~A299 & \new_[24864]_ ;
  assign \new_[24866]_  = \new_[24865]_  & \new_[24860]_ ;
  assign \new_[24870]_  = A199 & A166;
  assign \new_[24871]_  = A167 & \new_[24870]_ ;
  assign \new_[24875]_  = A203 & A201;
  assign \new_[24876]_  = ~A200 & \new_[24875]_ ;
  assign \new_[24877]_  = \new_[24876]_  & \new_[24871]_ ;
  assign \new_[24881]_  = A298 & A266;
  assign \new_[24882]_  = A265 & \new_[24881]_ ;
  assign \new_[24886]_  = A302 & A300;
  assign \new_[24887]_  = ~A299 & \new_[24886]_ ;
  assign \new_[24888]_  = \new_[24887]_  & \new_[24882]_ ;
  assign \new_[24892]_  = A199 & A166;
  assign \new_[24893]_  = A167 & \new_[24892]_ ;
  assign \new_[24897]_  = A203 & A201;
  assign \new_[24898]_  = ~A200 & \new_[24897]_ ;
  assign \new_[24899]_  = \new_[24898]_  & \new_[24893]_ ;
  assign \new_[24903]_  = ~A298 & A266;
  assign \new_[24904]_  = A265 & \new_[24903]_ ;
  assign \new_[24908]_  = A301 & A300;
  assign \new_[24909]_  = A299 & \new_[24908]_ ;
  assign \new_[24910]_  = \new_[24909]_  & \new_[24904]_ ;
  assign \new_[24914]_  = A199 & A166;
  assign \new_[24915]_  = A167 & \new_[24914]_ ;
  assign \new_[24919]_  = A203 & A201;
  assign \new_[24920]_  = ~A200 & \new_[24919]_ ;
  assign \new_[24921]_  = \new_[24920]_  & \new_[24915]_ ;
  assign \new_[24925]_  = ~A298 & A266;
  assign \new_[24926]_  = A265 & \new_[24925]_ ;
  assign \new_[24930]_  = A302 & A300;
  assign \new_[24931]_  = A299 & \new_[24930]_ ;
  assign \new_[24932]_  = \new_[24931]_  & \new_[24926]_ ;
  assign \new_[24936]_  = A199 & A166;
  assign \new_[24937]_  = A167 & \new_[24936]_ ;
  assign \new_[24941]_  = A203 & A201;
  assign \new_[24942]_  = ~A200 & \new_[24941]_ ;
  assign \new_[24943]_  = \new_[24942]_  & \new_[24937]_ ;
  assign \new_[24947]_  = A298 & ~A266;
  assign \new_[24948]_  = ~A265 & \new_[24947]_ ;
  assign \new_[24952]_  = A301 & A300;
  assign \new_[24953]_  = ~A299 & \new_[24952]_ ;
  assign \new_[24954]_  = \new_[24953]_  & \new_[24948]_ ;
  assign \new_[24958]_  = A199 & A166;
  assign \new_[24959]_  = A167 & \new_[24958]_ ;
  assign \new_[24963]_  = A203 & A201;
  assign \new_[24964]_  = ~A200 & \new_[24963]_ ;
  assign \new_[24965]_  = \new_[24964]_  & \new_[24959]_ ;
  assign \new_[24969]_  = A298 & ~A266;
  assign \new_[24970]_  = ~A265 & \new_[24969]_ ;
  assign \new_[24974]_  = A302 & A300;
  assign \new_[24975]_  = ~A299 & \new_[24974]_ ;
  assign \new_[24976]_  = \new_[24975]_  & \new_[24970]_ ;
  assign \new_[24980]_  = A199 & A166;
  assign \new_[24981]_  = A167 & \new_[24980]_ ;
  assign \new_[24985]_  = A203 & A201;
  assign \new_[24986]_  = ~A200 & \new_[24985]_ ;
  assign \new_[24987]_  = \new_[24986]_  & \new_[24981]_ ;
  assign \new_[24991]_  = ~A298 & ~A266;
  assign \new_[24992]_  = ~A265 & \new_[24991]_ ;
  assign \new_[24996]_  = A301 & A300;
  assign \new_[24997]_  = A299 & \new_[24996]_ ;
  assign \new_[24998]_  = \new_[24997]_  & \new_[24992]_ ;
  assign \new_[25002]_  = A199 & A166;
  assign \new_[25003]_  = A167 & \new_[25002]_ ;
  assign \new_[25007]_  = A203 & A201;
  assign \new_[25008]_  = ~A200 & \new_[25007]_ ;
  assign \new_[25009]_  = \new_[25008]_  & \new_[25003]_ ;
  assign \new_[25013]_  = ~A298 & ~A266;
  assign \new_[25014]_  = ~A265 & \new_[25013]_ ;
  assign \new_[25018]_  = A302 & A300;
  assign \new_[25019]_  = A299 & \new_[25018]_ ;
  assign \new_[25020]_  = \new_[25019]_  & \new_[25014]_ ;
  assign \new_[25024]_  = ~A199 & A166;
  assign \new_[25025]_  = A167 & \new_[25024]_ ;
  assign \new_[25029]_  = A266 & ~A265;
  assign \new_[25030]_  = ~A200 & \new_[25029]_ ;
  assign \new_[25031]_  = \new_[25030]_  & \new_[25025]_ ;
  assign \new_[25035]_  = ~A269 & ~A268;
  assign \new_[25036]_  = ~A267 & \new_[25035]_ ;
  assign \new_[25040]_  = ~A302 & ~A301;
  assign \new_[25041]_  = A300 & \new_[25040]_ ;
  assign \new_[25042]_  = \new_[25041]_  & \new_[25036]_ ;
  assign \new_[25046]_  = ~A199 & A166;
  assign \new_[25047]_  = A167 & \new_[25046]_ ;
  assign \new_[25051]_  = ~A266 & A265;
  assign \new_[25052]_  = ~A200 & \new_[25051]_ ;
  assign \new_[25053]_  = \new_[25052]_  & \new_[25047]_ ;
  assign \new_[25057]_  = ~A269 & ~A268;
  assign \new_[25058]_  = ~A267 & \new_[25057]_ ;
  assign \new_[25062]_  = ~A302 & ~A301;
  assign \new_[25063]_  = A300 & \new_[25062]_ ;
  assign \new_[25064]_  = \new_[25063]_  & \new_[25058]_ ;
  assign \new_[25068]_  = A201 & ~A166;
  assign \new_[25069]_  = ~A167 & \new_[25068]_ ;
  assign \new_[25073]_  = ~A265 & ~A203;
  assign \new_[25074]_  = ~A202 & \new_[25073]_ ;
  assign \new_[25075]_  = \new_[25074]_  & \new_[25069]_ ;
  assign \new_[25079]_  = A268 & A267;
  assign \new_[25080]_  = A266 & \new_[25079]_ ;
  assign \new_[25084]_  = ~A302 & ~A301;
  assign \new_[25085]_  = A300 & \new_[25084]_ ;
  assign \new_[25086]_  = \new_[25085]_  & \new_[25080]_ ;
  assign \new_[25090]_  = A201 & ~A166;
  assign \new_[25091]_  = ~A167 & \new_[25090]_ ;
  assign \new_[25095]_  = ~A265 & ~A203;
  assign \new_[25096]_  = ~A202 & \new_[25095]_ ;
  assign \new_[25097]_  = \new_[25096]_  & \new_[25091]_ ;
  assign \new_[25101]_  = A269 & A267;
  assign \new_[25102]_  = A266 & \new_[25101]_ ;
  assign \new_[25106]_  = ~A302 & ~A301;
  assign \new_[25107]_  = A300 & \new_[25106]_ ;
  assign \new_[25108]_  = \new_[25107]_  & \new_[25102]_ ;
  assign \new_[25112]_  = A201 & ~A166;
  assign \new_[25113]_  = ~A167 & \new_[25112]_ ;
  assign \new_[25117]_  = ~A265 & ~A203;
  assign \new_[25118]_  = ~A202 & \new_[25117]_ ;
  assign \new_[25119]_  = \new_[25118]_  & \new_[25113]_ ;
  assign \new_[25123]_  = ~A268 & ~A267;
  assign \new_[25124]_  = A266 & \new_[25123]_ ;
  assign \new_[25128]_  = A301 & ~A300;
  assign \new_[25129]_  = ~A269 & \new_[25128]_ ;
  assign \new_[25130]_  = \new_[25129]_  & \new_[25124]_ ;
  assign \new_[25134]_  = A201 & ~A166;
  assign \new_[25135]_  = ~A167 & \new_[25134]_ ;
  assign \new_[25139]_  = ~A265 & ~A203;
  assign \new_[25140]_  = ~A202 & \new_[25139]_ ;
  assign \new_[25141]_  = \new_[25140]_  & \new_[25135]_ ;
  assign \new_[25145]_  = ~A268 & ~A267;
  assign \new_[25146]_  = A266 & \new_[25145]_ ;
  assign \new_[25150]_  = A302 & ~A300;
  assign \new_[25151]_  = ~A269 & \new_[25150]_ ;
  assign \new_[25152]_  = \new_[25151]_  & \new_[25146]_ ;
  assign \new_[25156]_  = A201 & ~A166;
  assign \new_[25157]_  = ~A167 & \new_[25156]_ ;
  assign \new_[25161]_  = ~A265 & ~A203;
  assign \new_[25162]_  = ~A202 & \new_[25161]_ ;
  assign \new_[25163]_  = \new_[25162]_  & \new_[25157]_ ;
  assign \new_[25167]_  = ~A268 & ~A267;
  assign \new_[25168]_  = A266 & \new_[25167]_ ;
  assign \new_[25172]_  = A299 & A298;
  assign \new_[25173]_  = ~A269 & \new_[25172]_ ;
  assign \new_[25174]_  = \new_[25173]_  & \new_[25168]_ ;
  assign \new_[25178]_  = A201 & ~A166;
  assign \new_[25179]_  = ~A167 & \new_[25178]_ ;
  assign \new_[25183]_  = ~A265 & ~A203;
  assign \new_[25184]_  = ~A202 & \new_[25183]_ ;
  assign \new_[25185]_  = \new_[25184]_  & \new_[25179]_ ;
  assign \new_[25189]_  = ~A268 & ~A267;
  assign \new_[25190]_  = A266 & \new_[25189]_ ;
  assign \new_[25194]_  = ~A299 & ~A298;
  assign \new_[25195]_  = ~A269 & \new_[25194]_ ;
  assign \new_[25196]_  = \new_[25195]_  & \new_[25190]_ ;
  assign \new_[25200]_  = A201 & ~A166;
  assign \new_[25201]_  = ~A167 & \new_[25200]_ ;
  assign \new_[25205]_  = A265 & ~A203;
  assign \new_[25206]_  = ~A202 & \new_[25205]_ ;
  assign \new_[25207]_  = \new_[25206]_  & \new_[25201]_ ;
  assign \new_[25211]_  = A268 & A267;
  assign \new_[25212]_  = ~A266 & \new_[25211]_ ;
  assign \new_[25216]_  = ~A302 & ~A301;
  assign \new_[25217]_  = A300 & \new_[25216]_ ;
  assign \new_[25218]_  = \new_[25217]_  & \new_[25212]_ ;
  assign \new_[25222]_  = A201 & ~A166;
  assign \new_[25223]_  = ~A167 & \new_[25222]_ ;
  assign \new_[25227]_  = A265 & ~A203;
  assign \new_[25228]_  = ~A202 & \new_[25227]_ ;
  assign \new_[25229]_  = \new_[25228]_  & \new_[25223]_ ;
  assign \new_[25233]_  = A269 & A267;
  assign \new_[25234]_  = ~A266 & \new_[25233]_ ;
  assign \new_[25238]_  = ~A302 & ~A301;
  assign \new_[25239]_  = A300 & \new_[25238]_ ;
  assign \new_[25240]_  = \new_[25239]_  & \new_[25234]_ ;
  assign \new_[25244]_  = A201 & ~A166;
  assign \new_[25245]_  = ~A167 & \new_[25244]_ ;
  assign \new_[25249]_  = A265 & ~A203;
  assign \new_[25250]_  = ~A202 & \new_[25249]_ ;
  assign \new_[25251]_  = \new_[25250]_  & \new_[25245]_ ;
  assign \new_[25255]_  = ~A268 & ~A267;
  assign \new_[25256]_  = ~A266 & \new_[25255]_ ;
  assign \new_[25260]_  = A301 & ~A300;
  assign \new_[25261]_  = ~A269 & \new_[25260]_ ;
  assign \new_[25262]_  = \new_[25261]_  & \new_[25256]_ ;
  assign \new_[25266]_  = A201 & ~A166;
  assign \new_[25267]_  = ~A167 & \new_[25266]_ ;
  assign \new_[25271]_  = A265 & ~A203;
  assign \new_[25272]_  = ~A202 & \new_[25271]_ ;
  assign \new_[25273]_  = \new_[25272]_  & \new_[25267]_ ;
  assign \new_[25277]_  = ~A268 & ~A267;
  assign \new_[25278]_  = ~A266 & \new_[25277]_ ;
  assign \new_[25282]_  = A302 & ~A300;
  assign \new_[25283]_  = ~A269 & \new_[25282]_ ;
  assign \new_[25284]_  = \new_[25283]_  & \new_[25278]_ ;
  assign \new_[25288]_  = A201 & ~A166;
  assign \new_[25289]_  = ~A167 & \new_[25288]_ ;
  assign \new_[25293]_  = A265 & ~A203;
  assign \new_[25294]_  = ~A202 & \new_[25293]_ ;
  assign \new_[25295]_  = \new_[25294]_  & \new_[25289]_ ;
  assign \new_[25299]_  = ~A268 & ~A267;
  assign \new_[25300]_  = ~A266 & \new_[25299]_ ;
  assign \new_[25304]_  = A299 & A298;
  assign \new_[25305]_  = ~A269 & \new_[25304]_ ;
  assign \new_[25306]_  = \new_[25305]_  & \new_[25300]_ ;
  assign \new_[25310]_  = A201 & ~A166;
  assign \new_[25311]_  = ~A167 & \new_[25310]_ ;
  assign \new_[25315]_  = A265 & ~A203;
  assign \new_[25316]_  = ~A202 & \new_[25315]_ ;
  assign \new_[25317]_  = \new_[25316]_  & \new_[25311]_ ;
  assign \new_[25321]_  = ~A268 & ~A267;
  assign \new_[25322]_  = ~A266 & \new_[25321]_ ;
  assign \new_[25326]_  = ~A299 & ~A298;
  assign \new_[25327]_  = ~A269 & \new_[25326]_ ;
  assign \new_[25328]_  = \new_[25327]_  & \new_[25322]_ ;
  assign \new_[25332]_  = ~A201 & ~A166;
  assign \new_[25333]_  = ~A167 & \new_[25332]_ ;
  assign \new_[25337]_  = A266 & ~A265;
  assign \new_[25338]_  = A202 & \new_[25337]_ ;
  assign \new_[25339]_  = \new_[25338]_  & \new_[25333]_ ;
  assign \new_[25343]_  = ~A269 & ~A268;
  assign \new_[25344]_  = ~A267 & \new_[25343]_ ;
  assign \new_[25348]_  = ~A302 & ~A301;
  assign \new_[25349]_  = A300 & \new_[25348]_ ;
  assign \new_[25350]_  = \new_[25349]_  & \new_[25344]_ ;
  assign \new_[25354]_  = ~A201 & ~A166;
  assign \new_[25355]_  = ~A167 & \new_[25354]_ ;
  assign \new_[25359]_  = ~A266 & A265;
  assign \new_[25360]_  = A202 & \new_[25359]_ ;
  assign \new_[25361]_  = \new_[25360]_  & \new_[25355]_ ;
  assign \new_[25365]_  = ~A269 & ~A268;
  assign \new_[25366]_  = ~A267 & \new_[25365]_ ;
  assign \new_[25370]_  = ~A302 & ~A301;
  assign \new_[25371]_  = A300 & \new_[25370]_ ;
  assign \new_[25372]_  = \new_[25371]_  & \new_[25366]_ ;
  assign \new_[25376]_  = ~A201 & ~A166;
  assign \new_[25377]_  = ~A167 & \new_[25376]_ ;
  assign \new_[25381]_  = A266 & ~A265;
  assign \new_[25382]_  = A203 & \new_[25381]_ ;
  assign \new_[25383]_  = \new_[25382]_  & \new_[25377]_ ;
  assign \new_[25387]_  = ~A269 & ~A268;
  assign \new_[25388]_  = ~A267 & \new_[25387]_ ;
  assign \new_[25392]_  = ~A302 & ~A301;
  assign \new_[25393]_  = A300 & \new_[25392]_ ;
  assign \new_[25394]_  = \new_[25393]_  & \new_[25388]_ ;
  assign \new_[25398]_  = ~A201 & ~A166;
  assign \new_[25399]_  = ~A167 & \new_[25398]_ ;
  assign \new_[25403]_  = ~A266 & A265;
  assign \new_[25404]_  = A203 & \new_[25403]_ ;
  assign \new_[25405]_  = \new_[25404]_  & \new_[25399]_ ;
  assign \new_[25409]_  = ~A269 & ~A268;
  assign \new_[25410]_  = ~A267 & \new_[25409]_ ;
  assign \new_[25414]_  = ~A302 & ~A301;
  assign \new_[25415]_  = A300 & \new_[25414]_ ;
  assign \new_[25416]_  = \new_[25415]_  & \new_[25410]_ ;
  assign \new_[25420]_  = A199 & ~A166;
  assign \new_[25421]_  = ~A167 & \new_[25420]_ ;
  assign \new_[25425]_  = A266 & ~A265;
  assign \new_[25426]_  = A200 & \new_[25425]_ ;
  assign \new_[25427]_  = \new_[25426]_  & \new_[25421]_ ;
  assign \new_[25431]_  = ~A269 & ~A268;
  assign \new_[25432]_  = ~A267 & \new_[25431]_ ;
  assign \new_[25436]_  = ~A302 & ~A301;
  assign \new_[25437]_  = A300 & \new_[25436]_ ;
  assign \new_[25438]_  = \new_[25437]_  & \new_[25432]_ ;
  assign \new_[25442]_  = A199 & ~A166;
  assign \new_[25443]_  = ~A167 & \new_[25442]_ ;
  assign \new_[25447]_  = ~A266 & A265;
  assign \new_[25448]_  = A200 & \new_[25447]_ ;
  assign \new_[25449]_  = \new_[25448]_  & \new_[25443]_ ;
  assign \new_[25453]_  = ~A269 & ~A268;
  assign \new_[25454]_  = ~A267 & \new_[25453]_ ;
  assign \new_[25458]_  = ~A302 & ~A301;
  assign \new_[25459]_  = A300 & \new_[25458]_ ;
  assign \new_[25460]_  = \new_[25459]_  & \new_[25454]_ ;
  assign \new_[25464]_  = ~A199 & ~A166;
  assign \new_[25465]_  = ~A167 & \new_[25464]_ ;
  assign \new_[25469]_  = A202 & A201;
  assign \new_[25470]_  = A200 & \new_[25469]_ ;
  assign \new_[25471]_  = \new_[25470]_  & \new_[25465]_ ;
  assign \new_[25475]_  = A298 & A268;
  assign \new_[25476]_  = ~A267 & \new_[25475]_ ;
  assign \new_[25480]_  = A301 & A300;
  assign \new_[25481]_  = ~A299 & \new_[25480]_ ;
  assign \new_[25482]_  = \new_[25481]_  & \new_[25476]_ ;
  assign \new_[25486]_  = ~A199 & ~A166;
  assign \new_[25487]_  = ~A167 & \new_[25486]_ ;
  assign \new_[25491]_  = A202 & A201;
  assign \new_[25492]_  = A200 & \new_[25491]_ ;
  assign \new_[25493]_  = \new_[25492]_  & \new_[25487]_ ;
  assign \new_[25497]_  = A298 & A268;
  assign \new_[25498]_  = ~A267 & \new_[25497]_ ;
  assign \new_[25502]_  = A302 & A300;
  assign \new_[25503]_  = ~A299 & \new_[25502]_ ;
  assign \new_[25504]_  = \new_[25503]_  & \new_[25498]_ ;
  assign \new_[25508]_  = ~A199 & ~A166;
  assign \new_[25509]_  = ~A167 & \new_[25508]_ ;
  assign \new_[25513]_  = A202 & A201;
  assign \new_[25514]_  = A200 & \new_[25513]_ ;
  assign \new_[25515]_  = \new_[25514]_  & \new_[25509]_ ;
  assign \new_[25519]_  = ~A298 & A268;
  assign \new_[25520]_  = ~A267 & \new_[25519]_ ;
  assign \new_[25524]_  = A301 & A300;
  assign \new_[25525]_  = A299 & \new_[25524]_ ;
  assign \new_[25526]_  = \new_[25525]_  & \new_[25520]_ ;
  assign \new_[25530]_  = ~A199 & ~A166;
  assign \new_[25531]_  = ~A167 & \new_[25530]_ ;
  assign \new_[25535]_  = A202 & A201;
  assign \new_[25536]_  = A200 & \new_[25535]_ ;
  assign \new_[25537]_  = \new_[25536]_  & \new_[25531]_ ;
  assign \new_[25541]_  = ~A298 & A268;
  assign \new_[25542]_  = ~A267 & \new_[25541]_ ;
  assign \new_[25546]_  = A302 & A300;
  assign \new_[25547]_  = A299 & \new_[25546]_ ;
  assign \new_[25548]_  = \new_[25547]_  & \new_[25542]_ ;
  assign \new_[25552]_  = ~A199 & ~A166;
  assign \new_[25553]_  = ~A167 & \new_[25552]_ ;
  assign \new_[25557]_  = A202 & A201;
  assign \new_[25558]_  = A200 & \new_[25557]_ ;
  assign \new_[25559]_  = \new_[25558]_  & \new_[25553]_ ;
  assign \new_[25563]_  = A298 & A269;
  assign \new_[25564]_  = ~A267 & \new_[25563]_ ;
  assign \new_[25568]_  = A301 & A300;
  assign \new_[25569]_  = ~A299 & \new_[25568]_ ;
  assign \new_[25570]_  = \new_[25569]_  & \new_[25564]_ ;
  assign \new_[25574]_  = ~A199 & ~A166;
  assign \new_[25575]_  = ~A167 & \new_[25574]_ ;
  assign \new_[25579]_  = A202 & A201;
  assign \new_[25580]_  = A200 & \new_[25579]_ ;
  assign \new_[25581]_  = \new_[25580]_  & \new_[25575]_ ;
  assign \new_[25585]_  = A298 & A269;
  assign \new_[25586]_  = ~A267 & \new_[25585]_ ;
  assign \new_[25590]_  = A302 & A300;
  assign \new_[25591]_  = ~A299 & \new_[25590]_ ;
  assign \new_[25592]_  = \new_[25591]_  & \new_[25586]_ ;
  assign \new_[25596]_  = ~A199 & ~A166;
  assign \new_[25597]_  = ~A167 & \new_[25596]_ ;
  assign \new_[25601]_  = A202 & A201;
  assign \new_[25602]_  = A200 & \new_[25601]_ ;
  assign \new_[25603]_  = \new_[25602]_  & \new_[25597]_ ;
  assign \new_[25607]_  = ~A298 & A269;
  assign \new_[25608]_  = ~A267 & \new_[25607]_ ;
  assign \new_[25612]_  = A301 & A300;
  assign \new_[25613]_  = A299 & \new_[25612]_ ;
  assign \new_[25614]_  = \new_[25613]_  & \new_[25608]_ ;
  assign \new_[25618]_  = ~A199 & ~A166;
  assign \new_[25619]_  = ~A167 & \new_[25618]_ ;
  assign \new_[25623]_  = A202 & A201;
  assign \new_[25624]_  = A200 & \new_[25623]_ ;
  assign \new_[25625]_  = \new_[25624]_  & \new_[25619]_ ;
  assign \new_[25629]_  = ~A298 & A269;
  assign \new_[25630]_  = ~A267 & \new_[25629]_ ;
  assign \new_[25634]_  = A302 & A300;
  assign \new_[25635]_  = A299 & \new_[25634]_ ;
  assign \new_[25636]_  = \new_[25635]_  & \new_[25630]_ ;
  assign \new_[25640]_  = ~A199 & ~A166;
  assign \new_[25641]_  = ~A167 & \new_[25640]_ ;
  assign \new_[25645]_  = A202 & A201;
  assign \new_[25646]_  = A200 & \new_[25645]_ ;
  assign \new_[25647]_  = \new_[25646]_  & \new_[25641]_ ;
  assign \new_[25651]_  = A298 & A266;
  assign \new_[25652]_  = A265 & \new_[25651]_ ;
  assign \new_[25656]_  = A301 & A300;
  assign \new_[25657]_  = ~A299 & \new_[25656]_ ;
  assign \new_[25658]_  = \new_[25657]_  & \new_[25652]_ ;
  assign \new_[25662]_  = ~A199 & ~A166;
  assign \new_[25663]_  = ~A167 & \new_[25662]_ ;
  assign \new_[25667]_  = A202 & A201;
  assign \new_[25668]_  = A200 & \new_[25667]_ ;
  assign \new_[25669]_  = \new_[25668]_  & \new_[25663]_ ;
  assign \new_[25673]_  = A298 & A266;
  assign \new_[25674]_  = A265 & \new_[25673]_ ;
  assign \new_[25678]_  = A302 & A300;
  assign \new_[25679]_  = ~A299 & \new_[25678]_ ;
  assign \new_[25680]_  = \new_[25679]_  & \new_[25674]_ ;
  assign \new_[25684]_  = ~A199 & ~A166;
  assign \new_[25685]_  = ~A167 & \new_[25684]_ ;
  assign \new_[25689]_  = A202 & A201;
  assign \new_[25690]_  = A200 & \new_[25689]_ ;
  assign \new_[25691]_  = \new_[25690]_  & \new_[25685]_ ;
  assign \new_[25695]_  = ~A298 & A266;
  assign \new_[25696]_  = A265 & \new_[25695]_ ;
  assign \new_[25700]_  = A301 & A300;
  assign \new_[25701]_  = A299 & \new_[25700]_ ;
  assign \new_[25702]_  = \new_[25701]_  & \new_[25696]_ ;
  assign \new_[25706]_  = ~A199 & ~A166;
  assign \new_[25707]_  = ~A167 & \new_[25706]_ ;
  assign \new_[25711]_  = A202 & A201;
  assign \new_[25712]_  = A200 & \new_[25711]_ ;
  assign \new_[25713]_  = \new_[25712]_  & \new_[25707]_ ;
  assign \new_[25717]_  = ~A298 & A266;
  assign \new_[25718]_  = A265 & \new_[25717]_ ;
  assign \new_[25722]_  = A302 & A300;
  assign \new_[25723]_  = A299 & \new_[25722]_ ;
  assign \new_[25724]_  = \new_[25723]_  & \new_[25718]_ ;
  assign \new_[25728]_  = ~A199 & ~A166;
  assign \new_[25729]_  = ~A167 & \new_[25728]_ ;
  assign \new_[25733]_  = A202 & A201;
  assign \new_[25734]_  = A200 & \new_[25733]_ ;
  assign \new_[25735]_  = \new_[25734]_  & \new_[25729]_ ;
  assign \new_[25739]_  = A298 & ~A266;
  assign \new_[25740]_  = ~A265 & \new_[25739]_ ;
  assign \new_[25744]_  = A301 & A300;
  assign \new_[25745]_  = ~A299 & \new_[25744]_ ;
  assign \new_[25746]_  = \new_[25745]_  & \new_[25740]_ ;
  assign \new_[25750]_  = ~A199 & ~A166;
  assign \new_[25751]_  = ~A167 & \new_[25750]_ ;
  assign \new_[25755]_  = A202 & A201;
  assign \new_[25756]_  = A200 & \new_[25755]_ ;
  assign \new_[25757]_  = \new_[25756]_  & \new_[25751]_ ;
  assign \new_[25761]_  = A298 & ~A266;
  assign \new_[25762]_  = ~A265 & \new_[25761]_ ;
  assign \new_[25766]_  = A302 & A300;
  assign \new_[25767]_  = ~A299 & \new_[25766]_ ;
  assign \new_[25768]_  = \new_[25767]_  & \new_[25762]_ ;
  assign \new_[25772]_  = ~A199 & ~A166;
  assign \new_[25773]_  = ~A167 & \new_[25772]_ ;
  assign \new_[25777]_  = A202 & A201;
  assign \new_[25778]_  = A200 & \new_[25777]_ ;
  assign \new_[25779]_  = \new_[25778]_  & \new_[25773]_ ;
  assign \new_[25783]_  = ~A298 & ~A266;
  assign \new_[25784]_  = ~A265 & \new_[25783]_ ;
  assign \new_[25788]_  = A301 & A300;
  assign \new_[25789]_  = A299 & \new_[25788]_ ;
  assign \new_[25790]_  = \new_[25789]_  & \new_[25784]_ ;
  assign \new_[25794]_  = ~A199 & ~A166;
  assign \new_[25795]_  = ~A167 & \new_[25794]_ ;
  assign \new_[25799]_  = A202 & A201;
  assign \new_[25800]_  = A200 & \new_[25799]_ ;
  assign \new_[25801]_  = \new_[25800]_  & \new_[25795]_ ;
  assign \new_[25805]_  = ~A298 & ~A266;
  assign \new_[25806]_  = ~A265 & \new_[25805]_ ;
  assign \new_[25810]_  = A302 & A300;
  assign \new_[25811]_  = A299 & \new_[25810]_ ;
  assign \new_[25812]_  = \new_[25811]_  & \new_[25806]_ ;
  assign \new_[25816]_  = ~A199 & ~A166;
  assign \new_[25817]_  = ~A167 & \new_[25816]_ ;
  assign \new_[25821]_  = A203 & A201;
  assign \new_[25822]_  = A200 & \new_[25821]_ ;
  assign \new_[25823]_  = \new_[25822]_  & \new_[25817]_ ;
  assign \new_[25827]_  = A298 & A268;
  assign \new_[25828]_  = ~A267 & \new_[25827]_ ;
  assign \new_[25832]_  = A301 & A300;
  assign \new_[25833]_  = ~A299 & \new_[25832]_ ;
  assign \new_[25834]_  = \new_[25833]_  & \new_[25828]_ ;
  assign \new_[25838]_  = ~A199 & ~A166;
  assign \new_[25839]_  = ~A167 & \new_[25838]_ ;
  assign \new_[25843]_  = A203 & A201;
  assign \new_[25844]_  = A200 & \new_[25843]_ ;
  assign \new_[25845]_  = \new_[25844]_  & \new_[25839]_ ;
  assign \new_[25849]_  = A298 & A268;
  assign \new_[25850]_  = ~A267 & \new_[25849]_ ;
  assign \new_[25854]_  = A302 & A300;
  assign \new_[25855]_  = ~A299 & \new_[25854]_ ;
  assign \new_[25856]_  = \new_[25855]_  & \new_[25850]_ ;
  assign \new_[25860]_  = ~A199 & ~A166;
  assign \new_[25861]_  = ~A167 & \new_[25860]_ ;
  assign \new_[25865]_  = A203 & A201;
  assign \new_[25866]_  = A200 & \new_[25865]_ ;
  assign \new_[25867]_  = \new_[25866]_  & \new_[25861]_ ;
  assign \new_[25871]_  = ~A298 & A268;
  assign \new_[25872]_  = ~A267 & \new_[25871]_ ;
  assign \new_[25876]_  = A301 & A300;
  assign \new_[25877]_  = A299 & \new_[25876]_ ;
  assign \new_[25878]_  = \new_[25877]_  & \new_[25872]_ ;
  assign \new_[25882]_  = ~A199 & ~A166;
  assign \new_[25883]_  = ~A167 & \new_[25882]_ ;
  assign \new_[25887]_  = A203 & A201;
  assign \new_[25888]_  = A200 & \new_[25887]_ ;
  assign \new_[25889]_  = \new_[25888]_  & \new_[25883]_ ;
  assign \new_[25893]_  = ~A298 & A268;
  assign \new_[25894]_  = ~A267 & \new_[25893]_ ;
  assign \new_[25898]_  = A302 & A300;
  assign \new_[25899]_  = A299 & \new_[25898]_ ;
  assign \new_[25900]_  = \new_[25899]_  & \new_[25894]_ ;
  assign \new_[25904]_  = ~A199 & ~A166;
  assign \new_[25905]_  = ~A167 & \new_[25904]_ ;
  assign \new_[25909]_  = A203 & A201;
  assign \new_[25910]_  = A200 & \new_[25909]_ ;
  assign \new_[25911]_  = \new_[25910]_  & \new_[25905]_ ;
  assign \new_[25915]_  = A298 & A269;
  assign \new_[25916]_  = ~A267 & \new_[25915]_ ;
  assign \new_[25920]_  = A301 & A300;
  assign \new_[25921]_  = ~A299 & \new_[25920]_ ;
  assign \new_[25922]_  = \new_[25921]_  & \new_[25916]_ ;
  assign \new_[25926]_  = ~A199 & ~A166;
  assign \new_[25927]_  = ~A167 & \new_[25926]_ ;
  assign \new_[25931]_  = A203 & A201;
  assign \new_[25932]_  = A200 & \new_[25931]_ ;
  assign \new_[25933]_  = \new_[25932]_  & \new_[25927]_ ;
  assign \new_[25937]_  = A298 & A269;
  assign \new_[25938]_  = ~A267 & \new_[25937]_ ;
  assign \new_[25942]_  = A302 & A300;
  assign \new_[25943]_  = ~A299 & \new_[25942]_ ;
  assign \new_[25944]_  = \new_[25943]_  & \new_[25938]_ ;
  assign \new_[25948]_  = ~A199 & ~A166;
  assign \new_[25949]_  = ~A167 & \new_[25948]_ ;
  assign \new_[25953]_  = A203 & A201;
  assign \new_[25954]_  = A200 & \new_[25953]_ ;
  assign \new_[25955]_  = \new_[25954]_  & \new_[25949]_ ;
  assign \new_[25959]_  = ~A298 & A269;
  assign \new_[25960]_  = ~A267 & \new_[25959]_ ;
  assign \new_[25964]_  = A301 & A300;
  assign \new_[25965]_  = A299 & \new_[25964]_ ;
  assign \new_[25966]_  = \new_[25965]_  & \new_[25960]_ ;
  assign \new_[25970]_  = ~A199 & ~A166;
  assign \new_[25971]_  = ~A167 & \new_[25970]_ ;
  assign \new_[25975]_  = A203 & A201;
  assign \new_[25976]_  = A200 & \new_[25975]_ ;
  assign \new_[25977]_  = \new_[25976]_  & \new_[25971]_ ;
  assign \new_[25981]_  = ~A298 & A269;
  assign \new_[25982]_  = ~A267 & \new_[25981]_ ;
  assign \new_[25986]_  = A302 & A300;
  assign \new_[25987]_  = A299 & \new_[25986]_ ;
  assign \new_[25988]_  = \new_[25987]_  & \new_[25982]_ ;
  assign \new_[25992]_  = ~A199 & ~A166;
  assign \new_[25993]_  = ~A167 & \new_[25992]_ ;
  assign \new_[25997]_  = A203 & A201;
  assign \new_[25998]_  = A200 & \new_[25997]_ ;
  assign \new_[25999]_  = \new_[25998]_  & \new_[25993]_ ;
  assign \new_[26003]_  = A298 & A266;
  assign \new_[26004]_  = A265 & \new_[26003]_ ;
  assign \new_[26008]_  = A301 & A300;
  assign \new_[26009]_  = ~A299 & \new_[26008]_ ;
  assign \new_[26010]_  = \new_[26009]_  & \new_[26004]_ ;
  assign \new_[26014]_  = ~A199 & ~A166;
  assign \new_[26015]_  = ~A167 & \new_[26014]_ ;
  assign \new_[26019]_  = A203 & A201;
  assign \new_[26020]_  = A200 & \new_[26019]_ ;
  assign \new_[26021]_  = \new_[26020]_  & \new_[26015]_ ;
  assign \new_[26025]_  = A298 & A266;
  assign \new_[26026]_  = A265 & \new_[26025]_ ;
  assign \new_[26030]_  = A302 & A300;
  assign \new_[26031]_  = ~A299 & \new_[26030]_ ;
  assign \new_[26032]_  = \new_[26031]_  & \new_[26026]_ ;
  assign \new_[26036]_  = ~A199 & ~A166;
  assign \new_[26037]_  = ~A167 & \new_[26036]_ ;
  assign \new_[26041]_  = A203 & A201;
  assign \new_[26042]_  = A200 & \new_[26041]_ ;
  assign \new_[26043]_  = \new_[26042]_  & \new_[26037]_ ;
  assign \new_[26047]_  = ~A298 & A266;
  assign \new_[26048]_  = A265 & \new_[26047]_ ;
  assign \new_[26052]_  = A301 & A300;
  assign \new_[26053]_  = A299 & \new_[26052]_ ;
  assign \new_[26054]_  = \new_[26053]_  & \new_[26048]_ ;
  assign \new_[26058]_  = ~A199 & ~A166;
  assign \new_[26059]_  = ~A167 & \new_[26058]_ ;
  assign \new_[26063]_  = A203 & A201;
  assign \new_[26064]_  = A200 & \new_[26063]_ ;
  assign \new_[26065]_  = \new_[26064]_  & \new_[26059]_ ;
  assign \new_[26069]_  = ~A298 & A266;
  assign \new_[26070]_  = A265 & \new_[26069]_ ;
  assign \new_[26074]_  = A302 & A300;
  assign \new_[26075]_  = A299 & \new_[26074]_ ;
  assign \new_[26076]_  = \new_[26075]_  & \new_[26070]_ ;
  assign \new_[26080]_  = ~A199 & ~A166;
  assign \new_[26081]_  = ~A167 & \new_[26080]_ ;
  assign \new_[26085]_  = A203 & A201;
  assign \new_[26086]_  = A200 & \new_[26085]_ ;
  assign \new_[26087]_  = \new_[26086]_  & \new_[26081]_ ;
  assign \new_[26091]_  = A298 & ~A266;
  assign \new_[26092]_  = ~A265 & \new_[26091]_ ;
  assign \new_[26096]_  = A301 & A300;
  assign \new_[26097]_  = ~A299 & \new_[26096]_ ;
  assign \new_[26098]_  = \new_[26097]_  & \new_[26092]_ ;
  assign \new_[26102]_  = ~A199 & ~A166;
  assign \new_[26103]_  = ~A167 & \new_[26102]_ ;
  assign \new_[26107]_  = A203 & A201;
  assign \new_[26108]_  = A200 & \new_[26107]_ ;
  assign \new_[26109]_  = \new_[26108]_  & \new_[26103]_ ;
  assign \new_[26113]_  = A298 & ~A266;
  assign \new_[26114]_  = ~A265 & \new_[26113]_ ;
  assign \new_[26118]_  = A302 & A300;
  assign \new_[26119]_  = ~A299 & \new_[26118]_ ;
  assign \new_[26120]_  = \new_[26119]_  & \new_[26114]_ ;
  assign \new_[26124]_  = ~A199 & ~A166;
  assign \new_[26125]_  = ~A167 & \new_[26124]_ ;
  assign \new_[26129]_  = A203 & A201;
  assign \new_[26130]_  = A200 & \new_[26129]_ ;
  assign \new_[26131]_  = \new_[26130]_  & \new_[26125]_ ;
  assign \new_[26135]_  = ~A298 & ~A266;
  assign \new_[26136]_  = ~A265 & \new_[26135]_ ;
  assign \new_[26140]_  = A301 & A300;
  assign \new_[26141]_  = A299 & \new_[26140]_ ;
  assign \new_[26142]_  = \new_[26141]_  & \new_[26136]_ ;
  assign \new_[26146]_  = ~A199 & ~A166;
  assign \new_[26147]_  = ~A167 & \new_[26146]_ ;
  assign \new_[26151]_  = A203 & A201;
  assign \new_[26152]_  = A200 & \new_[26151]_ ;
  assign \new_[26153]_  = \new_[26152]_  & \new_[26147]_ ;
  assign \new_[26157]_  = ~A298 & ~A266;
  assign \new_[26158]_  = ~A265 & \new_[26157]_ ;
  assign \new_[26162]_  = A302 & A300;
  assign \new_[26163]_  = A299 & \new_[26162]_ ;
  assign \new_[26164]_  = \new_[26163]_  & \new_[26158]_ ;
  assign \new_[26168]_  = A199 & ~A166;
  assign \new_[26169]_  = ~A167 & \new_[26168]_ ;
  assign \new_[26173]_  = A202 & A201;
  assign \new_[26174]_  = ~A200 & \new_[26173]_ ;
  assign \new_[26175]_  = \new_[26174]_  & \new_[26169]_ ;
  assign \new_[26179]_  = A298 & A268;
  assign \new_[26180]_  = ~A267 & \new_[26179]_ ;
  assign \new_[26184]_  = A301 & A300;
  assign \new_[26185]_  = ~A299 & \new_[26184]_ ;
  assign \new_[26186]_  = \new_[26185]_  & \new_[26180]_ ;
  assign \new_[26190]_  = A199 & ~A166;
  assign \new_[26191]_  = ~A167 & \new_[26190]_ ;
  assign \new_[26195]_  = A202 & A201;
  assign \new_[26196]_  = ~A200 & \new_[26195]_ ;
  assign \new_[26197]_  = \new_[26196]_  & \new_[26191]_ ;
  assign \new_[26201]_  = A298 & A268;
  assign \new_[26202]_  = ~A267 & \new_[26201]_ ;
  assign \new_[26206]_  = A302 & A300;
  assign \new_[26207]_  = ~A299 & \new_[26206]_ ;
  assign \new_[26208]_  = \new_[26207]_  & \new_[26202]_ ;
  assign \new_[26212]_  = A199 & ~A166;
  assign \new_[26213]_  = ~A167 & \new_[26212]_ ;
  assign \new_[26217]_  = A202 & A201;
  assign \new_[26218]_  = ~A200 & \new_[26217]_ ;
  assign \new_[26219]_  = \new_[26218]_  & \new_[26213]_ ;
  assign \new_[26223]_  = ~A298 & A268;
  assign \new_[26224]_  = ~A267 & \new_[26223]_ ;
  assign \new_[26228]_  = A301 & A300;
  assign \new_[26229]_  = A299 & \new_[26228]_ ;
  assign \new_[26230]_  = \new_[26229]_  & \new_[26224]_ ;
  assign \new_[26234]_  = A199 & ~A166;
  assign \new_[26235]_  = ~A167 & \new_[26234]_ ;
  assign \new_[26239]_  = A202 & A201;
  assign \new_[26240]_  = ~A200 & \new_[26239]_ ;
  assign \new_[26241]_  = \new_[26240]_  & \new_[26235]_ ;
  assign \new_[26245]_  = ~A298 & A268;
  assign \new_[26246]_  = ~A267 & \new_[26245]_ ;
  assign \new_[26250]_  = A302 & A300;
  assign \new_[26251]_  = A299 & \new_[26250]_ ;
  assign \new_[26252]_  = \new_[26251]_  & \new_[26246]_ ;
  assign \new_[26256]_  = A199 & ~A166;
  assign \new_[26257]_  = ~A167 & \new_[26256]_ ;
  assign \new_[26261]_  = A202 & A201;
  assign \new_[26262]_  = ~A200 & \new_[26261]_ ;
  assign \new_[26263]_  = \new_[26262]_  & \new_[26257]_ ;
  assign \new_[26267]_  = A298 & A269;
  assign \new_[26268]_  = ~A267 & \new_[26267]_ ;
  assign \new_[26272]_  = A301 & A300;
  assign \new_[26273]_  = ~A299 & \new_[26272]_ ;
  assign \new_[26274]_  = \new_[26273]_  & \new_[26268]_ ;
  assign \new_[26278]_  = A199 & ~A166;
  assign \new_[26279]_  = ~A167 & \new_[26278]_ ;
  assign \new_[26283]_  = A202 & A201;
  assign \new_[26284]_  = ~A200 & \new_[26283]_ ;
  assign \new_[26285]_  = \new_[26284]_  & \new_[26279]_ ;
  assign \new_[26289]_  = A298 & A269;
  assign \new_[26290]_  = ~A267 & \new_[26289]_ ;
  assign \new_[26294]_  = A302 & A300;
  assign \new_[26295]_  = ~A299 & \new_[26294]_ ;
  assign \new_[26296]_  = \new_[26295]_  & \new_[26290]_ ;
  assign \new_[26300]_  = A199 & ~A166;
  assign \new_[26301]_  = ~A167 & \new_[26300]_ ;
  assign \new_[26305]_  = A202 & A201;
  assign \new_[26306]_  = ~A200 & \new_[26305]_ ;
  assign \new_[26307]_  = \new_[26306]_  & \new_[26301]_ ;
  assign \new_[26311]_  = ~A298 & A269;
  assign \new_[26312]_  = ~A267 & \new_[26311]_ ;
  assign \new_[26316]_  = A301 & A300;
  assign \new_[26317]_  = A299 & \new_[26316]_ ;
  assign \new_[26318]_  = \new_[26317]_  & \new_[26312]_ ;
  assign \new_[26322]_  = A199 & ~A166;
  assign \new_[26323]_  = ~A167 & \new_[26322]_ ;
  assign \new_[26327]_  = A202 & A201;
  assign \new_[26328]_  = ~A200 & \new_[26327]_ ;
  assign \new_[26329]_  = \new_[26328]_  & \new_[26323]_ ;
  assign \new_[26333]_  = ~A298 & A269;
  assign \new_[26334]_  = ~A267 & \new_[26333]_ ;
  assign \new_[26338]_  = A302 & A300;
  assign \new_[26339]_  = A299 & \new_[26338]_ ;
  assign \new_[26340]_  = \new_[26339]_  & \new_[26334]_ ;
  assign \new_[26344]_  = A199 & ~A166;
  assign \new_[26345]_  = ~A167 & \new_[26344]_ ;
  assign \new_[26349]_  = A202 & A201;
  assign \new_[26350]_  = ~A200 & \new_[26349]_ ;
  assign \new_[26351]_  = \new_[26350]_  & \new_[26345]_ ;
  assign \new_[26355]_  = A298 & A266;
  assign \new_[26356]_  = A265 & \new_[26355]_ ;
  assign \new_[26360]_  = A301 & A300;
  assign \new_[26361]_  = ~A299 & \new_[26360]_ ;
  assign \new_[26362]_  = \new_[26361]_  & \new_[26356]_ ;
  assign \new_[26366]_  = A199 & ~A166;
  assign \new_[26367]_  = ~A167 & \new_[26366]_ ;
  assign \new_[26371]_  = A202 & A201;
  assign \new_[26372]_  = ~A200 & \new_[26371]_ ;
  assign \new_[26373]_  = \new_[26372]_  & \new_[26367]_ ;
  assign \new_[26377]_  = A298 & A266;
  assign \new_[26378]_  = A265 & \new_[26377]_ ;
  assign \new_[26382]_  = A302 & A300;
  assign \new_[26383]_  = ~A299 & \new_[26382]_ ;
  assign \new_[26384]_  = \new_[26383]_  & \new_[26378]_ ;
  assign \new_[26388]_  = A199 & ~A166;
  assign \new_[26389]_  = ~A167 & \new_[26388]_ ;
  assign \new_[26393]_  = A202 & A201;
  assign \new_[26394]_  = ~A200 & \new_[26393]_ ;
  assign \new_[26395]_  = \new_[26394]_  & \new_[26389]_ ;
  assign \new_[26399]_  = ~A298 & A266;
  assign \new_[26400]_  = A265 & \new_[26399]_ ;
  assign \new_[26404]_  = A301 & A300;
  assign \new_[26405]_  = A299 & \new_[26404]_ ;
  assign \new_[26406]_  = \new_[26405]_  & \new_[26400]_ ;
  assign \new_[26410]_  = A199 & ~A166;
  assign \new_[26411]_  = ~A167 & \new_[26410]_ ;
  assign \new_[26415]_  = A202 & A201;
  assign \new_[26416]_  = ~A200 & \new_[26415]_ ;
  assign \new_[26417]_  = \new_[26416]_  & \new_[26411]_ ;
  assign \new_[26421]_  = ~A298 & A266;
  assign \new_[26422]_  = A265 & \new_[26421]_ ;
  assign \new_[26426]_  = A302 & A300;
  assign \new_[26427]_  = A299 & \new_[26426]_ ;
  assign \new_[26428]_  = \new_[26427]_  & \new_[26422]_ ;
  assign \new_[26432]_  = A199 & ~A166;
  assign \new_[26433]_  = ~A167 & \new_[26432]_ ;
  assign \new_[26437]_  = A202 & A201;
  assign \new_[26438]_  = ~A200 & \new_[26437]_ ;
  assign \new_[26439]_  = \new_[26438]_  & \new_[26433]_ ;
  assign \new_[26443]_  = A298 & ~A266;
  assign \new_[26444]_  = ~A265 & \new_[26443]_ ;
  assign \new_[26448]_  = A301 & A300;
  assign \new_[26449]_  = ~A299 & \new_[26448]_ ;
  assign \new_[26450]_  = \new_[26449]_  & \new_[26444]_ ;
  assign \new_[26454]_  = A199 & ~A166;
  assign \new_[26455]_  = ~A167 & \new_[26454]_ ;
  assign \new_[26459]_  = A202 & A201;
  assign \new_[26460]_  = ~A200 & \new_[26459]_ ;
  assign \new_[26461]_  = \new_[26460]_  & \new_[26455]_ ;
  assign \new_[26465]_  = A298 & ~A266;
  assign \new_[26466]_  = ~A265 & \new_[26465]_ ;
  assign \new_[26470]_  = A302 & A300;
  assign \new_[26471]_  = ~A299 & \new_[26470]_ ;
  assign \new_[26472]_  = \new_[26471]_  & \new_[26466]_ ;
  assign \new_[26476]_  = A199 & ~A166;
  assign \new_[26477]_  = ~A167 & \new_[26476]_ ;
  assign \new_[26481]_  = A202 & A201;
  assign \new_[26482]_  = ~A200 & \new_[26481]_ ;
  assign \new_[26483]_  = \new_[26482]_  & \new_[26477]_ ;
  assign \new_[26487]_  = ~A298 & ~A266;
  assign \new_[26488]_  = ~A265 & \new_[26487]_ ;
  assign \new_[26492]_  = A301 & A300;
  assign \new_[26493]_  = A299 & \new_[26492]_ ;
  assign \new_[26494]_  = \new_[26493]_  & \new_[26488]_ ;
  assign \new_[26498]_  = A199 & ~A166;
  assign \new_[26499]_  = ~A167 & \new_[26498]_ ;
  assign \new_[26503]_  = A202 & A201;
  assign \new_[26504]_  = ~A200 & \new_[26503]_ ;
  assign \new_[26505]_  = \new_[26504]_  & \new_[26499]_ ;
  assign \new_[26509]_  = ~A298 & ~A266;
  assign \new_[26510]_  = ~A265 & \new_[26509]_ ;
  assign \new_[26514]_  = A302 & A300;
  assign \new_[26515]_  = A299 & \new_[26514]_ ;
  assign \new_[26516]_  = \new_[26515]_  & \new_[26510]_ ;
  assign \new_[26520]_  = A199 & ~A166;
  assign \new_[26521]_  = ~A167 & \new_[26520]_ ;
  assign \new_[26525]_  = A203 & A201;
  assign \new_[26526]_  = ~A200 & \new_[26525]_ ;
  assign \new_[26527]_  = \new_[26526]_  & \new_[26521]_ ;
  assign \new_[26531]_  = A298 & A268;
  assign \new_[26532]_  = ~A267 & \new_[26531]_ ;
  assign \new_[26536]_  = A301 & A300;
  assign \new_[26537]_  = ~A299 & \new_[26536]_ ;
  assign \new_[26538]_  = \new_[26537]_  & \new_[26532]_ ;
  assign \new_[26542]_  = A199 & ~A166;
  assign \new_[26543]_  = ~A167 & \new_[26542]_ ;
  assign \new_[26547]_  = A203 & A201;
  assign \new_[26548]_  = ~A200 & \new_[26547]_ ;
  assign \new_[26549]_  = \new_[26548]_  & \new_[26543]_ ;
  assign \new_[26553]_  = A298 & A268;
  assign \new_[26554]_  = ~A267 & \new_[26553]_ ;
  assign \new_[26558]_  = A302 & A300;
  assign \new_[26559]_  = ~A299 & \new_[26558]_ ;
  assign \new_[26560]_  = \new_[26559]_  & \new_[26554]_ ;
  assign \new_[26564]_  = A199 & ~A166;
  assign \new_[26565]_  = ~A167 & \new_[26564]_ ;
  assign \new_[26569]_  = A203 & A201;
  assign \new_[26570]_  = ~A200 & \new_[26569]_ ;
  assign \new_[26571]_  = \new_[26570]_  & \new_[26565]_ ;
  assign \new_[26575]_  = ~A298 & A268;
  assign \new_[26576]_  = ~A267 & \new_[26575]_ ;
  assign \new_[26580]_  = A301 & A300;
  assign \new_[26581]_  = A299 & \new_[26580]_ ;
  assign \new_[26582]_  = \new_[26581]_  & \new_[26576]_ ;
  assign \new_[26586]_  = A199 & ~A166;
  assign \new_[26587]_  = ~A167 & \new_[26586]_ ;
  assign \new_[26591]_  = A203 & A201;
  assign \new_[26592]_  = ~A200 & \new_[26591]_ ;
  assign \new_[26593]_  = \new_[26592]_  & \new_[26587]_ ;
  assign \new_[26597]_  = ~A298 & A268;
  assign \new_[26598]_  = ~A267 & \new_[26597]_ ;
  assign \new_[26602]_  = A302 & A300;
  assign \new_[26603]_  = A299 & \new_[26602]_ ;
  assign \new_[26604]_  = \new_[26603]_  & \new_[26598]_ ;
  assign \new_[26608]_  = A199 & ~A166;
  assign \new_[26609]_  = ~A167 & \new_[26608]_ ;
  assign \new_[26613]_  = A203 & A201;
  assign \new_[26614]_  = ~A200 & \new_[26613]_ ;
  assign \new_[26615]_  = \new_[26614]_  & \new_[26609]_ ;
  assign \new_[26619]_  = A298 & A269;
  assign \new_[26620]_  = ~A267 & \new_[26619]_ ;
  assign \new_[26624]_  = A301 & A300;
  assign \new_[26625]_  = ~A299 & \new_[26624]_ ;
  assign \new_[26626]_  = \new_[26625]_  & \new_[26620]_ ;
  assign \new_[26630]_  = A199 & ~A166;
  assign \new_[26631]_  = ~A167 & \new_[26630]_ ;
  assign \new_[26635]_  = A203 & A201;
  assign \new_[26636]_  = ~A200 & \new_[26635]_ ;
  assign \new_[26637]_  = \new_[26636]_  & \new_[26631]_ ;
  assign \new_[26641]_  = A298 & A269;
  assign \new_[26642]_  = ~A267 & \new_[26641]_ ;
  assign \new_[26646]_  = A302 & A300;
  assign \new_[26647]_  = ~A299 & \new_[26646]_ ;
  assign \new_[26648]_  = \new_[26647]_  & \new_[26642]_ ;
  assign \new_[26652]_  = A199 & ~A166;
  assign \new_[26653]_  = ~A167 & \new_[26652]_ ;
  assign \new_[26657]_  = A203 & A201;
  assign \new_[26658]_  = ~A200 & \new_[26657]_ ;
  assign \new_[26659]_  = \new_[26658]_  & \new_[26653]_ ;
  assign \new_[26663]_  = ~A298 & A269;
  assign \new_[26664]_  = ~A267 & \new_[26663]_ ;
  assign \new_[26668]_  = A301 & A300;
  assign \new_[26669]_  = A299 & \new_[26668]_ ;
  assign \new_[26670]_  = \new_[26669]_  & \new_[26664]_ ;
  assign \new_[26674]_  = A199 & ~A166;
  assign \new_[26675]_  = ~A167 & \new_[26674]_ ;
  assign \new_[26679]_  = A203 & A201;
  assign \new_[26680]_  = ~A200 & \new_[26679]_ ;
  assign \new_[26681]_  = \new_[26680]_  & \new_[26675]_ ;
  assign \new_[26685]_  = ~A298 & A269;
  assign \new_[26686]_  = ~A267 & \new_[26685]_ ;
  assign \new_[26690]_  = A302 & A300;
  assign \new_[26691]_  = A299 & \new_[26690]_ ;
  assign \new_[26692]_  = \new_[26691]_  & \new_[26686]_ ;
  assign \new_[26696]_  = A199 & ~A166;
  assign \new_[26697]_  = ~A167 & \new_[26696]_ ;
  assign \new_[26701]_  = A203 & A201;
  assign \new_[26702]_  = ~A200 & \new_[26701]_ ;
  assign \new_[26703]_  = \new_[26702]_  & \new_[26697]_ ;
  assign \new_[26707]_  = A298 & A266;
  assign \new_[26708]_  = A265 & \new_[26707]_ ;
  assign \new_[26712]_  = A301 & A300;
  assign \new_[26713]_  = ~A299 & \new_[26712]_ ;
  assign \new_[26714]_  = \new_[26713]_  & \new_[26708]_ ;
  assign \new_[26718]_  = A199 & ~A166;
  assign \new_[26719]_  = ~A167 & \new_[26718]_ ;
  assign \new_[26723]_  = A203 & A201;
  assign \new_[26724]_  = ~A200 & \new_[26723]_ ;
  assign \new_[26725]_  = \new_[26724]_  & \new_[26719]_ ;
  assign \new_[26729]_  = A298 & A266;
  assign \new_[26730]_  = A265 & \new_[26729]_ ;
  assign \new_[26734]_  = A302 & A300;
  assign \new_[26735]_  = ~A299 & \new_[26734]_ ;
  assign \new_[26736]_  = \new_[26735]_  & \new_[26730]_ ;
  assign \new_[26740]_  = A199 & ~A166;
  assign \new_[26741]_  = ~A167 & \new_[26740]_ ;
  assign \new_[26745]_  = A203 & A201;
  assign \new_[26746]_  = ~A200 & \new_[26745]_ ;
  assign \new_[26747]_  = \new_[26746]_  & \new_[26741]_ ;
  assign \new_[26751]_  = ~A298 & A266;
  assign \new_[26752]_  = A265 & \new_[26751]_ ;
  assign \new_[26756]_  = A301 & A300;
  assign \new_[26757]_  = A299 & \new_[26756]_ ;
  assign \new_[26758]_  = \new_[26757]_  & \new_[26752]_ ;
  assign \new_[26762]_  = A199 & ~A166;
  assign \new_[26763]_  = ~A167 & \new_[26762]_ ;
  assign \new_[26767]_  = A203 & A201;
  assign \new_[26768]_  = ~A200 & \new_[26767]_ ;
  assign \new_[26769]_  = \new_[26768]_  & \new_[26763]_ ;
  assign \new_[26773]_  = ~A298 & A266;
  assign \new_[26774]_  = A265 & \new_[26773]_ ;
  assign \new_[26778]_  = A302 & A300;
  assign \new_[26779]_  = A299 & \new_[26778]_ ;
  assign \new_[26780]_  = \new_[26779]_  & \new_[26774]_ ;
  assign \new_[26784]_  = A199 & ~A166;
  assign \new_[26785]_  = ~A167 & \new_[26784]_ ;
  assign \new_[26789]_  = A203 & A201;
  assign \new_[26790]_  = ~A200 & \new_[26789]_ ;
  assign \new_[26791]_  = \new_[26790]_  & \new_[26785]_ ;
  assign \new_[26795]_  = A298 & ~A266;
  assign \new_[26796]_  = ~A265 & \new_[26795]_ ;
  assign \new_[26800]_  = A301 & A300;
  assign \new_[26801]_  = ~A299 & \new_[26800]_ ;
  assign \new_[26802]_  = \new_[26801]_  & \new_[26796]_ ;
  assign \new_[26806]_  = A199 & ~A166;
  assign \new_[26807]_  = ~A167 & \new_[26806]_ ;
  assign \new_[26811]_  = A203 & A201;
  assign \new_[26812]_  = ~A200 & \new_[26811]_ ;
  assign \new_[26813]_  = \new_[26812]_  & \new_[26807]_ ;
  assign \new_[26817]_  = A298 & ~A266;
  assign \new_[26818]_  = ~A265 & \new_[26817]_ ;
  assign \new_[26822]_  = A302 & A300;
  assign \new_[26823]_  = ~A299 & \new_[26822]_ ;
  assign \new_[26824]_  = \new_[26823]_  & \new_[26818]_ ;
  assign \new_[26828]_  = A199 & ~A166;
  assign \new_[26829]_  = ~A167 & \new_[26828]_ ;
  assign \new_[26833]_  = A203 & A201;
  assign \new_[26834]_  = ~A200 & \new_[26833]_ ;
  assign \new_[26835]_  = \new_[26834]_  & \new_[26829]_ ;
  assign \new_[26839]_  = ~A298 & ~A266;
  assign \new_[26840]_  = ~A265 & \new_[26839]_ ;
  assign \new_[26844]_  = A301 & A300;
  assign \new_[26845]_  = A299 & \new_[26844]_ ;
  assign \new_[26846]_  = \new_[26845]_  & \new_[26840]_ ;
  assign \new_[26850]_  = A199 & ~A166;
  assign \new_[26851]_  = ~A167 & \new_[26850]_ ;
  assign \new_[26855]_  = A203 & A201;
  assign \new_[26856]_  = ~A200 & \new_[26855]_ ;
  assign \new_[26857]_  = \new_[26856]_  & \new_[26851]_ ;
  assign \new_[26861]_  = ~A298 & ~A266;
  assign \new_[26862]_  = ~A265 & \new_[26861]_ ;
  assign \new_[26866]_  = A302 & A300;
  assign \new_[26867]_  = A299 & \new_[26866]_ ;
  assign \new_[26868]_  = \new_[26867]_  & \new_[26862]_ ;
  assign \new_[26872]_  = ~A199 & ~A166;
  assign \new_[26873]_  = ~A167 & \new_[26872]_ ;
  assign \new_[26877]_  = A266 & ~A265;
  assign \new_[26878]_  = ~A200 & \new_[26877]_ ;
  assign \new_[26879]_  = \new_[26878]_  & \new_[26873]_ ;
  assign \new_[26883]_  = ~A269 & ~A268;
  assign \new_[26884]_  = ~A267 & \new_[26883]_ ;
  assign \new_[26888]_  = ~A302 & ~A301;
  assign \new_[26889]_  = A300 & \new_[26888]_ ;
  assign \new_[26890]_  = \new_[26889]_  & \new_[26884]_ ;
  assign \new_[26894]_  = ~A199 & ~A166;
  assign \new_[26895]_  = ~A167 & \new_[26894]_ ;
  assign \new_[26899]_  = ~A266 & A265;
  assign \new_[26900]_  = ~A200 & \new_[26899]_ ;
  assign \new_[26901]_  = \new_[26900]_  & \new_[26895]_ ;
  assign \new_[26905]_  = ~A269 & ~A268;
  assign \new_[26906]_  = ~A267 & \new_[26905]_ ;
  assign \new_[26910]_  = ~A302 & ~A301;
  assign \new_[26911]_  = A300 & \new_[26910]_ ;
  assign \new_[26912]_  = \new_[26911]_  & \new_[26906]_ ;
  assign \new_[26916]_  = A167 & A168;
  assign \new_[26917]_  = ~A170 & \new_[26916]_ ;
  assign \new_[26921]_  = A202 & ~A201;
  assign \new_[26922]_  = ~A166 & \new_[26921]_ ;
  assign \new_[26923]_  = \new_[26922]_  & \new_[26917]_ ;
  assign \new_[26927]_  = A298 & A268;
  assign \new_[26928]_  = ~A267 & \new_[26927]_ ;
  assign \new_[26932]_  = A301 & A300;
  assign \new_[26933]_  = ~A299 & \new_[26932]_ ;
  assign \new_[26934]_  = \new_[26933]_  & \new_[26928]_ ;
  assign \new_[26938]_  = A167 & A168;
  assign \new_[26939]_  = ~A170 & \new_[26938]_ ;
  assign \new_[26943]_  = A202 & ~A201;
  assign \new_[26944]_  = ~A166 & \new_[26943]_ ;
  assign \new_[26945]_  = \new_[26944]_  & \new_[26939]_ ;
  assign \new_[26949]_  = A298 & A268;
  assign \new_[26950]_  = ~A267 & \new_[26949]_ ;
  assign \new_[26954]_  = A302 & A300;
  assign \new_[26955]_  = ~A299 & \new_[26954]_ ;
  assign \new_[26956]_  = \new_[26955]_  & \new_[26950]_ ;
  assign \new_[26960]_  = A167 & A168;
  assign \new_[26961]_  = ~A170 & \new_[26960]_ ;
  assign \new_[26965]_  = A202 & ~A201;
  assign \new_[26966]_  = ~A166 & \new_[26965]_ ;
  assign \new_[26967]_  = \new_[26966]_  & \new_[26961]_ ;
  assign \new_[26971]_  = ~A298 & A268;
  assign \new_[26972]_  = ~A267 & \new_[26971]_ ;
  assign \new_[26976]_  = A301 & A300;
  assign \new_[26977]_  = A299 & \new_[26976]_ ;
  assign \new_[26978]_  = \new_[26977]_  & \new_[26972]_ ;
  assign \new_[26982]_  = A167 & A168;
  assign \new_[26983]_  = ~A170 & \new_[26982]_ ;
  assign \new_[26987]_  = A202 & ~A201;
  assign \new_[26988]_  = ~A166 & \new_[26987]_ ;
  assign \new_[26989]_  = \new_[26988]_  & \new_[26983]_ ;
  assign \new_[26993]_  = ~A298 & A268;
  assign \new_[26994]_  = ~A267 & \new_[26993]_ ;
  assign \new_[26998]_  = A302 & A300;
  assign \new_[26999]_  = A299 & \new_[26998]_ ;
  assign \new_[27000]_  = \new_[26999]_  & \new_[26994]_ ;
  assign \new_[27004]_  = A167 & A168;
  assign \new_[27005]_  = ~A170 & \new_[27004]_ ;
  assign \new_[27009]_  = A202 & ~A201;
  assign \new_[27010]_  = ~A166 & \new_[27009]_ ;
  assign \new_[27011]_  = \new_[27010]_  & \new_[27005]_ ;
  assign \new_[27015]_  = A298 & A269;
  assign \new_[27016]_  = ~A267 & \new_[27015]_ ;
  assign \new_[27020]_  = A301 & A300;
  assign \new_[27021]_  = ~A299 & \new_[27020]_ ;
  assign \new_[27022]_  = \new_[27021]_  & \new_[27016]_ ;
  assign \new_[27026]_  = A167 & A168;
  assign \new_[27027]_  = ~A170 & \new_[27026]_ ;
  assign \new_[27031]_  = A202 & ~A201;
  assign \new_[27032]_  = ~A166 & \new_[27031]_ ;
  assign \new_[27033]_  = \new_[27032]_  & \new_[27027]_ ;
  assign \new_[27037]_  = A298 & A269;
  assign \new_[27038]_  = ~A267 & \new_[27037]_ ;
  assign \new_[27042]_  = A302 & A300;
  assign \new_[27043]_  = ~A299 & \new_[27042]_ ;
  assign \new_[27044]_  = \new_[27043]_  & \new_[27038]_ ;
  assign \new_[27048]_  = A167 & A168;
  assign \new_[27049]_  = ~A170 & \new_[27048]_ ;
  assign \new_[27053]_  = A202 & ~A201;
  assign \new_[27054]_  = ~A166 & \new_[27053]_ ;
  assign \new_[27055]_  = \new_[27054]_  & \new_[27049]_ ;
  assign \new_[27059]_  = ~A298 & A269;
  assign \new_[27060]_  = ~A267 & \new_[27059]_ ;
  assign \new_[27064]_  = A301 & A300;
  assign \new_[27065]_  = A299 & \new_[27064]_ ;
  assign \new_[27066]_  = \new_[27065]_  & \new_[27060]_ ;
  assign \new_[27070]_  = A167 & A168;
  assign \new_[27071]_  = ~A170 & \new_[27070]_ ;
  assign \new_[27075]_  = A202 & ~A201;
  assign \new_[27076]_  = ~A166 & \new_[27075]_ ;
  assign \new_[27077]_  = \new_[27076]_  & \new_[27071]_ ;
  assign \new_[27081]_  = ~A298 & A269;
  assign \new_[27082]_  = ~A267 & \new_[27081]_ ;
  assign \new_[27086]_  = A302 & A300;
  assign \new_[27087]_  = A299 & \new_[27086]_ ;
  assign \new_[27088]_  = \new_[27087]_  & \new_[27082]_ ;
  assign \new_[27092]_  = A167 & A168;
  assign \new_[27093]_  = ~A170 & \new_[27092]_ ;
  assign \new_[27097]_  = A202 & ~A201;
  assign \new_[27098]_  = ~A166 & \new_[27097]_ ;
  assign \new_[27099]_  = \new_[27098]_  & \new_[27093]_ ;
  assign \new_[27103]_  = A298 & A266;
  assign \new_[27104]_  = A265 & \new_[27103]_ ;
  assign \new_[27108]_  = A301 & A300;
  assign \new_[27109]_  = ~A299 & \new_[27108]_ ;
  assign \new_[27110]_  = \new_[27109]_  & \new_[27104]_ ;
  assign \new_[27114]_  = A167 & A168;
  assign \new_[27115]_  = ~A170 & \new_[27114]_ ;
  assign \new_[27119]_  = A202 & ~A201;
  assign \new_[27120]_  = ~A166 & \new_[27119]_ ;
  assign \new_[27121]_  = \new_[27120]_  & \new_[27115]_ ;
  assign \new_[27125]_  = A298 & A266;
  assign \new_[27126]_  = A265 & \new_[27125]_ ;
  assign \new_[27130]_  = A302 & A300;
  assign \new_[27131]_  = ~A299 & \new_[27130]_ ;
  assign \new_[27132]_  = \new_[27131]_  & \new_[27126]_ ;
  assign \new_[27136]_  = A167 & A168;
  assign \new_[27137]_  = ~A170 & \new_[27136]_ ;
  assign \new_[27141]_  = A202 & ~A201;
  assign \new_[27142]_  = ~A166 & \new_[27141]_ ;
  assign \new_[27143]_  = \new_[27142]_  & \new_[27137]_ ;
  assign \new_[27147]_  = ~A298 & A266;
  assign \new_[27148]_  = A265 & \new_[27147]_ ;
  assign \new_[27152]_  = A301 & A300;
  assign \new_[27153]_  = A299 & \new_[27152]_ ;
  assign \new_[27154]_  = \new_[27153]_  & \new_[27148]_ ;
  assign \new_[27158]_  = A167 & A168;
  assign \new_[27159]_  = ~A170 & \new_[27158]_ ;
  assign \new_[27163]_  = A202 & ~A201;
  assign \new_[27164]_  = ~A166 & \new_[27163]_ ;
  assign \new_[27165]_  = \new_[27164]_  & \new_[27159]_ ;
  assign \new_[27169]_  = ~A298 & A266;
  assign \new_[27170]_  = A265 & \new_[27169]_ ;
  assign \new_[27174]_  = A302 & A300;
  assign \new_[27175]_  = A299 & \new_[27174]_ ;
  assign \new_[27176]_  = \new_[27175]_  & \new_[27170]_ ;
  assign \new_[27180]_  = A167 & A168;
  assign \new_[27181]_  = ~A170 & \new_[27180]_ ;
  assign \new_[27185]_  = A202 & ~A201;
  assign \new_[27186]_  = ~A166 & \new_[27185]_ ;
  assign \new_[27187]_  = \new_[27186]_  & \new_[27181]_ ;
  assign \new_[27191]_  = A298 & ~A266;
  assign \new_[27192]_  = ~A265 & \new_[27191]_ ;
  assign \new_[27196]_  = A301 & A300;
  assign \new_[27197]_  = ~A299 & \new_[27196]_ ;
  assign \new_[27198]_  = \new_[27197]_  & \new_[27192]_ ;
  assign \new_[27202]_  = A167 & A168;
  assign \new_[27203]_  = ~A170 & \new_[27202]_ ;
  assign \new_[27207]_  = A202 & ~A201;
  assign \new_[27208]_  = ~A166 & \new_[27207]_ ;
  assign \new_[27209]_  = \new_[27208]_  & \new_[27203]_ ;
  assign \new_[27213]_  = A298 & ~A266;
  assign \new_[27214]_  = ~A265 & \new_[27213]_ ;
  assign \new_[27218]_  = A302 & A300;
  assign \new_[27219]_  = ~A299 & \new_[27218]_ ;
  assign \new_[27220]_  = \new_[27219]_  & \new_[27214]_ ;
  assign \new_[27224]_  = A167 & A168;
  assign \new_[27225]_  = ~A170 & \new_[27224]_ ;
  assign \new_[27229]_  = A202 & ~A201;
  assign \new_[27230]_  = ~A166 & \new_[27229]_ ;
  assign \new_[27231]_  = \new_[27230]_  & \new_[27225]_ ;
  assign \new_[27235]_  = ~A298 & ~A266;
  assign \new_[27236]_  = ~A265 & \new_[27235]_ ;
  assign \new_[27240]_  = A301 & A300;
  assign \new_[27241]_  = A299 & \new_[27240]_ ;
  assign \new_[27242]_  = \new_[27241]_  & \new_[27236]_ ;
  assign \new_[27246]_  = A167 & A168;
  assign \new_[27247]_  = ~A170 & \new_[27246]_ ;
  assign \new_[27251]_  = A202 & ~A201;
  assign \new_[27252]_  = ~A166 & \new_[27251]_ ;
  assign \new_[27253]_  = \new_[27252]_  & \new_[27247]_ ;
  assign \new_[27257]_  = ~A298 & ~A266;
  assign \new_[27258]_  = ~A265 & \new_[27257]_ ;
  assign \new_[27262]_  = A302 & A300;
  assign \new_[27263]_  = A299 & \new_[27262]_ ;
  assign \new_[27264]_  = \new_[27263]_  & \new_[27258]_ ;
  assign \new_[27268]_  = A167 & A168;
  assign \new_[27269]_  = ~A170 & \new_[27268]_ ;
  assign \new_[27273]_  = A203 & ~A201;
  assign \new_[27274]_  = ~A166 & \new_[27273]_ ;
  assign \new_[27275]_  = \new_[27274]_  & \new_[27269]_ ;
  assign \new_[27279]_  = A298 & A268;
  assign \new_[27280]_  = ~A267 & \new_[27279]_ ;
  assign \new_[27284]_  = A301 & A300;
  assign \new_[27285]_  = ~A299 & \new_[27284]_ ;
  assign \new_[27286]_  = \new_[27285]_  & \new_[27280]_ ;
  assign \new_[27290]_  = A167 & A168;
  assign \new_[27291]_  = ~A170 & \new_[27290]_ ;
  assign \new_[27295]_  = A203 & ~A201;
  assign \new_[27296]_  = ~A166 & \new_[27295]_ ;
  assign \new_[27297]_  = \new_[27296]_  & \new_[27291]_ ;
  assign \new_[27301]_  = A298 & A268;
  assign \new_[27302]_  = ~A267 & \new_[27301]_ ;
  assign \new_[27306]_  = A302 & A300;
  assign \new_[27307]_  = ~A299 & \new_[27306]_ ;
  assign \new_[27308]_  = \new_[27307]_  & \new_[27302]_ ;
  assign \new_[27312]_  = A167 & A168;
  assign \new_[27313]_  = ~A170 & \new_[27312]_ ;
  assign \new_[27317]_  = A203 & ~A201;
  assign \new_[27318]_  = ~A166 & \new_[27317]_ ;
  assign \new_[27319]_  = \new_[27318]_  & \new_[27313]_ ;
  assign \new_[27323]_  = ~A298 & A268;
  assign \new_[27324]_  = ~A267 & \new_[27323]_ ;
  assign \new_[27328]_  = A301 & A300;
  assign \new_[27329]_  = A299 & \new_[27328]_ ;
  assign \new_[27330]_  = \new_[27329]_  & \new_[27324]_ ;
  assign \new_[27334]_  = A167 & A168;
  assign \new_[27335]_  = ~A170 & \new_[27334]_ ;
  assign \new_[27339]_  = A203 & ~A201;
  assign \new_[27340]_  = ~A166 & \new_[27339]_ ;
  assign \new_[27341]_  = \new_[27340]_  & \new_[27335]_ ;
  assign \new_[27345]_  = ~A298 & A268;
  assign \new_[27346]_  = ~A267 & \new_[27345]_ ;
  assign \new_[27350]_  = A302 & A300;
  assign \new_[27351]_  = A299 & \new_[27350]_ ;
  assign \new_[27352]_  = \new_[27351]_  & \new_[27346]_ ;
  assign \new_[27356]_  = A167 & A168;
  assign \new_[27357]_  = ~A170 & \new_[27356]_ ;
  assign \new_[27361]_  = A203 & ~A201;
  assign \new_[27362]_  = ~A166 & \new_[27361]_ ;
  assign \new_[27363]_  = \new_[27362]_  & \new_[27357]_ ;
  assign \new_[27367]_  = A298 & A269;
  assign \new_[27368]_  = ~A267 & \new_[27367]_ ;
  assign \new_[27372]_  = A301 & A300;
  assign \new_[27373]_  = ~A299 & \new_[27372]_ ;
  assign \new_[27374]_  = \new_[27373]_  & \new_[27368]_ ;
  assign \new_[27378]_  = A167 & A168;
  assign \new_[27379]_  = ~A170 & \new_[27378]_ ;
  assign \new_[27383]_  = A203 & ~A201;
  assign \new_[27384]_  = ~A166 & \new_[27383]_ ;
  assign \new_[27385]_  = \new_[27384]_  & \new_[27379]_ ;
  assign \new_[27389]_  = A298 & A269;
  assign \new_[27390]_  = ~A267 & \new_[27389]_ ;
  assign \new_[27394]_  = A302 & A300;
  assign \new_[27395]_  = ~A299 & \new_[27394]_ ;
  assign \new_[27396]_  = \new_[27395]_  & \new_[27390]_ ;
  assign \new_[27400]_  = A167 & A168;
  assign \new_[27401]_  = ~A170 & \new_[27400]_ ;
  assign \new_[27405]_  = A203 & ~A201;
  assign \new_[27406]_  = ~A166 & \new_[27405]_ ;
  assign \new_[27407]_  = \new_[27406]_  & \new_[27401]_ ;
  assign \new_[27411]_  = ~A298 & A269;
  assign \new_[27412]_  = ~A267 & \new_[27411]_ ;
  assign \new_[27416]_  = A301 & A300;
  assign \new_[27417]_  = A299 & \new_[27416]_ ;
  assign \new_[27418]_  = \new_[27417]_  & \new_[27412]_ ;
  assign \new_[27422]_  = A167 & A168;
  assign \new_[27423]_  = ~A170 & \new_[27422]_ ;
  assign \new_[27427]_  = A203 & ~A201;
  assign \new_[27428]_  = ~A166 & \new_[27427]_ ;
  assign \new_[27429]_  = \new_[27428]_  & \new_[27423]_ ;
  assign \new_[27433]_  = ~A298 & A269;
  assign \new_[27434]_  = ~A267 & \new_[27433]_ ;
  assign \new_[27438]_  = A302 & A300;
  assign \new_[27439]_  = A299 & \new_[27438]_ ;
  assign \new_[27440]_  = \new_[27439]_  & \new_[27434]_ ;
  assign \new_[27444]_  = A167 & A168;
  assign \new_[27445]_  = ~A170 & \new_[27444]_ ;
  assign \new_[27449]_  = A203 & ~A201;
  assign \new_[27450]_  = ~A166 & \new_[27449]_ ;
  assign \new_[27451]_  = \new_[27450]_  & \new_[27445]_ ;
  assign \new_[27455]_  = A298 & A266;
  assign \new_[27456]_  = A265 & \new_[27455]_ ;
  assign \new_[27460]_  = A301 & A300;
  assign \new_[27461]_  = ~A299 & \new_[27460]_ ;
  assign \new_[27462]_  = \new_[27461]_  & \new_[27456]_ ;
  assign \new_[27466]_  = A167 & A168;
  assign \new_[27467]_  = ~A170 & \new_[27466]_ ;
  assign \new_[27471]_  = A203 & ~A201;
  assign \new_[27472]_  = ~A166 & \new_[27471]_ ;
  assign \new_[27473]_  = \new_[27472]_  & \new_[27467]_ ;
  assign \new_[27477]_  = A298 & A266;
  assign \new_[27478]_  = A265 & \new_[27477]_ ;
  assign \new_[27482]_  = A302 & A300;
  assign \new_[27483]_  = ~A299 & \new_[27482]_ ;
  assign \new_[27484]_  = \new_[27483]_  & \new_[27478]_ ;
  assign \new_[27488]_  = A167 & A168;
  assign \new_[27489]_  = ~A170 & \new_[27488]_ ;
  assign \new_[27493]_  = A203 & ~A201;
  assign \new_[27494]_  = ~A166 & \new_[27493]_ ;
  assign \new_[27495]_  = \new_[27494]_  & \new_[27489]_ ;
  assign \new_[27499]_  = ~A298 & A266;
  assign \new_[27500]_  = A265 & \new_[27499]_ ;
  assign \new_[27504]_  = A301 & A300;
  assign \new_[27505]_  = A299 & \new_[27504]_ ;
  assign \new_[27506]_  = \new_[27505]_  & \new_[27500]_ ;
  assign \new_[27510]_  = A167 & A168;
  assign \new_[27511]_  = ~A170 & \new_[27510]_ ;
  assign \new_[27515]_  = A203 & ~A201;
  assign \new_[27516]_  = ~A166 & \new_[27515]_ ;
  assign \new_[27517]_  = \new_[27516]_  & \new_[27511]_ ;
  assign \new_[27521]_  = ~A298 & A266;
  assign \new_[27522]_  = A265 & \new_[27521]_ ;
  assign \new_[27526]_  = A302 & A300;
  assign \new_[27527]_  = A299 & \new_[27526]_ ;
  assign \new_[27528]_  = \new_[27527]_  & \new_[27522]_ ;
  assign \new_[27532]_  = A167 & A168;
  assign \new_[27533]_  = ~A170 & \new_[27532]_ ;
  assign \new_[27537]_  = A203 & ~A201;
  assign \new_[27538]_  = ~A166 & \new_[27537]_ ;
  assign \new_[27539]_  = \new_[27538]_  & \new_[27533]_ ;
  assign \new_[27543]_  = A298 & ~A266;
  assign \new_[27544]_  = ~A265 & \new_[27543]_ ;
  assign \new_[27548]_  = A301 & A300;
  assign \new_[27549]_  = ~A299 & \new_[27548]_ ;
  assign \new_[27550]_  = \new_[27549]_  & \new_[27544]_ ;
  assign \new_[27554]_  = A167 & A168;
  assign \new_[27555]_  = ~A170 & \new_[27554]_ ;
  assign \new_[27559]_  = A203 & ~A201;
  assign \new_[27560]_  = ~A166 & \new_[27559]_ ;
  assign \new_[27561]_  = \new_[27560]_  & \new_[27555]_ ;
  assign \new_[27565]_  = A298 & ~A266;
  assign \new_[27566]_  = ~A265 & \new_[27565]_ ;
  assign \new_[27570]_  = A302 & A300;
  assign \new_[27571]_  = ~A299 & \new_[27570]_ ;
  assign \new_[27572]_  = \new_[27571]_  & \new_[27566]_ ;
  assign \new_[27576]_  = A167 & A168;
  assign \new_[27577]_  = ~A170 & \new_[27576]_ ;
  assign \new_[27581]_  = A203 & ~A201;
  assign \new_[27582]_  = ~A166 & \new_[27581]_ ;
  assign \new_[27583]_  = \new_[27582]_  & \new_[27577]_ ;
  assign \new_[27587]_  = ~A298 & ~A266;
  assign \new_[27588]_  = ~A265 & \new_[27587]_ ;
  assign \new_[27592]_  = A301 & A300;
  assign \new_[27593]_  = A299 & \new_[27592]_ ;
  assign \new_[27594]_  = \new_[27593]_  & \new_[27588]_ ;
  assign \new_[27598]_  = A167 & A168;
  assign \new_[27599]_  = ~A170 & \new_[27598]_ ;
  assign \new_[27603]_  = A203 & ~A201;
  assign \new_[27604]_  = ~A166 & \new_[27603]_ ;
  assign \new_[27605]_  = \new_[27604]_  & \new_[27599]_ ;
  assign \new_[27609]_  = ~A298 & ~A266;
  assign \new_[27610]_  = ~A265 & \new_[27609]_ ;
  assign \new_[27614]_  = A302 & A300;
  assign \new_[27615]_  = A299 & \new_[27614]_ ;
  assign \new_[27616]_  = \new_[27615]_  & \new_[27610]_ ;
  assign \new_[27620]_  = A167 & A168;
  assign \new_[27621]_  = ~A170 & \new_[27620]_ ;
  assign \new_[27625]_  = A200 & A199;
  assign \new_[27626]_  = ~A166 & \new_[27625]_ ;
  assign \new_[27627]_  = \new_[27626]_  & \new_[27621]_ ;
  assign \new_[27631]_  = A298 & A268;
  assign \new_[27632]_  = ~A267 & \new_[27631]_ ;
  assign \new_[27636]_  = A301 & A300;
  assign \new_[27637]_  = ~A299 & \new_[27636]_ ;
  assign \new_[27638]_  = \new_[27637]_  & \new_[27632]_ ;
  assign \new_[27642]_  = A167 & A168;
  assign \new_[27643]_  = ~A170 & \new_[27642]_ ;
  assign \new_[27647]_  = A200 & A199;
  assign \new_[27648]_  = ~A166 & \new_[27647]_ ;
  assign \new_[27649]_  = \new_[27648]_  & \new_[27643]_ ;
  assign \new_[27653]_  = A298 & A268;
  assign \new_[27654]_  = ~A267 & \new_[27653]_ ;
  assign \new_[27658]_  = A302 & A300;
  assign \new_[27659]_  = ~A299 & \new_[27658]_ ;
  assign \new_[27660]_  = \new_[27659]_  & \new_[27654]_ ;
  assign \new_[27664]_  = A167 & A168;
  assign \new_[27665]_  = ~A170 & \new_[27664]_ ;
  assign \new_[27669]_  = A200 & A199;
  assign \new_[27670]_  = ~A166 & \new_[27669]_ ;
  assign \new_[27671]_  = \new_[27670]_  & \new_[27665]_ ;
  assign \new_[27675]_  = ~A298 & A268;
  assign \new_[27676]_  = ~A267 & \new_[27675]_ ;
  assign \new_[27680]_  = A301 & A300;
  assign \new_[27681]_  = A299 & \new_[27680]_ ;
  assign \new_[27682]_  = \new_[27681]_  & \new_[27676]_ ;
  assign \new_[27686]_  = A167 & A168;
  assign \new_[27687]_  = ~A170 & \new_[27686]_ ;
  assign \new_[27691]_  = A200 & A199;
  assign \new_[27692]_  = ~A166 & \new_[27691]_ ;
  assign \new_[27693]_  = \new_[27692]_  & \new_[27687]_ ;
  assign \new_[27697]_  = ~A298 & A268;
  assign \new_[27698]_  = ~A267 & \new_[27697]_ ;
  assign \new_[27702]_  = A302 & A300;
  assign \new_[27703]_  = A299 & \new_[27702]_ ;
  assign \new_[27704]_  = \new_[27703]_  & \new_[27698]_ ;
  assign \new_[27708]_  = A167 & A168;
  assign \new_[27709]_  = ~A170 & \new_[27708]_ ;
  assign \new_[27713]_  = A200 & A199;
  assign \new_[27714]_  = ~A166 & \new_[27713]_ ;
  assign \new_[27715]_  = \new_[27714]_  & \new_[27709]_ ;
  assign \new_[27719]_  = A298 & A269;
  assign \new_[27720]_  = ~A267 & \new_[27719]_ ;
  assign \new_[27724]_  = A301 & A300;
  assign \new_[27725]_  = ~A299 & \new_[27724]_ ;
  assign \new_[27726]_  = \new_[27725]_  & \new_[27720]_ ;
  assign \new_[27730]_  = A167 & A168;
  assign \new_[27731]_  = ~A170 & \new_[27730]_ ;
  assign \new_[27735]_  = A200 & A199;
  assign \new_[27736]_  = ~A166 & \new_[27735]_ ;
  assign \new_[27737]_  = \new_[27736]_  & \new_[27731]_ ;
  assign \new_[27741]_  = A298 & A269;
  assign \new_[27742]_  = ~A267 & \new_[27741]_ ;
  assign \new_[27746]_  = A302 & A300;
  assign \new_[27747]_  = ~A299 & \new_[27746]_ ;
  assign \new_[27748]_  = \new_[27747]_  & \new_[27742]_ ;
  assign \new_[27752]_  = A167 & A168;
  assign \new_[27753]_  = ~A170 & \new_[27752]_ ;
  assign \new_[27757]_  = A200 & A199;
  assign \new_[27758]_  = ~A166 & \new_[27757]_ ;
  assign \new_[27759]_  = \new_[27758]_  & \new_[27753]_ ;
  assign \new_[27763]_  = ~A298 & A269;
  assign \new_[27764]_  = ~A267 & \new_[27763]_ ;
  assign \new_[27768]_  = A301 & A300;
  assign \new_[27769]_  = A299 & \new_[27768]_ ;
  assign \new_[27770]_  = \new_[27769]_  & \new_[27764]_ ;
  assign \new_[27774]_  = A167 & A168;
  assign \new_[27775]_  = ~A170 & \new_[27774]_ ;
  assign \new_[27779]_  = A200 & A199;
  assign \new_[27780]_  = ~A166 & \new_[27779]_ ;
  assign \new_[27781]_  = \new_[27780]_  & \new_[27775]_ ;
  assign \new_[27785]_  = ~A298 & A269;
  assign \new_[27786]_  = ~A267 & \new_[27785]_ ;
  assign \new_[27790]_  = A302 & A300;
  assign \new_[27791]_  = A299 & \new_[27790]_ ;
  assign \new_[27792]_  = \new_[27791]_  & \new_[27786]_ ;
  assign \new_[27796]_  = A167 & A168;
  assign \new_[27797]_  = ~A170 & \new_[27796]_ ;
  assign \new_[27801]_  = A200 & A199;
  assign \new_[27802]_  = ~A166 & \new_[27801]_ ;
  assign \new_[27803]_  = \new_[27802]_  & \new_[27797]_ ;
  assign \new_[27807]_  = A298 & A266;
  assign \new_[27808]_  = A265 & \new_[27807]_ ;
  assign \new_[27812]_  = A301 & A300;
  assign \new_[27813]_  = ~A299 & \new_[27812]_ ;
  assign \new_[27814]_  = \new_[27813]_  & \new_[27808]_ ;
  assign \new_[27818]_  = A167 & A168;
  assign \new_[27819]_  = ~A170 & \new_[27818]_ ;
  assign \new_[27823]_  = A200 & A199;
  assign \new_[27824]_  = ~A166 & \new_[27823]_ ;
  assign \new_[27825]_  = \new_[27824]_  & \new_[27819]_ ;
  assign \new_[27829]_  = A298 & A266;
  assign \new_[27830]_  = A265 & \new_[27829]_ ;
  assign \new_[27834]_  = A302 & A300;
  assign \new_[27835]_  = ~A299 & \new_[27834]_ ;
  assign \new_[27836]_  = \new_[27835]_  & \new_[27830]_ ;
  assign \new_[27840]_  = A167 & A168;
  assign \new_[27841]_  = ~A170 & \new_[27840]_ ;
  assign \new_[27845]_  = A200 & A199;
  assign \new_[27846]_  = ~A166 & \new_[27845]_ ;
  assign \new_[27847]_  = \new_[27846]_  & \new_[27841]_ ;
  assign \new_[27851]_  = ~A298 & A266;
  assign \new_[27852]_  = A265 & \new_[27851]_ ;
  assign \new_[27856]_  = A301 & A300;
  assign \new_[27857]_  = A299 & \new_[27856]_ ;
  assign \new_[27858]_  = \new_[27857]_  & \new_[27852]_ ;
  assign \new_[27862]_  = A167 & A168;
  assign \new_[27863]_  = ~A170 & \new_[27862]_ ;
  assign \new_[27867]_  = A200 & A199;
  assign \new_[27868]_  = ~A166 & \new_[27867]_ ;
  assign \new_[27869]_  = \new_[27868]_  & \new_[27863]_ ;
  assign \new_[27873]_  = ~A298 & A266;
  assign \new_[27874]_  = A265 & \new_[27873]_ ;
  assign \new_[27878]_  = A302 & A300;
  assign \new_[27879]_  = A299 & \new_[27878]_ ;
  assign \new_[27880]_  = \new_[27879]_  & \new_[27874]_ ;
  assign \new_[27884]_  = A167 & A168;
  assign \new_[27885]_  = ~A170 & \new_[27884]_ ;
  assign \new_[27889]_  = A200 & A199;
  assign \new_[27890]_  = ~A166 & \new_[27889]_ ;
  assign \new_[27891]_  = \new_[27890]_  & \new_[27885]_ ;
  assign \new_[27895]_  = A298 & ~A266;
  assign \new_[27896]_  = ~A265 & \new_[27895]_ ;
  assign \new_[27900]_  = A301 & A300;
  assign \new_[27901]_  = ~A299 & \new_[27900]_ ;
  assign \new_[27902]_  = \new_[27901]_  & \new_[27896]_ ;
  assign \new_[27906]_  = A167 & A168;
  assign \new_[27907]_  = ~A170 & \new_[27906]_ ;
  assign \new_[27911]_  = A200 & A199;
  assign \new_[27912]_  = ~A166 & \new_[27911]_ ;
  assign \new_[27913]_  = \new_[27912]_  & \new_[27907]_ ;
  assign \new_[27917]_  = A298 & ~A266;
  assign \new_[27918]_  = ~A265 & \new_[27917]_ ;
  assign \new_[27922]_  = A302 & A300;
  assign \new_[27923]_  = ~A299 & \new_[27922]_ ;
  assign \new_[27924]_  = \new_[27923]_  & \new_[27918]_ ;
  assign \new_[27928]_  = A167 & A168;
  assign \new_[27929]_  = ~A170 & \new_[27928]_ ;
  assign \new_[27933]_  = A200 & A199;
  assign \new_[27934]_  = ~A166 & \new_[27933]_ ;
  assign \new_[27935]_  = \new_[27934]_  & \new_[27929]_ ;
  assign \new_[27939]_  = ~A298 & ~A266;
  assign \new_[27940]_  = ~A265 & \new_[27939]_ ;
  assign \new_[27944]_  = A301 & A300;
  assign \new_[27945]_  = A299 & \new_[27944]_ ;
  assign \new_[27946]_  = \new_[27945]_  & \new_[27940]_ ;
  assign \new_[27950]_  = A167 & A168;
  assign \new_[27951]_  = ~A170 & \new_[27950]_ ;
  assign \new_[27955]_  = A200 & A199;
  assign \new_[27956]_  = ~A166 & \new_[27955]_ ;
  assign \new_[27957]_  = \new_[27956]_  & \new_[27951]_ ;
  assign \new_[27961]_  = ~A298 & ~A266;
  assign \new_[27962]_  = ~A265 & \new_[27961]_ ;
  assign \new_[27966]_  = A302 & A300;
  assign \new_[27967]_  = A299 & \new_[27966]_ ;
  assign \new_[27968]_  = \new_[27967]_  & \new_[27962]_ ;
  assign \new_[27972]_  = A167 & A168;
  assign \new_[27973]_  = ~A170 & \new_[27972]_ ;
  assign \new_[27977]_  = ~A200 & ~A199;
  assign \new_[27978]_  = ~A166 & \new_[27977]_ ;
  assign \new_[27979]_  = \new_[27978]_  & \new_[27973]_ ;
  assign \new_[27983]_  = A298 & A268;
  assign \new_[27984]_  = ~A267 & \new_[27983]_ ;
  assign \new_[27988]_  = A301 & A300;
  assign \new_[27989]_  = ~A299 & \new_[27988]_ ;
  assign \new_[27990]_  = \new_[27989]_  & \new_[27984]_ ;
  assign \new_[27994]_  = A167 & A168;
  assign \new_[27995]_  = ~A170 & \new_[27994]_ ;
  assign \new_[27999]_  = ~A200 & ~A199;
  assign \new_[28000]_  = ~A166 & \new_[27999]_ ;
  assign \new_[28001]_  = \new_[28000]_  & \new_[27995]_ ;
  assign \new_[28005]_  = A298 & A268;
  assign \new_[28006]_  = ~A267 & \new_[28005]_ ;
  assign \new_[28010]_  = A302 & A300;
  assign \new_[28011]_  = ~A299 & \new_[28010]_ ;
  assign \new_[28012]_  = \new_[28011]_  & \new_[28006]_ ;
  assign \new_[28016]_  = A167 & A168;
  assign \new_[28017]_  = ~A170 & \new_[28016]_ ;
  assign \new_[28021]_  = ~A200 & ~A199;
  assign \new_[28022]_  = ~A166 & \new_[28021]_ ;
  assign \new_[28023]_  = \new_[28022]_  & \new_[28017]_ ;
  assign \new_[28027]_  = ~A298 & A268;
  assign \new_[28028]_  = ~A267 & \new_[28027]_ ;
  assign \new_[28032]_  = A301 & A300;
  assign \new_[28033]_  = A299 & \new_[28032]_ ;
  assign \new_[28034]_  = \new_[28033]_  & \new_[28028]_ ;
  assign \new_[28038]_  = A167 & A168;
  assign \new_[28039]_  = ~A170 & \new_[28038]_ ;
  assign \new_[28043]_  = ~A200 & ~A199;
  assign \new_[28044]_  = ~A166 & \new_[28043]_ ;
  assign \new_[28045]_  = \new_[28044]_  & \new_[28039]_ ;
  assign \new_[28049]_  = ~A298 & A268;
  assign \new_[28050]_  = ~A267 & \new_[28049]_ ;
  assign \new_[28054]_  = A302 & A300;
  assign \new_[28055]_  = A299 & \new_[28054]_ ;
  assign \new_[28056]_  = \new_[28055]_  & \new_[28050]_ ;
  assign \new_[28060]_  = A167 & A168;
  assign \new_[28061]_  = ~A170 & \new_[28060]_ ;
  assign \new_[28065]_  = ~A200 & ~A199;
  assign \new_[28066]_  = ~A166 & \new_[28065]_ ;
  assign \new_[28067]_  = \new_[28066]_  & \new_[28061]_ ;
  assign \new_[28071]_  = A298 & A269;
  assign \new_[28072]_  = ~A267 & \new_[28071]_ ;
  assign \new_[28076]_  = A301 & A300;
  assign \new_[28077]_  = ~A299 & \new_[28076]_ ;
  assign \new_[28078]_  = \new_[28077]_  & \new_[28072]_ ;
  assign \new_[28082]_  = A167 & A168;
  assign \new_[28083]_  = ~A170 & \new_[28082]_ ;
  assign \new_[28087]_  = ~A200 & ~A199;
  assign \new_[28088]_  = ~A166 & \new_[28087]_ ;
  assign \new_[28089]_  = \new_[28088]_  & \new_[28083]_ ;
  assign \new_[28093]_  = A298 & A269;
  assign \new_[28094]_  = ~A267 & \new_[28093]_ ;
  assign \new_[28098]_  = A302 & A300;
  assign \new_[28099]_  = ~A299 & \new_[28098]_ ;
  assign \new_[28100]_  = \new_[28099]_  & \new_[28094]_ ;
  assign \new_[28104]_  = A167 & A168;
  assign \new_[28105]_  = ~A170 & \new_[28104]_ ;
  assign \new_[28109]_  = ~A200 & ~A199;
  assign \new_[28110]_  = ~A166 & \new_[28109]_ ;
  assign \new_[28111]_  = \new_[28110]_  & \new_[28105]_ ;
  assign \new_[28115]_  = ~A298 & A269;
  assign \new_[28116]_  = ~A267 & \new_[28115]_ ;
  assign \new_[28120]_  = A301 & A300;
  assign \new_[28121]_  = A299 & \new_[28120]_ ;
  assign \new_[28122]_  = \new_[28121]_  & \new_[28116]_ ;
  assign \new_[28126]_  = A167 & A168;
  assign \new_[28127]_  = ~A170 & \new_[28126]_ ;
  assign \new_[28131]_  = ~A200 & ~A199;
  assign \new_[28132]_  = ~A166 & \new_[28131]_ ;
  assign \new_[28133]_  = \new_[28132]_  & \new_[28127]_ ;
  assign \new_[28137]_  = ~A298 & A269;
  assign \new_[28138]_  = ~A267 & \new_[28137]_ ;
  assign \new_[28142]_  = A302 & A300;
  assign \new_[28143]_  = A299 & \new_[28142]_ ;
  assign \new_[28144]_  = \new_[28143]_  & \new_[28138]_ ;
  assign \new_[28148]_  = A167 & A168;
  assign \new_[28149]_  = ~A170 & \new_[28148]_ ;
  assign \new_[28153]_  = ~A200 & ~A199;
  assign \new_[28154]_  = ~A166 & \new_[28153]_ ;
  assign \new_[28155]_  = \new_[28154]_  & \new_[28149]_ ;
  assign \new_[28159]_  = A298 & A266;
  assign \new_[28160]_  = A265 & \new_[28159]_ ;
  assign \new_[28164]_  = A301 & A300;
  assign \new_[28165]_  = ~A299 & \new_[28164]_ ;
  assign \new_[28166]_  = \new_[28165]_  & \new_[28160]_ ;
  assign \new_[28170]_  = A167 & A168;
  assign \new_[28171]_  = ~A170 & \new_[28170]_ ;
  assign \new_[28175]_  = ~A200 & ~A199;
  assign \new_[28176]_  = ~A166 & \new_[28175]_ ;
  assign \new_[28177]_  = \new_[28176]_  & \new_[28171]_ ;
  assign \new_[28181]_  = A298 & A266;
  assign \new_[28182]_  = A265 & \new_[28181]_ ;
  assign \new_[28186]_  = A302 & A300;
  assign \new_[28187]_  = ~A299 & \new_[28186]_ ;
  assign \new_[28188]_  = \new_[28187]_  & \new_[28182]_ ;
  assign \new_[28192]_  = A167 & A168;
  assign \new_[28193]_  = ~A170 & \new_[28192]_ ;
  assign \new_[28197]_  = ~A200 & ~A199;
  assign \new_[28198]_  = ~A166 & \new_[28197]_ ;
  assign \new_[28199]_  = \new_[28198]_  & \new_[28193]_ ;
  assign \new_[28203]_  = ~A298 & A266;
  assign \new_[28204]_  = A265 & \new_[28203]_ ;
  assign \new_[28208]_  = A301 & A300;
  assign \new_[28209]_  = A299 & \new_[28208]_ ;
  assign \new_[28210]_  = \new_[28209]_  & \new_[28204]_ ;
  assign \new_[28214]_  = A167 & A168;
  assign \new_[28215]_  = ~A170 & \new_[28214]_ ;
  assign \new_[28219]_  = ~A200 & ~A199;
  assign \new_[28220]_  = ~A166 & \new_[28219]_ ;
  assign \new_[28221]_  = \new_[28220]_  & \new_[28215]_ ;
  assign \new_[28225]_  = ~A298 & A266;
  assign \new_[28226]_  = A265 & \new_[28225]_ ;
  assign \new_[28230]_  = A302 & A300;
  assign \new_[28231]_  = A299 & \new_[28230]_ ;
  assign \new_[28232]_  = \new_[28231]_  & \new_[28226]_ ;
  assign \new_[28236]_  = A167 & A168;
  assign \new_[28237]_  = ~A170 & \new_[28236]_ ;
  assign \new_[28241]_  = ~A200 & ~A199;
  assign \new_[28242]_  = ~A166 & \new_[28241]_ ;
  assign \new_[28243]_  = \new_[28242]_  & \new_[28237]_ ;
  assign \new_[28247]_  = A298 & ~A266;
  assign \new_[28248]_  = ~A265 & \new_[28247]_ ;
  assign \new_[28252]_  = A301 & A300;
  assign \new_[28253]_  = ~A299 & \new_[28252]_ ;
  assign \new_[28254]_  = \new_[28253]_  & \new_[28248]_ ;
  assign \new_[28258]_  = A167 & A168;
  assign \new_[28259]_  = ~A170 & \new_[28258]_ ;
  assign \new_[28263]_  = ~A200 & ~A199;
  assign \new_[28264]_  = ~A166 & \new_[28263]_ ;
  assign \new_[28265]_  = \new_[28264]_  & \new_[28259]_ ;
  assign \new_[28269]_  = A298 & ~A266;
  assign \new_[28270]_  = ~A265 & \new_[28269]_ ;
  assign \new_[28274]_  = A302 & A300;
  assign \new_[28275]_  = ~A299 & \new_[28274]_ ;
  assign \new_[28276]_  = \new_[28275]_  & \new_[28270]_ ;
  assign \new_[28280]_  = A167 & A168;
  assign \new_[28281]_  = ~A170 & \new_[28280]_ ;
  assign \new_[28285]_  = ~A200 & ~A199;
  assign \new_[28286]_  = ~A166 & \new_[28285]_ ;
  assign \new_[28287]_  = \new_[28286]_  & \new_[28281]_ ;
  assign \new_[28291]_  = ~A298 & ~A266;
  assign \new_[28292]_  = ~A265 & \new_[28291]_ ;
  assign \new_[28296]_  = A301 & A300;
  assign \new_[28297]_  = A299 & \new_[28296]_ ;
  assign \new_[28298]_  = \new_[28297]_  & \new_[28292]_ ;
  assign \new_[28302]_  = A167 & A168;
  assign \new_[28303]_  = ~A170 & \new_[28302]_ ;
  assign \new_[28307]_  = ~A200 & ~A199;
  assign \new_[28308]_  = ~A166 & \new_[28307]_ ;
  assign \new_[28309]_  = \new_[28308]_  & \new_[28303]_ ;
  assign \new_[28313]_  = ~A298 & ~A266;
  assign \new_[28314]_  = ~A265 & \new_[28313]_ ;
  assign \new_[28318]_  = A302 & A300;
  assign \new_[28319]_  = A299 & \new_[28318]_ ;
  assign \new_[28320]_  = \new_[28319]_  & \new_[28314]_ ;
  assign \new_[28324]_  = ~A167 & A168;
  assign \new_[28325]_  = ~A170 & \new_[28324]_ ;
  assign \new_[28329]_  = A202 & ~A201;
  assign \new_[28330]_  = A166 & \new_[28329]_ ;
  assign \new_[28331]_  = \new_[28330]_  & \new_[28325]_ ;
  assign \new_[28335]_  = A298 & A268;
  assign \new_[28336]_  = ~A267 & \new_[28335]_ ;
  assign \new_[28340]_  = A301 & A300;
  assign \new_[28341]_  = ~A299 & \new_[28340]_ ;
  assign \new_[28342]_  = \new_[28341]_  & \new_[28336]_ ;
  assign \new_[28346]_  = ~A167 & A168;
  assign \new_[28347]_  = ~A170 & \new_[28346]_ ;
  assign \new_[28351]_  = A202 & ~A201;
  assign \new_[28352]_  = A166 & \new_[28351]_ ;
  assign \new_[28353]_  = \new_[28352]_  & \new_[28347]_ ;
  assign \new_[28357]_  = A298 & A268;
  assign \new_[28358]_  = ~A267 & \new_[28357]_ ;
  assign \new_[28362]_  = A302 & A300;
  assign \new_[28363]_  = ~A299 & \new_[28362]_ ;
  assign \new_[28364]_  = \new_[28363]_  & \new_[28358]_ ;
  assign \new_[28368]_  = ~A167 & A168;
  assign \new_[28369]_  = ~A170 & \new_[28368]_ ;
  assign \new_[28373]_  = A202 & ~A201;
  assign \new_[28374]_  = A166 & \new_[28373]_ ;
  assign \new_[28375]_  = \new_[28374]_  & \new_[28369]_ ;
  assign \new_[28379]_  = ~A298 & A268;
  assign \new_[28380]_  = ~A267 & \new_[28379]_ ;
  assign \new_[28384]_  = A301 & A300;
  assign \new_[28385]_  = A299 & \new_[28384]_ ;
  assign \new_[28386]_  = \new_[28385]_  & \new_[28380]_ ;
  assign \new_[28390]_  = ~A167 & A168;
  assign \new_[28391]_  = ~A170 & \new_[28390]_ ;
  assign \new_[28395]_  = A202 & ~A201;
  assign \new_[28396]_  = A166 & \new_[28395]_ ;
  assign \new_[28397]_  = \new_[28396]_  & \new_[28391]_ ;
  assign \new_[28401]_  = ~A298 & A268;
  assign \new_[28402]_  = ~A267 & \new_[28401]_ ;
  assign \new_[28406]_  = A302 & A300;
  assign \new_[28407]_  = A299 & \new_[28406]_ ;
  assign \new_[28408]_  = \new_[28407]_  & \new_[28402]_ ;
  assign \new_[28412]_  = ~A167 & A168;
  assign \new_[28413]_  = ~A170 & \new_[28412]_ ;
  assign \new_[28417]_  = A202 & ~A201;
  assign \new_[28418]_  = A166 & \new_[28417]_ ;
  assign \new_[28419]_  = \new_[28418]_  & \new_[28413]_ ;
  assign \new_[28423]_  = A298 & A269;
  assign \new_[28424]_  = ~A267 & \new_[28423]_ ;
  assign \new_[28428]_  = A301 & A300;
  assign \new_[28429]_  = ~A299 & \new_[28428]_ ;
  assign \new_[28430]_  = \new_[28429]_  & \new_[28424]_ ;
  assign \new_[28434]_  = ~A167 & A168;
  assign \new_[28435]_  = ~A170 & \new_[28434]_ ;
  assign \new_[28439]_  = A202 & ~A201;
  assign \new_[28440]_  = A166 & \new_[28439]_ ;
  assign \new_[28441]_  = \new_[28440]_  & \new_[28435]_ ;
  assign \new_[28445]_  = A298 & A269;
  assign \new_[28446]_  = ~A267 & \new_[28445]_ ;
  assign \new_[28450]_  = A302 & A300;
  assign \new_[28451]_  = ~A299 & \new_[28450]_ ;
  assign \new_[28452]_  = \new_[28451]_  & \new_[28446]_ ;
  assign \new_[28456]_  = ~A167 & A168;
  assign \new_[28457]_  = ~A170 & \new_[28456]_ ;
  assign \new_[28461]_  = A202 & ~A201;
  assign \new_[28462]_  = A166 & \new_[28461]_ ;
  assign \new_[28463]_  = \new_[28462]_  & \new_[28457]_ ;
  assign \new_[28467]_  = ~A298 & A269;
  assign \new_[28468]_  = ~A267 & \new_[28467]_ ;
  assign \new_[28472]_  = A301 & A300;
  assign \new_[28473]_  = A299 & \new_[28472]_ ;
  assign \new_[28474]_  = \new_[28473]_  & \new_[28468]_ ;
  assign \new_[28478]_  = ~A167 & A168;
  assign \new_[28479]_  = ~A170 & \new_[28478]_ ;
  assign \new_[28483]_  = A202 & ~A201;
  assign \new_[28484]_  = A166 & \new_[28483]_ ;
  assign \new_[28485]_  = \new_[28484]_  & \new_[28479]_ ;
  assign \new_[28489]_  = ~A298 & A269;
  assign \new_[28490]_  = ~A267 & \new_[28489]_ ;
  assign \new_[28494]_  = A302 & A300;
  assign \new_[28495]_  = A299 & \new_[28494]_ ;
  assign \new_[28496]_  = \new_[28495]_  & \new_[28490]_ ;
  assign \new_[28500]_  = ~A167 & A168;
  assign \new_[28501]_  = ~A170 & \new_[28500]_ ;
  assign \new_[28505]_  = A202 & ~A201;
  assign \new_[28506]_  = A166 & \new_[28505]_ ;
  assign \new_[28507]_  = \new_[28506]_  & \new_[28501]_ ;
  assign \new_[28511]_  = A298 & A266;
  assign \new_[28512]_  = A265 & \new_[28511]_ ;
  assign \new_[28516]_  = A301 & A300;
  assign \new_[28517]_  = ~A299 & \new_[28516]_ ;
  assign \new_[28518]_  = \new_[28517]_  & \new_[28512]_ ;
  assign \new_[28522]_  = ~A167 & A168;
  assign \new_[28523]_  = ~A170 & \new_[28522]_ ;
  assign \new_[28527]_  = A202 & ~A201;
  assign \new_[28528]_  = A166 & \new_[28527]_ ;
  assign \new_[28529]_  = \new_[28528]_  & \new_[28523]_ ;
  assign \new_[28533]_  = A298 & A266;
  assign \new_[28534]_  = A265 & \new_[28533]_ ;
  assign \new_[28538]_  = A302 & A300;
  assign \new_[28539]_  = ~A299 & \new_[28538]_ ;
  assign \new_[28540]_  = \new_[28539]_  & \new_[28534]_ ;
  assign \new_[28544]_  = ~A167 & A168;
  assign \new_[28545]_  = ~A170 & \new_[28544]_ ;
  assign \new_[28549]_  = A202 & ~A201;
  assign \new_[28550]_  = A166 & \new_[28549]_ ;
  assign \new_[28551]_  = \new_[28550]_  & \new_[28545]_ ;
  assign \new_[28555]_  = ~A298 & A266;
  assign \new_[28556]_  = A265 & \new_[28555]_ ;
  assign \new_[28560]_  = A301 & A300;
  assign \new_[28561]_  = A299 & \new_[28560]_ ;
  assign \new_[28562]_  = \new_[28561]_  & \new_[28556]_ ;
  assign \new_[28566]_  = ~A167 & A168;
  assign \new_[28567]_  = ~A170 & \new_[28566]_ ;
  assign \new_[28571]_  = A202 & ~A201;
  assign \new_[28572]_  = A166 & \new_[28571]_ ;
  assign \new_[28573]_  = \new_[28572]_  & \new_[28567]_ ;
  assign \new_[28577]_  = ~A298 & A266;
  assign \new_[28578]_  = A265 & \new_[28577]_ ;
  assign \new_[28582]_  = A302 & A300;
  assign \new_[28583]_  = A299 & \new_[28582]_ ;
  assign \new_[28584]_  = \new_[28583]_  & \new_[28578]_ ;
  assign \new_[28588]_  = ~A167 & A168;
  assign \new_[28589]_  = ~A170 & \new_[28588]_ ;
  assign \new_[28593]_  = A202 & ~A201;
  assign \new_[28594]_  = A166 & \new_[28593]_ ;
  assign \new_[28595]_  = \new_[28594]_  & \new_[28589]_ ;
  assign \new_[28599]_  = A298 & ~A266;
  assign \new_[28600]_  = ~A265 & \new_[28599]_ ;
  assign \new_[28604]_  = A301 & A300;
  assign \new_[28605]_  = ~A299 & \new_[28604]_ ;
  assign \new_[28606]_  = \new_[28605]_  & \new_[28600]_ ;
  assign \new_[28610]_  = ~A167 & A168;
  assign \new_[28611]_  = ~A170 & \new_[28610]_ ;
  assign \new_[28615]_  = A202 & ~A201;
  assign \new_[28616]_  = A166 & \new_[28615]_ ;
  assign \new_[28617]_  = \new_[28616]_  & \new_[28611]_ ;
  assign \new_[28621]_  = A298 & ~A266;
  assign \new_[28622]_  = ~A265 & \new_[28621]_ ;
  assign \new_[28626]_  = A302 & A300;
  assign \new_[28627]_  = ~A299 & \new_[28626]_ ;
  assign \new_[28628]_  = \new_[28627]_  & \new_[28622]_ ;
  assign \new_[28632]_  = ~A167 & A168;
  assign \new_[28633]_  = ~A170 & \new_[28632]_ ;
  assign \new_[28637]_  = A202 & ~A201;
  assign \new_[28638]_  = A166 & \new_[28637]_ ;
  assign \new_[28639]_  = \new_[28638]_  & \new_[28633]_ ;
  assign \new_[28643]_  = ~A298 & ~A266;
  assign \new_[28644]_  = ~A265 & \new_[28643]_ ;
  assign \new_[28648]_  = A301 & A300;
  assign \new_[28649]_  = A299 & \new_[28648]_ ;
  assign \new_[28650]_  = \new_[28649]_  & \new_[28644]_ ;
  assign \new_[28654]_  = ~A167 & A168;
  assign \new_[28655]_  = ~A170 & \new_[28654]_ ;
  assign \new_[28659]_  = A202 & ~A201;
  assign \new_[28660]_  = A166 & \new_[28659]_ ;
  assign \new_[28661]_  = \new_[28660]_  & \new_[28655]_ ;
  assign \new_[28665]_  = ~A298 & ~A266;
  assign \new_[28666]_  = ~A265 & \new_[28665]_ ;
  assign \new_[28670]_  = A302 & A300;
  assign \new_[28671]_  = A299 & \new_[28670]_ ;
  assign \new_[28672]_  = \new_[28671]_  & \new_[28666]_ ;
  assign \new_[28676]_  = ~A167 & A168;
  assign \new_[28677]_  = ~A170 & \new_[28676]_ ;
  assign \new_[28681]_  = A203 & ~A201;
  assign \new_[28682]_  = A166 & \new_[28681]_ ;
  assign \new_[28683]_  = \new_[28682]_  & \new_[28677]_ ;
  assign \new_[28687]_  = A298 & A268;
  assign \new_[28688]_  = ~A267 & \new_[28687]_ ;
  assign \new_[28692]_  = A301 & A300;
  assign \new_[28693]_  = ~A299 & \new_[28692]_ ;
  assign \new_[28694]_  = \new_[28693]_  & \new_[28688]_ ;
  assign \new_[28698]_  = ~A167 & A168;
  assign \new_[28699]_  = ~A170 & \new_[28698]_ ;
  assign \new_[28703]_  = A203 & ~A201;
  assign \new_[28704]_  = A166 & \new_[28703]_ ;
  assign \new_[28705]_  = \new_[28704]_  & \new_[28699]_ ;
  assign \new_[28709]_  = A298 & A268;
  assign \new_[28710]_  = ~A267 & \new_[28709]_ ;
  assign \new_[28714]_  = A302 & A300;
  assign \new_[28715]_  = ~A299 & \new_[28714]_ ;
  assign \new_[28716]_  = \new_[28715]_  & \new_[28710]_ ;
  assign \new_[28720]_  = ~A167 & A168;
  assign \new_[28721]_  = ~A170 & \new_[28720]_ ;
  assign \new_[28725]_  = A203 & ~A201;
  assign \new_[28726]_  = A166 & \new_[28725]_ ;
  assign \new_[28727]_  = \new_[28726]_  & \new_[28721]_ ;
  assign \new_[28731]_  = ~A298 & A268;
  assign \new_[28732]_  = ~A267 & \new_[28731]_ ;
  assign \new_[28736]_  = A301 & A300;
  assign \new_[28737]_  = A299 & \new_[28736]_ ;
  assign \new_[28738]_  = \new_[28737]_  & \new_[28732]_ ;
  assign \new_[28742]_  = ~A167 & A168;
  assign \new_[28743]_  = ~A170 & \new_[28742]_ ;
  assign \new_[28747]_  = A203 & ~A201;
  assign \new_[28748]_  = A166 & \new_[28747]_ ;
  assign \new_[28749]_  = \new_[28748]_  & \new_[28743]_ ;
  assign \new_[28753]_  = ~A298 & A268;
  assign \new_[28754]_  = ~A267 & \new_[28753]_ ;
  assign \new_[28758]_  = A302 & A300;
  assign \new_[28759]_  = A299 & \new_[28758]_ ;
  assign \new_[28760]_  = \new_[28759]_  & \new_[28754]_ ;
  assign \new_[28764]_  = ~A167 & A168;
  assign \new_[28765]_  = ~A170 & \new_[28764]_ ;
  assign \new_[28769]_  = A203 & ~A201;
  assign \new_[28770]_  = A166 & \new_[28769]_ ;
  assign \new_[28771]_  = \new_[28770]_  & \new_[28765]_ ;
  assign \new_[28775]_  = A298 & A269;
  assign \new_[28776]_  = ~A267 & \new_[28775]_ ;
  assign \new_[28780]_  = A301 & A300;
  assign \new_[28781]_  = ~A299 & \new_[28780]_ ;
  assign \new_[28782]_  = \new_[28781]_  & \new_[28776]_ ;
  assign \new_[28786]_  = ~A167 & A168;
  assign \new_[28787]_  = ~A170 & \new_[28786]_ ;
  assign \new_[28791]_  = A203 & ~A201;
  assign \new_[28792]_  = A166 & \new_[28791]_ ;
  assign \new_[28793]_  = \new_[28792]_  & \new_[28787]_ ;
  assign \new_[28797]_  = A298 & A269;
  assign \new_[28798]_  = ~A267 & \new_[28797]_ ;
  assign \new_[28802]_  = A302 & A300;
  assign \new_[28803]_  = ~A299 & \new_[28802]_ ;
  assign \new_[28804]_  = \new_[28803]_  & \new_[28798]_ ;
  assign \new_[28808]_  = ~A167 & A168;
  assign \new_[28809]_  = ~A170 & \new_[28808]_ ;
  assign \new_[28813]_  = A203 & ~A201;
  assign \new_[28814]_  = A166 & \new_[28813]_ ;
  assign \new_[28815]_  = \new_[28814]_  & \new_[28809]_ ;
  assign \new_[28819]_  = ~A298 & A269;
  assign \new_[28820]_  = ~A267 & \new_[28819]_ ;
  assign \new_[28824]_  = A301 & A300;
  assign \new_[28825]_  = A299 & \new_[28824]_ ;
  assign \new_[28826]_  = \new_[28825]_  & \new_[28820]_ ;
  assign \new_[28830]_  = ~A167 & A168;
  assign \new_[28831]_  = ~A170 & \new_[28830]_ ;
  assign \new_[28835]_  = A203 & ~A201;
  assign \new_[28836]_  = A166 & \new_[28835]_ ;
  assign \new_[28837]_  = \new_[28836]_  & \new_[28831]_ ;
  assign \new_[28841]_  = ~A298 & A269;
  assign \new_[28842]_  = ~A267 & \new_[28841]_ ;
  assign \new_[28846]_  = A302 & A300;
  assign \new_[28847]_  = A299 & \new_[28846]_ ;
  assign \new_[28848]_  = \new_[28847]_  & \new_[28842]_ ;
  assign \new_[28852]_  = ~A167 & A168;
  assign \new_[28853]_  = ~A170 & \new_[28852]_ ;
  assign \new_[28857]_  = A203 & ~A201;
  assign \new_[28858]_  = A166 & \new_[28857]_ ;
  assign \new_[28859]_  = \new_[28858]_  & \new_[28853]_ ;
  assign \new_[28863]_  = A298 & A266;
  assign \new_[28864]_  = A265 & \new_[28863]_ ;
  assign \new_[28868]_  = A301 & A300;
  assign \new_[28869]_  = ~A299 & \new_[28868]_ ;
  assign \new_[28870]_  = \new_[28869]_  & \new_[28864]_ ;
  assign \new_[28874]_  = ~A167 & A168;
  assign \new_[28875]_  = ~A170 & \new_[28874]_ ;
  assign \new_[28879]_  = A203 & ~A201;
  assign \new_[28880]_  = A166 & \new_[28879]_ ;
  assign \new_[28881]_  = \new_[28880]_  & \new_[28875]_ ;
  assign \new_[28885]_  = A298 & A266;
  assign \new_[28886]_  = A265 & \new_[28885]_ ;
  assign \new_[28890]_  = A302 & A300;
  assign \new_[28891]_  = ~A299 & \new_[28890]_ ;
  assign \new_[28892]_  = \new_[28891]_  & \new_[28886]_ ;
  assign \new_[28896]_  = ~A167 & A168;
  assign \new_[28897]_  = ~A170 & \new_[28896]_ ;
  assign \new_[28901]_  = A203 & ~A201;
  assign \new_[28902]_  = A166 & \new_[28901]_ ;
  assign \new_[28903]_  = \new_[28902]_  & \new_[28897]_ ;
  assign \new_[28907]_  = ~A298 & A266;
  assign \new_[28908]_  = A265 & \new_[28907]_ ;
  assign \new_[28912]_  = A301 & A300;
  assign \new_[28913]_  = A299 & \new_[28912]_ ;
  assign \new_[28914]_  = \new_[28913]_  & \new_[28908]_ ;
  assign \new_[28918]_  = ~A167 & A168;
  assign \new_[28919]_  = ~A170 & \new_[28918]_ ;
  assign \new_[28923]_  = A203 & ~A201;
  assign \new_[28924]_  = A166 & \new_[28923]_ ;
  assign \new_[28925]_  = \new_[28924]_  & \new_[28919]_ ;
  assign \new_[28929]_  = ~A298 & A266;
  assign \new_[28930]_  = A265 & \new_[28929]_ ;
  assign \new_[28934]_  = A302 & A300;
  assign \new_[28935]_  = A299 & \new_[28934]_ ;
  assign \new_[28936]_  = \new_[28935]_  & \new_[28930]_ ;
  assign \new_[28940]_  = ~A167 & A168;
  assign \new_[28941]_  = ~A170 & \new_[28940]_ ;
  assign \new_[28945]_  = A203 & ~A201;
  assign \new_[28946]_  = A166 & \new_[28945]_ ;
  assign \new_[28947]_  = \new_[28946]_  & \new_[28941]_ ;
  assign \new_[28951]_  = A298 & ~A266;
  assign \new_[28952]_  = ~A265 & \new_[28951]_ ;
  assign \new_[28956]_  = A301 & A300;
  assign \new_[28957]_  = ~A299 & \new_[28956]_ ;
  assign \new_[28958]_  = \new_[28957]_  & \new_[28952]_ ;
  assign \new_[28962]_  = ~A167 & A168;
  assign \new_[28963]_  = ~A170 & \new_[28962]_ ;
  assign \new_[28967]_  = A203 & ~A201;
  assign \new_[28968]_  = A166 & \new_[28967]_ ;
  assign \new_[28969]_  = \new_[28968]_  & \new_[28963]_ ;
  assign \new_[28973]_  = A298 & ~A266;
  assign \new_[28974]_  = ~A265 & \new_[28973]_ ;
  assign \new_[28978]_  = A302 & A300;
  assign \new_[28979]_  = ~A299 & \new_[28978]_ ;
  assign \new_[28980]_  = \new_[28979]_  & \new_[28974]_ ;
  assign \new_[28984]_  = ~A167 & A168;
  assign \new_[28985]_  = ~A170 & \new_[28984]_ ;
  assign \new_[28989]_  = A203 & ~A201;
  assign \new_[28990]_  = A166 & \new_[28989]_ ;
  assign \new_[28991]_  = \new_[28990]_  & \new_[28985]_ ;
  assign \new_[28995]_  = ~A298 & ~A266;
  assign \new_[28996]_  = ~A265 & \new_[28995]_ ;
  assign \new_[29000]_  = A301 & A300;
  assign \new_[29001]_  = A299 & \new_[29000]_ ;
  assign \new_[29002]_  = \new_[29001]_  & \new_[28996]_ ;
  assign \new_[29006]_  = ~A167 & A168;
  assign \new_[29007]_  = ~A170 & \new_[29006]_ ;
  assign \new_[29011]_  = A203 & ~A201;
  assign \new_[29012]_  = A166 & \new_[29011]_ ;
  assign \new_[29013]_  = \new_[29012]_  & \new_[29007]_ ;
  assign \new_[29017]_  = ~A298 & ~A266;
  assign \new_[29018]_  = ~A265 & \new_[29017]_ ;
  assign \new_[29022]_  = A302 & A300;
  assign \new_[29023]_  = A299 & \new_[29022]_ ;
  assign \new_[29024]_  = \new_[29023]_  & \new_[29018]_ ;
  assign \new_[29028]_  = ~A167 & A168;
  assign \new_[29029]_  = ~A170 & \new_[29028]_ ;
  assign \new_[29033]_  = A200 & A199;
  assign \new_[29034]_  = A166 & \new_[29033]_ ;
  assign \new_[29035]_  = \new_[29034]_  & \new_[29029]_ ;
  assign \new_[29039]_  = A298 & A268;
  assign \new_[29040]_  = ~A267 & \new_[29039]_ ;
  assign \new_[29044]_  = A301 & A300;
  assign \new_[29045]_  = ~A299 & \new_[29044]_ ;
  assign \new_[29046]_  = \new_[29045]_  & \new_[29040]_ ;
  assign \new_[29050]_  = ~A167 & A168;
  assign \new_[29051]_  = ~A170 & \new_[29050]_ ;
  assign \new_[29055]_  = A200 & A199;
  assign \new_[29056]_  = A166 & \new_[29055]_ ;
  assign \new_[29057]_  = \new_[29056]_  & \new_[29051]_ ;
  assign \new_[29061]_  = A298 & A268;
  assign \new_[29062]_  = ~A267 & \new_[29061]_ ;
  assign \new_[29066]_  = A302 & A300;
  assign \new_[29067]_  = ~A299 & \new_[29066]_ ;
  assign \new_[29068]_  = \new_[29067]_  & \new_[29062]_ ;
  assign \new_[29072]_  = ~A167 & A168;
  assign \new_[29073]_  = ~A170 & \new_[29072]_ ;
  assign \new_[29077]_  = A200 & A199;
  assign \new_[29078]_  = A166 & \new_[29077]_ ;
  assign \new_[29079]_  = \new_[29078]_  & \new_[29073]_ ;
  assign \new_[29083]_  = ~A298 & A268;
  assign \new_[29084]_  = ~A267 & \new_[29083]_ ;
  assign \new_[29088]_  = A301 & A300;
  assign \new_[29089]_  = A299 & \new_[29088]_ ;
  assign \new_[29090]_  = \new_[29089]_  & \new_[29084]_ ;
  assign \new_[29094]_  = ~A167 & A168;
  assign \new_[29095]_  = ~A170 & \new_[29094]_ ;
  assign \new_[29099]_  = A200 & A199;
  assign \new_[29100]_  = A166 & \new_[29099]_ ;
  assign \new_[29101]_  = \new_[29100]_  & \new_[29095]_ ;
  assign \new_[29105]_  = ~A298 & A268;
  assign \new_[29106]_  = ~A267 & \new_[29105]_ ;
  assign \new_[29110]_  = A302 & A300;
  assign \new_[29111]_  = A299 & \new_[29110]_ ;
  assign \new_[29112]_  = \new_[29111]_  & \new_[29106]_ ;
  assign \new_[29116]_  = ~A167 & A168;
  assign \new_[29117]_  = ~A170 & \new_[29116]_ ;
  assign \new_[29121]_  = A200 & A199;
  assign \new_[29122]_  = A166 & \new_[29121]_ ;
  assign \new_[29123]_  = \new_[29122]_  & \new_[29117]_ ;
  assign \new_[29127]_  = A298 & A269;
  assign \new_[29128]_  = ~A267 & \new_[29127]_ ;
  assign \new_[29132]_  = A301 & A300;
  assign \new_[29133]_  = ~A299 & \new_[29132]_ ;
  assign \new_[29134]_  = \new_[29133]_  & \new_[29128]_ ;
  assign \new_[29138]_  = ~A167 & A168;
  assign \new_[29139]_  = ~A170 & \new_[29138]_ ;
  assign \new_[29143]_  = A200 & A199;
  assign \new_[29144]_  = A166 & \new_[29143]_ ;
  assign \new_[29145]_  = \new_[29144]_  & \new_[29139]_ ;
  assign \new_[29149]_  = A298 & A269;
  assign \new_[29150]_  = ~A267 & \new_[29149]_ ;
  assign \new_[29154]_  = A302 & A300;
  assign \new_[29155]_  = ~A299 & \new_[29154]_ ;
  assign \new_[29156]_  = \new_[29155]_  & \new_[29150]_ ;
  assign \new_[29160]_  = ~A167 & A168;
  assign \new_[29161]_  = ~A170 & \new_[29160]_ ;
  assign \new_[29165]_  = A200 & A199;
  assign \new_[29166]_  = A166 & \new_[29165]_ ;
  assign \new_[29167]_  = \new_[29166]_  & \new_[29161]_ ;
  assign \new_[29171]_  = ~A298 & A269;
  assign \new_[29172]_  = ~A267 & \new_[29171]_ ;
  assign \new_[29176]_  = A301 & A300;
  assign \new_[29177]_  = A299 & \new_[29176]_ ;
  assign \new_[29178]_  = \new_[29177]_  & \new_[29172]_ ;
  assign \new_[29182]_  = ~A167 & A168;
  assign \new_[29183]_  = ~A170 & \new_[29182]_ ;
  assign \new_[29187]_  = A200 & A199;
  assign \new_[29188]_  = A166 & \new_[29187]_ ;
  assign \new_[29189]_  = \new_[29188]_  & \new_[29183]_ ;
  assign \new_[29193]_  = ~A298 & A269;
  assign \new_[29194]_  = ~A267 & \new_[29193]_ ;
  assign \new_[29198]_  = A302 & A300;
  assign \new_[29199]_  = A299 & \new_[29198]_ ;
  assign \new_[29200]_  = \new_[29199]_  & \new_[29194]_ ;
  assign \new_[29204]_  = ~A167 & A168;
  assign \new_[29205]_  = ~A170 & \new_[29204]_ ;
  assign \new_[29209]_  = A200 & A199;
  assign \new_[29210]_  = A166 & \new_[29209]_ ;
  assign \new_[29211]_  = \new_[29210]_  & \new_[29205]_ ;
  assign \new_[29215]_  = A298 & A266;
  assign \new_[29216]_  = A265 & \new_[29215]_ ;
  assign \new_[29220]_  = A301 & A300;
  assign \new_[29221]_  = ~A299 & \new_[29220]_ ;
  assign \new_[29222]_  = \new_[29221]_  & \new_[29216]_ ;
  assign \new_[29226]_  = ~A167 & A168;
  assign \new_[29227]_  = ~A170 & \new_[29226]_ ;
  assign \new_[29231]_  = A200 & A199;
  assign \new_[29232]_  = A166 & \new_[29231]_ ;
  assign \new_[29233]_  = \new_[29232]_  & \new_[29227]_ ;
  assign \new_[29237]_  = A298 & A266;
  assign \new_[29238]_  = A265 & \new_[29237]_ ;
  assign \new_[29242]_  = A302 & A300;
  assign \new_[29243]_  = ~A299 & \new_[29242]_ ;
  assign \new_[29244]_  = \new_[29243]_  & \new_[29238]_ ;
  assign \new_[29248]_  = ~A167 & A168;
  assign \new_[29249]_  = ~A170 & \new_[29248]_ ;
  assign \new_[29253]_  = A200 & A199;
  assign \new_[29254]_  = A166 & \new_[29253]_ ;
  assign \new_[29255]_  = \new_[29254]_  & \new_[29249]_ ;
  assign \new_[29259]_  = ~A298 & A266;
  assign \new_[29260]_  = A265 & \new_[29259]_ ;
  assign \new_[29264]_  = A301 & A300;
  assign \new_[29265]_  = A299 & \new_[29264]_ ;
  assign \new_[29266]_  = \new_[29265]_  & \new_[29260]_ ;
  assign \new_[29270]_  = ~A167 & A168;
  assign \new_[29271]_  = ~A170 & \new_[29270]_ ;
  assign \new_[29275]_  = A200 & A199;
  assign \new_[29276]_  = A166 & \new_[29275]_ ;
  assign \new_[29277]_  = \new_[29276]_  & \new_[29271]_ ;
  assign \new_[29281]_  = ~A298 & A266;
  assign \new_[29282]_  = A265 & \new_[29281]_ ;
  assign \new_[29286]_  = A302 & A300;
  assign \new_[29287]_  = A299 & \new_[29286]_ ;
  assign \new_[29288]_  = \new_[29287]_  & \new_[29282]_ ;
  assign \new_[29292]_  = ~A167 & A168;
  assign \new_[29293]_  = ~A170 & \new_[29292]_ ;
  assign \new_[29297]_  = A200 & A199;
  assign \new_[29298]_  = A166 & \new_[29297]_ ;
  assign \new_[29299]_  = \new_[29298]_  & \new_[29293]_ ;
  assign \new_[29303]_  = A298 & ~A266;
  assign \new_[29304]_  = ~A265 & \new_[29303]_ ;
  assign \new_[29308]_  = A301 & A300;
  assign \new_[29309]_  = ~A299 & \new_[29308]_ ;
  assign \new_[29310]_  = \new_[29309]_  & \new_[29304]_ ;
  assign \new_[29314]_  = ~A167 & A168;
  assign \new_[29315]_  = ~A170 & \new_[29314]_ ;
  assign \new_[29319]_  = A200 & A199;
  assign \new_[29320]_  = A166 & \new_[29319]_ ;
  assign \new_[29321]_  = \new_[29320]_  & \new_[29315]_ ;
  assign \new_[29325]_  = A298 & ~A266;
  assign \new_[29326]_  = ~A265 & \new_[29325]_ ;
  assign \new_[29330]_  = A302 & A300;
  assign \new_[29331]_  = ~A299 & \new_[29330]_ ;
  assign \new_[29332]_  = \new_[29331]_  & \new_[29326]_ ;
  assign \new_[29336]_  = ~A167 & A168;
  assign \new_[29337]_  = ~A170 & \new_[29336]_ ;
  assign \new_[29341]_  = A200 & A199;
  assign \new_[29342]_  = A166 & \new_[29341]_ ;
  assign \new_[29343]_  = \new_[29342]_  & \new_[29337]_ ;
  assign \new_[29347]_  = ~A298 & ~A266;
  assign \new_[29348]_  = ~A265 & \new_[29347]_ ;
  assign \new_[29352]_  = A301 & A300;
  assign \new_[29353]_  = A299 & \new_[29352]_ ;
  assign \new_[29354]_  = \new_[29353]_  & \new_[29348]_ ;
  assign \new_[29358]_  = ~A167 & A168;
  assign \new_[29359]_  = ~A170 & \new_[29358]_ ;
  assign \new_[29363]_  = A200 & A199;
  assign \new_[29364]_  = A166 & \new_[29363]_ ;
  assign \new_[29365]_  = \new_[29364]_  & \new_[29359]_ ;
  assign \new_[29369]_  = ~A298 & ~A266;
  assign \new_[29370]_  = ~A265 & \new_[29369]_ ;
  assign \new_[29374]_  = A302 & A300;
  assign \new_[29375]_  = A299 & \new_[29374]_ ;
  assign \new_[29376]_  = \new_[29375]_  & \new_[29370]_ ;
  assign \new_[29380]_  = ~A167 & A168;
  assign \new_[29381]_  = ~A170 & \new_[29380]_ ;
  assign \new_[29385]_  = ~A200 & ~A199;
  assign \new_[29386]_  = A166 & \new_[29385]_ ;
  assign \new_[29387]_  = \new_[29386]_  & \new_[29381]_ ;
  assign \new_[29391]_  = A298 & A268;
  assign \new_[29392]_  = ~A267 & \new_[29391]_ ;
  assign \new_[29396]_  = A301 & A300;
  assign \new_[29397]_  = ~A299 & \new_[29396]_ ;
  assign \new_[29398]_  = \new_[29397]_  & \new_[29392]_ ;
  assign \new_[29402]_  = ~A167 & A168;
  assign \new_[29403]_  = ~A170 & \new_[29402]_ ;
  assign \new_[29407]_  = ~A200 & ~A199;
  assign \new_[29408]_  = A166 & \new_[29407]_ ;
  assign \new_[29409]_  = \new_[29408]_  & \new_[29403]_ ;
  assign \new_[29413]_  = A298 & A268;
  assign \new_[29414]_  = ~A267 & \new_[29413]_ ;
  assign \new_[29418]_  = A302 & A300;
  assign \new_[29419]_  = ~A299 & \new_[29418]_ ;
  assign \new_[29420]_  = \new_[29419]_  & \new_[29414]_ ;
  assign \new_[29424]_  = ~A167 & A168;
  assign \new_[29425]_  = ~A170 & \new_[29424]_ ;
  assign \new_[29429]_  = ~A200 & ~A199;
  assign \new_[29430]_  = A166 & \new_[29429]_ ;
  assign \new_[29431]_  = \new_[29430]_  & \new_[29425]_ ;
  assign \new_[29435]_  = ~A298 & A268;
  assign \new_[29436]_  = ~A267 & \new_[29435]_ ;
  assign \new_[29440]_  = A301 & A300;
  assign \new_[29441]_  = A299 & \new_[29440]_ ;
  assign \new_[29442]_  = \new_[29441]_  & \new_[29436]_ ;
  assign \new_[29446]_  = ~A167 & A168;
  assign \new_[29447]_  = ~A170 & \new_[29446]_ ;
  assign \new_[29451]_  = ~A200 & ~A199;
  assign \new_[29452]_  = A166 & \new_[29451]_ ;
  assign \new_[29453]_  = \new_[29452]_  & \new_[29447]_ ;
  assign \new_[29457]_  = ~A298 & A268;
  assign \new_[29458]_  = ~A267 & \new_[29457]_ ;
  assign \new_[29462]_  = A302 & A300;
  assign \new_[29463]_  = A299 & \new_[29462]_ ;
  assign \new_[29464]_  = \new_[29463]_  & \new_[29458]_ ;
  assign \new_[29468]_  = ~A167 & A168;
  assign \new_[29469]_  = ~A170 & \new_[29468]_ ;
  assign \new_[29473]_  = ~A200 & ~A199;
  assign \new_[29474]_  = A166 & \new_[29473]_ ;
  assign \new_[29475]_  = \new_[29474]_  & \new_[29469]_ ;
  assign \new_[29479]_  = A298 & A269;
  assign \new_[29480]_  = ~A267 & \new_[29479]_ ;
  assign \new_[29484]_  = A301 & A300;
  assign \new_[29485]_  = ~A299 & \new_[29484]_ ;
  assign \new_[29486]_  = \new_[29485]_  & \new_[29480]_ ;
  assign \new_[29490]_  = ~A167 & A168;
  assign \new_[29491]_  = ~A170 & \new_[29490]_ ;
  assign \new_[29495]_  = ~A200 & ~A199;
  assign \new_[29496]_  = A166 & \new_[29495]_ ;
  assign \new_[29497]_  = \new_[29496]_  & \new_[29491]_ ;
  assign \new_[29501]_  = A298 & A269;
  assign \new_[29502]_  = ~A267 & \new_[29501]_ ;
  assign \new_[29506]_  = A302 & A300;
  assign \new_[29507]_  = ~A299 & \new_[29506]_ ;
  assign \new_[29508]_  = \new_[29507]_  & \new_[29502]_ ;
  assign \new_[29512]_  = ~A167 & A168;
  assign \new_[29513]_  = ~A170 & \new_[29512]_ ;
  assign \new_[29517]_  = ~A200 & ~A199;
  assign \new_[29518]_  = A166 & \new_[29517]_ ;
  assign \new_[29519]_  = \new_[29518]_  & \new_[29513]_ ;
  assign \new_[29523]_  = ~A298 & A269;
  assign \new_[29524]_  = ~A267 & \new_[29523]_ ;
  assign \new_[29528]_  = A301 & A300;
  assign \new_[29529]_  = A299 & \new_[29528]_ ;
  assign \new_[29530]_  = \new_[29529]_  & \new_[29524]_ ;
  assign \new_[29534]_  = ~A167 & A168;
  assign \new_[29535]_  = ~A170 & \new_[29534]_ ;
  assign \new_[29539]_  = ~A200 & ~A199;
  assign \new_[29540]_  = A166 & \new_[29539]_ ;
  assign \new_[29541]_  = \new_[29540]_  & \new_[29535]_ ;
  assign \new_[29545]_  = ~A298 & A269;
  assign \new_[29546]_  = ~A267 & \new_[29545]_ ;
  assign \new_[29550]_  = A302 & A300;
  assign \new_[29551]_  = A299 & \new_[29550]_ ;
  assign \new_[29552]_  = \new_[29551]_  & \new_[29546]_ ;
  assign \new_[29556]_  = ~A167 & A168;
  assign \new_[29557]_  = ~A170 & \new_[29556]_ ;
  assign \new_[29561]_  = ~A200 & ~A199;
  assign \new_[29562]_  = A166 & \new_[29561]_ ;
  assign \new_[29563]_  = \new_[29562]_  & \new_[29557]_ ;
  assign \new_[29567]_  = A298 & A266;
  assign \new_[29568]_  = A265 & \new_[29567]_ ;
  assign \new_[29572]_  = A301 & A300;
  assign \new_[29573]_  = ~A299 & \new_[29572]_ ;
  assign \new_[29574]_  = \new_[29573]_  & \new_[29568]_ ;
  assign \new_[29578]_  = ~A167 & A168;
  assign \new_[29579]_  = ~A170 & \new_[29578]_ ;
  assign \new_[29583]_  = ~A200 & ~A199;
  assign \new_[29584]_  = A166 & \new_[29583]_ ;
  assign \new_[29585]_  = \new_[29584]_  & \new_[29579]_ ;
  assign \new_[29589]_  = A298 & A266;
  assign \new_[29590]_  = A265 & \new_[29589]_ ;
  assign \new_[29594]_  = A302 & A300;
  assign \new_[29595]_  = ~A299 & \new_[29594]_ ;
  assign \new_[29596]_  = \new_[29595]_  & \new_[29590]_ ;
  assign \new_[29600]_  = ~A167 & A168;
  assign \new_[29601]_  = ~A170 & \new_[29600]_ ;
  assign \new_[29605]_  = ~A200 & ~A199;
  assign \new_[29606]_  = A166 & \new_[29605]_ ;
  assign \new_[29607]_  = \new_[29606]_  & \new_[29601]_ ;
  assign \new_[29611]_  = ~A298 & A266;
  assign \new_[29612]_  = A265 & \new_[29611]_ ;
  assign \new_[29616]_  = A301 & A300;
  assign \new_[29617]_  = A299 & \new_[29616]_ ;
  assign \new_[29618]_  = \new_[29617]_  & \new_[29612]_ ;
  assign \new_[29622]_  = ~A167 & A168;
  assign \new_[29623]_  = ~A170 & \new_[29622]_ ;
  assign \new_[29627]_  = ~A200 & ~A199;
  assign \new_[29628]_  = A166 & \new_[29627]_ ;
  assign \new_[29629]_  = \new_[29628]_  & \new_[29623]_ ;
  assign \new_[29633]_  = ~A298 & A266;
  assign \new_[29634]_  = A265 & \new_[29633]_ ;
  assign \new_[29638]_  = A302 & A300;
  assign \new_[29639]_  = A299 & \new_[29638]_ ;
  assign \new_[29640]_  = \new_[29639]_  & \new_[29634]_ ;
  assign \new_[29644]_  = ~A167 & A168;
  assign \new_[29645]_  = ~A170 & \new_[29644]_ ;
  assign \new_[29649]_  = ~A200 & ~A199;
  assign \new_[29650]_  = A166 & \new_[29649]_ ;
  assign \new_[29651]_  = \new_[29650]_  & \new_[29645]_ ;
  assign \new_[29655]_  = A298 & ~A266;
  assign \new_[29656]_  = ~A265 & \new_[29655]_ ;
  assign \new_[29660]_  = A301 & A300;
  assign \new_[29661]_  = ~A299 & \new_[29660]_ ;
  assign \new_[29662]_  = \new_[29661]_  & \new_[29656]_ ;
  assign \new_[29666]_  = ~A167 & A168;
  assign \new_[29667]_  = ~A170 & \new_[29666]_ ;
  assign \new_[29671]_  = ~A200 & ~A199;
  assign \new_[29672]_  = A166 & \new_[29671]_ ;
  assign \new_[29673]_  = \new_[29672]_  & \new_[29667]_ ;
  assign \new_[29677]_  = A298 & ~A266;
  assign \new_[29678]_  = ~A265 & \new_[29677]_ ;
  assign \new_[29682]_  = A302 & A300;
  assign \new_[29683]_  = ~A299 & \new_[29682]_ ;
  assign \new_[29684]_  = \new_[29683]_  & \new_[29678]_ ;
  assign \new_[29688]_  = ~A167 & A168;
  assign \new_[29689]_  = ~A170 & \new_[29688]_ ;
  assign \new_[29693]_  = ~A200 & ~A199;
  assign \new_[29694]_  = A166 & \new_[29693]_ ;
  assign \new_[29695]_  = \new_[29694]_  & \new_[29689]_ ;
  assign \new_[29699]_  = ~A298 & ~A266;
  assign \new_[29700]_  = ~A265 & \new_[29699]_ ;
  assign \new_[29704]_  = A301 & A300;
  assign \new_[29705]_  = A299 & \new_[29704]_ ;
  assign \new_[29706]_  = \new_[29705]_  & \new_[29700]_ ;
  assign \new_[29710]_  = ~A167 & A168;
  assign \new_[29711]_  = ~A170 & \new_[29710]_ ;
  assign \new_[29715]_  = ~A200 & ~A199;
  assign \new_[29716]_  = A166 & \new_[29715]_ ;
  assign \new_[29717]_  = \new_[29716]_  & \new_[29711]_ ;
  assign \new_[29721]_  = ~A298 & ~A266;
  assign \new_[29722]_  = ~A265 & \new_[29721]_ ;
  assign \new_[29726]_  = A302 & A300;
  assign \new_[29727]_  = A299 & \new_[29726]_ ;
  assign \new_[29728]_  = \new_[29727]_  & \new_[29722]_ ;
  assign \new_[29732]_  = A201 & ~A168;
  assign \new_[29733]_  = ~A170 & \new_[29732]_ ;
  assign \new_[29737]_  = ~A265 & ~A203;
  assign \new_[29738]_  = ~A202 & \new_[29737]_ ;
  assign \new_[29739]_  = \new_[29738]_  & \new_[29733]_ ;
  assign \new_[29743]_  = A268 & A267;
  assign \new_[29744]_  = A266 & \new_[29743]_ ;
  assign \new_[29748]_  = ~A302 & ~A301;
  assign \new_[29749]_  = A300 & \new_[29748]_ ;
  assign \new_[29750]_  = \new_[29749]_  & \new_[29744]_ ;
  assign \new_[29754]_  = A201 & ~A168;
  assign \new_[29755]_  = ~A170 & \new_[29754]_ ;
  assign \new_[29759]_  = ~A265 & ~A203;
  assign \new_[29760]_  = ~A202 & \new_[29759]_ ;
  assign \new_[29761]_  = \new_[29760]_  & \new_[29755]_ ;
  assign \new_[29765]_  = A269 & A267;
  assign \new_[29766]_  = A266 & \new_[29765]_ ;
  assign \new_[29770]_  = ~A302 & ~A301;
  assign \new_[29771]_  = A300 & \new_[29770]_ ;
  assign \new_[29772]_  = \new_[29771]_  & \new_[29766]_ ;
  assign \new_[29776]_  = A201 & ~A168;
  assign \new_[29777]_  = ~A170 & \new_[29776]_ ;
  assign \new_[29781]_  = ~A265 & ~A203;
  assign \new_[29782]_  = ~A202 & \new_[29781]_ ;
  assign \new_[29783]_  = \new_[29782]_  & \new_[29777]_ ;
  assign \new_[29787]_  = ~A268 & ~A267;
  assign \new_[29788]_  = A266 & \new_[29787]_ ;
  assign \new_[29792]_  = A301 & ~A300;
  assign \new_[29793]_  = ~A269 & \new_[29792]_ ;
  assign \new_[29794]_  = \new_[29793]_  & \new_[29788]_ ;
  assign \new_[29798]_  = A201 & ~A168;
  assign \new_[29799]_  = ~A170 & \new_[29798]_ ;
  assign \new_[29803]_  = ~A265 & ~A203;
  assign \new_[29804]_  = ~A202 & \new_[29803]_ ;
  assign \new_[29805]_  = \new_[29804]_  & \new_[29799]_ ;
  assign \new_[29809]_  = ~A268 & ~A267;
  assign \new_[29810]_  = A266 & \new_[29809]_ ;
  assign \new_[29814]_  = A302 & ~A300;
  assign \new_[29815]_  = ~A269 & \new_[29814]_ ;
  assign \new_[29816]_  = \new_[29815]_  & \new_[29810]_ ;
  assign \new_[29820]_  = A201 & ~A168;
  assign \new_[29821]_  = ~A170 & \new_[29820]_ ;
  assign \new_[29825]_  = ~A265 & ~A203;
  assign \new_[29826]_  = ~A202 & \new_[29825]_ ;
  assign \new_[29827]_  = \new_[29826]_  & \new_[29821]_ ;
  assign \new_[29831]_  = ~A268 & ~A267;
  assign \new_[29832]_  = A266 & \new_[29831]_ ;
  assign \new_[29836]_  = A299 & A298;
  assign \new_[29837]_  = ~A269 & \new_[29836]_ ;
  assign \new_[29838]_  = \new_[29837]_  & \new_[29832]_ ;
  assign \new_[29842]_  = A201 & ~A168;
  assign \new_[29843]_  = ~A170 & \new_[29842]_ ;
  assign \new_[29847]_  = ~A265 & ~A203;
  assign \new_[29848]_  = ~A202 & \new_[29847]_ ;
  assign \new_[29849]_  = \new_[29848]_  & \new_[29843]_ ;
  assign \new_[29853]_  = ~A268 & ~A267;
  assign \new_[29854]_  = A266 & \new_[29853]_ ;
  assign \new_[29858]_  = ~A299 & ~A298;
  assign \new_[29859]_  = ~A269 & \new_[29858]_ ;
  assign \new_[29860]_  = \new_[29859]_  & \new_[29854]_ ;
  assign \new_[29864]_  = A201 & ~A168;
  assign \new_[29865]_  = ~A170 & \new_[29864]_ ;
  assign \new_[29869]_  = A265 & ~A203;
  assign \new_[29870]_  = ~A202 & \new_[29869]_ ;
  assign \new_[29871]_  = \new_[29870]_  & \new_[29865]_ ;
  assign \new_[29875]_  = A268 & A267;
  assign \new_[29876]_  = ~A266 & \new_[29875]_ ;
  assign \new_[29880]_  = ~A302 & ~A301;
  assign \new_[29881]_  = A300 & \new_[29880]_ ;
  assign \new_[29882]_  = \new_[29881]_  & \new_[29876]_ ;
  assign \new_[29886]_  = A201 & ~A168;
  assign \new_[29887]_  = ~A170 & \new_[29886]_ ;
  assign \new_[29891]_  = A265 & ~A203;
  assign \new_[29892]_  = ~A202 & \new_[29891]_ ;
  assign \new_[29893]_  = \new_[29892]_  & \new_[29887]_ ;
  assign \new_[29897]_  = A269 & A267;
  assign \new_[29898]_  = ~A266 & \new_[29897]_ ;
  assign \new_[29902]_  = ~A302 & ~A301;
  assign \new_[29903]_  = A300 & \new_[29902]_ ;
  assign \new_[29904]_  = \new_[29903]_  & \new_[29898]_ ;
  assign \new_[29908]_  = A201 & ~A168;
  assign \new_[29909]_  = ~A170 & \new_[29908]_ ;
  assign \new_[29913]_  = A265 & ~A203;
  assign \new_[29914]_  = ~A202 & \new_[29913]_ ;
  assign \new_[29915]_  = \new_[29914]_  & \new_[29909]_ ;
  assign \new_[29919]_  = ~A268 & ~A267;
  assign \new_[29920]_  = ~A266 & \new_[29919]_ ;
  assign \new_[29924]_  = A301 & ~A300;
  assign \new_[29925]_  = ~A269 & \new_[29924]_ ;
  assign \new_[29926]_  = \new_[29925]_  & \new_[29920]_ ;
  assign \new_[29930]_  = A201 & ~A168;
  assign \new_[29931]_  = ~A170 & \new_[29930]_ ;
  assign \new_[29935]_  = A265 & ~A203;
  assign \new_[29936]_  = ~A202 & \new_[29935]_ ;
  assign \new_[29937]_  = \new_[29936]_  & \new_[29931]_ ;
  assign \new_[29941]_  = ~A268 & ~A267;
  assign \new_[29942]_  = ~A266 & \new_[29941]_ ;
  assign \new_[29946]_  = A302 & ~A300;
  assign \new_[29947]_  = ~A269 & \new_[29946]_ ;
  assign \new_[29948]_  = \new_[29947]_  & \new_[29942]_ ;
  assign \new_[29952]_  = A201 & ~A168;
  assign \new_[29953]_  = ~A170 & \new_[29952]_ ;
  assign \new_[29957]_  = A265 & ~A203;
  assign \new_[29958]_  = ~A202 & \new_[29957]_ ;
  assign \new_[29959]_  = \new_[29958]_  & \new_[29953]_ ;
  assign \new_[29963]_  = ~A268 & ~A267;
  assign \new_[29964]_  = ~A266 & \new_[29963]_ ;
  assign \new_[29968]_  = A299 & A298;
  assign \new_[29969]_  = ~A269 & \new_[29968]_ ;
  assign \new_[29970]_  = \new_[29969]_  & \new_[29964]_ ;
  assign \new_[29974]_  = A201 & ~A168;
  assign \new_[29975]_  = ~A170 & \new_[29974]_ ;
  assign \new_[29979]_  = A265 & ~A203;
  assign \new_[29980]_  = ~A202 & \new_[29979]_ ;
  assign \new_[29981]_  = \new_[29980]_  & \new_[29975]_ ;
  assign \new_[29985]_  = ~A268 & ~A267;
  assign \new_[29986]_  = ~A266 & \new_[29985]_ ;
  assign \new_[29990]_  = ~A299 & ~A298;
  assign \new_[29991]_  = ~A269 & \new_[29990]_ ;
  assign \new_[29992]_  = \new_[29991]_  & \new_[29986]_ ;
  assign \new_[29996]_  = ~A201 & ~A168;
  assign \new_[29997]_  = ~A170 & \new_[29996]_ ;
  assign \new_[30001]_  = A266 & ~A265;
  assign \new_[30002]_  = A202 & \new_[30001]_ ;
  assign \new_[30003]_  = \new_[30002]_  & \new_[29997]_ ;
  assign \new_[30007]_  = ~A269 & ~A268;
  assign \new_[30008]_  = ~A267 & \new_[30007]_ ;
  assign \new_[30012]_  = ~A302 & ~A301;
  assign \new_[30013]_  = A300 & \new_[30012]_ ;
  assign \new_[30014]_  = \new_[30013]_  & \new_[30008]_ ;
  assign \new_[30018]_  = ~A201 & ~A168;
  assign \new_[30019]_  = ~A170 & \new_[30018]_ ;
  assign \new_[30023]_  = ~A266 & A265;
  assign \new_[30024]_  = A202 & \new_[30023]_ ;
  assign \new_[30025]_  = \new_[30024]_  & \new_[30019]_ ;
  assign \new_[30029]_  = ~A269 & ~A268;
  assign \new_[30030]_  = ~A267 & \new_[30029]_ ;
  assign \new_[30034]_  = ~A302 & ~A301;
  assign \new_[30035]_  = A300 & \new_[30034]_ ;
  assign \new_[30036]_  = \new_[30035]_  & \new_[30030]_ ;
  assign \new_[30040]_  = ~A201 & ~A168;
  assign \new_[30041]_  = ~A170 & \new_[30040]_ ;
  assign \new_[30045]_  = A266 & ~A265;
  assign \new_[30046]_  = A203 & \new_[30045]_ ;
  assign \new_[30047]_  = \new_[30046]_  & \new_[30041]_ ;
  assign \new_[30051]_  = ~A269 & ~A268;
  assign \new_[30052]_  = ~A267 & \new_[30051]_ ;
  assign \new_[30056]_  = ~A302 & ~A301;
  assign \new_[30057]_  = A300 & \new_[30056]_ ;
  assign \new_[30058]_  = \new_[30057]_  & \new_[30052]_ ;
  assign \new_[30062]_  = ~A201 & ~A168;
  assign \new_[30063]_  = ~A170 & \new_[30062]_ ;
  assign \new_[30067]_  = ~A266 & A265;
  assign \new_[30068]_  = A203 & \new_[30067]_ ;
  assign \new_[30069]_  = \new_[30068]_  & \new_[30063]_ ;
  assign \new_[30073]_  = ~A269 & ~A268;
  assign \new_[30074]_  = ~A267 & \new_[30073]_ ;
  assign \new_[30078]_  = ~A302 & ~A301;
  assign \new_[30079]_  = A300 & \new_[30078]_ ;
  assign \new_[30080]_  = \new_[30079]_  & \new_[30074]_ ;
  assign \new_[30084]_  = A199 & ~A168;
  assign \new_[30085]_  = ~A170 & \new_[30084]_ ;
  assign \new_[30089]_  = A266 & ~A265;
  assign \new_[30090]_  = A200 & \new_[30089]_ ;
  assign \new_[30091]_  = \new_[30090]_  & \new_[30085]_ ;
  assign \new_[30095]_  = ~A269 & ~A268;
  assign \new_[30096]_  = ~A267 & \new_[30095]_ ;
  assign \new_[30100]_  = ~A302 & ~A301;
  assign \new_[30101]_  = A300 & \new_[30100]_ ;
  assign \new_[30102]_  = \new_[30101]_  & \new_[30096]_ ;
  assign \new_[30106]_  = A199 & ~A168;
  assign \new_[30107]_  = ~A170 & \new_[30106]_ ;
  assign \new_[30111]_  = ~A266 & A265;
  assign \new_[30112]_  = A200 & \new_[30111]_ ;
  assign \new_[30113]_  = \new_[30112]_  & \new_[30107]_ ;
  assign \new_[30117]_  = ~A269 & ~A268;
  assign \new_[30118]_  = ~A267 & \new_[30117]_ ;
  assign \new_[30122]_  = ~A302 & ~A301;
  assign \new_[30123]_  = A300 & \new_[30122]_ ;
  assign \new_[30124]_  = \new_[30123]_  & \new_[30118]_ ;
  assign \new_[30128]_  = ~A199 & ~A168;
  assign \new_[30129]_  = ~A170 & \new_[30128]_ ;
  assign \new_[30133]_  = A202 & A201;
  assign \new_[30134]_  = A200 & \new_[30133]_ ;
  assign \new_[30135]_  = \new_[30134]_  & \new_[30129]_ ;
  assign \new_[30139]_  = A298 & A268;
  assign \new_[30140]_  = ~A267 & \new_[30139]_ ;
  assign \new_[30144]_  = A301 & A300;
  assign \new_[30145]_  = ~A299 & \new_[30144]_ ;
  assign \new_[30146]_  = \new_[30145]_  & \new_[30140]_ ;
  assign \new_[30150]_  = ~A199 & ~A168;
  assign \new_[30151]_  = ~A170 & \new_[30150]_ ;
  assign \new_[30155]_  = A202 & A201;
  assign \new_[30156]_  = A200 & \new_[30155]_ ;
  assign \new_[30157]_  = \new_[30156]_  & \new_[30151]_ ;
  assign \new_[30161]_  = A298 & A268;
  assign \new_[30162]_  = ~A267 & \new_[30161]_ ;
  assign \new_[30166]_  = A302 & A300;
  assign \new_[30167]_  = ~A299 & \new_[30166]_ ;
  assign \new_[30168]_  = \new_[30167]_  & \new_[30162]_ ;
  assign \new_[30172]_  = ~A199 & ~A168;
  assign \new_[30173]_  = ~A170 & \new_[30172]_ ;
  assign \new_[30177]_  = A202 & A201;
  assign \new_[30178]_  = A200 & \new_[30177]_ ;
  assign \new_[30179]_  = \new_[30178]_  & \new_[30173]_ ;
  assign \new_[30183]_  = ~A298 & A268;
  assign \new_[30184]_  = ~A267 & \new_[30183]_ ;
  assign \new_[30188]_  = A301 & A300;
  assign \new_[30189]_  = A299 & \new_[30188]_ ;
  assign \new_[30190]_  = \new_[30189]_  & \new_[30184]_ ;
  assign \new_[30194]_  = ~A199 & ~A168;
  assign \new_[30195]_  = ~A170 & \new_[30194]_ ;
  assign \new_[30199]_  = A202 & A201;
  assign \new_[30200]_  = A200 & \new_[30199]_ ;
  assign \new_[30201]_  = \new_[30200]_  & \new_[30195]_ ;
  assign \new_[30205]_  = ~A298 & A268;
  assign \new_[30206]_  = ~A267 & \new_[30205]_ ;
  assign \new_[30210]_  = A302 & A300;
  assign \new_[30211]_  = A299 & \new_[30210]_ ;
  assign \new_[30212]_  = \new_[30211]_  & \new_[30206]_ ;
  assign \new_[30216]_  = ~A199 & ~A168;
  assign \new_[30217]_  = ~A170 & \new_[30216]_ ;
  assign \new_[30221]_  = A202 & A201;
  assign \new_[30222]_  = A200 & \new_[30221]_ ;
  assign \new_[30223]_  = \new_[30222]_  & \new_[30217]_ ;
  assign \new_[30227]_  = A298 & A269;
  assign \new_[30228]_  = ~A267 & \new_[30227]_ ;
  assign \new_[30232]_  = A301 & A300;
  assign \new_[30233]_  = ~A299 & \new_[30232]_ ;
  assign \new_[30234]_  = \new_[30233]_  & \new_[30228]_ ;
  assign \new_[30238]_  = ~A199 & ~A168;
  assign \new_[30239]_  = ~A170 & \new_[30238]_ ;
  assign \new_[30243]_  = A202 & A201;
  assign \new_[30244]_  = A200 & \new_[30243]_ ;
  assign \new_[30245]_  = \new_[30244]_  & \new_[30239]_ ;
  assign \new_[30249]_  = A298 & A269;
  assign \new_[30250]_  = ~A267 & \new_[30249]_ ;
  assign \new_[30254]_  = A302 & A300;
  assign \new_[30255]_  = ~A299 & \new_[30254]_ ;
  assign \new_[30256]_  = \new_[30255]_  & \new_[30250]_ ;
  assign \new_[30260]_  = ~A199 & ~A168;
  assign \new_[30261]_  = ~A170 & \new_[30260]_ ;
  assign \new_[30265]_  = A202 & A201;
  assign \new_[30266]_  = A200 & \new_[30265]_ ;
  assign \new_[30267]_  = \new_[30266]_  & \new_[30261]_ ;
  assign \new_[30271]_  = ~A298 & A269;
  assign \new_[30272]_  = ~A267 & \new_[30271]_ ;
  assign \new_[30276]_  = A301 & A300;
  assign \new_[30277]_  = A299 & \new_[30276]_ ;
  assign \new_[30278]_  = \new_[30277]_  & \new_[30272]_ ;
  assign \new_[30282]_  = ~A199 & ~A168;
  assign \new_[30283]_  = ~A170 & \new_[30282]_ ;
  assign \new_[30287]_  = A202 & A201;
  assign \new_[30288]_  = A200 & \new_[30287]_ ;
  assign \new_[30289]_  = \new_[30288]_  & \new_[30283]_ ;
  assign \new_[30293]_  = ~A298 & A269;
  assign \new_[30294]_  = ~A267 & \new_[30293]_ ;
  assign \new_[30298]_  = A302 & A300;
  assign \new_[30299]_  = A299 & \new_[30298]_ ;
  assign \new_[30300]_  = \new_[30299]_  & \new_[30294]_ ;
  assign \new_[30304]_  = ~A199 & ~A168;
  assign \new_[30305]_  = ~A170 & \new_[30304]_ ;
  assign \new_[30309]_  = A202 & A201;
  assign \new_[30310]_  = A200 & \new_[30309]_ ;
  assign \new_[30311]_  = \new_[30310]_  & \new_[30305]_ ;
  assign \new_[30315]_  = A298 & A266;
  assign \new_[30316]_  = A265 & \new_[30315]_ ;
  assign \new_[30320]_  = A301 & A300;
  assign \new_[30321]_  = ~A299 & \new_[30320]_ ;
  assign \new_[30322]_  = \new_[30321]_  & \new_[30316]_ ;
  assign \new_[30326]_  = ~A199 & ~A168;
  assign \new_[30327]_  = ~A170 & \new_[30326]_ ;
  assign \new_[30331]_  = A202 & A201;
  assign \new_[30332]_  = A200 & \new_[30331]_ ;
  assign \new_[30333]_  = \new_[30332]_  & \new_[30327]_ ;
  assign \new_[30337]_  = A298 & A266;
  assign \new_[30338]_  = A265 & \new_[30337]_ ;
  assign \new_[30342]_  = A302 & A300;
  assign \new_[30343]_  = ~A299 & \new_[30342]_ ;
  assign \new_[30344]_  = \new_[30343]_  & \new_[30338]_ ;
  assign \new_[30348]_  = ~A199 & ~A168;
  assign \new_[30349]_  = ~A170 & \new_[30348]_ ;
  assign \new_[30353]_  = A202 & A201;
  assign \new_[30354]_  = A200 & \new_[30353]_ ;
  assign \new_[30355]_  = \new_[30354]_  & \new_[30349]_ ;
  assign \new_[30359]_  = ~A298 & A266;
  assign \new_[30360]_  = A265 & \new_[30359]_ ;
  assign \new_[30364]_  = A301 & A300;
  assign \new_[30365]_  = A299 & \new_[30364]_ ;
  assign \new_[30366]_  = \new_[30365]_  & \new_[30360]_ ;
  assign \new_[30370]_  = ~A199 & ~A168;
  assign \new_[30371]_  = ~A170 & \new_[30370]_ ;
  assign \new_[30375]_  = A202 & A201;
  assign \new_[30376]_  = A200 & \new_[30375]_ ;
  assign \new_[30377]_  = \new_[30376]_  & \new_[30371]_ ;
  assign \new_[30381]_  = ~A298 & A266;
  assign \new_[30382]_  = A265 & \new_[30381]_ ;
  assign \new_[30386]_  = A302 & A300;
  assign \new_[30387]_  = A299 & \new_[30386]_ ;
  assign \new_[30388]_  = \new_[30387]_  & \new_[30382]_ ;
  assign \new_[30392]_  = ~A199 & ~A168;
  assign \new_[30393]_  = ~A170 & \new_[30392]_ ;
  assign \new_[30397]_  = A202 & A201;
  assign \new_[30398]_  = A200 & \new_[30397]_ ;
  assign \new_[30399]_  = \new_[30398]_  & \new_[30393]_ ;
  assign \new_[30403]_  = A298 & ~A266;
  assign \new_[30404]_  = ~A265 & \new_[30403]_ ;
  assign \new_[30408]_  = A301 & A300;
  assign \new_[30409]_  = ~A299 & \new_[30408]_ ;
  assign \new_[30410]_  = \new_[30409]_  & \new_[30404]_ ;
  assign \new_[30414]_  = ~A199 & ~A168;
  assign \new_[30415]_  = ~A170 & \new_[30414]_ ;
  assign \new_[30419]_  = A202 & A201;
  assign \new_[30420]_  = A200 & \new_[30419]_ ;
  assign \new_[30421]_  = \new_[30420]_  & \new_[30415]_ ;
  assign \new_[30425]_  = A298 & ~A266;
  assign \new_[30426]_  = ~A265 & \new_[30425]_ ;
  assign \new_[30430]_  = A302 & A300;
  assign \new_[30431]_  = ~A299 & \new_[30430]_ ;
  assign \new_[30432]_  = \new_[30431]_  & \new_[30426]_ ;
  assign \new_[30436]_  = ~A199 & ~A168;
  assign \new_[30437]_  = ~A170 & \new_[30436]_ ;
  assign \new_[30441]_  = A202 & A201;
  assign \new_[30442]_  = A200 & \new_[30441]_ ;
  assign \new_[30443]_  = \new_[30442]_  & \new_[30437]_ ;
  assign \new_[30447]_  = ~A298 & ~A266;
  assign \new_[30448]_  = ~A265 & \new_[30447]_ ;
  assign \new_[30452]_  = A301 & A300;
  assign \new_[30453]_  = A299 & \new_[30452]_ ;
  assign \new_[30454]_  = \new_[30453]_  & \new_[30448]_ ;
  assign \new_[30458]_  = ~A199 & ~A168;
  assign \new_[30459]_  = ~A170 & \new_[30458]_ ;
  assign \new_[30463]_  = A202 & A201;
  assign \new_[30464]_  = A200 & \new_[30463]_ ;
  assign \new_[30465]_  = \new_[30464]_  & \new_[30459]_ ;
  assign \new_[30469]_  = ~A298 & ~A266;
  assign \new_[30470]_  = ~A265 & \new_[30469]_ ;
  assign \new_[30474]_  = A302 & A300;
  assign \new_[30475]_  = A299 & \new_[30474]_ ;
  assign \new_[30476]_  = \new_[30475]_  & \new_[30470]_ ;
  assign \new_[30480]_  = ~A199 & ~A168;
  assign \new_[30481]_  = ~A170 & \new_[30480]_ ;
  assign \new_[30485]_  = A203 & A201;
  assign \new_[30486]_  = A200 & \new_[30485]_ ;
  assign \new_[30487]_  = \new_[30486]_  & \new_[30481]_ ;
  assign \new_[30491]_  = A298 & A268;
  assign \new_[30492]_  = ~A267 & \new_[30491]_ ;
  assign \new_[30496]_  = A301 & A300;
  assign \new_[30497]_  = ~A299 & \new_[30496]_ ;
  assign \new_[30498]_  = \new_[30497]_  & \new_[30492]_ ;
  assign \new_[30502]_  = ~A199 & ~A168;
  assign \new_[30503]_  = ~A170 & \new_[30502]_ ;
  assign \new_[30507]_  = A203 & A201;
  assign \new_[30508]_  = A200 & \new_[30507]_ ;
  assign \new_[30509]_  = \new_[30508]_  & \new_[30503]_ ;
  assign \new_[30513]_  = A298 & A268;
  assign \new_[30514]_  = ~A267 & \new_[30513]_ ;
  assign \new_[30518]_  = A302 & A300;
  assign \new_[30519]_  = ~A299 & \new_[30518]_ ;
  assign \new_[30520]_  = \new_[30519]_  & \new_[30514]_ ;
  assign \new_[30524]_  = ~A199 & ~A168;
  assign \new_[30525]_  = ~A170 & \new_[30524]_ ;
  assign \new_[30529]_  = A203 & A201;
  assign \new_[30530]_  = A200 & \new_[30529]_ ;
  assign \new_[30531]_  = \new_[30530]_  & \new_[30525]_ ;
  assign \new_[30535]_  = ~A298 & A268;
  assign \new_[30536]_  = ~A267 & \new_[30535]_ ;
  assign \new_[30540]_  = A301 & A300;
  assign \new_[30541]_  = A299 & \new_[30540]_ ;
  assign \new_[30542]_  = \new_[30541]_  & \new_[30536]_ ;
  assign \new_[30546]_  = ~A199 & ~A168;
  assign \new_[30547]_  = ~A170 & \new_[30546]_ ;
  assign \new_[30551]_  = A203 & A201;
  assign \new_[30552]_  = A200 & \new_[30551]_ ;
  assign \new_[30553]_  = \new_[30552]_  & \new_[30547]_ ;
  assign \new_[30557]_  = ~A298 & A268;
  assign \new_[30558]_  = ~A267 & \new_[30557]_ ;
  assign \new_[30562]_  = A302 & A300;
  assign \new_[30563]_  = A299 & \new_[30562]_ ;
  assign \new_[30564]_  = \new_[30563]_  & \new_[30558]_ ;
  assign \new_[30568]_  = ~A199 & ~A168;
  assign \new_[30569]_  = ~A170 & \new_[30568]_ ;
  assign \new_[30573]_  = A203 & A201;
  assign \new_[30574]_  = A200 & \new_[30573]_ ;
  assign \new_[30575]_  = \new_[30574]_  & \new_[30569]_ ;
  assign \new_[30579]_  = A298 & A269;
  assign \new_[30580]_  = ~A267 & \new_[30579]_ ;
  assign \new_[30584]_  = A301 & A300;
  assign \new_[30585]_  = ~A299 & \new_[30584]_ ;
  assign \new_[30586]_  = \new_[30585]_  & \new_[30580]_ ;
  assign \new_[30590]_  = ~A199 & ~A168;
  assign \new_[30591]_  = ~A170 & \new_[30590]_ ;
  assign \new_[30595]_  = A203 & A201;
  assign \new_[30596]_  = A200 & \new_[30595]_ ;
  assign \new_[30597]_  = \new_[30596]_  & \new_[30591]_ ;
  assign \new_[30601]_  = A298 & A269;
  assign \new_[30602]_  = ~A267 & \new_[30601]_ ;
  assign \new_[30606]_  = A302 & A300;
  assign \new_[30607]_  = ~A299 & \new_[30606]_ ;
  assign \new_[30608]_  = \new_[30607]_  & \new_[30602]_ ;
  assign \new_[30612]_  = ~A199 & ~A168;
  assign \new_[30613]_  = ~A170 & \new_[30612]_ ;
  assign \new_[30617]_  = A203 & A201;
  assign \new_[30618]_  = A200 & \new_[30617]_ ;
  assign \new_[30619]_  = \new_[30618]_  & \new_[30613]_ ;
  assign \new_[30623]_  = ~A298 & A269;
  assign \new_[30624]_  = ~A267 & \new_[30623]_ ;
  assign \new_[30628]_  = A301 & A300;
  assign \new_[30629]_  = A299 & \new_[30628]_ ;
  assign \new_[30630]_  = \new_[30629]_  & \new_[30624]_ ;
  assign \new_[30634]_  = ~A199 & ~A168;
  assign \new_[30635]_  = ~A170 & \new_[30634]_ ;
  assign \new_[30639]_  = A203 & A201;
  assign \new_[30640]_  = A200 & \new_[30639]_ ;
  assign \new_[30641]_  = \new_[30640]_  & \new_[30635]_ ;
  assign \new_[30645]_  = ~A298 & A269;
  assign \new_[30646]_  = ~A267 & \new_[30645]_ ;
  assign \new_[30650]_  = A302 & A300;
  assign \new_[30651]_  = A299 & \new_[30650]_ ;
  assign \new_[30652]_  = \new_[30651]_  & \new_[30646]_ ;
  assign \new_[30656]_  = ~A199 & ~A168;
  assign \new_[30657]_  = ~A170 & \new_[30656]_ ;
  assign \new_[30661]_  = A203 & A201;
  assign \new_[30662]_  = A200 & \new_[30661]_ ;
  assign \new_[30663]_  = \new_[30662]_  & \new_[30657]_ ;
  assign \new_[30667]_  = A298 & A266;
  assign \new_[30668]_  = A265 & \new_[30667]_ ;
  assign \new_[30672]_  = A301 & A300;
  assign \new_[30673]_  = ~A299 & \new_[30672]_ ;
  assign \new_[30674]_  = \new_[30673]_  & \new_[30668]_ ;
  assign \new_[30678]_  = ~A199 & ~A168;
  assign \new_[30679]_  = ~A170 & \new_[30678]_ ;
  assign \new_[30683]_  = A203 & A201;
  assign \new_[30684]_  = A200 & \new_[30683]_ ;
  assign \new_[30685]_  = \new_[30684]_  & \new_[30679]_ ;
  assign \new_[30689]_  = A298 & A266;
  assign \new_[30690]_  = A265 & \new_[30689]_ ;
  assign \new_[30694]_  = A302 & A300;
  assign \new_[30695]_  = ~A299 & \new_[30694]_ ;
  assign \new_[30696]_  = \new_[30695]_  & \new_[30690]_ ;
  assign \new_[30700]_  = ~A199 & ~A168;
  assign \new_[30701]_  = ~A170 & \new_[30700]_ ;
  assign \new_[30705]_  = A203 & A201;
  assign \new_[30706]_  = A200 & \new_[30705]_ ;
  assign \new_[30707]_  = \new_[30706]_  & \new_[30701]_ ;
  assign \new_[30711]_  = ~A298 & A266;
  assign \new_[30712]_  = A265 & \new_[30711]_ ;
  assign \new_[30716]_  = A301 & A300;
  assign \new_[30717]_  = A299 & \new_[30716]_ ;
  assign \new_[30718]_  = \new_[30717]_  & \new_[30712]_ ;
  assign \new_[30722]_  = ~A199 & ~A168;
  assign \new_[30723]_  = ~A170 & \new_[30722]_ ;
  assign \new_[30727]_  = A203 & A201;
  assign \new_[30728]_  = A200 & \new_[30727]_ ;
  assign \new_[30729]_  = \new_[30728]_  & \new_[30723]_ ;
  assign \new_[30733]_  = ~A298 & A266;
  assign \new_[30734]_  = A265 & \new_[30733]_ ;
  assign \new_[30738]_  = A302 & A300;
  assign \new_[30739]_  = A299 & \new_[30738]_ ;
  assign \new_[30740]_  = \new_[30739]_  & \new_[30734]_ ;
  assign \new_[30744]_  = ~A199 & ~A168;
  assign \new_[30745]_  = ~A170 & \new_[30744]_ ;
  assign \new_[30749]_  = A203 & A201;
  assign \new_[30750]_  = A200 & \new_[30749]_ ;
  assign \new_[30751]_  = \new_[30750]_  & \new_[30745]_ ;
  assign \new_[30755]_  = A298 & ~A266;
  assign \new_[30756]_  = ~A265 & \new_[30755]_ ;
  assign \new_[30760]_  = A301 & A300;
  assign \new_[30761]_  = ~A299 & \new_[30760]_ ;
  assign \new_[30762]_  = \new_[30761]_  & \new_[30756]_ ;
  assign \new_[30766]_  = ~A199 & ~A168;
  assign \new_[30767]_  = ~A170 & \new_[30766]_ ;
  assign \new_[30771]_  = A203 & A201;
  assign \new_[30772]_  = A200 & \new_[30771]_ ;
  assign \new_[30773]_  = \new_[30772]_  & \new_[30767]_ ;
  assign \new_[30777]_  = A298 & ~A266;
  assign \new_[30778]_  = ~A265 & \new_[30777]_ ;
  assign \new_[30782]_  = A302 & A300;
  assign \new_[30783]_  = ~A299 & \new_[30782]_ ;
  assign \new_[30784]_  = \new_[30783]_  & \new_[30778]_ ;
  assign \new_[30788]_  = ~A199 & ~A168;
  assign \new_[30789]_  = ~A170 & \new_[30788]_ ;
  assign \new_[30793]_  = A203 & A201;
  assign \new_[30794]_  = A200 & \new_[30793]_ ;
  assign \new_[30795]_  = \new_[30794]_  & \new_[30789]_ ;
  assign \new_[30799]_  = ~A298 & ~A266;
  assign \new_[30800]_  = ~A265 & \new_[30799]_ ;
  assign \new_[30804]_  = A301 & A300;
  assign \new_[30805]_  = A299 & \new_[30804]_ ;
  assign \new_[30806]_  = \new_[30805]_  & \new_[30800]_ ;
  assign \new_[30810]_  = ~A199 & ~A168;
  assign \new_[30811]_  = ~A170 & \new_[30810]_ ;
  assign \new_[30815]_  = A203 & A201;
  assign \new_[30816]_  = A200 & \new_[30815]_ ;
  assign \new_[30817]_  = \new_[30816]_  & \new_[30811]_ ;
  assign \new_[30821]_  = ~A298 & ~A266;
  assign \new_[30822]_  = ~A265 & \new_[30821]_ ;
  assign \new_[30826]_  = A302 & A300;
  assign \new_[30827]_  = A299 & \new_[30826]_ ;
  assign \new_[30828]_  = \new_[30827]_  & \new_[30822]_ ;
  assign \new_[30832]_  = A199 & ~A168;
  assign \new_[30833]_  = ~A170 & \new_[30832]_ ;
  assign \new_[30837]_  = A202 & A201;
  assign \new_[30838]_  = ~A200 & \new_[30837]_ ;
  assign \new_[30839]_  = \new_[30838]_  & \new_[30833]_ ;
  assign \new_[30843]_  = A298 & A268;
  assign \new_[30844]_  = ~A267 & \new_[30843]_ ;
  assign \new_[30848]_  = A301 & A300;
  assign \new_[30849]_  = ~A299 & \new_[30848]_ ;
  assign \new_[30850]_  = \new_[30849]_  & \new_[30844]_ ;
  assign \new_[30854]_  = A199 & ~A168;
  assign \new_[30855]_  = ~A170 & \new_[30854]_ ;
  assign \new_[30859]_  = A202 & A201;
  assign \new_[30860]_  = ~A200 & \new_[30859]_ ;
  assign \new_[30861]_  = \new_[30860]_  & \new_[30855]_ ;
  assign \new_[30865]_  = A298 & A268;
  assign \new_[30866]_  = ~A267 & \new_[30865]_ ;
  assign \new_[30870]_  = A302 & A300;
  assign \new_[30871]_  = ~A299 & \new_[30870]_ ;
  assign \new_[30872]_  = \new_[30871]_  & \new_[30866]_ ;
  assign \new_[30876]_  = A199 & ~A168;
  assign \new_[30877]_  = ~A170 & \new_[30876]_ ;
  assign \new_[30881]_  = A202 & A201;
  assign \new_[30882]_  = ~A200 & \new_[30881]_ ;
  assign \new_[30883]_  = \new_[30882]_  & \new_[30877]_ ;
  assign \new_[30887]_  = ~A298 & A268;
  assign \new_[30888]_  = ~A267 & \new_[30887]_ ;
  assign \new_[30892]_  = A301 & A300;
  assign \new_[30893]_  = A299 & \new_[30892]_ ;
  assign \new_[30894]_  = \new_[30893]_  & \new_[30888]_ ;
  assign \new_[30898]_  = A199 & ~A168;
  assign \new_[30899]_  = ~A170 & \new_[30898]_ ;
  assign \new_[30903]_  = A202 & A201;
  assign \new_[30904]_  = ~A200 & \new_[30903]_ ;
  assign \new_[30905]_  = \new_[30904]_  & \new_[30899]_ ;
  assign \new_[30909]_  = ~A298 & A268;
  assign \new_[30910]_  = ~A267 & \new_[30909]_ ;
  assign \new_[30914]_  = A302 & A300;
  assign \new_[30915]_  = A299 & \new_[30914]_ ;
  assign \new_[30916]_  = \new_[30915]_  & \new_[30910]_ ;
  assign \new_[30920]_  = A199 & ~A168;
  assign \new_[30921]_  = ~A170 & \new_[30920]_ ;
  assign \new_[30925]_  = A202 & A201;
  assign \new_[30926]_  = ~A200 & \new_[30925]_ ;
  assign \new_[30927]_  = \new_[30926]_  & \new_[30921]_ ;
  assign \new_[30931]_  = A298 & A269;
  assign \new_[30932]_  = ~A267 & \new_[30931]_ ;
  assign \new_[30936]_  = A301 & A300;
  assign \new_[30937]_  = ~A299 & \new_[30936]_ ;
  assign \new_[30938]_  = \new_[30937]_  & \new_[30932]_ ;
  assign \new_[30942]_  = A199 & ~A168;
  assign \new_[30943]_  = ~A170 & \new_[30942]_ ;
  assign \new_[30947]_  = A202 & A201;
  assign \new_[30948]_  = ~A200 & \new_[30947]_ ;
  assign \new_[30949]_  = \new_[30948]_  & \new_[30943]_ ;
  assign \new_[30953]_  = A298 & A269;
  assign \new_[30954]_  = ~A267 & \new_[30953]_ ;
  assign \new_[30958]_  = A302 & A300;
  assign \new_[30959]_  = ~A299 & \new_[30958]_ ;
  assign \new_[30960]_  = \new_[30959]_  & \new_[30954]_ ;
  assign \new_[30964]_  = A199 & ~A168;
  assign \new_[30965]_  = ~A170 & \new_[30964]_ ;
  assign \new_[30969]_  = A202 & A201;
  assign \new_[30970]_  = ~A200 & \new_[30969]_ ;
  assign \new_[30971]_  = \new_[30970]_  & \new_[30965]_ ;
  assign \new_[30975]_  = ~A298 & A269;
  assign \new_[30976]_  = ~A267 & \new_[30975]_ ;
  assign \new_[30980]_  = A301 & A300;
  assign \new_[30981]_  = A299 & \new_[30980]_ ;
  assign \new_[30982]_  = \new_[30981]_  & \new_[30976]_ ;
  assign \new_[30986]_  = A199 & ~A168;
  assign \new_[30987]_  = ~A170 & \new_[30986]_ ;
  assign \new_[30991]_  = A202 & A201;
  assign \new_[30992]_  = ~A200 & \new_[30991]_ ;
  assign \new_[30993]_  = \new_[30992]_  & \new_[30987]_ ;
  assign \new_[30997]_  = ~A298 & A269;
  assign \new_[30998]_  = ~A267 & \new_[30997]_ ;
  assign \new_[31002]_  = A302 & A300;
  assign \new_[31003]_  = A299 & \new_[31002]_ ;
  assign \new_[31004]_  = \new_[31003]_  & \new_[30998]_ ;
  assign \new_[31008]_  = A199 & ~A168;
  assign \new_[31009]_  = ~A170 & \new_[31008]_ ;
  assign \new_[31013]_  = A202 & A201;
  assign \new_[31014]_  = ~A200 & \new_[31013]_ ;
  assign \new_[31015]_  = \new_[31014]_  & \new_[31009]_ ;
  assign \new_[31019]_  = A298 & A266;
  assign \new_[31020]_  = A265 & \new_[31019]_ ;
  assign \new_[31024]_  = A301 & A300;
  assign \new_[31025]_  = ~A299 & \new_[31024]_ ;
  assign \new_[31026]_  = \new_[31025]_  & \new_[31020]_ ;
  assign \new_[31030]_  = A199 & ~A168;
  assign \new_[31031]_  = ~A170 & \new_[31030]_ ;
  assign \new_[31035]_  = A202 & A201;
  assign \new_[31036]_  = ~A200 & \new_[31035]_ ;
  assign \new_[31037]_  = \new_[31036]_  & \new_[31031]_ ;
  assign \new_[31041]_  = A298 & A266;
  assign \new_[31042]_  = A265 & \new_[31041]_ ;
  assign \new_[31046]_  = A302 & A300;
  assign \new_[31047]_  = ~A299 & \new_[31046]_ ;
  assign \new_[31048]_  = \new_[31047]_  & \new_[31042]_ ;
  assign \new_[31052]_  = A199 & ~A168;
  assign \new_[31053]_  = ~A170 & \new_[31052]_ ;
  assign \new_[31057]_  = A202 & A201;
  assign \new_[31058]_  = ~A200 & \new_[31057]_ ;
  assign \new_[31059]_  = \new_[31058]_  & \new_[31053]_ ;
  assign \new_[31063]_  = ~A298 & A266;
  assign \new_[31064]_  = A265 & \new_[31063]_ ;
  assign \new_[31068]_  = A301 & A300;
  assign \new_[31069]_  = A299 & \new_[31068]_ ;
  assign \new_[31070]_  = \new_[31069]_  & \new_[31064]_ ;
  assign \new_[31074]_  = A199 & ~A168;
  assign \new_[31075]_  = ~A170 & \new_[31074]_ ;
  assign \new_[31079]_  = A202 & A201;
  assign \new_[31080]_  = ~A200 & \new_[31079]_ ;
  assign \new_[31081]_  = \new_[31080]_  & \new_[31075]_ ;
  assign \new_[31085]_  = ~A298 & A266;
  assign \new_[31086]_  = A265 & \new_[31085]_ ;
  assign \new_[31090]_  = A302 & A300;
  assign \new_[31091]_  = A299 & \new_[31090]_ ;
  assign \new_[31092]_  = \new_[31091]_  & \new_[31086]_ ;
  assign \new_[31096]_  = A199 & ~A168;
  assign \new_[31097]_  = ~A170 & \new_[31096]_ ;
  assign \new_[31101]_  = A202 & A201;
  assign \new_[31102]_  = ~A200 & \new_[31101]_ ;
  assign \new_[31103]_  = \new_[31102]_  & \new_[31097]_ ;
  assign \new_[31107]_  = A298 & ~A266;
  assign \new_[31108]_  = ~A265 & \new_[31107]_ ;
  assign \new_[31112]_  = A301 & A300;
  assign \new_[31113]_  = ~A299 & \new_[31112]_ ;
  assign \new_[31114]_  = \new_[31113]_  & \new_[31108]_ ;
  assign \new_[31118]_  = A199 & ~A168;
  assign \new_[31119]_  = ~A170 & \new_[31118]_ ;
  assign \new_[31123]_  = A202 & A201;
  assign \new_[31124]_  = ~A200 & \new_[31123]_ ;
  assign \new_[31125]_  = \new_[31124]_  & \new_[31119]_ ;
  assign \new_[31129]_  = A298 & ~A266;
  assign \new_[31130]_  = ~A265 & \new_[31129]_ ;
  assign \new_[31134]_  = A302 & A300;
  assign \new_[31135]_  = ~A299 & \new_[31134]_ ;
  assign \new_[31136]_  = \new_[31135]_  & \new_[31130]_ ;
  assign \new_[31140]_  = A199 & ~A168;
  assign \new_[31141]_  = ~A170 & \new_[31140]_ ;
  assign \new_[31145]_  = A202 & A201;
  assign \new_[31146]_  = ~A200 & \new_[31145]_ ;
  assign \new_[31147]_  = \new_[31146]_  & \new_[31141]_ ;
  assign \new_[31151]_  = ~A298 & ~A266;
  assign \new_[31152]_  = ~A265 & \new_[31151]_ ;
  assign \new_[31156]_  = A301 & A300;
  assign \new_[31157]_  = A299 & \new_[31156]_ ;
  assign \new_[31158]_  = \new_[31157]_  & \new_[31152]_ ;
  assign \new_[31162]_  = A199 & ~A168;
  assign \new_[31163]_  = ~A170 & \new_[31162]_ ;
  assign \new_[31167]_  = A202 & A201;
  assign \new_[31168]_  = ~A200 & \new_[31167]_ ;
  assign \new_[31169]_  = \new_[31168]_  & \new_[31163]_ ;
  assign \new_[31173]_  = ~A298 & ~A266;
  assign \new_[31174]_  = ~A265 & \new_[31173]_ ;
  assign \new_[31178]_  = A302 & A300;
  assign \new_[31179]_  = A299 & \new_[31178]_ ;
  assign \new_[31180]_  = \new_[31179]_  & \new_[31174]_ ;
  assign \new_[31184]_  = A199 & ~A168;
  assign \new_[31185]_  = ~A170 & \new_[31184]_ ;
  assign \new_[31189]_  = A203 & A201;
  assign \new_[31190]_  = ~A200 & \new_[31189]_ ;
  assign \new_[31191]_  = \new_[31190]_  & \new_[31185]_ ;
  assign \new_[31195]_  = A298 & A268;
  assign \new_[31196]_  = ~A267 & \new_[31195]_ ;
  assign \new_[31200]_  = A301 & A300;
  assign \new_[31201]_  = ~A299 & \new_[31200]_ ;
  assign \new_[31202]_  = \new_[31201]_  & \new_[31196]_ ;
  assign \new_[31206]_  = A199 & ~A168;
  assign \new_[31207]_  = ~A170 & \new_[31206]_ ;
  assign \new_[31211]_  = A203 & A201;
  assign \new_[31212]_  = ~A200 & \new_[31211]_ ;
  assign \new_[31213]_  = \new_[31212]_  & \new_[31207]_ ;
  assign \new_[31217]_  = A298 & A268;
  assign \new_[31218]_  = ~A267 & \new_[31217]_ ;
  assign \new_[31222]_  = A302 & A300;
  assign \new_[31223]_  = ~A299 & \new_[31222]_ ;
  assign \new_[31224]_  = \new_[31223]_  & \new_[31218]_ ;
  assign \new_[31228]_  = A199 & ~A168;
  assign \new_[31229]_  = ~A170 & \new_[31228]_ ;
  assign \new_[31233]_  = A203 & A201;
  assign \new_[31234]_  = ~A200 & \new_[31233]_ ;
  assign \new_[31235]_  = \new_[31234]_  & \new_[31229]_ ;
  assign \new_[31239]_  = ~A298 & A268;
  assign \new_[31240]_  = ~A267 & \new_[31239]_ ;
  assign \new_[31244]_  = A301 & A300;
  assign \new_[31245]_  = A299 & \new_[31244]_ ;
  assign \new_[31246]_  = \new_[31245]_  & \new_[31240]_ ;
  assign \new_[31250]_  = A199 & ~A168;
  assign \new_[31251]_  = ~A170 & \new_[31250]_ ;
  assign \new_[31255]_  = A203 & A201;
  assign \new_[31256]_  = ~A200 & \new_[31255]_ ;
  assign \new_[31257]_  = \new_[31256]_  & \new_[31251]_ ;
  assign \new_[31261]_  = ~A298 & A268;
  assign \new_[31262]_  = ~A267 & \new_[31261]_ ;
  assign \new_[31266]_  = A302 & A300;
  assign \new_[31267]_  = A299 & \new_[31266]_ ;
  assign \new_[31268]_  = \new_[31267]_  & \new_[31262]_ ;
  assign \new_[31272]_  = A199 & ~A168;
  assign \new_[31273]_  = ~A170 & \new_[31272]_ ;
  assign \new_[31277]_  = A203 & A201;
  assign \new_[31278]_  = ~A200 & \new_[31277]_ ;
  assign \new_[31279]_  = \new_[31278]_  & \new_[31273]_ ;
  assign \new_[31283]_  = A298 & A269;
  assign \new_[31284]_  = ~A267 & \new_[31283]_ ;
  assign \new_[31288]_  = A301 & A300;
  assign \new_[31289]_  = ~A299 & \new_[31288]_ ;
  assign \new_[31290]_  = \new_[31289]_  & \new_[31284]_ ;
  assign \new_[31294]_  = A199 & ~A168;
  assign \new_[31295]_  = ~A170 & \new_[31294]_ ;
  assign \new_[31299]_  = A203 & A201;
  assign \new_[31300]_  = ~A200 & \new_[31299]_ ;
  assign \new_[31301]_  = \new_[31300]_  & \new_[31295]_ ;
  assign \new_[31305]_  = A298 & A269;
  assign \new_[31306]_  = ~A267 & \new_[31305]_ ;
  assign \new_[31310]_  = A302 & A300;
  assign \new_[31311]_  = ~A299 & \new_[31310]_ ;
  assign \new_[31312]_  = \new_[31311]_  & \new_[31306]_ ;
  assign \new_[31316]_  = A199 & ~A168;
  assign \new_[31317]_  = ~A170 & \new_[31316]_ ;
  assign \new_[31321]_  = A203 & A201;
  assign \new_[31322]_  = ~A200 & \new_[31321]_ ;
  assign \new_[31323]_  = \new_[31322]_  & \new_[31317]_ ;
  assign \new_[31327]_  = ~A298 & A269;
  assign \new_[31328]_  = ~A267 & \new_[31327]_ ;
  assign \new_[31332]_  = A301 & A300;
  assign \new_[31333]_  = A299 & \new_[31332]_ ;
  assign \new_[31334]_  = \new_[31333]_  & \new_[31328]_ ;
  assign \new_[31338]_  = A199 & ~A168;
  assign \new_[31339]_  = ~A170 & \new_[31338]_ ;
  assign \new_[31343]_  = A203 & A201;
  assign \new_[31344]_  = ~A200 & \new_[31343]_ ;
  assign \new_[31345]_  = \new_[31344]_  & \new_[31339]_ ;
  assign \new_[31349]_  = ~A298 & A269;
  assign \new_[31350]_  = ~A267 & \new_[31349]_ ;
  assign \new_[31354]_  = A302 & A300;
  assign \new_[31355]_  = A299 & \new_[31354]_ ;
  assign \new_[31356]_  = \new_[31355]_  & \new_[31350]_ ;
  assign \new_[31360]_  = A199 & ~A168;
  assign \new_[31361]_  = ~A170 & \new_[31360]_ ;
  assign \new_[31365]_  = A203 & A201;
  assign \new_[31366]_  = ~A200 & \new_[31365]_ ;
  assign \new_[31367]_  = \new_[31366]_  & \new_[31361]_ ;
  assign \new_[31371]_  = A298 & A266;
  assign \new_[31372]_  = A265 & \new_[31371]_ ;
  assign \new_[31376]_  = A301 & A300;
  assign \new_[31377]_  = ~A299 & \new_[31376]_ ;
  assign \new_[31378]_  = \new_[31377]_  & \new_[31372]_ ;
  assign \new_[31382]_  = A199 & ~A168;
  assign \new_[31383]_  = ~A170 & \new_[31382]_ ;
  assign \new_[31387]_  = A203 & A201;
  assign \new_[31388]_  = ~A200 & \new_[31387]_ ;
  assign \new_[31389]_  = \new_[31388]_  & \new_[31383]_ ;
  assign \new_[31393]_  = A298 & A266;
  assign \new_[31394]_  = A265 & \new_[31393]_ ;
  assign \new_[31398]_  = A302 & A300;
  assign \new_[31399]_  = ~A299 & \new_[31398]_ ;
  assign \new_[31400]_  = \new_[31399]_  & \new_[31394]_ ;
  assign \new_[31404]_  = A199 & ~A168;
  assign \new_[31405]_  = ~A170 & \new_[31404]_ ;
  assign \new_[31409]_  = A203 & A201;
  assign \new_[31410]_  = ~A200 & \new_[31409]_ ;
  assign \new_[31411]_  = \new_[31410]_  & \new_[31405]_ ;
  assign \new_[31415]_  = ~A298 & A266;
  assign \new_[31416]_  = A265 & \new_[31415]_ ;
  assign \new_[31420]_  = A301 & A300;
  assign \new_[31421]_  = A299 & \new_[31420]_ ;
  assign \new_[31422]_  = \new_[31421]_  & \new_[31416]_ ;
  assign \new_[31426]_  = A199 & ~A168;
  assign \new_[31427]_  = ~A170 & \new_[31426]_ ;
  assign \new_[31431]_  = A203 & A201;
  assign \new_[31432]_  = ~A200 & \new_[31431]_ ;
  assign \new_[31433]_  = \new_[31432]_  & \new_[31427]_ ;
  assign \new_[31437]_  = ~A298 & A266;
  assign \new_[31438]_  = A265 & \new_[31437]_ ;
  assign \new_[31442]_  = A302 & A300;
  assign \new_[31443]_  = A299 & \new_[31442]_ ;
  assign \new_[31444]_  = \new_[31443]_  & \new_[31438]_ ;
  assign \new_[31448]_  = A199 & ~A168;
  assign \new_[31449]_  = ~A170 & \new_[31448]_ ;
  assign \new_[31453]_  = A203 & A201;
  assign \new_[31454]_  = ~A200 & \new_[31453]_ ;
  assign \new_[31455]_  = \new_[31454]_  & \new_[31449]_ ;
  assign \new_[31459]_  = A298 & ~A266;
  assign \new_[31460]_  = ~A265 & \new_[31459]_ ;
  assign \new_[31464]_  = A301 & A300;
  assign \new_[31465]_  = ~A299 & \new_[31464]_ ;
  assign \new_[31466]_  = \new_[31465]_  & \new_[31460]_ ;
  assign \new_[31470]_  = A199 & ~A168;
  assign \new_[31471]_  = ~A170 & \new_[31470]_ ;
  assign \new_[31475]_  = A203 & A201;
  assign \new_[31476]_  = ~A200 & \new_[31475]_ ;
  assign \new_[31477]_  = \new_[31476]_  & \new_[31471]_ ;
  assign \new_[31481]_  = A298 & ~A266;
  assign \new_[31482]_  = ~A265 & \new_[31481]_ ;
  assign \new_[31486]_  = A302 & A300;
  assign \new_[31487]_  = ~A299 & \new_[31486]_ ;
  assign \new_[31488]_  = \new_[31487]_  & \new_[31482]_ ;
  assign \new_[31492]_  = A199 & ~A168;
  assign \new_[31493]_  = ~A170 & \new_[31492]_ ;
  assign \new_[31497]_  = A203 & A201;
  assign \new_[31498]_  = ~A200 & \new_[31497]_ ;
  assign \new_[31499]_  = \new_[31498]_  & \new_[31493]_ ;
  assign \new_[31503]_  = ~A298 & ~A266;
  assign \new_[31504]_  = ~A265 & \new_[31503]_ ;
  assign \new_[31508]_  = A301 & A300;
  assign \new_[31509]_  = A299 & \new_[31508]_ ;
  assign \new_[31510]_  = \new_[31509]_  & \new_[31504]_ ;
  assign \new_[31514]_  = A199 & ~A168;
  assign \new_[31515]_  = ~A170 & \new_[31514]_ ;
  assign \new_[31519]_  = A203 & A201;
  assign \new_[31520]_  = ~A200 & \new_[31519]_ ;
  assign \new_[31521]_  = \new_[31520]_  & \new_[31515]_ ;
  assign \new_[31525]_  = ~A298 & ~A266;
  assign \new_[31526]_  = ~A265 & \new_[31525]_ ;
  assign \new_[31530]_  = A302 & A300;
  assign \new_[31531]_  = A299 & \new_[31530]_ ;
  assign \new_[31532]_  = \new_[31531]_  & \new_[31526]_ ;
  assign \new_[31536]_  = ~A199 & ~A168;
  assign \new_[31537]_  = ~A170 & \new_[31536]_ ;
  assign \new_[31541]_  = A266 & ~A265;
  assign \new_[31542]_  = ~A200 & \new_[31541]_ ;
  assign \new_[31543]_  = \new_[31542]_  & \new_[31537]_ ;
  assign \new_[31547]_  = ~A269 & ~A268;
  assign \new_[31548]_  = ~A267 & \new_[31547]_ ;
  assign \new_[31552]_  = ~A302 & ~A301;
  assign \new_[31553]_  = A300 & \new_[31552]_ ;
  assign \new_[31554]_  = \new_[31553]_  & \new_[31548]_ ;
  assign \new_[31558]_  = ~A199 & ~A168;
  assign \new_[31559]_  = ~A170 & \new_[31558]_ ;
  assign \new_[31563]_  = ~A266 & A265;
  assign \new_[31564]_  = ~A200 & \new_[31563]_ ;
  assign \new_[31565]_  = \new_[31564]_  & \new_[31559]_ ;
  assign \new_[31569]_  = ~A269 & ~A268;
  assign \new_[31570]_  = ~A267 & \new_[31569]_ ;
  assign \new_[31574]_  = ~A302 & ~A301;
  assign \new_[31575]_  = A300 & \new_[31574]_ ;
  assign \new_[31576]_  = \new_[31575]_  & \new_[31570]_ ;
  assign \new_[31580]_  = A167 & A168;
  assign \new_[31581]_  = A169 & \new_[31580]_ ;
  assign \new_[31585]_  = A202 & ~A201;
  assign \new_[31586]_  = ~A166 & \new_[31585]_ ;
  assign \new_[31587]_  = \new_[31586]_  & \new_[31581]_ ;
  assign \new_[31591]_  = A298 & A268;
  assign \new_[31592]_  = ~A267 & \new_[31591]_ ;
  assign \new_[31596]_  = A301 & A300;
  assign \new_[31597]_  = ~A299 & \new_[31596]_ ;
  assign \new_[31598]_  = \new_[31597]_  & \new_[31592]_ ;
  assign \new_[31602]_  = A167 & A168;
  assign \new_[31603]_  = A169 & \new_[31602]_ ;
  assign \new_[31607]_  = A202 & ~A201;
  assign \new_[31608]_  = ~A166 & \new_[31607]_ ;
  assign \new_[31609]_  = \new_[31608]_  & \new_[31603]_ ;
  assign \new_[31613]_  = A298 & A268;
  assign \new_[31614]_  = ~A267 & \new_[31613]_ ;
  assign \new_[31618]_  = A302 & A300;
  assign \new_[31619]_  = ~A299 & \new_[31618]_ ;
  assign \new_[31620]_  = \new_[31619]_  & \new_[31614]_ ;
  assign \new_[31624]_  = A167 & A168;
  assign \new_[31625]_  = A169 & \new_[31624]_ ;
  assign \new_[31629]_  = A202 & ~A201;
  assign \new_[31630]_  = ~A166 & \new_[31629]_ ;
  assign \new_[31631]_  = \new_[31630]_  & \new_[31625]_ ;
  assign \new_[31635]_  = ~A298 & A268;
  assign \new_[31636]_  = ~A267 & \new_[31635]_ ;
  assign \new_[31640]_  = A301 & A300;
  assign \new_[31641]_  = A299 & \new_[31640]_ ;
  assign \new_[31642]_  = \new_[31641]_  & \new_[31636]_ ;
  assign \new_[31646]_  = A167 & A168;
  assign \new_[31647]_  = A169 & \new_[31646]_ ;
  assign \new_[31651]_  = A202 & ~A201;
  assign \new_[31652]_  = ~A166 & \new_[31651]_ ;
  assign \new_[31653]_  = \new_[31652]_  & \new_[31647]_ ;
  assign \new_[31657]_  = ~A298 & A268;
  assign \new_[31658]_  = ~A267 & \new_[31657]_ ;
  assign \new_[31662]_  = A302 & A300;
  assign \new_[31663]_  = A299 & \new_[31662]_ ;
  assign \new_[31664]_  = \new_[31663]_  & \new_[31658]_ ;
  assign \new_[31668]_  = A167 & A168;
  assign \new_[31669]_  = A169 & \new_[31668]_ ;
  assign \new_[31673]_  = A202 & ~A201;
  assign \new_[31674]_  = ~A166 & \new_[31673]_ ;
  assign \new_[31675]_  = \new_[31674]_  & \new_[31669]_ ;
  assign \new_[31679]_  = A298 & A269;
  assign \new_[31680]_  = ~A267 & \new_[31679]_ ;
  assign \new_[31684]_  = A301 & A300;
  assign \new_[31685]_  = ~A299 & \new_[31684]_ ;
  assign \new_[31686]_  = \new_[31685]_  & \new_[31680]_ ;
  assign \new_[31690]_  = A167 & A168;
  assign \new_[31691]_  = A169 & \new_[31690]_ ;
  assign \new_[31695]_  = A202 & ~A201;
  assign \new_[31696]_  = ~A166 & \new_[31695]_ ;
  assign \new_[31697]_  = \new_[31696]_  & \new_[31691]_ ;
  assign \new_[31701]_  = A298 & A269;
  assign \new_[31702]_  = ~A267 & \new_[31701]_ ;
  assign \new_[31706]_  = A302 & A300;
  assign \new_[31707]_  = ~A299 & \new_[31706]_ ;
  assign \new_[31708]_  = \new_[31707]_  & \new_[31702]_ ;
  assign \new_[31712]_  = A167 & A168;
  assign \new_[31713]_  = A169 & \new_[31712]_ ;
  assign \new_[31717]_  = A202 & ~A201;
  assign \new_[31718]_  = ~A166 & \new_[31717]_ ;
  assign \new_[31719]_  = \new_[31718]_  & \new_[31713]_ ;
  assign \new_[31723]_  = ~A298 & A269;
  assign \new_[31724]_  = ~A267 & \new_[31723]_ ;
  assign \new_[31728]_  = A301 & A300;
  assign \new_[31729]_  = A299 & \new_[31728]_ ;
  assign \new_[31730]_  = \new_[31729]_  & \new_[31724]_ ;
  assign \new_[31734]_  = A167 & A168;
  assign \new_[31735]_  = A169 & \new_[31734]_ ;
  assign \new_[31739]_  = A202 & ~A201;
  assign \new_[31740]_  = ~A166 & \new_[31739]_ ;
  assign \new_[31741]_  = \new_[31740]_  & \new_[31735]_ ;
  assign \new_[31745]_  = ~A298 & A269;
  assign \new_[31746]_  = ~A267 & \new_[31745]_ ;
  assign \new_[31750]_  = A302 & A300;
  assign \new_[31751]_  = A299 & \new_[31750]_ ;
  assign \new_[31752]_  = \new_[31751]_  & \new_[31746]_ ;
  assign \new_[31756]_  = A167 & A168;
  assign \new_[31757]_  = A169 & \new_[31756]_ ;
  assign \new_[31761]_  = A202 & ~A201;
  assign \new_[31762]_  = ~A166 & \new_[31761]_ ;
  assign \new_[31763]_  = \new_[31762]_  & \new_[31757]_ ;
  assign \new_[31767]_  = A298 & A266;
  assign \new_[31768]_  = A265 & \new_[31767]_ ;
  assign \new_[31772]_  = A301 & A300;
  assign \new_[31773]_  = ~A299 & \new_[31772]_ ;
  assign \new_[31774]_  = \new_[31773]_  & \new_[31768]_ ;
  assign \new_[31778]_  = A167 & A168;
  assign \new_[31779]_  = A169 & \new_[31778]_ ;
  assign \new_[31783]_  = A202 & ~A201;
  assign \new_[31784]_  = ~A166 & \new_[31783]_ ;
  assign \new_[31785]_  = \new_[31784]_  & \new_[31779]_ ;
  assign \new_[31789]_  = A298 & A266;
  assign \new_[31790]_  = A265 & \new_[31789]_ ;
  assign \new_[31794]_  = A302 & A300;
  assign \new_[31795]_  = ~A299 & \new_[31794]_ ;
  assign \new_[31796]_  = \new_[31795]_  & \new_[31790]_ ;
  assign \new_[31800]_  = A167 & A168;
  assign \new_[31801]_  = A169 & \new_[31800]_ ;
  assign \new_[31805]_  = A202 & ~A201;
  assign \new_[31806]_  = ~A166 & \new_[31805]_ ;
  assign \new_[31807]_  = \new_[31806]_  & \new_[31801]_ ;
  assign \new_[31811]_  = ~A298 & A266;
  assign \new_[31812]_  = A265 & \new_[31811]_ ;
  assign \new_[31816]_  = A301 & A300;
  assign \new_[31817]_  = A299 & \new_[31816]_ ;
  assign \new_[31818]_  = \new_[31817]_  & \new_[31812]_ ;
  assign \new_[31822]_  = A167 & A168;
  assign \new_[31823]_  = A169 & \new_[31822]_ ;
  assign \new_[31827]_  = A202 & ~A201;
  assign \new_[31828]_  = ~A166 & \new_[31827]_ ;
  assign \new_[31829]_  = \new_[31828]_  & \new_[31823]_ ;
  assign \new_[31833]_  = ~A298 & A266;
  assign \new_[31834]_  = A265 & \new_[31833]_ ;
  assign \new_[31838]_  = A302 & A300;
  assign \new_[31839]_  = A299 & \new_[31838]_ ;
  assign \new_[31840]_  = \new_[31839]_  & \new_[31834]_ ;
  assign \new_[31844]_  = A167 & A168;
  assign \new_[31845]_  = A169 & \new_[31844]_ ;
  assign \new_[31849]_  = A202 & ~A201;
  assign \new_[31850]_  = ~A166 & \new_[31849]_ ;
  assign \new_[31851]_  = \new_[31850]_  & \new_[31845]_ ;
  assign \new_[31855]_  = A298 & ~A266;
  assign \new_[31856]_  = ~A265 & \new_[31855]_ ;
  assign \new_[31860]_  = A301 & A300;
  assign \new_[31861]_  = ~A299 & \new_[31860]_ ;
  assign \new_[31862]_  = \new_[31861]_  & \new_[31856]_ ;
  assign \new_[31866]_  = A167 & A168;
  assign \new_[31867]_  = A169 & \new_[31866]_ ;
  assign \new_[31871]_  = A202 & ~A201;
  assign \new_[31872]_  = ~A166 & \new_[31871]_ ;
  assign \new_[31873]_  = \new_[31872]_  & \new_[31867]_ ;
  assign \new_[31877]_  = A298 & ~A266;
  assign \new_[31878]_  = ~A265 & \new_[31877]_ ;
  assign \new_[31882]_  = A302 & A300;
  assign \new_[31883]_  = ~A299 & \new_[31882]_ ;
  assign \new_[31884]_  = \new_[31883]_  & \new_[31878]_ ;
  assign \new_[31888]_  = A167 & A168;
  assign \new_[31889]_  = A169 & \new_[31888]_ ;
  assign \new_[31893]_  = A202 & ~A201;
  assign \new_[31894]_  = ~A166 & \new_[31893]_ ;
  assign \new_[31895]_  = \new_[31894]_  & \new_[31889]_ ;
  assign \new_[31899]_  = ~A298 & ~A266;
  assign \new_[31900]_  = ~A265 & \new_[31899]_ ;
  assign \new_[31904]_  = A301 & A300;
  assign \new_[31905]_  = A299 & \new_[31904]_ ;
  assign \new_[31906]_  = \new_[31905]_  & \new_[31900]_ ;
  assign \new_[31910]_  = A167 & A168;
  assign \new_[31911]_  = A169 & \new_[31910]_ ;
  assign \new_[31915]_  = A202 & ~A201;
  assign \new_[31916]_  = ~A166 & \new_[31915]_ ;
  assign \new_[31917]_  = \new_[31916]_  & \new_[31911]_ ;
  assign \new_[31921]_  = ~A298 & ~A266;
  assign \new_[31922]_  = ~A265 & \new_[31921]_ ;
  assign \new_[31926]_  = A302 & A300;
  assign \new_[31927]_  = A299 & \new_[31926]_ ;
  assign \new_[31928]_  = \new_[31927]_  & \new_[31922]_ ;
  assign \new_[31932]_  = A167 & A168;
  assign \new_[31933]_  = A169 & \new_[31932]_ ;
  assign \new_[31937]_  = A203 & ~A201;
  assign \new_[31938]_  = ~A166 & \new_[31937]_ ;
  assign \new_[31939]_  = \new_[31938]_  & \new_[31933]_ ;
  assign \new_[31943]_  = A298 & A268;
  assign \new_[31944]_  = ~A267 & \new_[31943]_ ;
  assign \new_[31948]_  = A301 & A300;
  assign \new_[31949]_  = ~A299 & \new_[31948]_ ;
  assign \new_[31950]_  = \new_[31949]_  & \new_[31944]_ ;
  assign \new_[31954]_  = A167 & A168;
  assign \new_[31955]_  = A169 & \new_[31954]_ ;
  assign \new_[31959]_  = A203 & ~A201;
  assign \new_[31960]_  = ~A166 & \new_[31959]_ ;
  assign \new_[31961]_  = \new_[31960]_  & \new_[31955]_ ;
  assign \new_[31965]_  = A298 & A268;
  assign \new_[31966]_  = ~A267 & \new_[31965]_ ;
  assign \new_[31970]_  = A302 & A300;
  assign \new_[31971]_  = ~A299 & \new_[31970]_ ;
  assign \new_[31972]_  = \new_[31971]_  & \new_[31966]_ ;
  assign \new_[31976]_  = A167 & A168;
  assign \new_[31977]_  = A169 & \new_[31976]_ ;
  assign \new_[31981]_  = A203 & ~A201;
  assign \new_[31982]_  = ~A166 & \new_[31981]_ ;
  assign \new_[31983]_  = \new_[31982]_  & \new_[31977]_ ;
  assign \new_[31987]_  = ~A298 & A268;
  assign \new_[31988]_  = ~A267 & \new_[31987]_ ;
  assign \new_[31992]_  = A301 & A300;
  assign \new_[31993]_  = A299 & \new_[31992]_ ;
  assign \new_[31994]_  = \new_[31993]_  & \new_[31988]_ ;
  assign \new_[31998]_  = A167 & A168;
  assign \new_[31999]_  = A169 & \new_[31998]_ ;
  assign \new_[32003]_  = A203 & ~A201;
  assign \new_[32004]_  = ~A166 & \new_[32003]_ ;
  assign \new_[32005]_  = \new_[32004]_  & \new_[31999]_ ;
  assign \new_[32009]_  = ~A298 & A268;
  assign \new_[32010]_  = ~A267 & \new_[32009]_ ;
  assign \new_[32014]_  = A302 & A300;
  assign \new_[32015]_  = A299 & \new_[32014]_ ;
  assign \new_[32016]_  = \new_[32015]_  & \new_[32010]_ ;
  assign \new_[32020]_  = A167 & A168;
  assign \new_[32021]_  = A169 & \new_[32020]_ ;
  assign \new_[32025]_  = A203 & ~A201;
  assign \new_[32026]_  = ~A166 & \new_[32025]_ ;
  assign \new_[32027]_  = \new_[32026]_  & \new_[32021]_ ;
  assign \new_[32031]_  = A298 & A269;
  assign \new_[32032]_  = ~A267 & \new_[32031]_ ;
  assign \new_[32036]_  = A301 & A300;
  assign \new_[32037]_  = ~A299 & \new_[32036]_ ;
  assign \new_[32038]_  = \new_[32037]_  & \new_[32032]_ ;
  assign \new_[32042]_  = A167 & A168;
  assign \new_[32043]_  = A169 & \new_[32042]_ ;
  assign \new_[32047]_  = A203 & ~A201;
  assign \new_[32048]_  = ~A166 & \new_[32047]_ ;
  assign \new_[32049]_  = \new_[32048]_  & \new_[32043]_ ;
  assign \new_[32053]_  = A298 & A269;
  assign \new_[32054]_  = ~A267 & \new_[32053]_ ;
  assign \new_[32058]_  = A302 & A300;
  assign \new_[32059]_  = ~A299 & \new_[32058]_ ;
  assign \new_[32060]_  = \new_[32059]_  & \new_[32054]_ ;
  assign \new_[32064]_  = A167 & A168;
  assign \new_[32065]_  = A169 & \new_[32064]_ ;
  assign \new_[32069]_  = A203 & ~A201;
  assign \new_[32070]_  = ~A166 & \new_[32069]_ ;
  assign \new_[32071]_  = \new_[32070]_  & \new_[32065]_ ;
  assign \new_[32075]_  = ~A298 & A269;
  assign \new_[32076]_  = ~A267 & \new_[32075]_ ;
  assign \new_[32080]_  = A301 & A300;
  assign \new_[32081]_  = A299 & \new_[32080]_ ;
  assign \new_[32082]_  = \new_[32081]_  & \new_[32076]_ ;
  assign \new_[32086]_  = A167 & A168;
  assign \new_[32087]_  = A169 & \new_[32086]_ ;
  assign \new_[32091]_  = A203 & ~A201;
  assign \new_[32092]_  = ~A166 & \new_[32091]_ ;
  assign \new_[32093]_  = \new_[32092]_  & \new_[32087]_ ;
  assign \new_[32097]_  = ~A298 & A269;
  assign \new_[32098]_  = ~A267 & \new_[32097]_ ;
  assign \new_[32102]_  = A302 & A300;
  assign \new_[32103]_  = A299 & \new_[32102]_ ;
  assign \new_[32104]_  = \new_[32103]_  & \new_[32098]_ ;
  assign \new_[32108]_  = A167 & A168;
  assign \new_[32109]_  = A169 & \new_[32108]_ ;
  assign \new_[32113]_  = A203 & ~A201;
  assign \new_[32114]_  = ~A166 & \new_[32113]_ ;
  assign \new_[32115]_  = \new_[32114]_  & \new_[32109]_ ;
  assign \new_[32119]_  = A298 & A266;
  assign \new_[32120]_  = A265 & \new_[32119]_ ;
  assign \new_[32124]_  = A301 & A300;
  assign \new_[32125]_  = ~A299 & \new_[32124]_ ;
  assign \new_[32126]_  = \new_[32125]_  & \new_[32120]_ ;
  assign \new_[32130]_  = A167 & A168;
  assign \new_[32131]_  = A169 & \new_[32130]_ ;
  assign \new_[32135]_  = A203 & ~A201;
  assign \new_[32136]_  = ~A166 & \new_[32135]_ ;
  assign \new_[32137]_  = \new_[32136]_  & \new_[32131]_ ;
  assign \new_[32141]_  = A298 & A266;
  assign \new_[32142]_  = A265 & \new_[32141]_ ;
  assign \new_[32146]_  = A302 & A300;
  assign \new_[32147]_  = ~A299 & \new_[32146]_ ;
  assign \new_[32148]_  = \new_[32147]_  & \new_[32142]_ ;
  assign \new_[32152]_  = A167 & A168;
  assign \new_[32153]_  = A169 & \new_[32152]_ ;
  assign \new_[32157]_  = A203 & ~A201;
  assign \new_[32158]_  = ~A166 & \new_[32157]_ ;
  assign \new_[32159]_  = \new_[32158]_  & \new_[32153]_ ;
  assign \new_[32163]_  = ~A298 & A266;
  assign \new_[32164]_  = A265 & \new_[32163]_ ;
  assign \new_[32168]_  = A301 & A300;
  assign \new_[32169]_  = A299 & \new_[32168]_ ;
  assign \new_[32170]_  = \new_[32169]_  & \new_[32164]_ ;
  assign \new_[32174]_  = A167 & A168;
  assign \new_[32175]_  = A169 & \new_[32174]_ ;
  assign \new_[32179]_  = A203 & ~A201;
  assign \new_[32180]_  = ~A166 & \new_[32179]_ ;
  assign \new_[32181]_  = \new_[32180]_  & \new_[32175]_ ;
  assign \new_[32185]_  = ~A298 & A266;
  assign \new_[32186]_  = A265 & \new_[32185]_ ;
  assign \new_[32190]_  = A302 & A300;
  assign \new_[32191]_  = A299 & \new_[32190]_ ;
  assign \new_[32192]_  = \new_[32191]_  & \new_[32186]_ ;
  assign \new_[32196]_  = A167 & A168;
  assign \new_[32197]_  = A169 & \new_[32196]_ ;
  assign \new_[32201]_  = A203 & ~A201;
  assign \new_[32202]_  = ~A166 & \new_[32201]_ ;
  assign \new_[32203]_  = \new_[32202]_  & \new_[32197]_ ;
  assign \new_[32207]_  = A298 & ~A266;
  assign \new_[32208]_  = ~A265 & \new_[32207]_ ;
  assign \new_[32212]_  = A301 & A300;
  assign \new_[32213]_  = ~A299 & \new_[32212]_ ;
  assign \new_[32214]_  = \new_[32213]_  & \new_[32208]_ ;
  assign \new_[32218]_  = A167 & A168;
  assign \new_[32219]_  = A169 & \new_[32218]_ ;
  assign \new_[32223]_  = A203 & ~A201;
  assign \new_[32224]_  = ~A166 & \new_[32223]_ ;
  assign \new_[32225]_  = \new_[32224]_  & \new_[32219]_ ;
  assign \new_[32229]_  = A298 & ~A266;
  assign \new_[32230]_  = ~A265 & \new_[32229]_ ;
  assign \new_[32234]_  = A302 & A300;
  assign \new_[32235]_  = ~A299 & \new_[32234]_ ;
  assign \new_[32236]_  = \new_[32235]_  & \new_[32230]_ ;
  assign \new_[32240]_  = A167 & A168;
  assign \new_[32241]_  = A169 & \new_[32240]_ ;
  assign \new_[32245]_  = A203 & ~A201;
  assign \new_[32246]_  = ~A166 & \new_[32245]_ ;
  assign \new_[32247]_  = \new_[32246]_  & \new_[32241]_ ;
  assign \new_[32251]_  = ~A298 & ~A266;
  assign \new_[32252]_  = ~A265 & \new_[32251]_ ;
  assign \new_[32256]_  = A301 & A300;
  assign \new_[32257]_  = A299 & \new_[32256]_ ;
  assign \new_[32258]_  = \new_[32257]_  & \new_[32252]_ ;
  assign \new_[32262]_  = A167 & A168;
  assign \new_[32263]_  = A169 & \new_[32262]_ ;
  assign \new_[32267]_  = A203 & ~A201;
  assign \new_[32268]_  = ~A166 & \new_[32267]_ ;
  assign \new_[32269]_  = \new_[32268]_  & \new_[32263]_ ;
  assign \new_[32273]_  = ~A298 & ~A266;
  assign \new_[32274]_  = ~A265 & \new_[32273]_ ;
  assign \new_[32278]_  = A302 & A300;
  assign \new_[32279]_  = A299 & \new_[32278]_ ;
  assign \new_[32280]_  = \new_[32279]_  & \new_[32274]_ ;
  assign \new_[32284]_  = A167 & A168;
  assign \new_[32285]_  = A169 & \new_[32284]_ ;
  assign \new_[32289]_  = A200 & A199;
  assign \new_[32290]_  = ~A166 & \new_[32289]_ ;
  assign \new_[32291]_  = \new_[32290]_  & \new_[32285]_ ;
  assign \new_[32295]_  = A298 & A268;
  assign \new_[32296]_  = ~A267 & \new_[32295]_ ;
  assign \new_[32300]_  = A301 & A300;
  assign \new_[32301]_  = ~A299 & \new_[32300]_ ;
  assign \new_[32302]_  = \new_[32301]_  & \new_[32296]_ ;
  assign \new_[32306]_  = A167 & A168;
  assign \new_[32307]_  = A169 & \new_[32306]_ ;
  assign \new_[32311]_  = A200 & A199;
  assign \new_[32312]_  = ~A166 & \new_[32311]_ ;
  assign \new_[32313]_  = \new_[32312]_  & \new_[32307]_ ;
  assign \new_[32317]_  = A298 & A268;
  assign \new_[32318]_  = ~A267 & \new_[32317]_ ;
  assign \new_[32322]_  = A302 & A300;
  assign \new_[32323]_  = ~A299 & \new_[32322]_ ;
  assign \new_[32324]_  = \new_[32323]_  & \new_[32318]_ ;
  assign \new_[32328]_  = A167 & A168;
  assign \new_[32329]_  = A169 & \new_[32328]_ ;
  assign \new_[32333]_  = A200 & A199;
  assign \new_[32334]_  = ~A166 & \new_[32333]_ ;
  assign \new_[32335]_  = \new_[32334]_  & \new_[32329]_ ;
  assign \new_[32339]_  = ~A298 & A268;
  assign \new_[32340]_  = ~A267 & \new_[32339]_ ;
  assign \new_[32344]_  = A301 & A300;
  assign \new_[32345]_  = A299 & \new_[32344]_ ;
  assign \new_[32346]_  = \new_[32345]_  & \new_[32340]_ ;
  assign \new_[32350]_  = A167 & A168;
  assign \new_[32351]_  = A169 & \new_[32350]_ ;
  assign \new_[32355]_  = A200 & A199;
  assign \new_[32356]_  = ~A166 & \new_[32355]_ ;
  assign \new_[32357]_  = \new_[32356]_  & \new_[32351]_ ;
  assign \new_[32361]_  = ~A298 & A268;
  assign \new_[32362]_  = ~A267 & \new_[32361]_ ;
  assign \new_[32366]_  = A302 & A300;
  assign \new_[32367]_  = A299 & \new_[32366]_ ;
  assign \new_[32368]_  = \new_[32367]_  & \new_[32362]_ ;
  assign \new_[32372]_  = A167 & A168;
  assign \new_[32373]_  = A169 & \new_[32372]_ ;
  assign \new_[32377]_  = A200 & A199;
  assign \new_[32378]_  = ~A166 & \new_[32377]_ ;
  assign \new_[32379]_  = \new_[32378]_  & \new_[32373]_ ;
  assign \new_[32383]_  = A298 & A269;
  assign \new_[32384]_  = ~A267 & \new_[32383]_ ;
  assign \new_[32388]_  = A301 & A300;
  assign \new_[32389]_  = ~A299 & \new_[32388]_ ;
  assign \new_[32390]_  = \new_[32389]_  & \new_[32384]_ ;
  assign \new_[32394]_  = A167 & A168;
  assign \new_[32395]_  = A169 & \new_[32394]_ ;
  assign \new_[32399]_  = A200 & A199;
  assign \new_[32400]_  = ~A166 & \new_[32399]_ ;
  assign \new_[32401]_  = \new_[32400]_  & \new_[32395]_ ;
  assign \new_[32405]_  = A298 & A269;
  assign \new_[32406]_  = ~A267 & \new_[32405]_ ;
  assign \new_[32410]_  = A302 & A300;
  assign \new_[32411]_  = ~A299 & \new_[32410]_ ;
  assign \new_[32412]_  = \new_[32411]_  & \new_[32406]_ ;
  assign \new_[32416]_  = A167 & A168;
  assign \new_[32417]_  = A169 & \new_[32416]_ ;
  assign \new_[32421]_  = A200 & A199;
  assign \new_[32422]_  = ~A166 & \new_[32421]_ ;
  assign \new_[32423]_  = \new_[32422]_  & \new_[32417]_ ;
  assign \new_[32427]_  = ~A298 & A269;
  assign \new_[32428]_  = ~A267 & \new_[32427]_ ;
  assign \new_[32432]_  = A301 & A300;
  assign \new_[32433]_  = A299 & \new_[32432]_ ;
  assign \new_[32434]_  = \new_[32433]_  & \new_[32428]_ ;
  assign \new_[32438]_  = A167 & A168;
  assign \new_[32439]_  = A169 & \new_[32438]_ ;
  assign \new_[32443]_  = A200 & A199;
  assign \new_[32444]_  = ~A166 & \new_[32443]_ ;
  assign \new_[32445]_  = \new_[32444]_  & \new_[32439]_ ;
  assign \new_[32449]_  = ~A298 & A269;
  assign \new_[32450]_  = ~A267 & \new_[32449]_ ;
  assign \new_[32454]_  = A302 & A300;
  assign \new_[32455]_  = A299 & \new_[32454]_ ;
  assign \new_[32456]_  = \new_[32455]_  & \new_[32450]_ ;
  assign \new_[32460]_  = A167 & A168;
  assign \new_[32461]_  = A169 & \new_[32460]_ ;
  assign \new_[32465]_  = A200 & A199;
  assign \new_[32466]_  = ~A166 & \new_[32465]_ ;
  assign \new_[32467]_  = \new_[32466]_  & \new_[32461]_ ;
  assign \new_[32471]_  = A298 & A266;
  assign \new_[32472]_  = A265 & \new_[32471]_ ;
  assign \new_[32476]_  = A301 & A300;
  assign \new_[32477]_  = ~A299 & \new_[32476]_ ;
  assign \new_[32478]_  = \new_[32477]_  & \new_[32472]_ ;
  assign \new_[32482]_  = A167 & A168;
  assign \new_[32483]_  = A169 & \new_[32482]_ ;
  assign \new_[32487]_  = A200 & A199;
  assign \new_[32488]_  = ~A166 & \new_[32487]_ ;
  assign \new_[32489]_  = \new_[32488]_  & \new_[32483]_ ;
  assign \new_[32493]_  = A298 & A266;
  assign \new_[32494]_  = A265 & \new_[32493]_ ;
  assign \new_[32498]_  = A302 & A300;
  assign \new_[32499]_  = ~A299 & \new_[32498]_ ;
  assign \new_[32500]_  = \new_[32499]_  & \new_[32494]_ ;
  assign \new_[32504]_  = A167 & A168;
  assign \new_[32505]_  = A169 & \new_[32504]_ ;
  assign \new_[32509]_  = A200 & A199;
  assign \new_[32510]_  = ~A166 & \new_[32509]_ ;
  assign \new_[32511]_  = \new_[32510]_  & \new_[32505]_ ;
  assign \new_[32515]_  = ~A298 & A266;
  assign \new_[32516]_  = A265 & \new_[32515]_ ;
  assign \new_[32520]_  = A301 & A300;
  assign \new_[32521]_  = A299 & \new_[32520]_ ;
  assign \new_[32522]_  = \new_[32521]_  & \new_[32516]_ ;
  assign \new_[32526]_  = A167 & A168;
  assign \new_[32527]_  = A169 & \new_[32526]_ ;
  assign \new_[32531]_  = A200 & A199;
  assign \new_[32532]_  = ~A166 & \new_[32531]_ ;
  assign \new_[32533]_  = \new_[32532]_  & \new_[32527]_ ;
  assign \new_[32537]_  = ~A298 & A266;
  assign \new_[32538]_  = A265 & \new_[32537]_ ;
  assign \new_[32542]_  = A302 & A300;
  assign \new_[32543]_  = A299 & \new_[32542]_ ;
  assign \new_[32544]_  = \new_[32543]_  & \new_[32538]_ ;
  assign \new_[32548]_  = A167 & A168;
  assign \new_[32549]_  = A169 & \new_[32548]_ ;
  assign \new_[32553]_  = A200 & A199;
  assign \new_[32554]_  = ~A166 & \new_[32553]_ ;
  assign \new_[32555]_  = \new_[32554]_  & \new_[32549]_ ;
  assign \new_[32559]_  = A298 & ~A266;
  assign \new_[32560]_  = ~A265 & \new_[32559]_ ;
  assign \new_[32564]_  = A301 & A300;
  assign \new_[32565]_  = ~A299 & \new_[32564]_ ;
  assign \new_[32566]_  = \new_[32565]_  & \new_[32560]_ ;
  assign \new_[32570]_  = A167 & A168;
  assign \new_[32571]_  = A169 & \new_[32570]_ ;
  assign \new_[32575]_  = A200 & A199;
  assign \new_[32576]_  = ~A166 & \new_[32575]_ ;
  assign \new_[32577]_  = \new_[32576]_  & \new_[32571]_ ;
  assign \new_[32581]_  = A298 & ~A266;
  assign \new_[32582]_  = ~A265 & \new_[32581]_ ;
  assign \new_[32586]_  = A302 & A300;
  assign \new_[32587]_  = ~A299 & \new_[32586]_ ;
  assign \new_[32588]_  = \new_[32587]_  & \new_[32582]_ ;
  assign \new_[32592]_  = A167 & A168;
  assign \new_[32593]_  = A169 & \new_[32592]_ ;
  assign \new_[32597]_  = A200 & A199;
  assign \new_[32598]_  = ~A166 & \new_[32597]_ ;
  assign \new_[32599]_  = \new_[32598]_  & \new_[32593]_ ;
  assign \new_[32603]_  = ~A298 & ~A266;
  assign \new_[32604]_  = ~A265 & \new_[32603]_ ;
  assign \new_[32608]_  = A301 & A300;
  assign \new_[32609]_  = A299 & \new_[32608]_ ;
  assign \new_[32610]_  = \new_[32609]_  & \new_[32604]_ ;
  assign \new_[32614]_  = A167 & A168;
  assign \new_[32615]_  = A169 & \new_[32614]_ ;
  assign \new_[32619]_  = A200 & A199;
  assign \new_[32620]_  = ~A166 & \new_[32619]_ ;
  assign \new_[32621]_  = \new_[32620]_  & \new_[32615]_ ;
  assign \new_[32625]_  = ~A298 & ~A266;
  assign \new_[32626]_  = ~A265 & \new_[32625]_ ;
  assign \new_[32630]_  = A302 & A300;
  assign \new_[32631]_  = A299 & \new_[32630]_ ;
  assign \new_[32632]_  = \new_[32631]_  & \new_[32626]_ ;
  assign \new_[32636]_  = A167 & A168;
  assign \new_[32637]_  = A169 & \new_[32636]_ ;
  assign \new_[32641]_  = ~A200 & ~A199;
  assign \new_[32642]_  = ~A166 & \new_[32641]_ ;
  assign \new_[32643]_  = \new_[32642]_  & \new_[32637]_ ;
  assign \new_[32647]_  = A298 & A268;
  assign \new_[32648]_  = ~A267 & \new_[32647]_ ;
  assign \new_[32652]_  = A301 & A300;
  assign \new_[32653]_  = ~A299 & \new_[32652]_ ;
  assign \new_[32654]_  = \new_[32653]_  & \new_[32648]_ ;
  assign \new_[32658]_  = A167 & A168;
  assign \new_[32659]_  = A169 & \new_[32658]_ ;
  assign \new_[32663]_  = ~A200 & ~A199;
  assign \new_[32664]_  = ~A166 & \new_[32663]_ ;
  assign \new_[32665]_  = \new_[32664]_  & \new_[32659]_ ;
  assign \new_[32669]_  = A298 & A268;
  assign \new_[32670]_  = ~A267 & \new_[32669]_ ;
  assign \new_[32674]_  = A302 & A300;
  assign \new_[32675]_  = ~A299 & \new_[32674]_ ;
  assign \new_[32676]_  = \new_[32675]_  & \new_[32670]_ ;
  assign \new_[32680]_  = A167 & A168;
  assign \new_[32681]_  = A169 & \new_[32680]_ ;
  assign \new_[32685]_  = ~A200 & ~A199;
  assign \new_[32686]_  = ~A166 & \new_[32685]_ ;
  assign \new_[32687]_  = \new_[32686]_  & \new_[32681]_ ;
  assign \new_[32691]_  = ~A298 & A268;
  assign \new_[32692]_  = ~A267 & \new_[32691]_ ;
  assign \new_[32696]_  = A301 & A300;
  assign \new_[32697]_  = A299 & \new_[32696]_ ;
  assign \new_[32698]_  = \new_[32697]_  & \new_[32692]_ ;
  assign \new_[32702]_  = A167 & A168;
  assign \new_[32703]_  = A169 & \new_[32702]_ ;
  assign \new_[32707]_  = ~A200 & ~A199;
  assign \new_[32708]_  = ~A166 & \new_[32707]_ ;
  assign \new_[32709]_  = \new_[32708]_  & \new_[32703]_ ;
  assign \new_[32713]_  = ~A298 & A268;
  assign \new_[32714]_  = ~A267 & \new_[32713]_ ;
  assign \new_[32718]_  = A302 & A300;
  assign \new_[32719]_  = A299 & \new_[32718]_ ;
  assign \new_[32720]_  = \new_[32719]_  & \new_[32714]_ ;
  assign \new_[32724]_  = A167 & A168;
  assign \new_[32725]_  = A169 & \new_[32724]_ ;
  assign \new_[32729]_  = ~A200 & ~A199;
  assign \new_[32730]_  = ~A166 & \new_[32729]_ ;
  assign \new_[32731]_  = \new_[32730]_  & \new_[32725]_ ;
  assign \new_[32735]_  = A298 & A269;
  assign \new_[32736]_  = ~A267 & \new_[32735]_ ;
  assign \new_[32740]_  = A301 & A300;
  assign \new_[32741]_  = ~A299 & \new_[32740]_ ;
  assign \new_[32742]_  = \new_[32741]_  & \new_[32736]_ ;
  assign \new_[32746]_  = A167 & A168;
  assign \new_[32747]_  = A169 & \new_[32746]_ ;
  assign \new_[32751]_  = ~A200 & ~A199;
  assign \new_[32752]_  = ~A166 & \new_[32751]_ ;
  assign \new_[32753]_  = \new_[32752]_  & \new_[32747]_ ;
  assign \new_[32757]_  = A298 & A269;
  assign \new_[32758]_  = ~A267 & \new_[32757]_ ;
  assign \new_[32762]_  = A302 & A300;
  assign \new_[32763]_  = ~A299 & \new_[32762]_ ;
  assign \new_[32764]_  = \new_[32763]_  & \new_[32758]_ ;
  assign \new_[32768]_  = A167 & A168;
  assign \new_[32769]_  = A169 & \new_[32768]_ ;
  assign \new_[32773]_  = ~A200 & ~A199;
  assign \new_[32774]_  = ~A166 & \new_[32773]_ ;
  assign \new_[32775]_  = \new_[32774]_  & \new_[32769]_ ;
  assign \new_[32779]_  = ~A298 & A269;
  assign \new_[32780]_  = ~A267 & \new_[32779]_ ;
  assign \new_[32784]_  = A301 & A300;
  assign \new_[32785]_  = A299 & \new_[32784]_ ;
  assign \new_[32786]_  = \new_[32785]_  & \new_[32780]_ ;
  assign \new_[32790]_  = A167 & A168;
  assign \new_[32791]_  = A169 & \new_[32790]_ ;
  assign \new_[32795]_  = ~A200 & ~A199;
  assign \new_[32796]_  = ~A166 & \new_[32795]_ ;
  assign \new_[32797]_  = \new_[32796]_  & \new_[32791]_ ;
  assign \new_[32801]_  = ~A298 & A269;
  assign \new_[32802]_  = ~A267 & \new_[32801]_ ;
  assign \new_[32806]_  = A302 & A300;
  assign \new_[32807]_  = A299 & \new_[32806]_ ;
  assign \new_[32808]_  = \new_[32807]_  & \new_[32802]_ ;
  assign \new_[32812]_  = A167 & A168;
  assign \new_[32813]_  = A169 & \new_[32812]_ ;
  assign \new_[32817]_  = ~A200 & ~A199;
  assign \new_[32818]_  = ~A166 & \new_[32817]_ ;
  assign \new_[32819]_  = \new_[32818]_  & \new_[32813]_ ;
  assign \new_[32823]_  = A298 & A266;
  assign \new_[32824]_  = A265 & \new_[32823]_ ;
  assign \new_[32828]_  = A301 & A300;
  assign \new_[32829]_  = ~A299 & \new_[32828]_ ;
  assign \new_[32830]_  = \new_[32829]_  & \new_[32824]_ ;
  assign \new_[32834]_  = A167 & A168;
  assign \new_[32835]_  = A169 & \new_[32834]_ ;
  assign \new_[32839]_  = ~A200 & ~A199;
  assign \new_[32840]_  = ~A166 & \new_[32839]_ ;
  assign \new_[32841]_  = \new_[32840]_  & \new_[32835]_ ;
  assign \new_[32845]_  = A298 & A266;
  assign \new_[32846]_  = A265 & \new_[32845]_ ;
  assign \new_[32850]_  = A302 & A300;
  assign \new_[32851]_  = ~A299 & \new_[32850]_ ;
  assign \new_[32852]_  = \new_[32851]_  & \new_[32846]_ ;
  assign \new_[32856]_  = A167 & A168;
  assign \new_[32857]_  = A169 & \new_[32856]_ ;
  assign \new_[32861]_  = ~A200 & ~A199;
  assign \new_[32862]_  = ~A166 & \new_[32861]_ ;
  assign \new_[32863]_  = \new_[32862]_  & \new_[32857]_ ;
  assign \new_[32867]_  = ~A298 & A266;
  assign \new_[32868]_  = A265 & \new_[32867]_ ;
  assign \new_[32872]_  = A301 & A300;
  assign \new_[32873]_  = A299 & \new_[32872]_ ;
  assign \new_[32874]_  = \new_[32873]_  & \new_[32868]_ ;
  assign \new_[32878]_  = A167 & A168;
  assign \new_[32879]_  = A169 & \new_[32878]_ ;
  assign \new_[32883]_  = ~A200 & ~A199;
  assign \new_[32884]_  = ~A166 & \new_[32883]_ ;
  assign \new_[32885]_  = \new_[32884]_  & \new_[32879]_ ;
  assign \new_[32889]_  = ~A298 & A266;
  assign \new_[32890]_  = A265 & \new_[32889]_ ;
  assign \new_[32894]_  = A302 & A300;
  assign \new_[32895]_  = A299 & \new_[32894]_ ;
  assign \new_[32896]_  = \new_[32895]_  & \new_[32890]_ ;
  assign \new_[32900]_  = A167 & A168;
  assign \new_[32901]_  = A169 & \new_[32900]_ ;
  assign \new_[32905]_  = ~A200 & ~A199;
  assign \new_[32906]_  = ~A166 & \new_[32905]_ ;
  assign \new_[32907]_  = \new_[32906]_  & \new_[32901]_ ;
  assign \new_[32911]_  = A298 & ~A266;
  assign \new_[32912]_  = ~A265 & \new_[32911]_ ;
  assign \new_[32916]_  = A301 & A300;
  assign \new_[32917]_  = ~A299 & \new_[32916]_ ;
  assign \new_[32918]_  = \new_[32917]_  & \new_[32912]_ ;
  assign \new_[32922]_  = A167 & A168;
  assign \new_[32923]_  = A169 & \new_[32922]_ ;
  assign \new_[32927]_  = ~A200 & ~A199;
  assign \new_[32928]_  = ~A166 & \new_[32927]_ ;
  assign \new_[32929]_  = \new_[32928]_  & \new_[32923]_ ;
  assign \new_[32933]_  = A298 & ~A266;
  assign \new_[32934]_  = ~A265 & \new_[32933]_ ;
  assign \new_[32938]_  = A302 & A300;
  assign \new_[32939]_  = ~A299 & \new_[32938]_ ;
  assign \new_[32940]_  = \new_[32939]_  & \new_[32934]_ ;
  assign \new_[32944]_  = A167 & A168;
  assign \new_[32945]_  = A169 & \new_[32944]_ ;
  assign \new_[32949]_  = ~A200 & ~A199;
  assign \new_[32950]_  = ~A166 & \new_[32949]_ ;
  assign \new_[32951]_  = \new_[32950]_  & \new_[32945]_ ;
  assign \new_[32955]_  = ~A298 & ~A266;
  assign \new_[32956]_  = ~A265 & \new_[32955]_ ;
  assign \new_[32960]_  = A301 & A300;
  assign \new_[32961]_  = A299 & \new_[32960]_ ;
  assign \new_[32962]_  = \new_[32961]_  & \new_[32956]_ ;
  assign \new_[32966]_  = A167 & A168;
  assign \new_[32967]_  = A169 & \new_[32966]_ ;
  assign \new_[32971]_  = ~A200 & ~A199;
  assign \new_[32972]_  = ~A166 & \new_[32971]_ ;
  assign \new_[32973]_  = \new_[32972]_  & \new_[32967]_ ;
  assign \new_[32977]_  = ~A298 & ~A266;
  assign \new_[32978]_  = ~A265 & \new_[32977]_ ;
  assign \new_[32982]_  = A302 & A300;
  assign \new_[32983]_  = A299 & \new_[32982]_ ;
  assign \new_[32984]_  = \new_[32983]_  & \new_[32978]_ ;
  assign \new_[32988]_  = ~A167 & A168;
  assign \new_[32989]_  = A169 & \new_[32988]_ ;
  assign \new_[32993]_  = A202 & ~A201;
  assign \new_[32994]_  = A166 & \new_[32993]_ ;
  assign \new_[32995]_  = \new_[32994]_  & \new_[32989]_ ;
  assign \new_[32999]_  = A298 & A268;
  assign \new_[33000]_  = ~A267 & \new_[32999]_ ;
  assign \new_[33004]_  = A301 & A300;
  assign \new_[33005]_  = ~A299 & \new_[33004]_ ;
  assign \new_[33006]_  = \new_[33005]_  & \new_[33000]_ ;
  assign \new_[33010]_  = ~A167 & A168;
  assign \new_[33011]_  = A169 & \new_[33010]_ ;
  assign \new_[33015]_  = A202 & ~A201;
  assign \new_[33016]_  = A166 & \new_[33015]_ ;
  assign \new_[33017]_  = \new_[33016]_  & \new_[33011]_ ;
  assign \new_[33021]_  = A298 & A268;
  assign \new_[33022]_  = ~A267 & \new_[33021]_ ;
  assign \new_[33026]_  = A302 & A300;
  assign \new_[33027]_  = ~A299 & \new_[33026]_ ;
  assign \new_[33028]_  = \new_[33027]_  & \new_[33022]_ ;
  assign \new_[33032]_  = ~A167 & A168;
  assign \new_[33033]_  = A169 & \new_[33032]_ ;
  assign \new_[33037]_  = A202 & ~A201;
  assign \new_[33038]_  = A166 & \new_[33037]_ ;
  assign \new_[33039]_  = \new_[33038]_  & \new_[33033]_ ;
  assign \new_[33043]_  = ~A298 & A268;
  assign \new_[33044]_  = ~A267 & \new_[33043]_ ;
  assign \new_[33048]_  = A301 & A300;
  assign \new_[33049]_  = A299 & \new_[33048]_ ;
  assign \new_[33050]_  = \new_[33049]_  & \new_[33044]_ ;
  assign \new_[33054]_  = ~A167 & A168;
  assign \new_[33055]_  = A169 & \new_[33054]_ ;
  assign \new_[33059]_  = A202 & ~A201;
  assign \new_[33060]_  = A166 & \new_[33059]_ ;
  assign \new_[33061]_  = \new_[33060]_  & \new_[33055]_ ;
  assign \new_[33065]_  = ~A298 & A268;
  assign \new_[33066]_  = ~A267 & \new_[33065]_ ;
  assign \new_[33070]_  = A302 & A300;
  assign \new_[33071]_  = A299 & \new_[33070]_ ;
  assign \new_[33072]_  = \new_[33071]_  & \new_[33066]_ ;
  assign \new_[33076]_  = ~A167 & A168;
  assign \new_[33077]_  = A169 & \new_[33076]_ ;
  assign \new_[33081]_  = A202 & ~A201;
  assign \new_[33082]_  = A166 & \new_[33081]_ ;
  assign \new_[33083]_  = \new_[33082]_  & \new_[33077]_ ;
  assign \new_[33087]_  = A298 & A269;
  assign \new_[33088]_  = ~A267 & \new_[33087]_ ;
  assign \new_[33092]_  = A301 & A300;
  assign \new_[33093]_  = ~A299 & \new_[33092]_ ;
  assign \new_[33094]_  = \new_[33093]_  & \new_[33088]_ ;
  assign \new_[33098]_  = ~A167 & A168;
  assign \new_[33099]_  = A169 & \new_[33098]_ ;
  assign \new_[33103]_  = A202 & ~A201;
  assign \new_[33104]_  = A166 & \new_[33103]_ ;
  assign \new_[33105]_  = \new_[33104]_  & \new_[33099]_ ;
  assign \new_[33109]_  = A298 & A269;
  assign \new_[33110]_  = ~A267 & \new_[33109]_ ;
  assign \new_[33114]_  = A302 & A300;
  assign \new_[33115]_  = ~A299 & \new_[33114]_ ;
  assign \new_[33116]_  = \new_[33115]_  & \new_[33110]_ ;
  assign \new_[33120]_  = ~A167 & A168;
  assign \new_[33121]_  = A169 & \new_[33120]_ ;
  assign \new_[33125]_  = A202 & ~A201;
  assign \new_[33126]_  = A166 & \new_[33125]_ ;
  assign \new_[33127]_  = \new_[33126]_  & \new_[33121]_ ;
  assign \new_[33131]_  = ~A298 & A269;
  assign \new_[33132]_  = ~A267 & \new_[33131]_ ;
  assign \new_[33136]_  = A301 & A300;
  assign \new_[33137]_  = A299 & \new_[33136]_ ;
  assign \new_[33138]_  = \new_[33137]_  & \new_[33132]_ ;
  assign \new_[33142]_  = ~A167 & A168;
  assign \new_[33143]_  = A169 & \new_[33142]_ ;
  assign \new_[33147]_  = A202 & ~A201;
  assign \new_[33148]_  = A166 & \new_[33147]_ ;
  assign \new_[33149]_  = \new_[33148]_  & \new_[33143]_ ;
  assign \new_[33153]_  = ~A298 & A269;
  assign \new_[33154]_  = ~A267 & \new_[33153]_ ;
  assign \new_[33158]_  = A302 & A300;
  assign \new_[33159]_  = A299 & \new_[33158]_ ;
  assign \new_[33160]_  = \new_[33159]_  & \new_[33154]_ ;
  assign \new_[33164]_  = ~A167 & A168;
  assign \new_[33165]_  = A169 & \new_[33164]_ ;
  assign \new_[33169]_  = A202 & ~A201;
  assign \new_[33170]_  = A166 & \new_[33169]_ ;
  assign \new_[33171]_  = \new_[33170]_  & \new_[33165]_ ;
  assign \new_[33175]_  = A298 & A266;
  assign \new_[33176]_  = A265 & \new_[33175]_ ;
  assign \new_[33180]_  = A301 & A300;
  assign \new_[33181]_  = ~A299 & \new_[33180]_ ;
  assign \new_[33182]_  = \new_[33181]_  & \new_[33176]_ ;
  assign \new_[33186]_  = ~A167 & A168;
  assign \new_[33187]_  = A169 & \new_[33186]_ ;
  assign \new_[33191]_  = A202 & ~A201;
  assign \new_[33192]_  = A166 & \new_[33191]_ ;
  assign \new_[33193]_  = \new_[33192]_  & \new_[33187]_ ;
  assign \new_[33197]_  = A298 & A266;
  assign \new_[33198]_  = A265 & \new_[33197]_ ;
  assign \new_[33202]_  = A302 & A300;
  assign \new_[33203]_  = ~A299 & \new_[33202]_ ;
  assign \new_[33204]_  = \new_[33203]_  & \new_[33198]_ ;
  assign \new_[33208]_  = ~A167 & A168;
  assign \new_[33209]_  = A169 & \new_[33208]_ ;
  assign \new_[33213]_  = A202 & ~A201;
  assign \new_[33214]_  = A166 & \new_[33213]_ ;
  assign \new_[33215]_  = \new_[33214]_  & \new_[33209]_ ;
  assign \new_[33219]_  = ~A298 & A266;
  assign \new_[33220]_  = A265 & \new_[33219]_ ;
  assign \new_[33224]_  = A301 & A300;
  assign \new_[33225]_  = A299 & \new_[33224]_ ;
  assign \new_[33226]_  = \new_[33225]_  & \new_[33220]_ ;
  assign \new_[33230]_  = ~A167 & A168;
  assign \new_[33231]_  = A169 & \new_[33230]_ ;
  assign \new_[33235]_  = A202 & ~A201;
  assign \new_[33236]_  = A166 & \new_[33235]_ ;
  assign \new_[33237]_  = \new_[33236]_  & \new_[33231]_ ;
  assign \new_[33241]_  = ~A298 & A266;
  assign \new_[33242]_  = A265 & \new_[33241]_ ;
  assign \new_[33246]_  = A302 & A300;
  assign \new_[33247]_  = A299 & \new_[33246]_ ;
  assign \new_[33248]_  = \new_[33247]_  & \new_[33242]_ ;
  assign \new_[33252]_  = ~A167 & A168;
  assign \new_[33253]_  = A169 & \new_[33252]_ ;
  assign \new_[33257]_  = A202 & ~A201;
  assign \new_[33258]_  = A166 & \new_[33257]_ ;
  assign \new_[33259]_  = \new_[33258]_  & \new_[33253]_ ;
  assign \new_[33263]_  = A298 & ~A266;
  assign \new_[33264]_  = ~A265 & \new_[33263]_ ;
  assign \new_[33268]_  = A301 & A300;
  assign \new_[33269]_  = ~A299 & \new_[33268]_ ;
  assign \new_[33270]_  = \new_[33269]_  & \new_[33264]_ ;
  assign \new_[33274]_  = ~A167 & A168;
  assign \new_[33275]_  = A169 & \new_[33274]_ ;
  assign \new_[33279]_  = A202 & ~A201;
  assign \new_[33280]_  = A166 & \new_[33279]_ ;
  assign \new_[33281]_  = \new_[33280]_  & \new_[33275]_ ;
  assign \new_[33285]_  = A298 & ~A266;
  assign \new_[33286]_  = ~A265 & \new_[33285]_ ;
  assign \new_[33290]_  = A302 & A300;
  assign \new_[33291]_  = ~A299 & \new_[33290]_ ;
  assign \new_[33292]_  = \new_[33291]_  & \new_[33286]_ ;
  assign \new_[33296]_  = ~A167 & A168;
  assign \new_[33297]_  = A169 & \new_[33296]_ ;
  assign \new_[33301]_  = A202 & ~A201;
  assign \new_[33302]_  = A166 & \new_[33301]_ ;
  assign \new_[33303]_  = \new_[33302]_  & \new_[33297]_ ;
  assign \new_[33307]_  = ~A298 & ~A266;
  assign \new_[33308]_  = ~A265 & \new_[33307]_ ;
  assign \new_[33312]_  = A301 & A300;
  assign \new_[33313]_  = A299 & \new_[33312]_ ;
  assign \new_[33314]_  = \new_[33313]_  & \new_[33308]_ ;
  assign \new_[33318]_  = ~A167 & A168;
  assign \new_[33319]_  = A169 & \new_[33318]_ ;
  assign \new_[33323]_  = A202 & ~A201;
  assign \new_[33324]_  = A166 & \new_[33323]_ ;
  assign \new_[33325]_  = \new_[33324]_  & \new_[33319]_ ;
  assign \new_[33329]_  = ~A298 & ~A266;
  assign \new_[33330]_  = ~A265 & \new_[33329]_ ;
  assign \new_[33334]_  = A302 & A300;
  assign \new_[33335]_  = A299 & \new_[33334]_ ;
  assign \new_[33336]_  = \new_[33335]_  & \new_[33330]_ ;
  assign \new_[33340]_  = ~A167 & A168;
  assign \new_[33341]_  = A169 & \new_[33340]_ ;
  assign \new_[33345]_  = A203 & ~A201;
  assign \new_[33346]_  = A166 & \new_[33345]_ ;
  assign \new_[33347]_  = \new_[33346]_  & \new_[33341]_ ;
  assign \new_[33351]_  = A298 & A268;
  assign \new_[33352]_  = ~A267 & \new_[33351]_ ;
  assign \new_[33356]_  = A301 & A300;
  assign \new_[33357]_  = ~A299 & \new_[33356]_ ;
  assign \new_[33358]_  = \new_[33357]_  & \new_[33352]_ ;
  assign \new_[33362]_  = ~A167 & A168;
  assign \new_[33363]_  = A169 & \new_[33362]_ ;
  assign \new_[33367]_  = A203 & ~A201;
  assign \new_[33368]_  = A166 & \new_[33367]_ ;
  assign \new_[33369]_  = \new_[33368]_  & \new_[33363]_ ;
  assign \new_[33373]_  = A298 & A268;
  assign \new_[33374]_  = ~A267 & \new_[33373]_ ;
  assign \new_[33378]_  = A302 & A300;
  assign \new_[33379]_  = ~A299 & \new_[33378]_ ;
  assign \new_[33380]_  = \new_[33379]_  & \new_[33374]_ ;
  assign \new_[33384]_  = ~A167 & A168;
  assign \new_[33385]_  = A169 & \new_[33384]_ ;
  assign \new_[33389]_  = A203 & ~A201;
  assign \new_[33390]_  = A166 & \new_[33389]_ ;
  assign \new_[33391]_  = \new_[33390]_  & \new_[33385]_ ;
  assign \new_[33395]_  = ~A298 & A268;
  assign \new_[33396]_  = ~A267 & \new_[33395]_ ;
  assign \new_[33400]_  = A301 & A300;
  assign \new_[33401]_  = A299 & \new_[33400]_ ;
  assign \new_[33402]_  = \new_[33401]_  & \new_[33396]_ ;
  assign \new_[33406]_  = ~A167 & A168;
  assign \new_[33407]_  = A169 & \new_[33406]_ ;
  assign \new_[33411]_  = A203 & ~A201;
  assign \new_[33412]_  = A166 & \new_[33411]_ ;
  assign \new_[33413]_  = \new_[33412]_  & \new_[33407]_ ;
  assign \new_[33417]_  = ~A298 & A268;
  assign \new_[33418]_  = ~A267 & \new_[33417]_ ;
  assign \new_[33422]_  = A302 & A300;
  assign \new_[33423]_  = A299 & \new_[33422]_ ;
  assign \new_[33424]_  = \new_[33423]_  & \new_[33418]_ ;
  assign \new_[33428]_  = ~A167 & A168;
  assign \new_[33429]_  = A169 & \new_[33428]_ ;
  assign \new_[33433]_  = A203 & ~A201;
  assign \new_[33434]_  = A166 & \new_[33433]_ ;
  assign \new_[33435]_  = \new_[33434]_  & \new_[33429]_ ;
  assign \new_[33439]_  = A298 & A269;
  assign \new_[33440]_  = ~A267 & \new_[33439]_ ;
  assign \new_[33444]_  = A301 & A300;
  assign \new_[33445]_  = ~A299 & \new_[33444]_ ;
  assign \new_[33446]_  = \new_[33445]_  & \new_[33440]_ ;
  assign \new_[33450]_  = ~A167 & A168;
  assign \new_[33451]_  = A169 & \new_[33450]_ ;
  assign \new_[33455]_  = A203 & ~A201;
  assign \new_[33456]_  = A166 & \new_[33455]_ ;
  assign \new_[33457]_  = \new_[33456]_  & \new_[33451]_ ;
  assign \new_[33461]_  = A298 & A269;
  assign \new_[33462]_  = ~A267 & \new_[33461]_ ;
  assign \new_[33466]_  = A302 & A300;
  assign \new_[33467]_  = ~A299 & \new_[33466]_ ;
  assign \new_[33468]_  = \new_[33467]_  & \new_[33462]_ ;
  assign \new_[33472]_  = ~A167 & A168;
  assign \new_[33473]_  = A169 & \new_[33472]_ ;
  assign \new_[33477]_  = A203 & ~A201;
  assign \new_[33478]_  = A166 & \new_[33477]_ ;
  assign \new_[33479]_  = \new_[33478]_  & \new_[33473]_ ;
  assign \new_[33483]_  = ~A298 & A269;
  assign \new_[33484]_  = ~A267 & \new_[33483]_ ;
  assign \new_[33488]_  = A301 & A300;
  assign \new_[33489]_  = A299 & \new_[33488]_ ;
  assign \new_[33490]_  = \new_[33489]_  & \new_[33484]_ ;
  assign \new_[33494]_  = ~A167 & A168;
  assign \new_[33495]_  = A169 & \new_[33494]_ ;
  assign \new_[33499]_  = A203 & ~A201;
  assign \new_[33500]_  = A166 & \new_[33499]_ ;
  assign \new_[33501]_  = \new_[33500]_  & \new_[33495]_ ;
  assign \new_[33505]_  = ~A298 & A269;
  assign \new_[33506]_  = ~A267 & \new_[33505]_ ;
  assign \new_[33510]_  = A302 & A300;
  assign \new_[33511]_  = A299 & \new_[33510]_ ;
  assign \new_[33512]_  = \new_[33511]_  & \new_[33506]_ ;
  assign \new_[33516]_  = ~A167 & A168;
  assign \new_[33517]_  = A169 & \new_[33516]_ ;
  assign \new_[33521]_  = A203 & ~A201;
  assign \new_[33522]_  = A166 & \new_[33521]_ ;
  assign \new_[33523]_  = \new_[33522]_  & \new_[33517]_ ;
  assign \new_[33527]_  = A298 & A266;
  assign \new_[33528]_  = A265 & \new_[33527]_ ;
  assign \new_[33532]_  = A301 & A300;
  assign \new_[33533]_  = ~A299 & \new_[33532]_ ;
  assign \new_[33534]_  = \new_[33533]_  & \new_[33528]_ ;
  assign \new_[33538]_  = ~A167 & A168;
  assign \new_[33539]_  = A169 & \new_[33538]_ ;
  assign \new_[33543]_  = A203 & ~A201;
  assign \new_[33544]_  = A166 & \new_[33543]_ ;
  assign \new_[33545]_  = \new_[33544]_  & \new_[33539]_ ;
  assign \new_[33549]_  = A298 & A266;
  assign \new_[33550]_  = A265 & \new_[33549]_ ;
  assign \new_[33554]_  = A302 & A300;
  assign \new_[33555]_  = ~A299 & \new_[33554]_ ;
  assign \new_[33556]_  = \new_[33555]_  & \new_[33550]_ ;
  assign \new_[33560]_  = ~A167 & A168;
  assign \new_[33561]_  = A169 & \new_[33560]_ ;
  assign \new_[33565]_  = A203 & ~A201;
  assign \new_[33566]_  = A166 & \new_[33565]_ ;
  assign \new_[33567]_  = \new_[33566]_  & \new_[33561]_ ;
  assign \new_[33571]_  = ~A298 & A266;
  assign \new_[33572]_  = A265 & \new_[33571]_ ;
  assign \new_[33576]_  = A301 & A300;
  assign \new_[33577]_  = A299 & \new_[33576]_ ;
  assign \new_[33578]_  = \new_[33577]_  & \new_[33572]_ ;
  assign \new_[33582]_  = ~A167 & A168;
  assign \new_[33583]_  = A169 & \new_[33582]_ ;
  assign \new_[33587]_  = A203 & ~A201;
  assign \new_[33588]_  = A166 & \new_[33587]_ ;
  assign \new_[33589]_  = \new_[33588]_  & \new_[33583]_ ;
  assign \new_[33593]_  = ~A298 & A266;
  assign \new_[33594]_  = A265 & \new_[33593]_ ;
  assign \new_[33598]_  = A302 & A300;
  assign \new_[33599]_  = A299 & \new_[33598]_ ;
  assign \new_[33600]_  = \new_[33599]_  & \new_[33594]_ ;
  assign \new_[33604]_  = ~A167 & A168;
  assign \new_[33605]_  = A169 & \new_[33604]_ ;
  assign \new_[33609]_  = A203 & ~A201;
  assign \new_[33610]_  = A166 & \new_[33609]_ ;
  assign \new_[33611]_  = \new_[33610]_  & \new_[33605]_ ;
  assign \new_[33615]_  = A298 & ~A266;
  assign \new_[33616]_  = ~A265 & \new_[33615]_ ;
  assign \new_[33620]_  = A301 & A300;
  assign \new_[33621]_  = ~A299 & \new_[33620]_ ;
  assign \new_[33622]_  = \new_[33621]_  & \new_[33616]_ ;
  assign \new_[33626]_  = ~A167 & A168;
  assign \new_[33627]_  = A169 & \new_[33626]_ ;
  assign \new_[33631]_  = A203 & ~A201;
  assign \new_[33632]_  = A166 & \new_[33631]_ ;
  assign \new_[33633]_  = \new_[33632]_  & \new_[33627]_ ;
  assign \new_[33637]_  = A298 & ~A266;
  assign \new_[33638]_  = ~A265 & \new_[33637]_ ;
  assign \new_[33642]_  = A302 & A300;
  assign \new_[33643]_  = ~A299 & \new_[33642]_ ;
  assign \new_[33644]_  = \new_[33643]_  & \new_[33638]_ ;
  assign \new_[33648]_  = ~A167 & A168;
  assign \new_[33649]_  = A169 & \new_[33648]_ ;
  assign \new_[33653]_  = A203 & ~A201;
  assign \new_[33654]_  = A166 & \new_[33653]_ ;
  assign \new_[33655]_  = \new_[33654]_  & \new_[33649]_ ;
  assign \new_[33659]_  = ~A298 & ~A266;
  assign \new_[33660]_  = ~A265 & \new_[33659]_ ;
  assign \new_[33664]_  = A301 & A300;
  assign \new_[33665]_  = A299 & \new_[33664]_ ;
  assign \new_[33666]_  = \new_[33665]_  & \new_[33660]_ ;
  assign \new_[33670]_  = ~A167 & A168;
  assign \new_[33671]_  = A169 & \new_[33670]_ ;
  assign \new_[33675]_  = A203 & ~A201;
  assign \new_[33676]_  = A166 & \new_[33675]_ ;
  assign \new_[33677]_  = \new_[33676]_  & \new_[33671]_ ;
  assign \new_[33681]_  = ~A298 & ~A266;
  assign \new_[33682]_  = ~A265 & \new_[33681]_ ;
  assign \new_[33686]_  = A302 & A300;
  assign \new_[33687]_  = A299 & \new_[33686]_ ;
  assign \new_[33688]_  = \new_[33687]_  & \new_[33682]_ ;
  assign \new_[33692]_  = ~A167 & A168;
  assign \new_[33693]_  = A169 & \new_[33692]_ ;
  assign \new_[33697]_  = A200 & A199;
  assign \new_[33698]_  = A166 & \new_[33697]_ ;
  assign \new_[33699]_  = \new_[33698]_  & \new_[33693]_ ;
  assign \new_[33703]_  = A298 & A268;
  assign \new_[33704]_  = ~A267 & \new_[33703]_ ;
  assign \new_[33708]_  = A301 & A300;
  assign \new_[33709]_  = ~A299 & \new_[33708]_ ;
  assign \new_[33710]_  = \new_[33709]_  & \new_[33704]_ ;
  assign \new_[33714]_  = ~A167 & A168;
  assign \new_[33715]_  = A169 & \new_[33714]_ ;
  assign \new_[33719]_  = A200 & A199;
  assign \new_[33720]_  = A166 & \new_[33719]_ ;
  assign \new_[33721]_  = \new_[33720]_  & \new_[33715]_ ;
  assign \new_[33725]_  = A298 & A268;
  assign \new_[33726]_  = ~A267 & \new_[33725]_ ;
  assign \new_[33730]_  = A302 & A300;
  assign \new_[33731]_  = ~A299 & \new_[33730]_ ;
  assign \new_[33732]_  = \new_[33731]_  & \new_[33726]_ ;
  assign \new_[33736]_  = ~A167 & A168;
  assign \new_[33737]_  = A169 & \new_[33736]_ ;
  assign \new_[33741]_  = A200 & A199;
  assign \new_[33742]_  = A166 & \new_[33741]_ ;
  assign \new_[33743]_  = \new_[33742]_  & \new_[33737]_ ;
  assign \new_[33747]_  = ~A298 & A268;
  assign \new_[33748]_  = ~A267 & \new_[33747]_ ;
  assign \new_[33752]_  = A301 & A300;
  assign \new_[33753]_  = A299 & \new_[33752]_ ;
  assign \new_[33754]_  = \new_[33753]_  & \new_[33748]_ ;
  assign \new_[33758]_  = ~A167 & A168;
  assign \new_[33759]_  = A169 & \new_[33758]_ ;
  assign \new_[33763]_  = A200 & A199;
  assign \new_[33764]_  = A166 & \new_[33763]_ ;
  assign \new_[33765]_  = \new_[33764]_  & \new_[33759]_ ;
  assign \new_[33769]_  = ~A298 & A268;
  assign \new_[33770]_  = ~A267 & \new_[33769]_ ;
  assign \new_[33774]_  = A302 & A300;
  assign \new_[33775]_  = A299 & \new_[33774]_ ;
  assign \new_[33776]_  = \new_[33775]_  & \new_[33770]_ ;
  assign \new_[33780]_  = ~A167 & A168;
  assign \new_[33781]_  = A169 & \new_[33780]_ ;
  assign \new_[33785]_  = A200 & A199;
  assign \new_[33786]_  = A166 & \new_[33785]_ ;
  assign \new_[33787]_  = \new_[33786]_  & \new_[33781]_ ;
  assign \new_[33791]_  = A298 & A269;
  assign \new_[33792]_  = ~A267 & \new_[33791]_ ;
  assign \new_[33796]_  = A301 & A300;
  assign \new_[33797]_  = ~A299 & \new_[33796]_ ;
  assign \new_[33798]_  = \new_[33797]_  & \new_[33792]_ ;
  assign \new_[33802]_  = ~A167 & A168;
  assign \new_[33803]_  = A169 & \new_[33802]_ ;
  assign \new_[33807]_  = A200 & A199;
  assign \new_[33808]_  = A166 & \new_[33807]_ ;
  assign \new_[33809]_  = \new_[33808]_  & \new_[33803]_ ;
  assign \new_[33813]_  = A298 & A269;
  assign \new_[33814]_  = ~A267 & \new_[33813]_ ;
  assign \new_[33818]_  = A302 & A300;
  assign \new_[33819]_  = ~A299 & \new_[33818]_ ;
  assign \new_[33820]_  = \new_[33819]_  & \new_[33814]_ ;
  assign \new_[33824]_  = ~A167 & A168;
  assign \new_[33825]_  = A169 & \new_[33824]_ ;
  assign \new_[33829]_  = A200 & A199;
  assign \new_[33830]_  = A166 & \new_[33829]_ ;
  assign \new_[33831]_  = \new_[33830]_  & \new_[33825]_ ;
  assign \new_[33835]_  = ~A298 & A269;
  assign \new_[33836]_  = ~A267 & \new_[33835]_ ;
  assign \new_[33840]_  = A301 & A300;
  assign \new_[33841]_  = A299 & \new_[33840]_ ;
  assign \new_[33842]_  = \new_[33841]_  & \new_[33836]_ ;
  assign \new_[33846]_  = ~A167 & A168;
  assign \new_[33847]_  = A169 & \new_[33846]_ ;
  assign \new_[33851]_  = A200 & A199;
  assign \new_[33852]_  = A166 & \new_[33851]_ ;
  assign \new_[33853]_  = \new_[33852]_  & \new_[33847]_ ;
  assign \new_[33857]_  = ~A298 & A269;
  assign \new_[33858]_  = ~A267 & \new_[33857]_ ;
  assign \new_[33862]_  = A302 & A300;
  assign \new_[33863]_  = A299 & \new_[33862]_ ;
  assign \new_[33864]_  = \new_[33863]_  & \new_[33858]_ ;
  assign \new_[33868]_  = ~A167 & A168;
  assign \new_[33869]_  = A169 & \new_[33868]_ ;
  assign \new_[33873]_  = A200 & A199;
  assign \new_[33874]_  = A166 & \new_[33873]_ ;
  assign \new_[33875]_  = \new_[33874]_  & \new_[33869]_ ;
  assign \new_[33879]_  = A298 & A266;
  assign \new_[33880]_  = A265 & \new_[33879]_ ;
  assign \new_[33884]_  = A301 & A300;
  assign \new_[33885]_  = ~A299 & \new_[33884]_ ;
  assign \new_[33886]_  = \new_[33885]_  & \new_[33880]_ ;
  assign \new_[33890]_  = ~A167 & A168;
  assign \new_[33891]_  = A169 & \new_[33890]_ ;
  assign \new_[33895]_  = A200 & A199;
  assign \new_[33896]_  = A166 & \new_[33895]_ ;
  assign \new_[33897]_  = \new_[33896]_  & \new_[33891]_ ;
  assign \new_[33901]_  = A298 & A266;
  assign \new_[33902]_  = A265 & \new_[33901]_ ;
  assign \new_[33906]_  = A302 & A300;
  assign \new_[33907]_  = ~A299 & \new_[33906]_ ;
  assign \new_[33908]_  = \new_[33907]_  & \new_[33902]_ ;
  assign \new_[33912]_  = ~A167 & A168;
  assign \new_[33913]_  = A169 & \new_[33912]_ ;
  assign \new_[33917]_  = A200 & A199;
  assign \new_[33918]_  = A166 & \new_[33917]_ ;
  assign \new_[33919]_  = \new_[33918]_  & \new_[33913]_ ;
  assign \new_[33923]_  = ~A298 & A266;
  assign \new_[33924]_  = A265 & \new_[33923]_ ;
  assign \new_[33928]_  = A301 & A300;
  assign \new_[33929]_  = A299 & \new_[33928]_ ;
  assign \new_[33930]_  = \new_[33929]_  & \new_[33924]_ ;
  assign \new_[33934]_  = ~A167 & A168;
  assign \new_[33935]_  = A169 & \new_[33934]_ ;
  assign \new_[33939]_  = A200 & A199;
  assign \new_[33940]_  = A166 & \new_[33939]_ ;
  assign \new_[33941]_  = \new_[33940]_  & \new_[33935]_ ;
  assign \new_[33945]_  = ~A298 & A266;
  assign \new_[33946]_  = A265 & \new_[33945]_ ;
  assign \new_[33950]_  = A302 & A300;
  assign \new_[33951]_  = A299 & \new_[33950]_ ;
  assign \new_[33952]_  = \new_[33951]_  & \new_[33946]_ ;
  assign \new_[33956]_  = ~A167 & A168;
  assign \new_[33957]_  = A169 & \new_[33956]_ ;
  assign \new_[33961]_  = A200 & A199;
  assign \new_[33962]_  = A166 & \new_[33961]_ ;
  assign \new_[33963]_  = \new_[33962]_  & \new_[33957]_ ;
  assign \new_[33967]_  = A298 & ~A266;
  assign \new_[33968]_  = ~A265 & \new_[33967]_ ;
  assign \new_[33972]_  = A301 & A300;
  assign \new_[33973]_  = ~A299 & \new_[33972]_ ;
  assign \new_[33974]_  = \new_[33973]_  & \new_[33968]_ ;
  assign \new_[33978]_  = ~A167 & A168;
  assign \new_[33979]_  = A169 & \new_[33978]_ ;
  assign \new_[33983]_  = A200 & A199;
  assign \new_[33984]_  = A166 & \new_[33983]_ ;
  assign \new_[33985]_  = \new_[33984]_  & \new_[33979]_ ;
  assign \new_[33989]_  = A298 & ~A266;
  assign \new_[33990]_  = ~A265 & \new_[33989]_ ;
  assign \new_[33994]_  = A302 & A300;
  assign \new_[33995]_  = ~A299 & \new_[33994]_ ;
  assign \new_[33996]_  = \new_[33995]_  & \new_[33990]_ ;
  assign \new_[34000]_  = ~A167 & A168;
  assign \new_[34001]_  = A169 & \new_[34000]_ ;
  assign \new_[34005]_  = A200 & A199;
  assign \new_[34006]_  = A166 & \new_[34005]_ ;
  assign \new_[34007]_  = \new_[34006]_  & \new_[34001]_ ;
  assign \new_[34011]_  = ~A298 & ~A266;
  assign \new_[34012]_  = ~A265 & \new_[34011]_ ;
  assign \new_[34016]_  = A301 & A300;
  assign \new_[34017]_  = A299 & \new_[34016]_ ;
  assign \new_[34018]_  = \new_[34017]_  & \new_[34012]_ ;
  assign \new_[34022]_  = ~A167 & A168;
  assign \new_[34023]_  = A169 & \new_[34022]_ ;
  assign \new_[34027]_  = A200 & A199;
  assign \new_[34028]_  = A166 & \new_[34027]_ ;
  assign \new_[34029]_  = \new_[34028]_  & \new_[34023]_ ;
  assign \new_[34033]_  = ~A298 & ~A266;
  assign \new_[34034]_  = ~A265 & \new_[34033]_ ;
  assign \new_[34038]_  = A302 & A300;
  assign \new_[34039]_  = A299 & \new_[34038]_ ;
  assign \new_[34040]_  = \new_[34039]_  & \new_[34034]_ ;
  assign \new_[34044]_  = ~A167 & A168;
  assign \new_[34045]_  = A169 & \new_[34044]_ ;
  assign \new_[34049]_  = ~A200 & ~A199;
  assign \new_[34050]_  = A166 & \new_[34049]_ ;
  assign \new_[34051]_  = \new_[34050]_  & \new_[34045]_ ;
  assign \new_[34055]_  = A298 & A268;
  assign \new_[34056]_  = ~A267 & \new_[34055]_ ;
  assign \new_[34060]_  = A301 & A300;
  assign \new_[34061]_  = ~A299 & \new_[34060]_ ;
  assign \new_[34062]_  = \new_[34061]_  & \new_[34056]_ ;
  assign \new_[34066]_  = ~A167 & A168;
  assign \new_[34067]_  = A169 & \new_[34066]_ ;
  assign \new_[34071]_  = ~A200 & ~A199;
  assign \new_[34072]_  = A166 & \new_[34071]_ ;
  assign \new_[34073]_  = \new_[34072]_  & \new_[34067]_ ;
  assign \new_[34077]_  = A298 & A268;
  assign \new_[34078]_  = ~A267 & \new_[34077]_ ;
  assign \new_[34082]_  = A302 & A300;
  assign \new_[34083]_  = ~A299 & \new_[34082]_ ;
  assign \new_[34084]_  = \new_[34083]_  & \new_[34078]_ ;
  assign \new_[34088]_  = ~A167 & A168;
  assign \new_[34089]_  = A169 & \new_[34088]_ ;
  assign \new_[34093]_  = ~A200 & ~A199;
  assign \new_[34094]_  = A166 & \new_[34093]_ ;
  assign \new_[34095]_  = \new_[34094]_  & \new_[34089]_ ;
  assign \new_[34099]_  = ~A298 & A268;
  assign \new_[34100]_  = ~A267 & \new_[34099]_ ;
  assign \new_[34104]_  = A301 & A300;
  assign \new_[34105]_  = A299 & \new_[34104]_ ;
  assign \new_[34106]_  = \new_[34105]_  & \new_[34100]_ ;
  assign \new_[34110]_  = ~A167 & A168;
  assign \new_[34111]_  = A169 & \new_[34110]_ ;
  assign \new_[34115]_  = ~A200 & ~A199;
  assign \new_[34116]_  = A166 & \new_[34115]_ ;
  assign \new_[34117]_  = \new_[34116]_  & \new_[34111]_ ;
  assign \new_[34121]_  = ~A298 & A268;
  assign \new_[34122]_  = ~A267 & \new_[34121]_ ;
  assign \new_[34126]_  = A302 & A300;
  assign \new_[34127]_  = A299 & \new_[34126]_ ;
  assign \new_[34128]_  = \new_[34127]_  & \new_[34122]_ ;
  assign \new_[34132]_  = ~A167 & A168;
  assign \new_[34133]_  = A169 & \new_[34132]_ ;
  assign \new_[34137]_  = ~A200 & ~A199;
  assign \new_[34138]_  = A166 & \new_[34137]_ ;
  assign \new_[34139]_  = \new_[34138]_  & \new_[34133]_ ;
  assign \new_[34143]_  = A298 & A269;
  assign \new_[34144]_  = ~A267 & \new_[34143]_ ;
  assign \new_[34148]_  = A301 & A300;
  assign \new_[34149]_  = ~A299 & \new_[34148]_ ;
  assign \new_[34150]_  = \new_[34149]_  & \new_[34144]_ ;
  assign \new_[34154]_  = ~A167 & A168;
  assign \new_[34155]_  = A169 & \new_[34154]_ ;
  assign \new_[34159]_  = ~A200 & ~A199;
  assign \new_[34160]_  = A166 & \new_[34159]_ ;
  assign \new_[34161]_  = \new_[34160]_  & \new_[34155]_ ;
  assign \new_[34165]_  = A298 & A269;
  assign \new_[34166]_  = ~A267 & \new_[34165]_ ;
  assign \new_[34170]_  = A302 & A300;
  assign \new_[34171]_  = ~A299 & \new_[34170]_ ;
  assign \new_[34172]_  = \new_[34171]_  & \new_[34166]_ ;
  assign \new_[34176]_  = ~A167 & A168;
  assign \new_[34177]_  = A169 & \new_[34176]_ ;
  assign \new_[34181]_  = ~A200 & ~A199;
  assign \new_[34182]_  = A166 & \new_[34181]_ ;
  assign \new_[34183]_  = \new_[34182]_  & \new_[34177]_ ;
  assign \new_[34187]_  = ~A298 & A269;
  assign \new_[34188]_  = ~A267 & \new_[34187]_ ;
  assign \new_[34192]_  = A301 & A300;
  assign \new_[34193]_  = A299 & \new_[34192]_ ;
  assign \new_[34194]_  = \new_[34193]_  & \new_[34188]_ ;
  assign \new_[34198]_  = ~A167 & A168;
  assign \new_[34199]_  = A169 & \new_[34198]_ ;
  assign \new_[34203]_  = ~A200 & ~A199;
  assign \new_[34204]_  = A166 & \new_[34203]_ ;
  assign \new_[34205]_  = \new_[34204]_  & \new_[34199]_ ;
  assign \new_[34209]_  = ~A298 & A269;
  assign \new_[34210]_  = ~A267 & \new_[34209]_ ;
  assign \new_[34214]_  = A302 & A300;
  assign \new_[34215]_  = A299 & \new_[34214]_ ;
  assign \new_[34216]_  = \new_[34215]_  & \new_[34210]_ ;
  assign \new_[34220]_  = ~A167 & A168;
  assign \new_[34221]_  = A169 & \new_[34220]_ ;
  assign \new_[34225]_  = ~A200 & ~A199;
  assign \new_[34226]_  = A166 & \new_[34225]_ ;
  assign \new_[34227]_  = \new_[34226]_  & \new_[34221]_ ;
  assign \new_[34231]_  = A298 & A266;
  assign \new_[34232]_  = A265 & \new_[34231]_ ;
  assign \new_[34236]_  = A301 & A300;
  assign \new_[34237]_  = ~A299 & \new_[34236]_ ;
  assign \new_[34238]_  = \new_[34237]_  & \new_[34232]_ ;
  assign \new_[34242]_  = ~A167 & A168;
  assign \new_[34243]_  = A169 & \new_[34242]_ ;
  assign \new_[34247]_  = ~A200 & ~A199;
  assign \new_[34248]_  = A166 & \new_[34247]_ ;
  assign \new_[34249]_  = \new_[34248]_  & \new_[34243]_ ;
  assign \new_[34253]_  = A298 & A266;
  assign \new_[34254]_  = A265 & \new_[34253]_ ;
  assign \new_[34258]_  = A302 & A300;
  assign \new_[34259]_  = ~A299 & \new_[34258]_ ;
  assign \new_[34260]_  = \new_[34259]_  & \new_[34254]_ ;
  assign \new_[34264]_  = ~A167 & A168;
  assign \new_[34265]_  = A169 & \new_[34264]_ ;
  assign \new_[34269]_  = ~A200 & ~A199;
  assign \new_[34270]_  = A166 & \new_[34269]_ ;
  assign \new_[34271]_  = \new_[34270]_  & \new_[34265]_ ;
  assign \new_[34275]_  = ~A298 & A266;
  assign \new_[34276]_  = A265 & \new_[34275]_ ;
  assign \new_[34280]_  = A301 & A300;
  assign \new_[34281]_  = A299 & \new_[34280]_ ;
  assign \new_[34282]_  = \new_[34281]_  & \new_[34276]_ ;
  assign \new_[34286]_  = ~A167 & A168;
  assign \new_[34287]_  = A169 & \new_[34286]_ ;
  assign \new_[34291]_  = ~A200 & ~A199;
  assign \new_[34292]_  = A166 & \new_[34291]_ ;
  assign \new_[34293]_  = \new_[34292]_  & \new_[34287]_ ;
  assign \new_[34297]_  = ~A298 & A266;
  assign \new_[34298]_  = A265 & \new_[34297]_ ;
  assign \new_[34302]_  = A302 & A300;
  assign \new_[34303]_  = A299 & \new_[34302]_ ;
  assign \new_[34304]_  = \new_[34303]_  & \new_[34298]_ ;
  assign \new_[34308]_  = ~A167 & A168;
  assign \new_[34309]_  = A169 & \new_[34308]_ ;
  assign \new_[34313]_  = ~A200 & ~A199;
  assign \new_[34314]_  = A166 & \new_[34313]_ ;
  assign \new_[34315]_  = \new_[34314]_  & \new_[34309]_ ;
  assign \new_[34319]_  = A298 & ~A266;
  assign \new_[34320]_  = ~A265 & \new_[34319]_ ;
  assign \new_[34324]_  = A301 & A300;
  assign \new_[34325]_  = ~A299 & \new_[34324]_ ;
  assign \new_[34326]_  = \new_[34325]_  & \new_[34320]_ ;
  assign \new_[34330]_  = ~A167 & A168;
  assign \new_[34331]_  = A169 & \new_[34330]_ ;
  assign \new_[34335]_  = ~A200 & ~A199;
  assign \new_[34336]_  = A166 & \new_[34335]_ ;
  assign \new_[34337]_  = \new_[34336]_  & \new_[34331]_ ;
  assign \new_[34341]_  = A298 & ~A266;
  assign \new_[34342]_  = ~A265 & \new_[34341]_ ;
  assign \new_[34346]_  = A302 & A300;
  assign \new_[34347]_  = ~A299 & \new_[34346]_ ;
  assign \new_[34348]_  = \new_[34347]_  & \new_[34342]_ ;
  assign \new_[34352]_  = ~A167 & A168;
  assign \new_[34353]_  = A169 & \new_[34352]_ ;
  assign \new_[34357]_  = ~A200 & ~A199;
  assign \new_[34358]_  = A166 & \new_[34357]_ ;
  assign \new_[34359]_  = \new_[34358]_  & \new_[34353]_ ;
  assign \new_[34363]_  = ~A298 & ~A266;
  assign \new_[34364]_  = ~A265 & \new_[34363]_ ;
  assign \new_[34368]_  = A301 & A300;
  assign \new_[34369]_  = A299 & \new_[34368]_ ;
  assign \new_[34370]_  = \new_[34369]_  & \new_[34364]_ ;
  assign \new_[34374]_  = ~A167 & A168;
  assign \new_[34375]_  = A169 & \new_[34374]_ ;
  assign \new_[34379]_  = ~A200 & ~A199;
  assign \new_[34380]_  = A166 & \new_[34379]_ ;
  assign \new_[34381]_  = \new_[34380]_  & \new_[34375]_ ;
  assign \new_[34385]_  = ~A298 & ~A266;
  assign \new_[34386]_  = ~A265 & \new_[34385]_ ;
  assign \new_[34390]_  = A302 & A300;
  assign \new_[34391]_  = A299 & \new_[34390]_ ;
  assign \new_[34392]_  = \new_[34391]_  & \new_[34386]_ ;
  assign \new_[34396]_  = A201 & ~A168;
  assign \new_[34397]_  = A169 & \new_[34396]_ ;
  assign \new_[34401]_  = ~A265 & ~A203;
  assign \new_[34402]_  = ~A202 & \new_[34401]_ ;
  assign \new_[34403]_  = \new_[34402]_  & \new_[34397]_ ;
  assign \new_[34407]_  = A268 & A267;
  assign \new_[34408]_  = A266 & \new_[34407]_ ;
  assign \new_[34412]_  = ~A302 & ~A301;
  assign \new_[34413]_  = A300 & \new_[34412]_ ;
  assign \new_[34414]_  = \new_[34413]_  & \new_[34408]_ ;
  assign \new_[34418]_  = A201 & ~A168;
  assign \new_[34419]_  = A169 & \new_[34418]_ ;
  assign \new_[34423]_  = ~A265 & ~A203;
  assign \new_[34424]_  = ~A202 & \new_[34423]_ ;
  assign \new_[34425]_  = \new_[34424]_  & \new_[34419]_ ;
  assign \new_[34429]_  = A269 & A267;
  assign \new_[34430]_  = A266 & \new_[34429]_ ;
  assign \new_[34434]_  = ~A302 & ~A301;
  assign \new_[34435]_  = A300 & \new_[34434]_ ;
  assign \new_[34436]_  = \new_[34435]_  & \new_[34430]_ ;
  assign \new_[34440]_  = A201 & ~A168;
  assign \new_[34441]_  = A169 & \new_[34440]_ ;
  assign \new_[34445]_  = ~A265 & ~A203;
  assign \new_[34446]_  = ~A202 & \new_[34445]_ ;
  assign \new_[34447]_  = \new_[34446]_  & \new_[34441]_ ;
  assign \new_[34451]_  = ~A268 & ~A267;
  assign \new_[34452]_  = A266 & \new_[34451]_ ;
  assign \new_[34456]_  = A301 & ~A300;
  assign \new_[34457]_  = ~A269 & \new_[34456]_ ;
  assign \new_[34458]_  = \new_[34457]_  & \new_[34452]_ ;
  assign \new_[34462]_  = A201 & ~A168;
  assign \new_[34463]_  = A169 & \new_[34462]_ ;
  assign \new_[34467]_  = ~A265 & ~A203;
  assign \new_[34468]_  = ~A202 & \new_[34467]_ ;
  assign \new_[34469]_  = \new_[34468]_  & \new_[34463]_ ;
  assign \new_[34473]_  = ~A268 & ~A267;
  assign \new_[34474]_  = A266 & \new_[34473]_ ;
  assign \new_[34478]_  = A302 & ~A300;
  assign \new_[34479]_  = ~A269 & \new_[34478]_ ;
  assign \new_[34480]_  = \new_[34479]_  & \new_[34474]_ ;
  assign \new_[34484]_  = A201 & ~A168;
  assign \new_[34485]_  = A169 & \new_[34484]_ ;
  assign \new_[34489]_  = ~A265 & ~A203;
  assign \new_[34490]_  = ~A202 & \new_[34489]_ ;
  assign \new_[34491]_  = \new_[34490]_  & \new_[34485]_ ;
  assign \new_[34495]_  = ~A268 & ~A267;
  assign \new_[34496]_  = A266 & \new_[34495]_ ;
  assign \new_[34500]_  = A299 & A298;
  assign \new_[34501]_  = ~A269 & \new_[34500]_ ;
  assign \new_[34502]_  = \new_[34501]_  & \new_[34496]_ ;
  assign \new_[34506]_  = A201 & ~A168;
  assign \new_[34507]_  = A169 & \new_[34506]_ ;
  assign \new_[34511]_  = ~A265 & ~A203;
  assign \new_[34512]_  = ~A202 & \new_[34511]_ ;
  assign \new_[34513]_  = \new_[34512]_  & \new_[34507]_ ;
  assign \new_[34517]_  = ~A268 & ~A267;
  assign \new_[34518]_  = A266 & \new_[34517]_ ;
  assign \new_[34522]_  = ~A299 & ~A298;
  assign \new_[34523]_  = ~A269 & \new_[34522]_ ;
  assign \new_[34524]_  = \new_[34523]_  & \new_[34518]_ ;
  assign \new_[34528]_  = A201 & ~A168;
  assign \new_[34529]_  = A169 & \new_[34528]_ ;
  assign \new_[34533]_  = A265 & ~A203;
  assign \new_[34534]_  = ~A202 & \new_[34533]_ ;
  assign \new_[34535]_  = \new_[34534]_  & \new_[34529]_ ;
  assign \new_[34539]_  = A268 & A267;
  assign \new_[34540]_  = ~A266 & \new_[34539]_ ;
  assign \new_[34544]_  = ~A302 & ~A301;
  assign \new_[34545]_  = A300 & \new_[34544]_ ;
  assign \new_[34546]_  = \new_[34545]_  & \new_[34540]_ ;
  assign \new_[34550]_  = A201 & ~A168;
  assign \new_[34551]_  = A169 & \new_[34550]_ ;
  assign \new_[34555]_  = A265 & ~A203;
  assign \new_[34556]_  = ~A202 & \new_[34555]_ ;
  assign \new_[34557]_  = \new_[34556]_  & \new_[34551]_ ;
  assign \new_[34561]_  = A269 & A267;
  assign \new_[34562]_  = ~A266 & \new_[34561]_ ;
  assign \new_[34566]_  = ~A302 & ~A301;
  assign \new_[34567]_  = A300 & \new_[34566]_ ;
  assign \new_[34568]_  = \new_[34567]_  & \new_[34562]_ ;
  assign \new_[34572]_  = A201 & ~A168;
  assign \new_[34573]_  = A169 & \new_[34572]_ ;
  assign \new_[34577]_  = A265 & ~A203;
  assign \new_[34578]_  = ~A202 & \new_[34577]_ ;
  assign \new_[34579]_  = \new_[34578]_  & \new_[34573]_ ;
  assign \new_[34583]_  = ~A268 & ~A267;
  assign \new_[34584]_  = ~A266 & \new_[34583]_ ;
  assign \new_[34588]_  = A301 & ~A300;
  assign \new_[34589]_  = ~A269 & \new_[34588]_ ;
  assign \new_[34590]_  = \new_[34589]_  & \new_[34584]_ ;
  assign \new_[34594]_  = A201 & ~A168;
  assign \new_[34595]_  = A169 & \new_[34594]_ ;
  assign \new_[34599]_  = A265 & ~A203;
  assign \new_[34600]_  = ~A202 & \new_[34599]_ ;
  assign \new_[34601]_  = \new_[34600]_  & \new_[34595]_ ;
  assign \new_[34605]_  = ~A268 & ~A267;
  assign \new_[34606]_  = ~A266 & \new_[34605]_ ;
  assign \new_[34610]_  = A302 & ~A300;
  assign \new_[34611]_  = ~A269 & \new_[34610]_ ;
  assign \new_[34612]_  = \new_[34611]_  & \new_[34606]_ ;
  assign \new_[34616]_  = A201 & ~A168;
  assign \new_[34617]_  = A169 & \new_[34616]_ ;
  assign \new_[34621]_  = A265 & ~A203;
  assign \new_[34622]_  = ~A202 & \new_[34621]_ ;
  assign \new_[34623]_  = \new_[34622]_  & \new_[34617]_ ;
  assign \new_[34627]_  = ~A268 & ~A267;
  assign \new_[34628]_  = ~A266 & \new_[34627]_ ;
  assign \new_[34632]_  = A299 & A298;
  assign \new_[34633]_  = ~A269 & \new_[34632]_ ;
  assign \new_[34634]_  = \new_[34633]_  & \new_[34628]_ ;
  assign \new_[34638]_  = A201 & ~A168;
  assign \new_[34639]_  = A169 & \new_[34638]_ ;
  assign \new_[34643]_  = A265 & ~A203;
  assign \new_[34644]_  = ~A202 & \new_[34643]_ ;
  assign \new_[34645]_  = \new_[34644]_  & \new_[34639]_ ;
  assign \new_[34649]_  = ~A268 & ~A267;
  assign \new_[34650]_  = ~A266 & \new_[34649]_ ;
  assign \new_[34654]_  = ~A299 & ~A298;
  assign \new_[34655]_  = ~A269 & \new_[34654]_ ;
  assign \new_[34656]_  = \new_[34655]_  & \new_[34650]_ ;
  assign \new_[34660]_  = ~A201 & ~A168;
  assign \new_[34661]_  = A169 & \new_[34660]_ ;
  assign \new_[34665]_  = A266 & ~A265;
  assign \new_[34666]_  = A202 & \new_[34665]_ ;
  assign \new_[34667]_  = \new_[34666]_  & \new_[34661]_ ;
  assign \new_[34671]_  = ~A269 & ~A268;
  assign \new_[34672]_  = ~A267 & \new_[34671]_ ;
  assign \new_[34676]_  = ~A302 & ~A301;
  assign \new_[34677]_  = A300 & \new_[34676]_ ;
  assign \new_[34678]_  = \new_[34677]_  & \new_[34672]_ ;
  assign \new_[34682]_  = ~A201 & ~A168;
  assign \new_[34683]_  = A169 & \new_[34682]_ ;
  assign \new_[34687]_  = ~A266 & A265;
  assign \new_[34688]_  = A202 & \new_[34687]_ ;
  assign \new_[34689]_  = \new_[34688]_  & \new_[34683]_ ;
  assign \new_[34693]_  = ~A269 & ~A268;
  assign \new_[34694]_  = ~A267 & \new_[34693]_ ;
  assign \new_[34698]_  = ~A302 & ~A301;
  assign \new_[34699]_  = A300 & \new_[34698]_ ;
  assign \new_[34700]_  = \new_[34699]_  & \new_[34694]_ ;
  assign \new_[34704]_  = ~A201 & ~A168;
  assign \new_[34705]_  = A169 & \new_[34704]_ ;
  assign \new_[34709]_  = A266 & ~A265;
  assign \new_[34710]_  = A203 & \new_[34709]_ ;
  assign \new_[34711]_  = \new_[34710]_  & \new_[34705]_ ;
  assign \new_[34715]_  = ~A269 & ~A268;
  assign \new_[34716]_  = ~A267 & \new_[34715]_ ;
  assign \new_[34720]_  = ~A302 & ~A301;
  assign \new_[34721]_  = A300 & \new_[34720]_ ;
  assign \new_[34722]_  = \new_[34721]_  & \new_[34716]_ ;
  assign \new_[34726]_  = ~A201 & ~A168;
  assign \new_[34727]_  = A169 & \new_[34726]_ ;
  assign \new_[34731]_  = ~A266 & A265;
  assign \new_[34732]_  = A203 & \new_[34731]_ ;
  assign \new_[34733]_  = \new_[34732]_  & \new_[34727]_ ;
  assign \new_[34737]_  = ~A269 & ~A268;
  assign \new_[34738]_  = ~A267 & \new_[34737]_ ;
  assign \new_[34742]_  = ~A302 & ~A301;
  assign \new_[34743]_  = A300 & \new_[34742]_ ;
  assign \new_[34744]_  = \new_[34743]_  & \new_[34738]_ ;
  assign \new_[34748]_  = A199 & ~A168;
  assign \new_[34749]_  = A169 & \new_[34748]_ ;
  assign \new_[34753]_  = A266 & ~A265;
  assign \new_[34754]_  = A200 & \new_[34753]_ ;
  assign \new_[34755]_  = \new_[34754]_  & \new_[34749]_ ;
  assign \new_[34759]_  = ~A269 & ~A268;
  assign \new_[34760]_  = ~A267 & \new_[34759]_ ;
  assign \new_[34764]_  = ~A302 & ~A301;
  assign \new_[34765]_  = A300 & \new_[34764]_ ;
  assign \new_[34766]_  = \new_[34765]_  & \new_[34760]_ ;
  assign \new_[34770]_  = A199 & ~A168;
  assign \new_[34771]_  = A169 & \new_[34770]_ ;
  assign \new_[34775]_  = ~A266 & A265;
  assign \new_[34776]_  = A200 & \new_[34775]_ ;
  assign \new_[34777]_  = \new_[34776]_  & \new_[34771]_ ;
  assign \new_[34781]_  = ~A269 & ~A268;
  assign \new_[34782]_  = ~A267 & \new_[34781]_ ;
  assign \new_[34786]_  = ~A302 & ~A301;
  assign \new_[34787]_  = A300 & \new_[34786]_ ;
  assign \new_[34788]_  = \new_[34787]_  & \new_[34782]_ ;
  assign \new_[34792]_  = ~A199 & ~A168;
  assign \new_[34793]_  = A169 & \new_[34792]_ ;
  assign \new_[34797]_  = A202 & A201;
  assign \new_[34798]_  = A200 & \new_[34797]_ ;
  assign \new_[34799]_  = \new_[34798]_  & \new_[34793]_ ;
  assign \new_[34803]_  = A298 & A268;
  assign \new_[34804]_  = ~A267 & \new_[34803]_ ;
  assign \new_[34808]_  = A301 & A300;
  assign \new_[34809]_  = ~A299 & \new_[34808]_ ;
  assign \new_[34810]_  = \new_[34809]_  & \new_[34804]_ ;
  assign \new_[34814]_  = ~A199 & ~A168;
  assign \new_[34815]_  = A169 & \new_[34814]_ ;
  assign \new_[34819]_  = A202 & A201;
  assign \new_[34820]_  = A200 & \new_[34819]_ ;
  assign \new_[34821]_  = \new_[34820]_  & \new_[34815]_ ;
  assign \new_[34825]_  = A298 & A268;
  assign \new_[34826]_  = ~A267 & \new_[34825]_ ;
  assign \new_[34830]_  = A302 & A300;
  assign \new_[34831]_  = ~A299 & \new_[34830]_ ;
  assign \new_[34832]_  = \new_[34831]_  & \new_[34826]_ ;
  assign \new_[34836]_  = ~A199 & ~A168;
  assign \new_[34837]_  = A169 & \new_[34836]_ ;
  assign \new_[34841]_  = A202 & A201;
  assign \new_[34842]_  = A200 & \new_[34841]_ ;
  assign \new_[34843]_  = \new_[34842]_  & \new_[34837]_ ;
  assign \new_[34847]_  = ~A298 & A268;
  assign \new_[34848]_  = ~A267 & \new_[34847]_ ;
  assign \new_[34852]_  = A301 & A300;
  assign \new_[34853]_  = A299 & \new_[34852]_ ;
  assign \new_[34854]_  = \new_[34853]_  & \new_[34848]_ ;
  assign \new_[34858]_  = ~A199 & ~A168;
  assign \new_[34859]_  = A169 & \new_[34858]_ ;
  assign \new_[34863]_  = A202 & A201;
  assign \new_[34864]_  = A200 & \new_[34863]_ ;
  assign \new_[34865]_  = \new_[34864]_  & \new_[34859]_ ;
  assign \new_[34869]_  = ~A298 & A268;
  assign \new_[34870]_  = ~A267 & \new_[34869]_ ;
  assign \new_[34874]_  = A302 & A300;
  assign \new_[34875]_  = A299 & \new_[34874]_ ;
  assign \new_[34876]_  = \new_[34875]_  & \new_[34870]_ ;
  assign \new_[34880]_  = ~A199 & ~A168;
  assign \new_[34881]_  = A169 & \new_[34880]_ ;
  assign \new_[34885]_  = A202 & A201;
  assign \new_[34886]_  = A200 & \new_[34885]_ ;
  assign \new_[34887]_  = \new_[34886]_  & \new_[34881]_ ;
  assign \new_[34891]_  = A298 & A269;
  assign \new_[34892]_  = ~A267 & \new_[34891]_ ;
  assign \new_[34896]_  = A301 & A300;
  assign \new_[34897]_  = ~A299 & \new_[34896]_ ;
  assign \new_[34898]_  = \new_[34897]_  & \new_[34892]_ ;
  assign \new_[34902]_  = ~A199 & ~A168;
  assign \new_[34903]_  = A169 & \new_[34902]_ ;
  assign \new_[34907]_  = A202 & A201;
  assign \new_[34908]_  = A200 & \new_[34907]_ ;
  assign \new_[34909]_  = \new_[34908]_  & \new_[34903]_ ;
  assign \new_[34913]_  = A298 & A269;
  assign \new_[34914]_  = ~A267 & \new_[34913]_ ;
  assign \new_[34918]_  = A302 & A300;
  assign \new_[34919]_  = ~A299 & \new_[34918]_ ;
  assign \new_[34920]_  = \new_[34919]_  & \new_[34914]_ ;
  assign \new_[34924]_  = ~A199 & ~A168;
  assign \new_[34925]_  = A169 & \new_[34924]_ ;
  assign \new_[34929]_  = A202 & A201;
  assign \new_[34930]_  = A200 & \new_[34929]_ ;
  assign \new_[34931]_  = \new_[34930]_  & \new_[34925]_ ;
  assign \new_[34935]_  = ~A298 & A269;
  assign \new_[34936]_  = ~A267 & \new_[34935]_ ;
  assign \new_[34940]_  = A301 & A300;
  assign \new_[34941]_  = A299 & \new_[34940]_ ;
  assign \new_[34942]_  = \new_[34941]_  & \new_[34936]_ ;
  assign \new_[34946]_  = ~A199 & ~A168;
  assign \new_[34947]_  = A169 & \new_[34946]_ ;
  assign \new_[34951]_  = A202 & A201;
  assign \new_[34952]_  = A200 & \new_[34951]_ ;
  assign \new_[34953]_  = \new_[34952]_  & \new_[34947]_ ;
  assign \new_[34957]_  = ~A298 & A269;
  assign \new_[34958]_  = ~A267 & \new_[34957]_ ;
  assign \new_[34962]_  = A302 & A300;
  assign \new_[34963]_  = A299 & \new_[34962]_ ;
  assign \new_[34964]_  = \new_[34963]_  & \new_[34958]_ ;
  assign \new_[34968]_  = ~A199 & ~A168;
  assign \new_[34969]_  = A169 & \new_[34968]_ ;
  assign \new_[34973]_  = A202 & A201;
  assign \new_[34974]_  = A200 & \new_[34973]_ ;
  assign \new_[34975]_  = \new_[34974]_  & \new_[34969]_ ;
  assign \new_[34979]_  = A298 & A266;
  assign \new_[34980]_  = A265 & \new_[34979]_ ;
  assign \new_[34984]_  = A301 & A300;
  assign \new_[34985]_  = ~A299 & \new_[34984]_ ;
  assign \new_[34986]_  = \new_[34985]_  & \new_[34980]_ ;
  assign \new_[34990]_  = ~A199 & ~A168;
  assign \new_[34991]_  = A169 & \new_[34990]_ ;
  assign \new_[34995]_  = A202 & A201;
  assign \new_[34996]_  = A200 & \new_[34995]_ ;
  assign \new_[34997]_  = \new_[34996]_  & \new_[34991]_ ;
  assign \new_[35001]_  = A298 & A266;
  assign \new_[35002]_  = A265 & \new_[35001]_ ;
  assign \new_[35006]_  = A302 & A300;
  assign \new_[35007]_  = ~A299 & \new_[35006]_ ;
  assign \new_[35008]_  = \new_[35007]_  & \new_[35002]_ ;
  assign \new_[35012]_  = ~A199 & ~A168;
  assign \new_[35013]_  = A169 & \new_[35012]_ ;
  assign \new_[35017]_  = A202 & A201;
  assign \new_[35018]_  = A200 & \new_[35017]_ ;
  assign \new_[35019]_  = \new_[35018]_  & \new_[35013]_ ;
  assign \new_[35023]_  = ~A298 & A266;
  assign \new_[35024]_  = A265 & \new_[35023]_ ;
  assign \new_[35028]_  = A301 & A300;
  assign \new_[35029]_  = A299 & \new_[35028]_ ;
  assign \new_[35030]_  = \new_[35029]_  & \new_[35024]_ ;
  assign \new_[35034]_  = ~A199 & ~A168;
  assign \new_[35035]_  = A169 & \new_[35034]_ ;
  assign \new_[35039]_  = A202 & A201;
  assign \new_[35040]_  = A200 & \new_[35039]_ ;
  assign \new_[35041]_  = \new_[35040]_  & \new_[35035]_ ;
  assign \new_[35045]_  = ~A298 & A266;
  assign \new_[35046]_  = A265 & \new_[35045]_ ;
  assign \new_[35050]_  = A302 & A300;
  assign \new_[35051]_  = A299 & \new_[35050]_ ;
  assign \new_[35052]_  = \new_[35051]_  & \new_[35046]_ ;
  assign \new_[35056]_  = ~A199 & ~A168;
  assign \new_[35057]_  = A169 & \new_[35056]_ ;
  assign \new_[35061]_  = A202 & A201;
  assign \new_[35062]_  = A200 & \new_[35061]_ ;
  assign \new_[35063]_  = \new_[35062]_  & \new_[35057]_ ;
  assign \new_[35067]_  = A298 & ~A266;
  assign \new_[35068]_  = ~A265 & \new_[35067]_ ;
  assign \new_[35072]_  = A301 & A300;
  assign \new_[35073]_  = ~A299 & \new_[35072]_ ;
  assign \new_[35074]_  = \new_[35073]_  & \new_[35068]_ ;
  assign \new_[35078]_  = ~A199 & ~A168;
  assign \new_[35079]_  = A169 & \new_[35078]_ ;
  assign \new_[35083]_  = A202 & A201;
  assign \new_[35084]_  = A200 & \new_[35083]_ ;
  assign \new_[35085]_  = \new_[35084]_  & \new_[35079]_ ;
  assign \new_[35089]_  = A298 & ~A266;
  assign \new_[35090]_  = ~A265 & \new_[35089]_ ;
  assign \new_[35094]_  = A302 & A300;
  assign \new_[35095]_  = ~A299 & \new_[35094]_ ;
  assign \new_[35096]_  = \new_[35095]_  & \new_[35090]_ ;
  assign \new_[35100]_  = ~A199 & ~A168;
  assign \new_[35101]_  = A169 & \new_[35100]_ ;
  assign \new_[35105]_  = A202 & A201;
  assign \new_[35106]_  = A200 & \new_[35105]_ ;
  assign \new_[35107]_  = \new_[35106]_  & \new_[35101]_ ;
  assign \new_[35111]_  = ~A298 & ~A266;
  assign \new_[35112]_  = ~A265 & \new_[35111]_ ;
  assign \new_[35116]_  = A301 & A300;
  assign \new_[35117]_  = A299 & \new_[35116]_ ;
  assign \new_[35118]_  = \new_[35117]_  & \new_[35112]_ ;
  assign \new_[35122]_  = ~A199 & ~A168;
  assign \new_[35123]_  = A169 & \new_[35122]_ ;
  assign \new_[35127]_  = A202 & A201;
  assign \new_[35128]_  = A200 & \new_[35127]_ ;
  assign \new_[35129]_  = \new_[35128]_  & \new_[35123]_ ;
  assign \new_[35133]_  = ~A298 & ~A266;
  assign \new_[35134]_  = ~A265 & \new_[35133]_ ;
  assign \new_[35138]_  = A302 & A300;
  assign \new_[35139]_  = A299 & \new_[35138]_ ;
  assign \new_[35140]_  = \new_[35139]_  & \new_[35134]_ ;
  assign \new_[35144]_  = ~A199 & ~A168;
  assign \new_[35145]_  = A169 & \new_[35144]_ ;
  assign \new_[35149]_  = A203 & A201;
  assign \new_[35150]_  = A200 & \new_[35149]_ ;
  assign \new_[35151]_  = \new_[35150]_  & \new_[35145]_ ;
  assign \new_[35155]_  = A298 & A268;
  assign \new_[35156]_  = ~A267 & \new_[35155]_ ;
  assign \new_[35160]_  = A301 & A300;
  assign \new_[35161]_  = ~A299 & \new_[35160]_ ;
  assign \new_[35162]_  = \new_[35161]_  & \new_[35156]_ ;
  assign \new_[35166]_  = ~A199 & ~A168;
  assign \new_[35167]_  = A169 & \new_[35166]_ ;
  assign \new_[35171]_  = A203 & A201;
  assign \new_[35172]_  = A200 & \new_[35171]_ ;
  assign \new_[35173]_  = \new_[35172]_  & \new_[35167]_ ;
  assign \new_[35177]_  = A298 & A268;
  assign \new_[35178]_  = ~A267 & \new_[35177]_ ;
  assign \new_[35182]_  = A302 & A300;
  assign \new_[35183]_  = ~A299 & \new_[35182]_ ;
  assign \new_[35184]_  = \new_[35183]_  & \new_[35178]_ ;
  assign \new_[35188]_  = ~A199 & ~A168;
  assign \new_[35189]_  = A169 & \new_[35188]_ ;
  assign \new_[35193]_  = A203 & A201;
  assign \new_[35194]_  = A200 & \new_[35193]_ ;
  assign \new_[35195]_  = \new_[35194]_  & \new_[35189]_ ;
  assign \new_[35199]_  = ~A298 & A268;
  assign \new_[35200]_  = ~A267 & \new_[35199]_ ;
  assign \new_[35204]_  = A301 & A300;
  assign \new_[35205]_  = A299 & \new_[35204]_ ;
  assign \new_[35206]_  = \new_[35205]_  & \new_[35200]_ ;
  assign \new_[35210]_  = ~A199 & ~A168;
  assign \new_[35211]_  = A169 & \new_[35210]_ ;
  assign \new_[35215]_  = A203 & A201;
  assign \new_[35216]_  = A200 & \new_[35215]_ ;
  assign \new_[35217]_  = \new_[35216]_  & \new_[35211]_ ;
  assign \new_[35221]_  = ~A298 & A268;
  assign \new_[35222]_  = ~A267 & \new_[35221]_ ;
  assign \new_[35226]_  = A302 & A300;
  assign \new_[35227]_  = A299 & \new_[35226]_ ;
  assign \new_[35228]_  = \new_[35227]_  & \new_[35222]_ ;
  assign \new_[35232]_  = ~A199 & ~A168;
  assign \new_[35233]_  = A169 & \new_[35232]_ ;
  assign \new_[35237]_  = A203 & A201;
  assign \new_[35238]_  = A200 & \new_[35237]_ ;
  assign \new_[35239]_  = \new_[35238]_  & \new_[35233]_ ;
  assign \new_[35243]_  = A298 & A269;
  assign \new_[35244]_  = ~A267 & \new_[35243]_ ;
  assign \new_[35248]_  = A301 & A300;
  assign \new_[35249]_  = ~A299 & \new_[35248]_ ;
  assign \new_[35250]_  = \new_[35249]_  & \new_[35244]_ ;
  assign \new_[35254]_  = ~A199 & ~A168;
  assign \new_[35255]_  = A169 & \new_[35254]_ ;
  assign \new_[35259]_  = A203 & A201;
  assign \new_[35260]_  = A200 & \new_[35259]_ ;
  assign \new_[35261]_  = \new_[35260]_  & \new_[35255]_ ;
  assign \new_[35265]_  = A298 & A269;
  assign \new_[35266]_  = ~A267 & \new_[35265]_ ;
  assign \new_[35270]_  = A302 & A300;
  assign \new_[35271]_  = ~A299 & \new_[35270]_ ;
  assign \new_[35272]_  = \new_[35271]_  & \new_[35266]_ ;
  assign \new_[35276]_  = ~A199 & ~A168;
  assign \new_[35277]_  = A169 & \new_[35276]_ ;
  assign \new_[35281]_  = A203 & A201;
  assign \new_[35282]_  = A200 & \new_[35281]_ ;
  assign \new_[35283]_  = \new_[35282]_  & \new_[35277]_ ;
  assign \new_[35287]_  = ~A298 & A269;
  assign \new_[35288]_  = ~A267 & \new_[35287]_ ;
  assign \new_[35292]_  = A301 & A300;
  assign \new_[35293]_  = A299 & \new_[35292]_ ;
  assign \new_[35294]_  = \new_[35293]_  & \new_[35288]_ ;
  assign \new_[35298]_  = ~A199 & ~A168;
  assign \new_[35299]_  = A169 & \new_[35298]_ ;
  assign \new_[35303]_  = A203 & A201;
  assign \new_[35304]_  = A200 & \new_[35303]_ ;
  assign \new_[35305]_  = \new_[35304]_  & \new_[35299]_ ;
  assign \new_[35309]_  = ~A298 & A269;
  assign \new_[35310]_  = ~A267 & \new_[35309]_ ;
  assign \new_[35314]_  = A302 & A300;
  assign \new_[35315]_  = A299 & \new_[35314]_ ;
  assign \new_[35316]_  = \new_[35315]_  & \new_[35310]_ ;
  assign \new_[35320]_  = ~A199 & ~A168;
  assign \new_[35321]_  = A169 & \new_[35320]_ ;
  assign \new_[35325]_  = A203 & A201;
  assign \new_[35326]_  = A200 & \new_[35325]_ ;
  assign \new_[35327]_  = \new_[35326]_  & \new_[35321]_ ;
  assign \new_[35331]_  = A298 & A266;
  assign \new_[35332]_  = A265 & \new_[35331]_ ;
  assign \new_[35336]_  = A301 & A300;
  assign \new_[35337]_  = ~A299 & \new_[35336]_ ;
  assign \new_[35338]_  = \new_[35337]_  & \new_[35332]_ ;
  assign \new_[35342]_  = ~A199 & ~A168;
  assign \new_[35343]_  = A169 & \new_[35342]_ ;
  assign \new_[35347]_  = A203 & A201;
  assign \new_[35348]_  = A200 & \new_[35347]_ ;
  assign \new_[35349]_  = \new_[35348]_  & \new_[35343]_ ;
  assign \new_[35353]_  = A298 & A266;
  assign \new_[35354]_  = A265 & \new_[35353]_ ;
  assign \new_[35358]_  = A302 & A300;
  assign \new_[35359]_  = ~A299 & \new_[35358]_ ;
  assign \new_[35360]_  = \new_[35359]_  & \new_[35354]_ ;
  assign \new_[35364]_  = ~A199 & ~A168;
  assign \new_[35365]_  = A169 & \new_[35364]_ ;
  assign \new_[35369]_  = A203 & A201;
  assign \new_[35370]_  = A200 & \new_[35369]_ ;
  assign \new_[35371]_  = \new_[35370]_  & \new_[35365]_ ;
  assign \new_[35375]_  = ~A298 & A266;
  assign \new_[35376]_  = A265 & \new_[35375]_ ;
  assign \new_[35380]_  = A301 & A300;
  assign \new_[35381]_  = A299 & \new_[35380]_ ;
  assign \new_[35382]_  = \new_[35381]_  & \new_[35376]_ ;
  assign \new_[35386]_  = ~A199 & ~A168;
  assign \new_[35387]_  = A169 & \new_[35386]_ ;
  assign \new_[35391]_  = A203 & A201;
  assign \new_[35392]_  = A200 & \new_[35391]_ ;
  assign \new_[35393]_  = \new_[35392]_  & \new_[35387]_ ;
  assign \new_[35397]_  = ~A298 & A266;
  assign \new_[35398]_  = A265 & \new_[35397]_ ;
  assign \new_[35402]_  = A302 & A300;
  assign \new_[35403]_  = A299 & \new_[35402]_ ;
  assign \new_[35404]_  = \new_[35403]_  & \new_[35398]_ ;
  assign \new_[35408]_  = ~A199 & ~A168;
  assign \new_[35409]_  = A169 & \new_[35408]_ ;
  assign \new_[35413]_  = A203 & A201;
  assign \new_[35414]_  = A200 & \new_[35413]_ ;
  assign \new_[35415]_  = \new_[35414]_  & \new_[35409]_ ;
  assign \new_[35419]_  = A298 & ~A266;
  assign \new_[35420]_  = ~A265 & \new_[35419]_ ;
  assign \new_[35424]_  = A301 & A300;
  assign \new_[35425]_  = ~A299 & \new_[35424]_ ;
  assign \new_[35426]_  = \new_[35425]_  & \new_[35420]_ ;
  assign \new_[35430]_  = ~A199 & ~A168;
  assign \new_[35431]_  = A169 & \new_[35430]_ ;
  assign \new_[35435]_  = A203 & A201;
  assign \new_[35436]_  = A200 & \new_[35435]_ ;
  assign \new_[35437]_  = \new_[35436]_  & \new_[35431]_ ;
  assign \new_[35441]_  = A298 & ~A266;
  assign \new_[35442]_  = ~A265 & \new_[35441]_ ;
  assign \new_[35446]_  = A302 & A300;
  assign \new_[35447]_  = ~A299 & \new_[35446]_ ;
  assign \new_[35448]_  = \new_[35447]_  & \new_[35442]_ ;
  assign \new_[35452]_  = ~A199 & ~A168;
  assign \new_[35453]_  = A169 & \new_[35452]_ ;
  assign \new_[35457]_  = A203 & A201;
  assign \new_[35458]_  = A200 & \new_[35457]_ ;
  assign \new_[35459]_  = \new_[35458]_  & \new_[35453]_ ;
  assign \new_[35463]_  = ~A298 & ~A266;
  assign \new_[35464]_  = ~A265 & \new_[35463]_ ;
  assign \new_[35468]_  = A301 & A300;
  assign \new_[35469]_  = A299 & \new_[35468]_ ;
  assign \new_[35470]_  = \new_[35469]_  & \new_[35464]_ ;
  assign \new_[35474]_  = ~A199 & ~A168;
  assign \new_[35475]_  = A169 & \new_[35474]_ ;
  assign \new_[35479]_  = A203 & A201;
  assign \new_[35480]_  = A200 & \new_[35479]_ ;
  assign \new_[35481]_  = \new_[35480]_  & \new_[35475]_ ;
  assign \new_[35485]_  = ~A298 & ~A266;
  assign \new_[35486]_  = ~A265 & \new_[35485]_ ;
  assign \new_[35490]_  = A302 & A300;
  assign \new_[35491]_  = A299 & \new_[35490]_ ;
  assign \new_[35492]_  = \new_[35491]_  & \new_[35486]_ ;
  assign \new_[35496]_  = A199 & ~A168;
  assign \new_[35497]_  = A169 & \new_[35496]_ ;
  assign \new_[35501]_  = A202 & A201;
  assign \new_[35502]_  = ~A200 & \new_[35501]_ ;
  assign \new_[35503]_  = \new_[35502]_  & \new_[35497]_ ;
  assign \new_[35507]_  = A298 & A268;
  assign \new_[35508]_  = ~A267 & \new_[35507]_ ;
  assign \new_[35512]_  = A301 & A300;
  assign \new_[35513]_  = ~A299 & \new_[35512]_ ;
  assign \new_[35514]_  = \new_[35513]_  & \new_[35508]_ ;
  assign \new_[35518]_  = A199 & ~A168;
  assign \new_[35519]_  = A169 & \new_[35518]_ ;
  assign \new_[35523]_  = A202 & A201;
  assign \new_[35524]_  = ~A200 & \new_[35523]_ ;
  assign \new_[35525]_  = \new_[35524]_  & \new_[35519]_ ;
  assign \new_[35529]_  = A298 & A268;
  assign \new_[35530]_  = ~A267 & \new_[35529]_ ;
  assign \new_[35534]_  = A302 & A300;
  assign \new_[35535]_  = ~A299 & \new_[35534]_ ;
  assign \new_[35536]_  = \new_[35535]_  & \new_[35530]_ ;
  assign \new_[35540]_  = A199 & ~A168;
  assign \new_[35541]_  = A169 & \new_[35540]_ ;
  assign \new_[35545]_  = A202 & A201;
  assign \new_[35546]_  = ~A200 & \new_[35545]_ ;
  assign \new_[35547]_  = \new_[35546]_  & \new_[35541]_ ;
  assign \new_[35551]_  = ~A298 & A268;
  assign \new_[35552]_  = ~A267 & \new_[35551]_ ;
  assign \new_[35556]_  = A301 & A300;
  assign \new_[35557]_  = A299 & \new_[35556]_ ;
  assign \new_[35558]_  = \new_[35557]_  & \new_[35552]_ ;
  assign \new_[35562]_  = A199 & ~A168;
  assign \new_[35563]_  = A169 & \new_[35562]_ ;
  assign \new_[35567]_  = A202 & A201;
  assign \new_[35568]_  = ~A200 & \new_[35567]_ ;
  assign \new_[35569]_  = \new_[35568]_  & \new_[35563]_ ;
  assign \new_[35573]_  = ~A298 & A268;
  assign \new_[35574]_  = ~A267 & \new_[35573]_ ;
  assign \new_[35578]_  = A302 & A300;
  assign \new_[35579]_  = A299 & \new_[35578]_ ;
  assign \new_[35580]_  = \new_[35579]_  & \new_[35574]_ ;
  assign \new_[35584]_  = A199 & ~A168;
  assign \new_[35585]_  = A169 & \new_[35584]_ ;
  assign \new_[35589]_  = A202 & A201;
  assign \new_[35590]_  = ~A200 & \new_[35589]_ ;
  assign \new_[35591]_  = \new_[35590]_  & \new_[35585]_ ;
  assign \new_[35595]_  = A298 & A269;
  assign \new_[35596]_  = ~A267 & \new_[35595]_ ;
  assign \new_[35600]_  = A301 & A300;
  assign \new_[35601]_  = ~A299 & \new_[35600]_ ;
  assign \new_[35602]_  = \new_[35601]_  & \new_[35596]_ ;
  assign \new_[35606]_  = A199 & ~A168;
  assign \new_[35607]_  = A169 & \new_[35606]_ ;
  assign \new_[35611]_  = A202 & A201;
  assign \new_[35612]_  = ~A200 & \new_[35611]_ ;
  assign \new_[35613]_  = \new_[35612]_  & \new_[35607]_ ;
  assign \new_[35617]_  = A298 & A269;
  assign \new_[35618]_  = ~A267 & \new_[35617]_ ;
  assign \new_[35622]_  = A302 & A300;
  assign \new_[35623]_  = ~A299 & \new_[35622]_ ;
  assign \new_[35624]_  = \new_[35623]_  & \new_[35618]_ ;
  assign \new_[35628]_  = A199 & ~A168;
  assign \new_[35629]_  = A169 & \new_[35628]_ ;
  assign \new_[35633]_  = A202 & A201;
  assign \new_[35634]_  = ~A200 & \new_[35633]_ ;
  assign \new_[35635]_  = \new_[35634]_  & \new_[35629]_ ;
  assign \new_[35639]_  = ~A298 & A269;
  assign \new_[35640]_  = ~A267 & \new_[35639]_ ;
  assign \new_[35644]_  = A301 & A300;
  assign \new_[35645]_  = A299 & \new_[35644]_ ;
  assign \new_[35646]_  = \new_[35645]_  & \new_[35640]_ ;
  assign \new_[35650]_  = A199 & ~A168;
  assign \new_[35651]_  = A169 & \new_[35650]_ ;
  assign \new_[35655]_  = A202 & A201;
  assign \new_[35656]_  = ~A200 & \new_[35655]_ ;
  assign \new_[35657]_  = \new_[35656]_  & \new_[35651]_ ;
  assign \new_[35661]_  = ~A298 & A269;
  assign \new_[35662]_  = ~A267 & \new_[35661]_ ;
  assign \new_[35666]_  = A302 & A300;
  assign \new_[35667]_  = A299 & \new_[35666]_ ;
  assign \new_[35668]_  = \new_[35667]_  & \new_[35662]_ ;
  assign \new_[35672]_  = A199 & ~A168;
  assign \new_[35673]_  = A169 & \new_[35672]_ ;
  assign \new_[35677]_  = A202 & A201;
  assign \new_[35678]_  = ~A200 & \new_[35677]_ ;
  assign \new_[35679]_  = \new_[35678]_  & \new_[35673]_ ;
  assign \new_[35683]_  = A298 & A266;
  assign \new_[35684]_  = A265 & \new_[35683]_ ;
  assign \new_[35688]_  = A301 & A300;
  assign \new_[35689]_  = ~A299 & \new_[35688]_ ;
  assign \new_[35690]_  = \new_[35689]_  & \new_[35684]_ ;
  assign \new_[35694]_  = A199 & ~A168;
  assign \new_[35695]_  = A169 & \new_[35694]_ ;
  assign \new_[35699]_  = A202 & A201;
  assign \new_[35700]_  = ~A200 & \new_[35699]_ ;
  assign \new_[35701]_  = \new_[35700]_  & \new_[35695]_ ;
  assign \new_[35705]_  = A298 & A266;
  assign \new_[35706]_  = A265 & \new_[35705]_ ;
  assign \new_[35710]_  = A302 & A300;
  assign \new_[35711]_  = ~A299 & \new_[35710]_ ;
  assign \new_[35712]_  = \new_[35711]_  & \new_[35706]_ ;
  assign \new_[35716]_  = A199 & ~A168;
  assign \new_[35717]_  = A169 & \new_[35716]_ ;
  assign \new_[35721]_  = A202 & A201;
  assign \new_[35722]_  = ~A200 & \new_[35721]_ ;
  assign \new_[35723]_  = \new_[35722]_  & \new_[35717]_ ;
  assign \new_[35727]_  = ~A298 & A266;
  assign \new_[35728]_  = A265 & \new_[35727]_ ;
  assign \new_[35732]_  = A301 & A300;
  assign \new_[35733]_  = A299 & \new_[35732]_ ;
  assign \new_[35734]_  = \new_[35733]_  & \new_[35728]_ ;
  assign \new_[35738]_  = A199 & ~A168;
  assign \new_[35739]_  = A169 & \new_[35738]_ ;
  assign \new_[35743]_  = A202 & A201;
  assign \new_[35744]_  = ~A200 & \new_[35743]_ ;
  assign \new_[35745]_  = \new_[35744]_  & \new_[35739]_ ;
  assign \new_[35749]_  = ~A298 & A266;
  assign \new_[35750]_  = A265 & \new_[35749]_ ;
  assign \new_[35754]_  = A302 & A300;
  assign \new_[35755]_  = A299 & \new_[35754]_ ;
  assign \new_[35756]_  = \new_[35755]_  & \new_[35750]_ ;
  assign \new_[35760]_  = A199 & ~A168;
  assign \new_[35761]_  = A169 & \new_[35760]_ ;
  assign \new_[35765]_  = A202 & A201;
  assign \new_[35766]_  = ~A200 & \new_[35765]_ ;
  assign \new_[35767]_  = \new_[35766]_  & \new_[35761]_ ;
  assign \new_[35771]_  = A298 & ~A266;
  assign \new_[35772]_  = ~A265 & \new_[35771]_ ;
  assign \new_[35776]_  = A301 & A300;
  assign \new_[35777]_  = ~A299 & \new_[35776]_ ;
  assign \new_[35778]_  = \new_[35777]_  & \new_[35772]_ ;
  assign \new_[35782]_  = A199 & ~A168;
  assign \new_[35783]_  = A169 & \new_[35782]_ ;
  assign \new_[35787]_  = A202 & A201;
  assign \new_[35788]_  = ~A200 & \new_[35787]_ ;
  assign \new_[35789]_  = \new_[35788]_  & \new_[35783]_ ;
  assign \new_[35793]_  = A298 & ~A266;
  assign \new_[35794]_  = ~A265 & \new_[35793]_ ;
  assign \new_[35798]_  = A302 & A300;
  assign \new_[35799]_  = ~A299 & \new_[35798]_ ;
  assign \new_[35800]_  = \new_[35799]_  & \new_[35794]_ ;
  assign \new_[35804]_  = A199 & ~A168;
  assign \new_[35805]_  = A169 & \new_[35804]_ ;
  assign \new_[35809]_  = A202 & A201;
  assign \new_[35810]_  = ~A200 & \new_[35809]_ ;
  assign \new_[35811]_  = \new_[35810]_  & \new_[35805]_ ;
  assign \new_[35815]_  = ~A298 & ~A266;
  assign \new_[35816]_  = ~A265 & \new_[35815]_ ;
  assign \new_[35820]_  = A301 & A300;
  assign \new_[35821]_  = A299 & \new_[35820]_ ;
  assign \new_[35822]_  = \new_[35821]_  & \new_[35816]_ ;
  assign \new_[35826]_  = A199 & ~A168;
  assign \new_[35827]_  = A169 & \new_[35826]_ ;
  assign \new_[35831]_  = A202 & A201;
  assign \new_[35832]_  = ~A200 & \new_[35831]_ ;
  assign \new_[35833]_  = \new_[35832]_  & \new_[35827]_ ;
  assign \new_[35837]_  = ~A298 & ~A266;
  assign \new_[35838]_  = ~A265 & \new_[35837]_ ;
  assign \new_[35842]_  = A302 & A300;
  assign \new_[35843]_  = A299 & \new_[35842]_ ;
  assign \new_[35844]_  = \new_[35843]_  & \new_[35838]_ ;
  assign \new_[35848]_  = A199 & ~A168;
  assign \new_[35849]_  = A169 & \new_[35848]_ ;
  assign \new_[35853]_  = A203 & A201;
  assign \new_[35854]_  = ~A200 & \new_[35853]_ ;
  assign \new_[35855]_  = \new_[35854]_  & \new_[35849]_ ;
  assign \new_[35859]_  = A298 & A268;
  assign \new_[35860]_  = ~A267 & \new_[35859]_ ;
  assign \new_[35864]_  = A301 & A300;
  assign \new_[35865]_  = ~A299 & \new_[35864]_ ;
  assign \new_[35866]_  = \new_[35865]_  & \new_[35860]_ ;
  assign \new_[35870]_  = A199 & ~A168;
  assign \new_[35871]_  = A169 & \new_[35870]_ ;
  assign \new_[35875]_  = A203 & A201;
  assign \new_[35876]_  = ~A200 & \new_[35875]_ ;
  assign \new_[35877]_  = \new_[35876]_  & \new_[35871]_ ;
  assign \new_[35881]_  = A298 & A268;
  assign \new_[35882]_  = ~A267 & \new_[35881]_ ;
  assign \new_[35886]_  = A302 & A300;
  assign \new_[35887]_  = ~A299 & \new_[35886]_ ;
  assign \new_[35888]_  = \new_[35887]_  & \new_[35882]_ ;
  assign \new_[35892]_  = A199 & ~A168;
  assign \new_[35893]_  = A169 & \new_[35892]_ ;
  assign \new_[35897]_  = A203 & A201;
  assign \new_[35898]_  = ~A200 & \new_[35897]_ ;
  assign \new_[35899]_  = \new_[35898]_  & \new_[35893]_ ;
  assign \new_[35903]_  = ~A298 & A268;
  assign \new_[35904]_  = ~A267 & \new_[35903]_ ;
  assign \new_[35908]_  = A301 & A300;
  assign \new_[35909]_  = A299 & \new_[35908]_ ;
  assign \new_[35910]_  = \new_[35909]_  & \new_[35904]_ ;
  assign \new_[35914]_  = A199 & ~A168;
  assign \new_[35915]_  = A169 & \new_[35914]_ ;
  assign \new_[35919]_  = A203 & A201;
  assign \new_[35920]_  = ~A200 & \new_[35919]_ ;
  assign \new_[35921]_  = \new_[35920]_  & \new_[35915]_ ;
  assign \new_[35925]_  = ~A298 & A268;
  assign \new_[35926]_  = ~A267 & \new_[35925]_ ;
  assign \new_[35930]_  = A302 & A300;
  assign \new_[35931]_  = A299 & \new_[35930]_ ;
  assign \new_[35932]_  = \new_[35931]_  & \new_[35926]_ ;
  assign \new_[35936]_  = A199 & ~A168;
  assign \new_[35937]_  = A169 & \new_[35936]_ ;
  assign \new_[35941]_  = A203 & A201;
  assign \new_[35942]_  = ~A200 & \new_[35941]_ ;
  assign \new_[35943]_  = \new_[35942]_  & \new_[35937]_ ;
  assign \new_[35947]_  = A298 & A269;
  assign \new_[35948]_  = ~A267 & \new_[35947]_ ;
  assign \new_[35952]_  = A301 & A300;
  assign \new_[35953]_  = ~A299 & \new_[35952]_ ;
  assign \new_[35954]_  = \new_[35953]_  & \new_[35948]_ ;
  assign \new_[35958]_  = A199 & ~A168;
  assign \new_[35959]_  = A169 & \new_[35958]_ ;
  assign \new_[35963]_  = A203 & A201;
  assign \new_[35964]_  = ~A200 & \new_[35963]_ ;
  assign \new_[35965]_  = \new_[35964]_  & \new_[35959]_ ;
  assign \new_[35969]_  = A298 & A269;
  assign \new_[35970]_  = ~A267 & \new_[35969]_ ;
  assign \new_[35974]_  = A302 & A300;
  assign \new_[35975]_  = ~A299 & \new_[35974]_ ;
  assign \new_[35976]_  = \new_[35975]_  & \new_[35970]_ ;
  assign \new_[35980]_  = A199 & ~A168;
  assign \new_[35981]_  = A169 & \new_[35980]_ ;
  assign \new_[35985]_  = A203 & A201;
  assign \new_[35986]_  = ~A200 & \new_[35985]_ ;
  assign \new_[35987]_  = \new_[35986]_  & \new_[35981]_ ;
  assign \new_[35991]_  = ~A298 & A269;
  assign \new_[35992]_  = ~A267 & \new_[35991]_ ;
  assign \new_[35996]_  = A301 & A300;
  assign \new_[35997]_  = A299 & \new_[35996]_ ;
  assign \new_[35998]_  = \new_[35997]_  & \new_[35992]_ ;
  assign \new_[36002]_  = A199 & ~A168;
  assign \new_[36003]_  = A169 & \new_[36002]_ ;
  assign \new_[36007]_  = A203 & A201;
  assign \new_[36008]_  = ~A200 & \new_[36007]_ ;
  assign \new_[36009]_  = \new_[36008]_  & \new_[36003]_ ;
  assign \new_[36013]_  = ~A298 & A269;
  assign \new_[36014]_  = ~A267 & \new_[36013]_ ;
  assign \new_[36018]_  = A302 & A300;
  assign \new_[36019]_  = A299 & \new_[36018]_ ;
  assign \new_[36020]_  = \new_[36019]_  & \new_[36014]_ ;
  assign \new_[36024]_  = A199 & ~A168;
  assign \new_[36025]_  = A169 & \new_[36024]_ ;
  assign \new_[36029]_  = A203 & A201;
  assign \new_[36030]_  = ~A200 & \new_[36029]_ ;
  assign \new_[36031]_  = \new_[36030]_  & \new_[36025]_ ;
  assign \new_[36035]_  = A298 & A266;
  assign \new_[36036]_  = A265 & \new_[36035]_ ;
  assign \new_[36040]_  = A301 & A300;
  assign \new_[36041]_  = ~A299 & \new_[36040]_ ;
  assign \new_[36042]_  = \new_[36041]_  & \new_[36036]_ ;
  assign \new_[36046]_  = A199 & ~A168;
  assign \new_[36047]_  = A169 & \new_[36046]_ ;
  assign \new_[36051]_  = A203 & A201;
  assign \new_[36052]_  = ~A200 & \new_[36051]_ ;
  assign \new_[36053]_  = \new_[36052]_  & \new_[36047]_ ;
  assign \new_[36057]_  = A298 & A266;
  assign \new_[36058]_  = A265 & \new_[36057]_ ;
  assign \new_[36062]_  = A302 & A300;
  assign \new_[36063]_  = ~A299 & \new_[36062]_ ;
  assign \new_[36064]_  = \new_[36063]_  & \new_[36058]_ ;
  assign \new_[36068]_  = A199 & ~A168;
  assign \new_[36069]_  = A169 & \new_[36068]_ ;
  assign \new_[36073]_  = A203 & A201;
  assign \new_[36074]_  = ~A200 & \new_[36073]_ ;
  assign \new_[36075]_  = \new_[36074]_  & \new_[36069]_ ;
  assign \new_[36079]_  = ~A298 & A266;
  assign \new_[36080]_  = A265 & \new_[36079]_ ;
  assign \new_[36084]_  = A301 & A300;
  assign \new_[36085]_  = A299 & \new_[36084]_ ;
  assign \new_[36086]_  = \new_[36085]_  & \new_[36080]_ ;
  assign \new_[36090]_  = A199 & ~A168;
  assign \new_[36091]_  = A169 & \new_[36090]_ ;
  assign \new_[36095]_  = A203 & A201;
  assign \new_[36096]_  = ~A200 & \new_[36095]_ ;
  assign \new_[36097]_  = \new_[36096]_  & \new_[36091]_ ;
  assign \new_[36101]_  = ~A298 & A266;
  assign \new_[36102]_  = A265 & \new_[36101]_ ;
  assign \new_[36106]_  = A302 & A300;
  assign \new_[36107]_  = A299 & \new_[36106]_ ;
  assign \new_[36108]_  = \new_[36107]_  & \new_[36102]_ ;
  assign \new_[36112]_  = A199 & ~A168;
  assign \new_[36113]_  = A169 & \new_[36112]_ ;
  assign \new_[36117]_  = A203 & A201;
  assign \new_[36118]_  = ~A200 & \new_[36117]_ ;
  assign \new_[36119]_  = \new_[36118]_  & \new_[36113]_ ;
  assign \new_[36123]_  = A298 & ~A266;
  assign \new_[36124]_  = ~A265 & \new_[36123]_ ;
  assign \new_[36128]_  = A301 & A300;
  assign \new_[36129]_  = ~A299 & \new_[36128]_ ;
  assign \new_[36130]_  = \new_[36129]_  & \new_[36124]_ ;
  assign \new_[36134]_  = A199 & ~A168;
  assign \new_[36135]_  = A169 & \new_[36134]_ ;
  assign \new_[36139]_  = A203 & A201;
  assign \new_[36140]_  = ~A200 & \new_[36139]_ ;
  assign \new_[36141]_  = \new_[36140]_  & \new_[36135]_ ;
  assign \new_[36145]_  = A298 & ~A266;
  assign \new_[36146]_  = ~A265 & \new_[36145]_ ;
  assign \new_[36150]_  = A302 & A300;
  assign \new_[36151]_  = ~A299 & \new_[36150]_ ;
  assign \new_[36152]_  = \new_[36151]_  & \new_[36146]_ ;
  assign \new_[36156]_  = A199 & ~A168;
  assign \new_[36157]_  = A169 & \new_[36156]_ ;
  assign \new_[36161]_  = A203 & A201;
  assign \new_[36162]_  = ~A200 & \new_[36161]_ ;
  assign \new_[36163]_  = \new_[36162]_  & \new_[36157]_ ;
  assign \new_[36167]_  = ~A298 & ~A266;
  assign \new_[36168]_  = ~A265 & \new_[36167]_ ;
  assign \new_[36172]_  = A301 & A300;
  assign \new_[36173]_  = A299 & \new_[36172]_ ;
  assign \new_[36174]_  = \new_[36173]_  & \new_[36168]_ ;
  assign \new_[36178]_  = A199 & ~A168;
  assign \new_[36179]_  = A169 & \new_[36178]_ ;
  assign \new_[36183]_  = A203 & A201;
  assign \new_[36184]_  = ~A200 & \new_[36183]_ ;
  assign \new_[36185]_  = \new_[36184]_  & \new_[36179]_ ;
  assign \new_[36189]_  = ~A298 & ~A266;
  assign \new_[36190]_  = ~A265 & \new_[36189]_ ;
  assign \new_[36194]_  = A302 & A300;
  assign \new_[36195]_  = A299 & \new_[36194]_ ;
  assign \new_[36196]_  = \new_[36195]_  & \new_[36190]_ ;
  assign \new_[36200]_  = ~A199 & ~A168;
  assign \new_[36201]_  = A169 & \new_[36200]_ ;
  assign \new_[36205]_  = A266 & ~A265;
  assign \new_[36206]_  = ~A200 & \new_[36205]_ ;
  assign \new_[36207]_  = \new_[36206]_  & \new_[36201]_ ;
  assign \new_[36211]_  = ~A269 & ~A268;
  assign \new_[36212]_  = ~A267 & \new_[36211]_ ;
  assign \new_[36216]_  = ~A302 & ~A301;
  assign \new_[36217]_  = A300 & \new_[36216]_ ;
  assign \new_[36218]_  = \new_[36217]_  & \new_[36212]_ ;
  assign \new_[36222]_  = ~A199 & ~A168;
  assign \new_[36223]_  = A169 & \new_[36222]_ ;
  assign \new_[36227]_  = ~A266 & A265;
  assign \new_[36228]_  = ~A200 & \new_[36227]_ ;
  assign \new_[36229]_  = \new_[36228]_  & \new_[36223]_ ;
  assign \new_[36233]_  = ~A269 & ~A268;
  assign \new_[36234]_  = ~A267 & \new_[36233]_ ;
  assign \new_[36238]_  = ~A302 & ~A301;
  assign \new_[36239]_  = A300 & \new_[36238]_ ;
  assign \new_[36240]_  = \new_[36239]_  & \new_[36234]_ ;
  assign \new_[36244]_  = A168 & ~A169;
  assign \new_[36245]_  = A170 & \new_[36244]_ ;
  assign \new_[36249]_  = ~A203 & ~A202;
  assign \new_[36250]_  = A201 & \new_[36249]_ ;
  assign \new_[36251]_  = \new_[36250]_  & \new_[36245]_ ;
  assign \new_[36255]_  = A267 & A266;
  assign \new_[36256]_  = ~A265 & \new_[36255]_ ;
  assign \new_[36260]_  = A301 & ~A300;
  assign \new_[36261]_  = A268 & \new_[36260]_ ;
  assign \new_[36262]_  = \new_[36261]_  & \new_[36256]_ ;
  assign \new_[36266]_  = A168 & ~A169;
  assign \new_[36267]_  = A170 & \new_[36266]_ ;
  assign \new_[36271]_  = ~A203 & ~A202;
  assign \new_[36272]_  = A201 & \new_[36271]_ ;
  assign \new_[36273]_  = \new_[36272]_  & \new_[36267]_ ;
  assign \new_[36277]_  = A267 & A266;
  assign \new_[36278]_  = ~A265 & \new_[36277]_ ;
  assign \new_[36282]_  = A302 & ~A300;
  assign \new_[36283]_  = A268 & \new_[36282]_ ;
  assign \new_[36284]_  = \new_[36283]_  & \new_[36278]_ ;
  assign \new_[36288]_  = A168 & ~A169;
  assign \new_[36289]_  = A170 & \new_[36288]_ ;
  assign \new_[36293]_  = ~A203 & ~A202;
  assign \new_[36294]_  = A201 & \new_[36293]_ ;
  assign \new_[36295]_  = \new_[36294]_  & \new_[36289]_ ;
  assign \new_[36299]_  = A267 & A266;
  assign \new_[36300]_  = ~A265 & \new_[36299]_ ;
  assign \new_[36304]_  = A299 & A298;
  assign \new_[36305]_  = A268 & \new_[36304]_ ;
  assign \new_[36306]_  = \new_[36305]_  & \new_[36300]_ ;
  assign \new_[36310]_  = A168 & ~A169;
  assign \new_[36311]_  = A170 & \new_[36310]_ ;
  assign \new_[36315]_  = ~A203 & ~A202;
  assign \new_[36316]_  = A201 & \new_[36315]_ ;
  assign \new_[36317]_  = \new_[36316]_  & \new_[36311]_ ;
  assign \new_[36321]_  = A267 & A266;
  assign \new_[36322]_  = ~A265 & \new_[36321]_ ;
  assign \new_[36326]_  = ~A299 & ~A298;
  assign \new_[36327]_  = A268 & \new_[36326]_ ;
  assign \new_[36328]_  = \new_[36327]_  & \new_[36322]_ ;
  assign \new_[36332]_  = A168 & ~A169;
  assign \new_[36333]_  = A170 & \new_[36332]_ ;
  assign \new_[36337]_  = ~A203 & ~A202;
  assign \new_[36338]_  = A201 & \new_[36337]_ ;
  assign \new_[36339]_  = \new_[36338]_  & \new_[36333]_ ;
  assign \new_[36343]_  = A267 & A266;
  assign \new_[36344]_  = ~A265 & \new_[36343]_ ;
  assign \new_[36348]_  = A301 & ~A300;
  assign \new_[36349]_  = A269 & \new_[36348]_ ;
  assign \new_[36350]_  = \new_[36349]_  & \new_[36344]_ ;
  assign \new_[36354]_  = A168 & ~A169;
  assign \new_[36355]_  = A170 & \new_[36354]_ ;
  assign \new_[36359]_  = ~A203 & ~A202;
  assign \new_[36360]_  = A201 & \new_[36359]_ ;
  assign \new_[36361]_  = \new_[36360]_  & \new_[36355]_ ;
  assign \new_[36365]_  = A267 & A266;
  assign \new_[36366]_  = ~A265 & \new_[36365]_ ;
  assign \new_[36370]_  = A302 & ~A300;
  assign \new_[36371]_  = A269 & \new_[36370]_ ;
  assign \new_[36372]_  = \new_[36371]_  & \new_[36366]_ ;
  assign \new_[36376]_  = A168 & ~A169;
  assign \new_[36377]_  = A170 & \new_[36376]_ ;
  assign \new_[36381]_  = ~A203 & ~A202;
  assign \new_[36382]_  = A201 & \new_[36381]_ ;
  assign \new_[36383]_  = \new_[36382]_  & \new_[36377]_ ;
  assign \new_[36387]_  = A267 & A266;
  assign \new_[36388]_  = ~A265 & \new_[36387]_ ;
  assign \new_[36392]_  = A299 & A298;
  assign \new_[36393]_  = A269 & \new_[36392]_ ;
  assign \new_[36394]_  = \new_[36393]_  & \new_[36388]_ ;
  assign \new_[36398]_  = A168 & ~A169;
  assign \new_[36399]_  = A170 & \new_[36398]_ ;
  assign \new_[36403]_  = ~A203 & ~A202;
  assign \new_[36404]_  = A201 & \new_[36403]_ ;
  assign \new_[36405]_  = \new_[36404]_  & \new_[36399]_ ;
  assign \new_[36409]_  = A267 & A266;
  assign \new_[36410]_  = ~A265 & \new_[36409]_ ;
  assign \new_[36414]_  = ~A299 & ~A298;
  assign \new_[36415]_  = A269 & \new_[36414]_ ;
  assign \new_[36416]_  = \new_[36415]_  & \new_[36410]_ ;
  assign \new_[36420]_  = A168 & ~A169;
  assign \new_[36421]_  = A170 & \new_[36420]_ ;
  assign \new_[36425]_  = ~A203 & ~A202;
  assign \new_[36426]_  = A201 & \new_[36425]_ ;
  assign \new_[36427]_  = \new_[36426]_  & \new_[36421]_ ;
  assign \new_[36431]_  = A267 & ~A266;
  assign \new_[36432]_  = A265 & \new_[36431]_ ;
  assign \new_[36436]_  = A301 & ~A300;
  assign \new_[36437]_  = A268 & \new_[36436]_ ;
  assign \new_[36438]_  = \new_[36437]_  & \new_[36432]_ ;
  assign \new_[36442]_  = A168 & ~A169;
  assign \new_[36443]_  = A170 & \new_[36442]_ ;
  assign \new_[36447]_  = ~A203 & ~A202;
  assign \new_[36448]_  = A201 & \new_[36447]_ ;
  assign \new_[36449]_  = \new_[36448]_  & \new_[36443]_ ;
  assign \new_[36453]_  = A267 & ~A266;
  assign \new_[36454]_  = A265 & \new_[36453]_ ;
  assign \new_[36458]_  = A302 & ~A300;
  assign \new_[36459]_  = A268 & \new_[36458]_ ;
  assign \new_[36460]_  = \new_[36459]_  & \new_[36454]_ ;
  assign \new_[36464]_  = A168 & ~A169;
  assign \new_[36465]_  = A170 & \new_[36464]_ ;
  assign \new_[36469]_  = ~A203 & ~A202;
  assign \new_[36470]_  = A201 & \new_[36469]_ ;
  assign \new_[36471]_  = \new_[36470]_  & \new_[36465]_ ;
  assign \new_[36475]_  = A267 & ~A266;
  assign \new_[36476]_  = A265 & \new_[36475]_ ;
  assign \new_[36480]_  = A299 & A298;
  assign \new_[36481]_  = A268 & \new_[36480]_ ;
  assign \new_[36482]_  = \new_[36481]_  & \new_[36476]_ ;
  assign \new_[36486]_  = A168 & ~A169;
  assign \new_[36487]_  = A170 & \new_[36486]_ ;
  assign \new_[36491]_  = ~A203 & ~A202;
  assign \new_[36492]_  = A201 & \new_[36491]_ ;
  assign \new_[36493]_  = \new_[36492]_  & \new_[36487]_ ;
  assign \new_[36497]_  = A267 & ~A266;
  assign \new_[36498]_  = A265 & \new_[36497]_ ;
  assign \new_[36502]_  = ~A299 & ~A298;
  assign \new_[36503]_  = A268 & \new_[36502]_ ;
  assign \new_[36504]_  = \new_[36503]_  & \new_[36498]_ ;
  assign \new_[36508]_  = A168 & ~A169;
  assign \new_[36509]_  = A170 & \new_[36508]_ ;
  assign \new_[36513]_  = ~A203 & ~A202;
  assign \new_[36514]_  = A201 & \new_[36513]_ ;
  assign \new_[36515]_  = \new_[36514]_  & \new_[36509]_ ;
  assign \new_[36519]_  = A267 & ~A266;
  assign \new_[36520]_  = A265 & \new_[36519]_ ;
  assign \new_[36524]_  = A301 & ~A300;
  assign \new_[36525]_  = A269 & \new_[36524]_ ;
  assign \new_[36526]_  = \new_[36525]_  & \new_[36520]_ ;
  assign \new_[36530]_  = A168 & ~A169;
  assign \new_[36531]_  = A170 & \new_[36530]_ ;
  assign \new_[36535]_  = ~A203 & ~A202;
  assign \new_[36536]_  = A201 & \new_[36535]_ ;
  assign \new_[36537]_  = \new_[36536]_  & \new_[36531]_ ;
  assign \new_[36541]_  = A267 & ~A266;
  assign \new_[36542]_  = A265 & \new_[36541]_ ;
  assign \new_[36546]_  = A302 & ~A300;
  assign \new_[36547]_  = A269 & \new_[36546]_ ;
  assign \new_[36548]_  = \new_[36547]_  & \new_[36542]_ ;
  assign \new_[36552]_  = A168 & ~A169;
  assign \new_[36553]_  = A170 & \new_[36552]_ ;
  assign \new_[36557]_  = ~A203 & ~A202;
  assign \new_[36558]_  = A201 & \new_[36557]_ ;
  assign \new_[36559]_  = \new_[36558]_  & \new_[36553]_ ;
  assign \new_[36563]_  = A267 & ~A266;
  assign \new_[36564]_  = A265 & \new_[36563]_ ;
  assign \new_[36568]_  = A299 & A298;
  assign \new_[36569]_  = A269 & \new_[36568]_ ;
  assign \new_[36570]_  = \new_[36569]_  & \new_[36564]_ ;
  assign \new_[36574]_  = A168 & ~A169;
  assign \new_[36575]_  = A170 & \new_[36574]_ ;
  assign \new_[36579]_  = ~A203 & ~A202;
  assign \new_[36580]_  = A201 & \new_[36579]_ ;
  assign \new_[36581]_  = \new_[36580]_  & \new_[36575]_ ;
  assign \new_[36585]_  = A267 & ~A266;
  assign \new_[36586]_  = A265 & \new_[36585]_ ;
  assign \new_[36590]_  = ~A299 & ~A298;
  assign \new_[36591]_  = A269 & \new_[36590]_ ;
  assign \new_[36592]_  = \new_[36591]_  & \new_[36586]_ ;
  assign \new_[36596]_  = A168 & ~A169;
  assign \new_[36597]_  = A170 & \new_[36596]_ ;
  assign \new_[36601]_  = ~A265 & A202;
  assign \new_[36602]_  = ~A201 & \new_[36601]_ ;
  assign \new_[36603]_  = \new_[36602]_  & \new_[36597]_ ;
  assign \new_[36607]_  = A268 & A267;
  assign \new_[36608]_  = A266 & \new_[36607]_ ;
  assign \new_[36612]_  = ~A302 & ~A301;
  assign \new_[36613]_  = A300 & \new_[36612]_ ;
  assign \new_[36614]_  = \new_[36613]_  & \new_[36608]_ ;
  assign \new_[36618]_  = A168 & ~A169;
  assign \new_[36619]_  = A170 & \new_[36618]_ ;
  assign \new_[36623]_  = ~A265 & A202;
  assign \new_[36624]_  = ~A201 & \new_[36623]_ ;
  assign \new_[36625]_  = \new_[36624]_  & \new_[36619]_ ;
  assign \new_[36629]_  = A269 & A267;
  assign \new_[36630]_  = A266 & \new_[36629]_ ;
  assign \new_[36634]_  = ~A302 & ~A301;
  assign \new_[36635]_  = A300 & \new_[36634]_ ;
  assign \new_[36636]_  = \new_[36635]_  & \new_[36630]_ ;
  assign \new_[36640]_  = A168 & ~A169;
  assign \new_[36641]_  = A170 & \new_[36640]_ ;
  assign \new_[36645]_  = ~A265 & A202;
  assign \new_[36646]_  = ~A201 & \new_[36645]_ ;
  assign \new_[36647]_  = \new_[36646]_  & \new_[36641]_ ;
  assign \new_[36651]_  = ~A268 & ~A267;
  assign \new_[36652]_  = A266 & \new_[36651]_ ;
  assign \new_[36656]_  = A301 & ~A300;
  assign \new_[36657]_  = ~A269 & \new_[36656]_ ;
  assign \new_[36658]_  = \new_[36657]_  & \new_[36652]_ ;
  assign \new_[36662]_  = A168 & ~A169;
  assign \new_[36663]_  = A170 & \new_[36662]_ ;
  assign \new_[36667]_  = ~A265 & A202;
  assign \new_[36668]_  = ~A201 & \new_[36667]_ ;
  assign \new_[36669]_  = \new_[36668]_  & \new_[36663]_ ;
  assign \new_[36673]_  = ~A268 & ~A267;
  assign \new_[36674]_  = A266 & \new_[36673]_ ;
  assign \new_[36678]_  = A302 & ~A300;
  assign \new_[36679]_  = ~A269 & \new_[36678]_ ;
  assign \new_[36680]_  = \new_[36679]_  & \new_[36674]_ ;
  assign \new_[36684]_  = A168 & ~A169;
  assign \new_[36685]_  = A170 & \new_[36684]_ ;
  assign \new_[36689]_  = ~A265 & A202;
  assign \new_[36690]_  = ~A201 & \new_[36689]_ ;
  assign \new_[36691]_  = \new_[36690]_  & \new_[36685]_ ;
  assign \new_[36695]_  = ~A268 & ~A267;
  assign \new_[36696]_  = A266 & \new_[36695]_ ;
  assign \new_[36700]_  = A299 & A298;
  assign \new_[36701]_  = ~A269 & \new_[36700]_ ;
  assign \new_[36702]_  = \new_[36701]_  & \new_[36696]_ ;
  assign \new_[36706]_  = A168 & ~A169;
  assign \new_[36707]_  = A170 & \new_[36706]_ ;
  assign \new_[36711]_  = ~A265 & A202;
  assign \new_[36712]_  = ~A201 & \new_[36711]_ ;
  assign \new_[36713]_  = \new_[36712]_  & \new_[36707]_ ;
  assign \new_[36717]_  = ~A268 & ~A267;
  assign \new_[36718]_  = A266 & \new_[36717]_ ;
  assign \new_[36722]_  = ~A299 & ~A298;
  assign \new_[36723]_  = ~A269 & \new_[36722]_ ;
  assign \new_[36724]_  = \new_[36723]_  & \new_[36718]_ ;
  assign \new_[36728]_  = A168 & ~A169;
  assign \new_[36729]_  = A170 & \new_[36728]_ ;
  assign \new_[36733]_  = A265 & A202;
  assign \new_[36734]_  = ~A201 & \new_[36733]_ ;
  assign \new_[36735]_  = \new_[36734]_  & \new_[36729]_ ;
  assign \new_[36739]_  = A268 & A267;
  assign \new_[36740]_  = ~A266 & \new_[36739]_ ;
  assign \new_[36744]_  = ~A302 & ~A301;
  assign \new_[36745]_  = A300 & \new_[36744]_ ;
  assign \new_[36746]_  = \new_[36745]_  & \new_[36740]_ ;
  assign \new_[36750]_  = A168 & ~A169;
  assign \new_[36751]_  = A170 & \new_[36750]_ ;
  assign \new_[36755]_  = A265 & A202;
  assign \new_[36756]_  = ~A201 & \new_[36755]_ ;
  assign \new_[36757]_  = \new_[36756]_  & \new_[36751]_ ;
  assign \new_[36761]_  = A269 & A267;
  assign \new_[36762]_  = ~A266 & \new_[36761]_ ;
  assign \new_[36766]_  = ~A302 & ~A301;
  assign \new_[36767]_  = A300 & \new_[36766]_ ;
  assign \new_[36768]_  = \new_[36767]_  & \new_[36762]_ ;
  assign \new_[36772]_  = A168 & ~A169;
  assign \new_[36773]_  = A170 & \new_[36772]_ ;
  assign \new_[36777]_  = A265 & A202;
  assign \new_[36778]_  = ~A201 & \new_[36777]_ ;
  assign \new_[36779]_  = \new_[36778]_  & \new_[36773]_ ;
  assign \new_[36783]_  = ~A268 & ~A267;
  assign \new_[36784]_  = ~A266 & \new_[36783]_ ;
  assign \new_[36788]_  = A301 & ~A300;
  assign \new_[36789]_  = ~A269 & \new_[36788]_ ;
  assign \new_[36790]_  = \new_[36789]_  & \new_[36784]_ ;
  assign \new_[36794]_  = A168 & ~A169;
  assign \new_[36795]_  = A170 & \new_[36794]_ ;
  assign \new_[36799]_  = A265 & A202;
  assign \new_[36800]_  = ~A201 & \new_[36799]_ ;
  assign \new_[36801]_  = \new_[36800]_  & \new_[36795]_ ;
  assign \new_[36805]_  = ~A268 & ~A267;
  assign \new_[36806]_  = ~A266 & \new_[36805]_ ;
  assign \new_[36810]_  = A302 & ~A300;
  assign \new_[36811]_  = ~A269 & \new_[36810]_ ;
  assign \new_[36812]_  = \new_[36811]_  & \new_[36806]_ ;
  assign \new_[36816]_  = A168 & ~A169;
  assign \new_[36817]_  = A170 & \new_[36816]_ ;
  assign \new_[36821]_  = A265 & A202;
  assign \new_[36822]_  = ~A201 & \new_[36821]_ ;
  assign \new_[36823]_  = \new_[36822]_  & \new_[36817]_ ;
  assign \new_[36827]_  = ~A268 & ~A267;
  assign \new_[36828]_  = ~A266 & \new_[36827]_ ;
  assign \new_[36832]_  = A299 & A298;
  assign \new_[36833]_  = ~A269 & \new_[36832]_ ;
  assign \new_[36834]_  = \new_[36833]_  & \new_[36828]_ ;
  assign \new_[36838]_  = A168 & ~A169;
  assign \new_[36839]_  = A170 & \new_[36838]_ ;
  assign \new_[36843]_  = A265 & A202;
  assign \new_[36844]_  = ~A201 & \new_[36843]_ ;
  assign \new_[36845]_  = \new_[36844]_  & \new_[36839]_ ;
  assign \new_[36849]_  = ~A268 & ~A267;
  assign \new_[36850]_  = ~A266 & \new_[36849]_ ;
  assign \new_[36854]_  = ~A299 & ~A298;
  assign \new_[36855]_  = ~A269 & \new_[36854]_ ;
  assign \new_[36856]_  = \new_[36855]_  & \new_[36850]_ ;
  assign \new_[36860]_  = A168 & ~A169;
  assign \new_[36861]_  = A170 & \new_[36860]_ ;
  assign \new_[36865]_  = ~A265 & A203;
  assign \new_[36866]_  = ~A201 & \new_[36865]_ ;
  assign \new_[36867]_  = \new_[36866]_  & \new_[36861]_ ;
  assign \new_[36871]_  = A268 & A267;
  assign \new_[36872]_  = A266 & \new_[36871]_ ;
  assign \new_[36876]_  = ~A302 & ~A301;
  assign \new_[36877]_  = A300 & \new_[36876]_ ;
  assign \new_[36878]_  = \new_[36877]_  & \new_[36872]_ ;
  assign \new_[36882]_  = A168 & ~A169;
  assign \new_[36883]_  = A170 & \new_[36882]_ ;
  assign \new_[36887]_  = ~A265 & A203;
  assign \new_[36888]_  = ~A201 & \new_[36887]_ ;
  assign \new_[36889]_  = \new_[36888]_  & \new_[36883]_ ;
  assign \new_[36893]_  = A269 & A267;
  assign \new_[36894]_  = A266 & \new_[36893]_ ;
  assign \new_[36898]_  = ~A302 & ~A301;
  assign \new_[36899]_  = A300 & \new_[36898]_ ;
  assign \new_[36900]_  = \new_[36899]_  & \new_[36894]_ ;
  assign \new_[36904]_  = A168 & ~A169;
  assign \new_[36905]_  = A170 & \new_[36904]_ ;
  assign \new_[36909]_  = ~A265 & A203;
  assign \new_[36910]_  = ~A201 & \new_[36909]_ ;
  assign \new_[36911]_  = \new_[36910]_  & \new_[36905]_ ;
  assign \new_[36915]_  = ~A268 & ~A267;
  assign \new_[36916]_  = A266 & \new_[36915]_ ;
  assign \new_[36920]_  = A301 & ~A300;
  assign \new_[36921]_  = ~A269 & \new_[36920]_ ;
  assign \new_[36922]_  = \new_[36921]_  & \new_[36916]_ ;
  assign \new_[36926]_  = A168 & ~A169;
  assign \new_[36927]_  = A170 & \new_[36926]_ ;
  assign \new_[36931]_  = ~A265 & A203;
  assign \new_[36932]_  = ~A201 & \new_[36931]_ ;
  assign \new_[36933]_  = \new_[36932]_  & \new_[36927]_ ;
  assign \new_[36937]_  = ~A268 & ~A267;
  assign \new_[36938]_  = A266 & \new_[36937]_ ;
  assign \new_[36942]_  = A302 & ~A300;
  assign \new_[36943]_  = ~A269 & \new_[36942]_ ;
  assign \new_[36944]_  = \new_[36943]_  & \new_[36938]_ ;
  assign \new_[36948]_  = A168 & ~A169;
  assign \new_[36949]_  = A170 & \new_[36948]_ ;
  assign \new_[36953]_  = ~A265 & A203;
  assign \new_[36954]_  = ~A201 & \new_[36953]_ ;
  assign \new_[36955]_  = \new_[36954]_  & \new_[36949]_ ;
  assign \new_[36959]_  = ~A268 & ~A267;
  assign \new_[36960]_  = A266 & \new_[36959]_ ;
  assign \new_[36964]_  = A299 & A298;
  assign \new_[36965]_  = ~A269 & \new_[36964]_ ;
  assign \new_[36966]_  = \new_[36965]_  & \new_[36960]_ ;
  assign \new_[36970]_  = A168 & ~A169;
  assign \new_[36971]_  = A170 & \new_[36970]_ ;
  assign \new_[36975]_  = ~A265 & A203;
  assign \new_[36976]_  = ~A201 & \new_[36975]_ ;
  assign \new_[36977]_  = \new_[36976]_  & \new_[36971]_ ;
  assign \new_[36981]_  = ~A268 & ~A267;
  assign \new_[36982]_  = A266 & \new_[36981]_ ;
  assign \new_[36986]_  = ~A299 & ~A298;
  assign \new_[36987]_  = ~A269 & \new_[36986]_ ;
  assign \new_[36988]_  = \new_[36987]_  & \new_[36982]_ ;
  assign \new_[36992]_  = A168 & ~A169;
  assign \new_[36993]_  = A170 & \new_[36992]_ ;
  assign \new_[36997]_  = A265 & A203;
  assign \new_[36998]_  = ~A201 & \new_[36997]_ ;
  assign \new_[36999]_  = \new_[36998]_  & \new_[36993]_ ;
  assign \new_[37003]_  = A268 & A267;
  assign \new_[37004]_  = ~A266 & \new_[37003]_ ;
  assign \new_[37008]_  = ~A302 & ~A301;
  assign \new_[37009]_  = A300 & \new_[37008]_ ;
  assign \new_[37010]_  = \new_[37009]_  & \new_[37004]_ ;
  assign \new_[37014]_  = A168 & ~A169;
  assign \new_[37015]_  = A170 & \new_[37014]_ ;
  assign \new_[37019]_  = A265 & A203;
  assign \new_[37020]_  = ~A201 & \new_[37019]_ ;
  assign \new_[37021]_  = \new_[37020]_  & \new_[37015]_ ;
  assign \new_[37025]_  = A269 & A267;
  assign \new_[37026]_  = ~A266 & \new_[37025]_ ;
  assign \new_[37030]_  = ~A302 & ~A301;
  assign \new_[37031]_  = A300 & \new_[37030]_ ;
  assign \new_[37032]_  = \new_[37031]_  & \new_[37026]_ ;
  assign \new_[37036]_  = A168 & ~A169;
  assign \new_[37037]_  = A170 & \new_[37036]_ ;
  assign \new_[37041]_  = A265 & A203;
  assign \new_[37042]_  = ~A201 & \new_[37041]_ ;
  assign \new_[37043]_  = \new_[37042]_  & \new_[37037]_ ;
  assign \new_[37047]_  = ~A268 & ~A267;
  assign \new_[37048]_  = ~A266 & \new_[37047]_ ;
  assign \new_[37052]_  = A301 & ~A300;
  assign \new_[37053]_  = ~A269 & \new_[37052]_ ;
  assign \new_[37054]_  = \new_[37053]_  & \new_[37048]_ ;
  assign \new_[37058]_  = A168 & ~A169;
  assign \new_[37059]_  = A170 & \new_[37058]_ ;
  assign \new_[37063]_  = A265 & A203;
  assign \new_[37064]_  = ~A201 & \new_[37063]_ ;
  assign \new_[37065]_  = \new_[37064]_  & \new_[37059]_ ;
  assign \new_[37069]_  = ~A268 & ~A267;
  assign \new_[37070]_  = ~A266 & \new_[37069]_ ;
  assign \new_[37074]_  = A302 & ~A300;
  assign \new_[37075]_  = ~A269 & \new_[37074]_ ;
  assign \new_[37076]_  = \new_[37075]_  & \new_[37070]_ ;
  assign \new_[37080]_  = A168 & ~A169;
  assign \new_[37081]_  = A170 & \new_[37080]_ ;
  assign \new_[37085]_  = A265 & A203;
  assign \new_[37086]_  = ~A201 & \new_[37085]_ ;
  assign \new_[37087]_  = \new_[37086]_  & \new_[37081]_ ;
  assign \new_[37091]_  = ~A268 & ~A267;
  assign \new_[37092]_  = ~A266 & \new_[37091]_ ;
  assign \new_[37096]_  = A299 & A298;
  assign \new_[37097]_  = ~A269 & \new_[37096]_ ;
  assign \new_[37098]_  = \new_[37097]_  & \new_[37092]_ ;
  assign \new_[37102]_  = A168 & ~A169;
  assign \new_[37103]_  = A170 & \new_[37102]_ ;
  assign \new_[37107]_  = A265 & A203;
  assign \new_[37108]_  = ~A201 & \new_[37107]_ ;
  assign \new_[37109]_  = \new_[37108]_  & \new_[37103]_ ;
  assign \new_[37113]_  = ~A268 & ~A267;
  assign \new_[37114]_  = ~A266 & \new_[37113]_ ;
  assign \new_[37118]_  = ~A299 & ~A298;
  assign \new_[37119]_  = ~A269 & \new_[37118]_ ;
  assign \new_[37120]_  = \new_[37119]_  & \new_[37114]_ ;
  assign \new_[37124]_  = A168 & ~A169;
  assign \new_[37125]_  = A170 & \new_[37124]_ ;
  assign \new_[37129]_  = ~A265 & A200;
  assign \new_[37130]_  = A199 & \new_[37129]_ ;
  assign \new_[37131]_  = \new_[37130]_  & \new_[37125]_ ;
  assign \new_[37135]_  = A268 & A267;
  assign \new_[37136]_  = A266 & \new_[37135]_ ;
  assign \new_[37140]_  = ~A302 & ~A301;
  assign \new_[37141]_  = A300 & \new_[37140]_ ;
  assign \new_[37142]_  = \new_[37141]_  & \new_[37136]_ ;
  assign \new_[37146]_  = A168 & ~A169;
  assign \new_[37147]_  = A170 & \new_[37146]_ ;
  assign \new_[37151]_  = ~A265 & A200;
  assign \new_[37152]_  = A199 & \new_[37151]_ ;
  assign \new_[37153]_  = \new_[37152]_  & \new_[37147]_ ;
  assign \new_[37157]_  = A269 & A267;
  assign \new_[37158]_  = A266 & \new_[37157]_ ;
  assign \new_[37162]_  = ~A302 & ~A301;
  assign \new_[37163]_  = A300 & \new_[37162]_ ;
  assign \new_[37164]_  = \new_[37163]_  & \new_[37158]_ ;
  assign \new_[37168]_  = A168 & ~A169;
  assign \new_[37169]_  = A170 & \new_[37168]_ ;
  assign \new_[37173]_  = ~A265 & A200;
  assign \new_[37174]_  = A199 & \new_[37173]_ ;
  assign \new_[37175]_  = \new_[37174]_  & \new_[37169]_ ;
  assign \new_[37179]_  = ~A268 & ~A267;
  assign \new_[37180]_  = A266 & \new_[37179]_ ;
  assign \new_[37184]_  = A301 & ~A300;
  assign \new_[37185]_  = ~A269 & \new_[37184]_ ;
  assign \new_[37186]_  = \new_[37185]_  & \new_[37180]_ ;
  assign \new_[37190]_  = A168 & ~A169;
  assign \new_[37191]_  = A170 & \new_[37190]_ ;
  assign \new_[37195]_  = ~A265 & A200;
  assign \new_[37196]_  = A199 & \new_[37195]_ ;
  assign \new_[37197]_  = \new_[37196]_  & \new_[37191]_ ;
  assign \new_[37201]_  = ~A268 & ~A267;
  assign \new_[37202]_  = A266 & \new_[37201]_ ;
  assign \new_[37206]_  = A302 & ~A300;
  assign \new_[37207]_  = ~A269 & \new_[37206]_ ;
  assign \new_[37208]_  = \new_[37207]_  & \new_[37202]_ ;
  assign \new_[37212]_  = A168 & ~A169;
  assign \new_[37213]_  = A170 & \new_[37212]_ ;
  assign \new_[37217]_  = ~A265 & A200;
  assign \new_[37218]_  = A199 & \new_[37217]_ ;
  assign \new_[37219]_  = \new_[37218]_  & \new_[37213]_ ;
  assign \new_[37223]_  = ~A268 & ~A267;
  assign \new_[37224]_  = A266 & \new_[37223]_ ;
  assign \new_[37228]_  = A299 & A298;
  assign \new_[37229]_  = ~A269 & \new_[37228]_ ;
  assign \new_[37230]_  = \new_[37229]_  & \new_[37224]_ ;
  assign \new_[37234]_  = A168 & ~A169;
  assign \new_[37235]_  = A170 & \new_[37234]_ ;
  assign \new_[37239]_  = ~A265 & A200;
  assign \new_[37240]_  = A199 & \new_[37239]_ ;
  assign \new_[37241]_  = \new_[37240]_  & \new_[37235]_ ;
  assign \new_[37245]_  = ~A268 & ~A267;
  assign \new_[37246]_  = A266 & \new_[37245]_ ;
  assign \new_[37250]_  = ~A299 & ~A298;
  assign \new_[37251]_  = ~A269 & \new_[37250]_ ;
  assign \new_[37252]_  = \new_[37251]_  & \new_[37246]_ ;
  assign \new_[37256]_  = A168 & ~A169;
  assign \new_[37257]_  = A170 & \new_[37256]_ ;
  assign \new_[37261]_  = A265 & A200;
  assign \new_[37262]_  = A199 & \new_[37261]_ ;
  assign \new_[37263]_  = \new_[37262]_  & \new_[37257]_ ;
  assign \new_[37267]_  = A268 & A267;
  assign \new_[37268]_  = ~A266 & \new_[37267]_ ;
  assign \new_[37272]_  = ~A302 & ~A301;
  assign \new_[37273]_  = A300 & \new_[37272]_ ;
  assign \new_[37274]_  = \new_[37273]_  & \new_[37268]_ ;
  assign \new_[37278]_  = A168 & ~A169;
  assign \new_[37279]_  = A170 & \new_[37278]_ ;
  assign \new_[37283]_  = A265 & A200;
  assign \new_[37284]_  = A199 & \new_[37283]_ ;
  assign \new_[37285]_  = \new_[37284]_  & \new_[37279]_ ;
  assign \new_[37289]_  = A269 & A267;
  assign \new_[37290]_  = ~A266 & \new_[37289]_ ;
  assign \new_[37294]_  = ~A302 & ~A301;
  assign \new_[37295]_  = A300 & \new_[37294]_ ;
  assign \new_[37296]_  = \new_[37295]_  & \new_[37290]_ ;
  assign \new_[37300]_  = A168 & ~A169;
  assign \new_[37301]_  = A170 & \new_[37300]_ ;
  assign \new_[37305]_  = A265 & A200;
  assign \new_[37306]_  = A199 & \new_[37305]_ ;
  assign \new_[37307]_  = \new_[37306]_  & \new_[37301]_ ;
  assign \new_[37311]_  = ~A268 & ~A267;
  assign \new_[37312]_  = ~A266 & \new_[37311]_ ;
  assign \new_[37316]_  = A301 & ~A300;
  assign \new_[37317]_  = ~A269 & \new_[37316]_ ;
  assign \new_[37318]_  = \new_[37317]_  & \new_[37312]_ ;
  assign \new_[37322]_  = A168 & ~A169;
  assign \new_[37323]_  = A170 & \new_[37322]_ ;
  assign \new_[37327]_  = A265 & A200;
  assign \new_[37328]_  = A199 & \new_[37327]_ ;
  assign \new_[37329]_  = \new_[37328]_  & \new_[37323]_ ;
  assign \new_[37333]_  = ~A268 & ~A267;
  assign \new_[37334]_  = ~A266 & \new_[37333]_ ;
  assign \new_[37338]_  = A302 & ~A300;
  assign \new_[37339]_  = ~A269 & \new_[37338]_ ;
  assign \new_[37340]_  = \new_[37339]_  & \new_[37334]_ ;
  assign \new_[37344]_  = A168 & ~A169;
  assign \new_[37345]_  = A170 & \new_[37344]_ ;
  assign \new_[37349]_  = A265 & A200;
  assign \new_[37350]_  = A199 & \new_[37349]_ ;
  assign \new_[37351]_  = \new_[37350]_  & \new_[37345]_ ;
  assign \new_[37355]_  = ~A268 & ~A267;
  assign \new_[37356]_  = ~A266 & \new_[37355]_ ;
  assign \new_[37360]_  = A299 & A298;
  assign \new_[37361]_  = ~A269 & \new_[37360]_ ;
  assign \new_[37362]_  = \new_[37361]_  & \new_[37356]_ ;
  assign \new_[37366]_  = A168 & ~A169;
  assign \new_[37367]_  = A170 & \new_[37366]_ ;
  assign \new_[37371]_  = A265 & A200;
  assign \new_[37372]_  = A199 & \new_[37371]_ ;
  assign \new_[37373]_  = \new_[37372]_  & \new_[37367]_ ;
  assign \new_[37377]_  = ~A268 & ~A267;
  assign \new_[37378]_  = ~A266 & \new_[37377]_ ;
  assign \new_[37382]_  = ~A299 & ~A298;
  assign \new_[37383]_  = ~A269 & \new_[37382]_ ;
  assign \new_[37384]_  = \new_[37383]_  & \new_[37378]_ ;
  assign \new_[37388]_  = A168 & ~A169;
  assign \new_[37389]_  = A170 & \new_[37388]_ ;
  assign \new_[37393]_  = ~A265 & ~A200;
  assign \new_[37394]_  = ~A199 & \new_[37393]_ ;
  assign \new_[37395]_  = \new_[37394]_  & \new_[37389]_ ;
  assign \new_[37399]_  = A268 & A267;
  assign \new_[37400]_  = A266 & \new_[37399]_ ;
  assign \new_[37404]_  = ~A302 & ~A301;
  assign \new_[37405]_  = A300 & \new_[37404]_ ;
  assign \new_[37406]_  = \new_[37405]_  & \new_[37400]_ ;
  assign \new_[37410]_  = A168 & ~A169;
  assign \new_[37411]_  = A170 & \new_[37410]_ ;
  assign \new_[37415]_  = ~A265 & ~A200;
  assign \new_[37416]_  = ~A199 & \new_[37415]_ ;
  assign \new_[37417]_  = \new_[37416]_  & \new_[37411]_ ;
  assign \new_[37421]_  = A269 & A267;
  assign \new_[37422]_  = A266 & \new_[37421]_ ;
  assign \new_[37426]_  = ~A302 & ~A301;
  assign \new_[37427]_  = A300 & \new_[37426]_ ;
  assign \new_[37428]_  = \new_[37427]_  & \new_[37422]_ ;
  assign \new_[37432]_  = A168 & ~A169;
  assign \new_[37433]_  = A170 & \new_[37432]_ ;
  assign \new_[37437]_  = ~A265 & ~A200;
  assign \new_[37438]_  = ~A199 & \new_[37437]_ ;
  assign \new_[37439]_  = \new_[37438]_  & \new_[37433]_ ;
  assign \new_[37443]_  = ~A268 & ~A267;
  assign \new_[37444]_  = A266 & \new_[37443]_ ;
  assign \new_[37448]_  = A301 & ~A300;
  assign \new_[37449]_  = ~A269 & \new_[37448]_ ;
  assign \new_[37450]_  = \new_[37449]_  & \new_[37444]_ ;
  assign \new_[37454]_  = A168 & ~A169;
  assign \new_[37455]_  = A170 & \new_[37454]_ ;
  assign \new_[37459]_  = ~A265 & ~A200;
  assign \new_[37460]_  = ~A199 & \new_[37459]_ ;
  assign \new_[37461]_  = \new_[37460]_  & \new_[37455]_ ;
  assign \new_[37465]_  = ~A268 & ~A267;
  assign \new_[37466]_  = A266 & \new_[37465]_ ;
  assign \new_[37470]_  = A302 & ~A300;
  assign \new_[37471]_  = ~A269 & \new_[37470]_ ;
  assign \new_[37472]_  = \new_[37471]_  & \new_[37466]_ ;
  assign \new_[37476]_  = A168 & ~A169;
  assign \new_[37477]_  = A170 & \new_[37476]_ ;
  assign \new_[37481]_  = ~A265 & ~A200;
  assign \new_[37482]_  = ~A199 & \new_[37481]_ ;
  assign \new_[37483]_  = \new_[37482]_  & \new_[37477]_ ;
  assign \new_[37487]_  = ~A268 & ~A267;
  assign \new_[37488]_  = A266 & \new_[37487]_ ;
  assign \new_[37492]_  = A299 & A298;
  assign \new_[37493]_  = ~A269 & \new_[37492]_ ;
  assign \new_[37494]_  = \new_[37493]_  & \new_[37488]_ ;
  assign \new_[37498]_  = A168 & ~A169;
  assign \new_[37499]_  = A170 & \new_[37498]_ ;
  assign \new_[37503]_  = ~A265 & ~A200;
  assign \new_[37504]_  = ~A199 & \new_[37503]_ ;
  assign \new_[37505]_  = \new_[37504]_  & \new_[37499]_ ;
  assign \new_[37509]_  = ~A268 & ~A267;
  assign \new_[37510]_  = A266 & \new_[37509]_ ;
  assign \new_[37514]_  = ~A299 & ~A298;
  assign \new_[37515]_  = ~A269 & \new_[37514]_ ;
  assign \new_[37516]_  = \new_[37515]_  & \new_[37510]_ ;
  assign \new_[37520]_  = A168 & ~A169;
  assign \new_[37521]_  = A170 & \new_[37520]_ ;
  assign \new_[37525]_  = A265 & ~A200;
  assign \new_[37526]_  = ~A199 & \new_[37525]_ ;
  assign \new_[37527]_  = \new_[37526]_  & \new_[37521]_ ;
  assign \new_[37531]_  = A268 & A267;
  assign \new_[37532]_  = ~A266 & \new_[37531]_ ;
  assign \new_[37536]_  = ~A302 & ~A301;
  assign \new_[37537]_  = A300 & \new_[37536]_ ;
  assign \new_[37538]_  = \new_[37537]_  & \new_[37532]_ ;
  assign \new_[37542]_  = A168 & ~A169;
  assign \new_[37543]_  = A170 & \new_[37542]_ ;
  assign \new_[37547]_  = A265 & ~A200;
  assign \new_[37548]_  = ~A199 & \new_[37547]_ ;
  assign \new_[37549]_  = \new_[37548]_  & \new_[37543]_ ;
  assign \new_[37553]_  = A269 & A267;
  assign \new_[37554]_  = ~A266 & \new_[37553]_ ;
  assign \new_[37558]_  = ~A302 & ~A301;
  assign \new_[37559]_  = A300 & \new_[37558]_ ;
  assign \new_[37560]_  = \new_[37559]_  & \new_[37554]_ ;
  assign \new_[37564]_  = A168 & ~A169;
  assign \new_[37565]_  = A170 & \new_[37564]_ ;
  assign \new_[37569]_  = A265 & ~A200;
  assign \new_[37570]_  = ~A199 & \new_[37569]_ ;
  assign \new_[37571]_  = \new_[37570]_  & \new_[37565]_ ;
  assign \new_[37575]_  = ~A268 & ~A267;
  assign \new_[37576]_  = ~A266 & \new_[37575]_ ;
  assign \new_[37580]_  = A301 & ~A300;
  assign \new_[37581]_  = ~A269 & \new_[37580]_ ;
  assign \new_[37582]_  = \new_[37581]_  & \new_[37576]_ ;
  assign \new_[37586]_  = A168 & ~A169;
  assign \new_[37587]_  = A170 & \new_[37586]_ ;
  assign \new_[37591]_  = A265 & ~A200;
  assign \new_[37592]_  = ~A199 & \new_[37591]_ ;
  assign \new_[37593]_  = \new_[37592]_  & \new_[37587]_ ;
  assign \new_[37597]_  = ~A268 & ~A267;
  assign \new_[37598]_  = ~A266 & \new_[37597]_ ;
  assign \new_[37602]_  = A302 & ~A300;
  assign \new_[37603]_  = ~A269 & \new_[37602]_ ;
  assign \new_[37604]_  = \new_[37603]_  & \new_[37598]_ ;
  assign \new_[37608]_  = A168 & ~A169;
  assign \new_[37609]_  = A170 & \new_[37608]_ ;
  assign \new_[37613]_  = A265 & ~A200;
  assign \new_[37614]_  = ~A199 & \new_[37613]_ ;
  assign \new_[37615]_  = \new_[37614]_  & \new_[37609]_ ;
  assign \new_[37619]_  = ~A268 & ~A267;
  assign \new_[37620]_  = ~A266 & \new_[37619]_ ;
  assign \new_[37624]_  = A299 & A298;
  assign \new_[37625]_  = ~A269 & \new_[37624]_ ;
  assign \new_[37626]_  = \new_[37625]_  & \new_[37620]_ ;
  assign \new_[37630]_  = A168 & ~A169;
  assign \new_[37631]_  = A170 & \new_[37630]_ ;
  assign \new_[37635]_  = A265 & ~A200;
  assign \new_[37636]_  = ~A199 & \new_[37635]_ ;
  assign \new_[37637]_  = \new_[37636]_  & \new_[37631]_ ;
  assign \new_[37641]_  = ~A268 & ~A267;
  assign \new_[37642]_  = ~A266 & \new_[37641]_ ;
  assign \new_[37646]_  = ~A299 & ~A298;
  assign \new_[37647]_  = ~A269 & \new_[37646]_ ;
  assign \new_[37648]_  = \new_[37647]_  & \new_[37642]_ ;
  assign \new_[37652]_  = A201 & A166;
  assign \new_[37653]_  = A167 & \new_[37652]_ ;
  assign \new_[37657]_  = ~A265 & ~A203;
  assign \new_[37658]_  = ~A202 & \new_[37657]_ ;
  assign \new_[37659]_  = \new_[37658]_  & \new_[37653]_ ;
  assign \new_[37663]_  = ~A268 & ~A267;
  assign \new_[37664]_  = A266 & \new_[37663]_ ;
  assign \new_[37667]_  = A300 & ~A269;
  assign \new_[37670]_  = ~A302 & ~A301;
  assign \new_[37671]_  = \new_[37670]_  & \new_[37667]_ ;
  assign \new_[37672]_  = \new_[37671]_  & \new_[37664]_ ;
  assign \new_[37676]_  = A201 & A166;
  assign \new_[37677]_  = A167 & \new_[37676]_ ;
  assign \new_[37681]_  = A265 & ~A203;
  assign \new_[37682]_  = ~A202 & \new_[37681]_ ;
  assign \new_[37683]_  = \new_[37682]_  & \new_[37677]_ ;
  assign \new_[37687]_  = ~A268 & ~A267;
  assign \new_[37688]_  = ~A266 & \new_[37687]_ ;
  assign \new_[37691]_  = A300 & ~A269;
  assign \new_[37694]_  = ~A302 & ~A301;
  assign \new_[37695]_  = \new_[37694]_  & \new_[37691]_ ;
  assign \new_[37696]_  = \new_[37695]_  & \new_[37688]_ ;
  assign \new_[37700]_  = ~A199 & A166;
  assign \new_[37701]_  = A167 & \new_[37700]_ ;
  assign \new_[37705]_  = A202 & A201;
  assign \new_[37706]_  = A200 & \new_[37705]_ ;
  assign \new_[37707]_  = \new_[37706]_  & \new_[37701]_ ;
  assign \new_[37711]_  = ~A269 & ~A268;
  assign \new_[37712]_  = A267 & \new_[37711]_ ;
  assign \new_[37715]_  = ~A299 & A298;
  assign \new_[37718]_  = A301 & A300;
  assign \new_[37719]_  = \new_[37718]_  & \new_[37715]_ ;
  assign \new_[37720]_  = \new_[37719]_  & \new_[37712]_ ;
  assign \new_[37724]_  = ~A199 & A166;
  assign \new_[37725]_  = A167 & \new_[37724]_ ;
  assign \new_[37729]_  = A202 & A201;
  assign \new_[37730]_  = A200 & \new_[37729]_ ;
  assign \new_[37731]_  = \new_[37730]_  & \new_[37725]_ ;
  assign \new_[37735]_  = ~A269 & ~A268;
  assign \new_[37736]_  = A267 & \new_[37735]_ ;
  assign \new_[37739]_  = ~A299 & A298;
  assign \new_[37742]_  = A302 & A300;
  assign \new_[37743]_  = \new_[37742]_  & \new_[37739]_ ;
  assign \new_[37744]_  = \new_[37743]_  & \new_[37736]_ ;
  assign \new_[37748]_  = ~A199 & A166;
  assign \new_[37749]_  = A167 & \new_[37748]_ ;
  assign \new_[37753]_  = A202 & A201;
  assign \new_[37754]_  = A200 & \new_[37753]_ ;
  assign \new_[37755]_  = \new_[37754]_  & \new_[37749]_ ;
  assign \new_[37759]_  = ~A269 & ~A268;
  assign \new_[37760]_  = A267 & \new_[37759]_ ;
  assign \new_[37763]_  = A299 & ~A298;
  assign \new_[37766]_  = A301 & A300;
  assign \new_[37767]_  = \new_[37766]_  & \new_[37763]_ ;
  assign \new_[37768]_  = \new_[37767]_  & \new_[37760]_ ;
  assign \new_[37772]_  = ~A199 & A166;
  assign \new_[37773]_  = A167 & \new_[37772]_ ;
  assign \new_[37777]_  = A202 & A201;
  assign \new_[37778]_  = A200 & \new_[37777]_ ;
  assign \new_[37779]_  = \new_[37778]_  & \new_[37773]_ ;
  assign \new_[37783]_  = ~A269 & ~A268;
  assign \new_[37784]_  = A267 & \new_[37783]_ ;
  assign \new_[37787]_  = A299 & ~A298;
  assign \new_[37790]_  = A302 & A300;
  assign \new_[37791]_  = \new_[37790]_  & \new_[37787]_ ;
  assign \new_[37792]_  = \new_[37791]_  & \new_[37784]_ ;
  assign \new_[37796]_  = ~A199 & A166;
  assign \new_[37797]_  = A167 & \new_[37796]_ ;
  assign \new_[37801]_  = A202 & A201;
  assign \new_[37802]_  = A200 & \new_[37801]_ ;
  assign \new_[37803]_  = \new_[37802]_  & \new_[37797]_ ;
  assign \new_[37807]_  = A298 & A268;
  assign \new_[37808]_  = ~A267 & \new_[37807]_ ;
  assign \new_[37811]_  = ~A300 & ~A299;
  assign \new_[37814]_  = ~A302 & ~A301;
  assign \new_[37815]_  = \new_[37814]_  & \new_[37811]_ ;
  assign \new_[37816]_  = \new_[37815]_  & \new_[37808]_ ;
  assign \new_[37820]_  = ~A199 & A166;
  assign \new_[37821]_  = A167 & \new_[37820]_ ;
  assign \new_[37825]_  = A202 & A201;
  assign \new_[37826]_  = A200 & \new_[37825]_ ;
  assign \new_[37827]_  = \new_[37826]_  & \new_[37821]_ ;
  assign \new_[37831]_  = ~A298 & A268;
  assign \new_[37832]_  = ~A267 & \new_[37831]_ ;
  assign \new_[37835]_  = ~A300 & A299;
  assign \new_[37838]_  = ~A302 & ~A301;
  assign \new_[37839]_  = \new_[37838]_  & \new_[37835]_ ;
  assign \new_[37840]_  = \new_[37839]_  & \new_[37832]_ ;
  assign \new_[37844]_  = ~A199 & A166;
  assign \new_[37845]_  = A167 & \new_[37844]_ ;
  assign \new_[37849]_  = A202 & A201;
  assign \new_[37850]_  = A200 & \new_[37849]_ ;
  assign \new_[37851]_  = \new_[37850]_  & \new_[37845]_ ;
  assign \new_[37855]_  = A298 & A269;
  assign \new_[37856]_  = ~A267 & \new_[37855]_ ;
  assign \new_[37859]_  = ~A300 & ~A299;
  assign \new_[37862]_  = ~A302 & ~A301;
  assign \new_[37863]_  = \new_[37862]_  & \new_[37859]_ ;
  assign \new_[37864]_  = \new_[37863]_  & \new_[37856]_ ;
  assign \new_[37868]_  = ~A199 & A166;
  assign \new_[37869]_  = A167 & \new_[37868]_ ;
  assign \new_[37873]_  = A202 & A201;
  assign \new_[37874]_  = A200 & \new_[37873]_ ;
  assign \new_[37875]_  = \new_[37874]_  & \new_[37869]_ ;
  assign \new_[37879]_  = ~A298 & A269;
  assign \new_[37880]_  = ~A267 & \new_[37879]_ ;
  assign \new_[37883]_  = ~A300 & A299;
  assign \new_[37886]_  = ~A302 & ~A301;
  assign \new_[37887]_  = \new_[37886]_  & \new_[37883]_ ;
  assign \new_[37888]_  = \new_[37887]_  & \new_[37880]_ ;
  assign \new_[37892]_  = ~A199 & A166;
  assign \new_[37893]_  = A167 & \new_[37892]_ ;
  assign \new_[37897]_  = A202 & A201;
  assign \new_[37898]_  = A200 & \new_[37897]_ ;
  assign \new_[37899]_  = \new_[37898]_  & \new_[37893]_ ;
  assign \new_[37903]_  = A298 & A266;
  assign \new_[37904]_  = A265 & \new_[37903]_ ;
  assign \new_[37907]_  = ~A300 & ~A299;
  assign \new_[37910]_  = ~A302 & ~A301;
  assign \new_[37911]_  = \new_[37910]_  & \new_[37907]_ ;
  assign \new_[37912]_  = \new_[37911]_  & \new_[37904]_ ;
  assign \new_[37916]_  = ~A199 & A166;
  assign \new_[37917]_  = A167 & \new_[37916]_ ;
  assign \new_[37921]_  = A202 & A201;
  assign \new_[37922]_  = A200 & \new_[37921]_ ;
  assign \new_[37923]_  = \new_[37922]_  & \new_[37917]_ ;
  assign \new_[37927]_  = ~A298 & A266;
  assign \new_[37928]_  = A265 & \new_[37927]_ ;
  assign \new_[37931]_  = ~A300 & A299;
  assign \new_[37934]_  = ~A302 & ~A301;
  assign \new_[37935]_  = \new_[37934]_  & \new_[37931]_ ;
  assign \new_[37936]_  = \new_[37935]_  & \new_[37928]_ ;
  assign \new_[37940]_  = ~A199 & A166;
  assign \new_[37941]_  = A167 & \new_[37940]_ ;
  assign \new_[37945]_  = A202 & A201;
  assign \new_[37946]_  = A200 & \new_[37945]_ ;
  assign \new_[37947]_  = \new_[37946]_  & \new_[37941]_ ;
  assign \new_[37951]_  = A298 & ~A266;
  assign \new_[37952]_  = ~A265 & \new_[37951]_ ;
  assign \new_[37955]_  = ~A300 & ~A299;
  assign \new_[37958]_  = ~A302 & ~A301;
  assign \new_[37959]_  = \new_[37958]_  & \new_[37955]_ ;
  assign \new_[37960]_  = \new_[37959]_  & \new_[37952]_ ;
  assign \new_[37964]_  = ~A199 & A166;
  assign \new_[37965]_  = A167 & \new_[37964]_ ;
  assign \new_[37969]_  = A202 & A201;
  assign \new_[37970]_  = A200 & \new_[37969]_ ;
  assign \new_[37971]_  = \new_[37970]_  & \new_[37965]_ ;
  assign \new_[37975]_  = ~A298 & ~A266;
  assign \new_[37976]_  = ~A265 & \new_[37975]_ ;
  assign \new_[37979]_  = ~A300 & A299;
  assign \new_[37982]_  = ~A302 & ~A301;
  assign \new_[37983]_  = \new_[37982]_  & \new_[37979]_ ;
  assign \new_[37984]_  = \new_[37983]_  & \new_[37976]_ ;
  assign \new_[37988]_  = ~A199 & A166;
  assign \new_[37989]_  = A167 & \new_[37988]_ ;
  assign \new_[37993]_  = A203 & A201;
  assign \new_[37994]_  = A200 & \new_[37993]_ ;
  assign \new_[37995]_  = \new_[37994]_  & \new_[37989]_ ;
  assign \new_[37999]_  = ~A269 & ~A268;
  assign \new_[38000]_  = A267 & \new_[37999]_ ;
  assign \new_[38003]_  = ~A299 & A298;
  assign \new_[38006]_  = A301 & A300;
  assign \new_[38007]_  = \new_[38006]_  & \new_[38003]_ ;
  assign \new_[38008]_  = \new_[38007]_  & \new_[38000]_ ;
  assign \new_[38012]_  = ~A199 & A166;
  assign \new_[38013]_  = A167 & \new_[38012]_ ;
  assign \new_[38017]_  = A203 & A201;
  assign \new_[38018]_  = A200 & \new_[38017]_ ;
  assign \new_[38019]_  = \new_[38018]_  & \new_[38013]_ ;
  assign \new_[38023]_  = ~A269 & ~A268;
  assign \new_[38024]_  = A267 & \new_[38023]_ ;
  assign \new_[38027]_  = ~A299 & A298;
  assign \new_[38030]_  = A302 & A300;
  assign \new_[38031]_  = \new_[38030]_  & \new_[38027]_ ;
  assign \new_[38032]_  = \new_[38031]_  & \new_[38024]_ ;
  assign \new_[38036]_  = ~A199 & A166;
  assign \new_[38037]_  = A167 & \new_[38036]_ ;
  assign \new_[38041]_  = A203 & A201;
  assign \new_[38042]_  = A200 & \new_[38041]_ ;
  assign \new_[38043]_  = \new_[38042]_  & \new_[38037]_ ;
  assign \new_[38047]_  = ~A269 & ~A268;
  assign \new_[38048]_  = A267 & \new_[38047]_ ;
  assign \new_[38051]_  = A299 & ~A298;
  assign \new_[38054]_  = A301 & A300;
  assign \new_[38055]_  = \new_[38054]_  & \new_[38051]_ ;
  assign \new_[38056]_  = \new_[38055]_  & \new_[38048]_ ;
  assign \new_[38060]_  = ~A199 & A166;
  assign \new_[38061]_  = A167 & \new_[38060]_ ;
  assign \new_[38065]_  = A203 & A201;
  assign \new_[38066]_  = A200 & \new_[38065]_ ;
  assign \new_[38067]_  = \new_[38066]_  & \new_[38061]_ ;
  assign \new_[38071]_  = ~A269 & ~A268;
  assign \new_[38072]_  = A267 & \new_[38071]_ ;
  assign \new_[38075]_  = A299 & ~A298;
  assign \new_[38078]_  = A302 & A300;
  assign \new_[38079]_  = \new_[38078]_  & \new_[38075]_ ;
  assign \new_[38080]_  = \new_[38079]_  & \new_[38072]_ ;
  assign \new_[38084]_  = ~A199 & A166;
  assign \new_[38085]_  = A167 & \new_[38084]_ ;
  assign \new_[38089]_  = A203 & A201;
  assign \new_[38090]_  = A200 & \new_[38089]_ ;
  assign \new_[38091]_  = \new_[38090]_  & \new_[38085]_ ;
  assign \new_[38095]_  = A298 & A268;
  assign \new_[38096]_  = ~A267 & \new_[38095]_ ;
  assign \new_[38099]_  = ~A300 & ~A299;
  assign \new_[38102]_  = ~A302 & ~A301;
  assign \new_[38103]_  = \new_[38102]_  & \new_[38099]_ ;
  assign \new_[38104]_  = \new_[38103]_  & \new_[38096]_ ;
  assign \new_[38108]_  = ~A199 & A166;
  assign \new_[38109]_  = A167 & \new_[38108]_ ;
  assign \new_[38113]_  = A203 & A201;
  assign \new_[38114]_  = A200 & \new_[38113]_ ;
  assign \new_[38115]_  = \new_[38114]_  & \new_[38109]_ ;
  assign \new_[38119]_  = ~A298 & A268;
  assign \new_[38120]_  = ~A267 & \new_[38119]_ ;
  assign \new_[38123]_  = ~A300 & A299;
  assign \new_[38126]_  = ~A302 & ~A301;
  assign \new_[38127]_  = \new_[38126]_  & \new_[38123]_ ;
  assign \new_[38128]_  = \new_[38127]_  & \new_[38120]_ ;
  assign \new_[38132]_  = ~A199 & A166;
  assign \new_[38133]_  = A167 & \new_[38132]_ ;
  assign \new_[38137]_  = A203 & A201;
  assign \new_[38138]_  = A200 & \new_[38137]_ ;
  assign \new_[38139]_  = \new_[38138]_  & \new_[38133]_ ;
  assign \new_[38143]_  = A298 & A269;
  assign \new_[38144]_  = ~A267 & \new_[38143]_ ;
  assign \new_[38147]_  = ~A300 & ~A299;
  assign \new_[38150]_  = ~A302 & ~A301;
  assign \new_[38151]_  = \new_[38150]_  & \new_[38147]_ ;
  assign \new_[38152]_  = \new_[38151]_  & \new_[38144]_ ;
  assign \new_[38156]_  = ~A199 & A166;
  assign \new_[38157]_  = A167 & \new_[38156]_ ;
  assign \new_[38161]_  = A203 & A201;
  assign \new_[38162]_  = A200 & \new_[38161]_ ;
  assign \new_[38163]_  = \new_[38162]_  & \new_[38157]_ ;
  assign \new_[38167]_  = ~A298 & A269;
  assign \new_[38168]_  = ~A267 & \new_[38167]_ ;
  assign \new_[38171]_  = ~A300 & A299;
  assign \new_[38174]_  = ~A302 & ~A301;
  assign \new_[38175]_  = \new_[38174]_  & \new_[38171]_ ;
  assign \new_[38176]_  = \new_[38175]_  & \new_[38168]_ ;
  assign \new_[38180]_  = ~A199 & A166;
  assign \new_[38181]_  = A167 & \new_[38180]_ ;
  assign \new_[38185]_  = A203 & A201;
  assign \new_[38186]_  = A200 & \new_[38185]_ ;
  assign \new_[38187]_  = \new_[38186]_  & \new_[38181]_ ;
  assign \new_[38191]_  = A298 & A266;
  assign \new_[38192]_  = A265 & \new_[38191]_ ;
  assign \new_[38195]_  = ~A300 & ~A299;
  assign \new_[38198]_  = ~A302 & ~A301;
  assign \new_[38199]_  = \new_[38198]_  & \new_[38195]_ ;
  assign \new_[38200]_  = \new_[38199]_  & \new_[38192]_ ;
  assign \new_[38204]_  = ~A199 & A166;
  assign \new_[38205]_  = A167 & \new_[38204]_ ;
  assign \new_[38209]_  = A203 & A201;
  assign \new_[38210]_  = A200 & \new_[38209]_ ;
  assign \new_[38211]_  = \new_[38210]_  & \new_[38205]_ ;
  assign \new_[38215]_  = ~A298 & A266;
  assign \new_[38216]_  = A265 & \new_[38215]_ ;
  assign \new_[38219]_  = ~A300 & A299;
  assign \new_[38222]_  = ~A302 & ~A301;
  assign \new_[38223]_  = \new_[38222]_  & \new_[38219]_ ;
  assign \new_[38224]_  = \new_[38223]_  & \new_[38216]_ ;
  assign \new_[38228]_  = ~A199 & A166;
  assign \new_[38229]_  = A167 & \new_[38228]_ ;
  assign \new_[38233]_  = A203 & A201;
  assign \new_[38234]_  = A200 & \new_[38233]_ ;
  assign \new_[38235]_  = \new_[38234]_  & \new_[38229]_ ;
  assign \new_[38239]_  = A298 & ~A266;
  assign \new_[38240]_  = ~A265 & \new_[38239]_ ;
  assign \new_[38243]_  = ~A300 & ~A299;
  assign \new_[38246]_  = ~A302 & ~A301;
  assign \new_[38247]_  = \new_[38246]_  & \new_[38243]_ ;
  assign \new_[38248]_  = \new_[38247]_  & \new_[38240]_ ;
  assign \new_[38252]_  = ~A199 & A166;
  assign \new_[38253]_  = A167 & \new_[38252]_ ;
  assign \new_[38257]_  = A203 & A201;
  assign \new_[38258]_  = A200 & \new_[38257]_ ;
  assign \new_[38259]_  = \new_[38258]_  & \new_[38253]_ ;
  assign \new_[38263]_  = ~A298 & ~A266;
  assign \new_[38264]_  = ~A265 & \new_[38263]_ ;
  assign \new_[38267]_  = ~A300 & A299;
  assign \new_[38270]_  = ~A302 & ~A301;
  assign \new_[38271]_  = \new_[38270]_  & \new_[38267]_ ;
  assign \new_[38272]_  = \new_[38271]_  & \new_[38264]_ ;
  assign \new_[38276]_  = ~A199 & A166;
  assign \new_[38277]_  = A167 & \new_[38276]_ ;
  assign \new_[38281]_  = ~A202 & ~A201;
  assign \new_[38282]_  = A200 & \new_[38281]_ ;
  assign \new_[38283]_  = \new_[38282]_  & \new_[38277]_ ;
  assign \new_[38287]_  = A268 & ~A267;
  assign \new_[38288]_  = ~A203 & \new_[38287]_ ;
  assign \new_[38291]_  = ~A299 & A298;
  assign \new_[38294]_  = A301 & A300;
  assign \new_[38295]_  = \new_[38294]_  & \new_[38291]_ ;
  assign \new_[38296]_  = \new_[38295]_  & \new_[38288]_ ;
  assign \new_[38300]_  = ~A199 & A166;
  assign \new_[38301]_  = A167 & \new_[38300]_ ;
  assign \new_[38305]_  = ~A202 & ~A201;
  assign \new_[38306]_  = A200 & \new_[38305]_ ;
  assign \new_[38307]_  = \new_[38306]_  & \new_[38301]_ ;
  assign \new_[38311]_  = A268 & ~A267;
  assign \new_[38312]_  = ~A203 & \new_[38311]_ ;
  assign \new_[38315]_  = ~A299 & A298;
  assign \new_[38318]_  = A302 & A300;
  assign \new_[38319]_  = \new_[38318]_  & \new_[38315]_ ;
  assign \new_[38320]_  = \new_[38319]_  & \new_[38312]_ ;
  assign \new_[38324]_  = ~A199 & A166;
  assign \new_[38325]_  = A167 & \new_[38324]_ ;
  assign \new_[38329]_  = ~A202 & ~A201;
  assign \new_[38330]_  = A200 & \new_[38329]_ ;
  assign \new_[38331]_  = \new_[38330]_  & \new_[38325]_ ;
  assign \new_[38335]_  = A268 & ~A267;
  assign \new_[38336]_  = ~A203 & \new_[38335]_ ;
  assign \new_[38339]_  = A299 & ~A298;
  assign \new_[38342]_  = A301 & A300;
  assign \new_[38343]_  = \new_[38342]_  & \new_[38339]_ ;
  assign \new_[38344]_  = \new_[38343]_  & \new_[38336]_ ;
  assign \new_[38348]_  = ~A199 & A166;
  assign \new_[38349]_  = A167 & \new_[38348]_ ;
  assign \new_[38353]_  = ~A202 & ~A201;
  assign \new_[38354]_  = A200 & \new_[38353]_ ;
  assign \new_[38355]_  = \new_[38354]_  & \new_[38349]_ ;
  assign \new_[38359]_  = A268 & ~A267;
  assign \new_[38360]_  = ~A203 & \new_[38359]_ ;
  assign \new_[38363]_  = A299 & ~A298;
  assign \new_[38366]_  = A302 & A300;
  assign \new_[38367]_  = \new_[38366]_  & \new_[38363]_ ;
  assign \new_[38368]_  = \new_[38367]_  & \new_[38360]_ ;
  assign \new_[38372]_  = ~A199 & A166;
  assign \new_[38373]_  = A167 & \new_[38372]_ ;
  assign \new_[38377]_  = ~A202 & ~A201;
  assign \new_[38378]_  = A200 & \new_[38377]_ ;
  assign \new_[38379]_  = \new_[38378]_  & \new_[38373]_ ;
  assign \new_[38383]_  = A269 & ~A267;
  assign \new_[38384]_  = ~A203 & \new_[38383]_ ;
  assign \new_[38387]_  = ~A299 & A298;
  assign \new_[38390]_  = A301 & A300;
  assign \new_[38391]_  = \new_[38390]_  & \new_[38387]_ ;
  assign \new_[38392]_  = \new_[38391]_  & \new_[38384]_ ;
  assign \new_[38396]_  = ~A199 & A166;
  assign \new_[38397]_  = A167 & \new_[38396]_ ;
  assign \new_[38401]_  = ~A202 & ~A201;
  assign \new_[38402]_  = A200 & \new_[38401]_ ;
  assign \new_[38403]_  = \new_[38402]_  & \new_[38397]_ ;
  assign \new_[38407]_  = A269 & ~A267;
  assign \new_[38408]_  = ~A203 & \new_[38407]_ ;
  assign \new_[38411]_  = ~A299 & A298;
  assign \new_[38414]_  = A302 & A300;
  assign \new_[38415]_  = \new_[38414]_  & \new_[38411]_ ;
  assign \new_[38416]_  = \new_[38415]_  & \new_[38408]_ ;
  assign \new_[38420]_  = ~A199 & A166;
  assign \new_[38421]_  = A167 & \new_[38420]_ ;
  assign \new_[38425]_  = ~A202 & ~A201;
  assign \new_[38426]_  = A200 & \new_[38425]_ ;
  assign \new_[38427]_  = \new_[38426]_  & \new_[38421]_ ;
  assign \new_[38431]_  = A269 & ~A267;
  assign \new_[38432]_  = ~A203 & \new_[38431]_ ;
  assign \new_[38435]_  = A299 & ~A298;
  assign \new_[38438]_  = A301 & A300;
  assign \new_[38439]_  = \new_[38438]_  & \new_[38435]_ ;
  assign \new_[38440]_  = \new_[38439]_  & \new_[38432]_ ;
  assign \new_[38444]_  = ~A199 & A166;
  assign \new_[38445]_  = A167 & \new_[38444]_ ;
  assign \new_[38449]_  = ~A202 & ~A201;
  assign \new_[38450]_  = A200 & \new_[38449]_ ;
  assign \new_[38451]_  = \new_[38450]_  & \new_[38445]_ ;
  assign \new_[38455]_  = A269 & ~A267;
  assign \new_[38456]_  = ~A203 & \new_[38455]_ ;
  assign \new_[38459]_  = A299 & ~A298;
  assign \new_[38462]_  = A302 & A300;
  assign \new_[38463]_  = \new_[38462]_  & \new_[38459]_ ;
  assign \new_[38464]_  = \new_[38463]_  & \new_[38456]_ ;
  assign \new_[38468]_  = ~A199 & A166;
  assign \new_[38469]_  = A167 & \new_[38468]_ ;
  assign \new_[38473]_  = ~A202 & ~A201;
  assign \new_[38474]_  = A200 & \new_[38473]_ ;
  assign \new_[38475]_  = \new_[38474]_  & \new_[38469]_ ;
  assign \new_[38479]_  = A266 & A265;
  assign \new_[38480]_  = ~A203 & \new_[38479]_ ;
  assign \new_[38483]_  = ~A299 & A298;
  assign \new_[38486]_  = A301 & A300;
  assign \new_[38487]_  = \new_[38486]_  & \new_[38483]_ ;
  assign \new_[38488]_  = \new_[38487]_  & \new_[38480]_ ;
  assign \new_[38492]_  = ~A199 & A166;
  assign \new_[38493]_  = A167 & \new_[38492]_ ;
  assign \new_[38497]_  = ~A202 & ~A201;
  assign \new_[38498]_  = A200 & \new_[38497]_ ;
  assign \new_[38499]_  = \new_[38498]_  & \new_[38493]_ ;
  assign \new_[38503]_  = A266 & A265;
  assign \new_[38504]_  = ~A203 & \new_[38503]_ ;
  assign \new_[38507]_  = ~A299 & A298;
  assign \new_[38510]_  = A302 & A300;
  assign \new_[38511]_  = \new_[38510]_  & \new_[38507]_ ;
  assign \new_[38512]_  = \new_[38511]_  & \new_[38504]_ ;
  assign \new_[38516]_  = ~A199 & A166;
  assign \new_[38517]_  = A167 & \new_[38516]_ ;
  assign \new_[38521]_  = ~A202 & ~A201;
  assign \new_[38522]_  = A200 & \new_[38521]_ ;
  assign \new_[38523]_  = \new_[38522]_  & \new_[38517]_ ;
  assign \new_[38527]_  = A266 & A265;
  assign \new_[38528]_  = ~A203 & \new_[38527]_ ;
  assign \new_[38531]_  = A299 & ~A298;
  assign \new_[38534]_  = A301 & A300;
  assign \new_[38535]_  = \new_[38534]_  & \new_[38531]_ ;
  assign \new_[38536]_  = \new_[38535]_  & \new_[38528]_ ;
  assign \new_[38540]_  = ~A199 & A166;
  assign \new_[38541]_  = A167 & \new_[38540]_ ;
  assign \new_[38545]_  = ~A202 & ~A201;
  assign \new_[38546]_  = A200 & \new_[38545]_ ;
  assign \new_[38547]_  = \new_[38546]_  & \new_[38541]_ ;
  assign \new_[38551]_  = A266 & A265;
  assign \new_[38552]_  = ~A203 & \new_[38551]_ ;
  assign \new_[38555]_  = A299 & ~A298;
  assign \new_[38558]_  = A302 & A300;
  assign \new_[38559]_  = \new_[38558]_  & \new_[38555]_ ;
  assign \new_[38560]_  = \new_[38559]_  & \new_[38552]_ ;
  assign \new_[38564]_  = ~A199 & A166;
  assign \new_[38565]_  = A167 & \new_[38564]_ ;
  assign \new_[38569]_  = ~A202 & ~A201;
  assign \new_[38570]_  = A200 & \new_[38569]_ ;
  assign \new_[38571]_  = \new_[38570]_  & \new_[38565]_ ;
  assign \new_[38575]_  = ~A266 & ~A265;
  assign \new_[38576]_  = ~A203 & \new_[38575]_ ;
  assign \new_[38579]_  = ~A299 & A298;
  assign \new_[38582]_  = A301 & A300;
  assign \new_[38583]_  = \new_[38582]_  & \new_[38579]_ ;
  assign \new_[38584]_  = \new_[38583]_  & \new_[38576]_ ;
  assign \new_[38588]_  = ~A199 & A166;
  assign \new_[38589]_  = A167 & \new_[38588]_ ;
  assign \new_[38593]_  = ~A202 & ~A201;
  assign \new_[38594]_  = A200 & \new_[38593]_ ;
  assign \new_[38595]_  = \new_[38594]_  & \new_[38589]_ ;
  assign \new_[38599]_  = ~A266 & ~A265;
  assign \new_[38600]_  = ~A203 & \new_[38599]_ ;
  assign \new_[38603]_  = ~A299 & A298;
  assign \new_[38606]_  = A302 & A300;
  assign \new_[38607]_  = \new_[38606]_  & \new_[38603]_ ;
  assign \new_[38608]_  = \new_[38607]_  & \new_[38600]_ ;
  assign \new_[38612]_  = ~A199 & A166;
  assign \new_[38613]_  = A167 & \new_[38612]_ ;
  assign \new_[38617]_  = ~A202 & ~A201;
  assign \new_[38618]_  = A200 & \new_[38617]_ ;
  assign \new_[38619]_  = \new_[38618]_  & \new_[38613]_ ;
  assign \new_[38623]_  = ~A266 & ~A265;
  assign \new_[38624]_  = ~A203 & \new_[38623]_ ;
  assign \new_[38627]_  = A299 & ~A298;
  assign \new_[38630]_  = A301 & A300;
  assign \new_[38631]_  = \new_[38630]_  & \new_[38627]_ ;
  assign \new_[38632]_  = \new_[38631]_  & \new_[38624]_ ;
  assign \new_[38636]_  = ~A199 & A166;
  assign \new_[38637]_  = A167 & \new_[38636]_ ;
  assign \new_[38641]_  = ~A202 & ~A201;
  assign \new_[38642]_  = A200 & \new_[38641]_ ;
  assign \new_[38643]_  = \new_[38642]_  & \new_[38637]_ ;
  assign \new_[38647]_  = ~A266 & ~A265;
  assign \new_[38648]_  = ~A203 & \new_[38647]_ ;
  assign \new_[38651]_  = A299 & ~A298;
  assign \new_[38654]_  = A302 & A300;
  assign \new_[38655]_  = \new_[38654]_  & \new_[38651]_ ;
  assign \new_[38656]_  = \new_[38655]_  & \new_[38648]_ ;
  assign \new_[38660]_  = A199 & A166;
  assign \new_[38661]_  = A167 & \new_[38660]_ ;
  assign \new_[38665]_  = A202 & A201;
  assign \new_[38666]_  = ~A200 & \new_[38665]_ ;
  assign \new_[38667]_  = \new_[38666]_  & \new_[38661]_ ;
  assign \new_[38671]_  = ~A269 & ~A268;
  assign \new_[38672]_  = A267 & \new_[38671]_ ;
  assign \new_[38675]_  = ~A299 & A298;
  assign \new_[38678]_  = A301 & A300;
  assign \new_[38679]_  = \new_[38678]_  & \new_[38675]_ ;
  assign \new_[38680]_  = \new_[38679]_  & \new_[38672]_ ;
  assign \new_[38684]_  = A199 & A166;
  assign \new_[38685]_  = A167 & \new_[38684]_ ;
  assign \new_[38689]_  = A202 & A201;
  assign \new_[38690]_  = ~A200 & \new_[38689]_ ;
  assign \new_[38691]_  = \new_[38690]_  & \new_[38685]_ ;
  assign \new_[38695]_  = ~A269 & ~A268;
  assign \new_[38696]_  = A267 & \new_[38695]_ ;
  assign \new_[38699]_  = ~A299 & A298;
  assign \new_[38702]_  = A302 & A300;
  assign \new_[38703]_  = \new_[38702]_  & \new_[38699]_ ;
  assign \new_[38704]_  = \new_[38703]_  & \new_[38696]_ ;
  assign \new_[38708]_  = A199 & A166;
  assign \new_[38709]_  = A167 & \new_[38708]_ ;
  assign \new_[38713]_  = A202 & A201;
  assign \new_[38714]_  = ~A200 & \new_[38713]_ ;
  assign \new_[38715]_  = \new_[38714]_  & \new_[38709]_ ;
  assign \new_[38719]_  = ~A269 & ~A268;
  assign \new_[38720]_  = A267 & \new_[38719]_ ;
  assign \new_[38723]_  = A299 & ~A298;
  assign \new_[38726]_  = A301 & A300;
  assign \new_[38727]_  = \new_[38726]_  & \new_[38723]_ ;
  assign \new_[38728]_  = \new_[38727]_  & \new_[38720]_ ;
  assign \new_[38732]_  = A199 & A166;
  assign \new_[38733]_  = A167 & \new_[38732]_ ;
  assign \new_[38737]_  = A202 & A201;
  assign \new_[38738]_  = ~A200 & \new_[38737]_ ;
  assign \new_[38739]_  = \new_[38738]_  & \new_[38733]_ ;
  assign \new_[38743]_  = ~A269 & ~A268;
  assign \new_[38744]_  = A267 & \new_[38743]_ ;
  assign \new_[38747]_  = A299 & ~A298;
  assign \new_[38750]_  = A302 & A300;
  assign \new_[38751]_  = \new_[38750]_  & \new_[38747]_ ;
  assign \new_[38752]_  = \new_[38751]_  & \new_[38744]_ ;
  assign \new_[38756]_  = A199 & A166;
  assign \new_[38757]_  = A167 & \new_[38756]_ ;
  assign \new_[38761]_  = A202 & A201;
  assign \new_[38762]_  = ~A200 & \new_[38761]_ ;
  assign \new_[38763]_  = \new_[38762]_  & \new_[38757]_ ;
  assign \new_[38767]_  = A298 & A268;
  assign \new_[38768]_  = ~A267 & \new_[38767]_ ;
  assign \new_[38771]_  = ~A300 & ~A299;
  assign \new_[38774]_  = ~A302 & ~A301;
  assign \new_[38775]_  = \new_[38774]_  & \new_[38771]_ ;
  assign \new_[38776]_  = \new_[38775]_  & \new_[38768]_ ;
  assign \new_[38780]_  = A199 & A166;
  assign \new_[38781]_  = A167 & \new_[38780]_ ;
  assign \new_[38785]_  = A202 & A201;
  assign \new_[38786]_  = ~A200 & \new_[38785]_ ;
  assign \new_[38787]_  = \new_[38786]_  & \new_[38781]_ ;
  assign \new_[38791]_  = ~A298 & A268;
  assign \new_[38792]_  = ~A267 & \new_[38791]_ ;
  assign \new_[38795]_  = ~A300 & A299;
  assign \new_[38798]_  = ~A302 & ~A301;
  assign \new_[38799]_  = \new_[38798]_  & \new_[38795]_ ;
  assign \new_[38800]_  = \new_[38799]_  & \new_[38792]_ ;
  assign \new_[38804]_  = A199 & A166;
  assign \new_[38805]_  = A167 & \new_[38804]_ ;
  assign \new_[38809]_  = A202 & A201;
  assign \new_[38810]_  = ~A200 & \new_[38809]_ ;
  assign \new_[38811]_  = \new_[38810]_  & \new_[38805]_ ;
  assign \new_[38815]_  = A298 & A269;
  assign \new_[38816]_  = ~A267 & \new_[38815]_ ;
  assign \new_[38819]_  = ~A300 & ~A299;
  assign \new_[38822]_  = ~A302 & ~A301;
  assign \new_[38823]_  = \new_[38822]_  & \new_[38819]_ ;
  assign \new_[38824]_  = \new_[38823]_  & \new_[38816]_ ;
  assign \new_[38828]_  = A199 & A166;
  assign \new_[38829]_  = A167 & \new_[38828]_ ;
  assign \new_[38833]_  = A202 & A201;
  assign \new_[38834]_  = ~A200 & \new_[38833]_ ;
  assign \new_[38835]_  = \new_[38834]_  & \new_[38829]_ ;
  assign \new_[38839]_  = ~A298 & A269;
  assign \new_[38840]_  = ~A267 & \new_[38839]_ ;
  assign \new_[38843]_  = ~A300 & A299;
  assign \new_[38846]_  = ~A302 & ~A301;
  assign \new_[38847]_  = \new_[38846]_  & \new_[38843]_ ;
  assign \new_[38848]_  = \new_[38847]_  & \new_[38840]_ ;
  assign \new_[38852]_  = A199 & A166;
  assign \new_[38853]_  = A167 & \new_[38852]_ ;
  assign \new_[38857]_  = A202 & A201;
  assign \new_[38858]_  = ~A200 & \new_[38857]_ ;
  assign \new_[38859]_  = \new_[38858]_  & \new_[38853]_ ;
  assign \new_[38863]_  = A298 & A266;
  assign \new_[38864]_  = A265 & \new_[38863]_ ;
  assign \new_[38867]_  = ~A300 & ~A299;
  assign \new_[38870]_  = ~A302 & ~A301;
  assign \new_[38871]_  = \new_[38870]_  & \new_[38867]_ ;
  assign \new_[38872]_  = \new_[38871]_  & \new_[38864]_ ;
  assign \new_[38876]_  = A199 & A166;
  assign \new_[38877]_  = A167 & \new_[38876]_ ;
  assign \new_[38881]_  = A202 & A201;
  assign \new_[38882]_  = ~A200 & \new_[38881]_ ;
  assign \new_[38883]_  = \new_[38882]_  & \new_[38877]_ ;
  assign \new_[38887]_  = ~A298 & A266;
  assign \new_[38888]_  = A265 & \new_[38887]_ ;
  assign \new_[38891]_  = ~A300 & A299;
  assign \new_[38894]_  = ~A302 & ~A301;
  assign \new_[38895]_  = \new_[38894]_  & \new_[38891]_ ;
  assign \new_[38896]_  = \new_[38895]_  & \new_[38888]_ ;
  assign \new_[38900]_  = A199 & A166;
  assign \new_[38901]_  = A167 & \new_[38900]_ ;
  assign \new_[38905]_  = A202 & A201;
  assign \new_[38906]_  = ~A200 & \new_[38905]_ ;
  assign \new_[38907]_  = \new_[38906]_  & \new_[38901]_ ;
  assign \new_[38911]_  = A298 & ~A266;
  assign \new_[38912]_  = ~A265 & \new_[38911]_ ;
  assign \new_[38915]_  = ~A300 & ~A299;
  assign \new_[38918]_  = ~A302 & ~A301;
  assign \new_[38919]_  = \new_[38918]_  & \new_[38915]_ ;
  assign \new_[38920]_  = \new_[38919]_  & \new_[38912]_ ;
  assign \new_[38924]_  = A199 & A166;
  assign \new_[38925]_  = A167 & \new_[38924]_ ;
  assign \new_[38929]_  = A202 & A201;
  assign \new_[38930]_  = ~A200 & \new_[38929]_ ;
  assign \new_[38931]_  = \new_[38930]_  & \new_[38925]_ ;
  assign \new_[38935]_  = ~A298 & ~A266;
  assign \new_[38936]_  = ~A265 & \new_[38935]_ ;
  assign \new_[38939]_  = ~A300 & A299;
  assign \new_[38942]_  = ~A302 & ~A301;
  assign \new_[38943]_  = \new_[38942]_  & \new_[38939]_ ;
  assign \new_[38944]_  = \new_[38943]_  & \new_[38936]_ ;
  assign \new_[38948]_  = A199 & A166;
  assign \new_[38949]_  = A167 & \new_[38948]_ ;
  assign \new_[38953]_  = A203 & A201;
  assign \new_[38954]_  = ~A200 & \new_[38953]_ ;
  assign \new_[38955]_  = \new_[38954]_  & \new_[38949]_ ;
  assign \new_[38959]_  = ~A269 & ~A268;
  assign \new_[38960]_  = A267 & \new_[38959]_ ;
  assign \new_[38963]_  = ~A299 & A298;
  assign \new_[38966]_  = A301 & A300;
  assign \new_[38967]_  = \new_[38966]_  & \new_[38963]_ ;
  assign \new_[38968]_  = \new_[38967]_  & \new_[38960]_ ;
  assign \new_[38972]_  = A199 & A166;
  assign \new_[38973]_  = A167 & \new_[38972]_ ;
  assign \new_[38977]_  = A203 & A201;
  assign \new_[38978]_  = ~A200 & \new_[38977]_ ;
  assign \new_[38979]_  = \new_[38978]_  & \new_[38973]_ ;
  assign \new_[38983]_  = ~A269 & ~A268;
  assign \new_[38984]_  = A267 & \new_[38983]_ ;
  assign \new_[38987]_  = ~A299 & A298;
  assign \new_[38990]_  = A302 & A300;
  assign \new_[38991]_  = \new_[38990]_  & \new_[38987]_ ;
  assign \new_[38992]_  = \new_[38991]_  & \new_[38984]_ ;
  assign \new_[38996]_  = A199 & A166;
  assign \new_[38997]_  = A167 & \new_[38996]_ ;
  assign \new_[39001]_  = A203 & A201;
  assign \new_[39002]_  = ~A200 & \new_[39001]_ ;
  assign \new_[39003]_  = \new_[39002]_  & \new_[38997]_ ;
  assign \new_[39007]_  = ~A269 & ~A268;
  assign \new_[39008]_  = A267 & \new_[39007]_ ;
  assign \new_[39011]_  = A299 & ~A298;
  assign \new_[39014]_  = A301 & A300;
  assign \new_[39015]_  = \new_[39014]_  & \new_[39011]_ ;
  assign \new_[39016]_  = \new_[39015]_  & \new_[39008]_ ;
  assign \new_[39020]_  = A199 & A166;
  assign \new_[39021]_  = A167 & \new_[39020]_ ;
  assign \new_[39025]_  = A203 & A201;
  assign \new_[39026]_  = ~A200 & \new_[39025]_ ;
  assign \new_[39027]_  = \new_[39026]_  & \new_[39021]_ ;
  assign \new_[39031]_  = ~A269 & ~A268;
  assign \new_[39032]_  = A267 & \new_[39031]_ ;
  assign \new_[39035]_  = A299 & ~A298;
  assign \new_[39038]_  = A302 & A300;
  assign \new_[39039]_  = \new_[39038]_  & \new_[39035]_ ;
  assign \new_[39040]_  = \new_[39039]_  & \new_[39032]_ ;
  assign \new_[39044]_  = A199 & A166;
  assign \new_[39045]_  = A167 & \new_[39044]_ ;
  assign \new_[39049]_  = A203 & A201;
  assign \new_[39050]_  = ~A200 & \new_[39049]_ ;
  assign \new_[39051]_  = \new_[39050]_  & \new_[39045]_ ;
  assign \new_[39055]_  = A298 & A268;
  assign \new_[39056]_  = ~A267 & \new_[39055]_ ;
  assign \new_[39059]_  = ~A300 & ~A299;
  assign \new_[39062]_  = ~A302 & ~A301;
  assign \new_[39063]_  = \new_[39062]_  & \new_[39059]_ ;
  assign \new_[39064]_  = \new_[39063]_  & \new_[39056]_ ;
  assign \new_[39068]_  = A199 & A166;
  assign \new_[39069]_  = A167 & \new_[39068]_ ;
  assign \new_[39073]_  = A203 & A201;
  assign \new_[39074]_  = ~A200 & \new_[39073]_ ;
  assign \new_[39075]_  = \new_[39074]_  & \new_[39069]_ ;
  assign \new_[39079]_  = ~A298 & A268;
  assign \new_[39080]_  = ~A267 & \new_[39079]_ ;
  assign \new_[39083]_  = ~A300 & A299;
  assign \new_[39086]_  = ~A302 & ~A301;
  assign \new_[39087]_  = \new_[39086]_  & \new_[39083]_ ;
  assign \new_[39088]_  = \new_[39087]_  & \new_[39080]_ ;
  assign \new_[39092]_  = A199 & A166;
  assign \new_[39093]_  = A167 & \new_[39092]_ ;
  assign \new_[39097]_  = A203 & A201;
  assign \new_[39098]_  = ~A200 & \new_[39097]_ ;
  assign \new_[39099]_  = \new_[39098]_  & \new_[39093]_ ;
  assign \new_[39103]_  = A298 & A269;
  assign \new_[39104]_  = ~A267 & \new_[39103]_ ;
  assign \new_[39107]_  = ~A300 & ~A299;
  assign \new_[39110]_  = ~A302 & ~A301;
  assign \new_[39111]_  = \new_[39110]_  & \new_[39107]_ ;
  assign \new_[39112]_  = \new_[39111]_  & \new_[39104]_ ;
  assign \new_[39116]_  = A199 & A166;
  assign \new_[39117]_  = A167 & \new_[39116]_ ;
  assign \new_[39121]_  = A203 & A201;
  assign \new_[39122]_  = ~A200 & \new_[39121]_ ;
  assign \new_[39123]_  = \new_[39122]_  & \new_[39117]_ ;
  assign \new_[39127]_  = ~A298 & A269;
  assign \new_[39128]_  = ~A267 & \new_[39127]_ ;
  assign \new_[39131]_  = ~A300 & A299;
  assign \new_[39134]_  = ~A302 & ~A301;
  assign \new_[39135]_  = \new_[39134]_  & \new_[39131]_ ;
  assign \new_[39136]_  = \new_[39135]_  & \new_[39128]_ ;
  assign \new_[39140]_  = A199 & A166;
  assign \new_[39141]_  = A167 & \new_[39140]_ ;
  assign \new_[39145]_  = A203 & A201;
  assign \new_[39146]_  = ~A200 & \new_[39145]_ ;
  assign \new_[39147]_  = \new_[39146]_  & \new_[39141]_ ;
  assign \new_[39151]_  = A298 & A266;
  assign \new_[39152]_  = A265 & \new_[39151]_ ;
  assign \new_[39155]_  = ~A300 & ~A299;
  assign \new_[39158]_  = ~A302 & ~A301;
  assign \new_[39159]_  = \new_[39158]_  & \new_[39155]_ ;
  assign \new_[39160]_  = \new_[39159]_  & \new_[39152]_ ;
  assign \new_[39164]_  = A199 & A166;
  assign \new_[39165]_  = A167 & \new_[39164]_ ;
  assign \new_[39169]_  = A203 & A201;
  assign \new_[39170]_  = ~A200 & \new_[39169]_ ;
  assign \new_[39171]_  = \new_[39170]_  & \new_[39165]_ ;
  assign \new_[39175]_  = ~A298 & A266;
  assign \new_[39176]_  = A265 & \new_[39175]_ ;
  assign \new_[39179]_  = ~A300 & A299;
  assign \new_[39182]_  = ~A302 & ~A301;
  assign \new_[39183]_  = \new_[39182]_  & \new_[39179]_ ;
  assign \new_[39184]_  = \new_[39183]_  & \new_[39176]_ ;
  assign \new_[39188]_  = A199 & A166;
  assign \new_[39189]_  = A167 & \new_[39188]_ ;
  assign \new_[39193]_  = A203 & A201;
  assign \new_[39194]_  = ~A200 & \new_[39193]_ ;
  assign \new_[39195]_  = \new_[39194]_  & \new_[39189]_ ;
  assign \new_[39199]_  = A298 & ~A266;
  assign \new_[39200]_  = ~A265 & \new_[39199]_ ;
  assign \new_[39203]_  = ~A300 & ~A299;
  assign \new_[39206]_  = ~A302 & ~A301;
  assign \new_[39207]_  = \new_[39206]_  & \new_[39203]_ ;
  assign \new_[39208]_  = \new_[39207]_  & \new_[39200]_ ;
  assign \new_[39212]_  = A199 & A166;
  assign \new_[39213]_  = A167 & \new_[39212]_ ;
  assign \new_[39217]_  = A203 & A201;
  assign \new_[39218]_  = ~A200 & \new_[39217]_ ;
  assign \new_[39219]_  = \new_[39218]_  & \new_[39213]_ ;
  assign \new_[39223]_  = ~A298 & ~A266;
  assign \new_[39224]_  = ~A265 & \new_[39223]_ ;
  assign \new_[39227]_  = ~A300 & A299;
  assign \new_[39230]_  = ~A302 & ~A301;
  assign \new_[39231]_  = \new_[39230]_  & \new_[39227]_ ;
  assign \new_[39232]_  = \new_[39231]_  & \new_[39224]_ ;
  assign \new_[39236]_  = A199 & A166;
  assign \new_[39237]_  = A167 & \new_[39236]_ ;
  assign \new_[39241]_  = ~A202 & ~A201;
  assign \new_[39242]_  = ~A200 & \new_[39241]_ ;
  assign \new_[39243]_  = \new_[39242]_  & \new_[39237]_ ;
  assign \new_[39247]_  = A268 & ~A267;
  assign \new_[39248]_  = ~A203 & \new_[39247]_ ;
  assign \new_[39251]_  = ~A299 & A298;
  assign \new_[39254]_  = A301 & A300;
  assign \new_[39255]_  = \new_[39254]_  & \new_[39251]_ ;
  assign \new_[39256]_  = \new_[39255]_  & \new_[39248]_ ;
  assign \new_[39260]_  = A199 & A166;
  assign \new_[39261]_  = A167 & \new_[39260]_ ;
  assign \new_[39265]_  = ~A202 & ~A201;
  assign \new_[39266]_  = ~A200 & \new_[39265]_ ;
  assign \new_[39267]_  = \new_[39266]_  & \new_[39261]_ ;
  assign \new_[39271]_  = A268 & ~A267;
  assign \new_[39272]_  = ~A203 & \new_[39271]_ ;
  assign \new_[39275]_  = ~A299 & A298;
  assign \new_[39278]_  = A302 & A300;
  assign \new_[39279]_  = \new_[39278]_  & \new_[39275]_ ;
  assign \new_[39280]_  = \new_[39279]_  & \new_[39272]_ ;
  assign \new_[39284]_  = A199 & A166;
  assign \new_[39285]_  = A167 & \new_[39284]_ ;
  assign \new_[39289]_  = ~A202 & ~A201;
  assign \new_[39290]_  = ~A200 & \new_[39289]_ ;
  assign \new_[39291]_  = \new_[39290]_  & \new_[39285]_ ;
  assign \new_[39295]_  = A268 & ~A267;
  assign \new_[39296]_  = ~A203 & \new_[39295]_ ;
  assign \new_[39299]_  = A299 & ~A298;
  assign \new_[39302]_  = A301 & A300;
  assign \new_[39303]_  = \new_[39302]_  & \new_[39299]_ ;
  assign \new_[39304]_  = \new_[39303]_  & \new_[39296]_ ;
  assign \new_[39308]_  = A199 & A166;
  assign \new_[39309]_  = A167 & \new_[39308]_ ;
  assign \new_[39313]_  = ~A202 & ~A201;
  assign \new_[39314]_  = ~A200 & \new_[39313]_ ;
  assign \new_[39315]_  = \new_[39314]_  & \new_[39309]_ ;
  assign \new_[39319]_  = A268 & ~A267;
  assign \new_[39320]_  = ~A203 & \new_[39319]_ ;
  assign \new_[39323]_  = A299 & ~A298;
  assign \new_[39326]_  = A302 & A300;
  assign \new_[39327]_  = \new_[39326]_  & \new_[39323]_ ;
  assign \new_[39328]_  = \new_[39327]_  & \new_[39320]_ ;
  assign \new_[39332]_  = A199 & A166;
  assign \new_[39333]_  = A167 & \new_[39332]_ ;
  assign \new_[39337]_  = ~A202 & ~A201;
  assign \new_[39338]_  = ~A200 & \new_[39337]_ ;
  assign \new_[39339]_  = \new_[39338]_  & \new_[39333]_ ;
  assign \new_[39343]_  = A269 & ~A267;
  assign \new_[39344]_  = ~A203 & \new_[39343]_ ;
  assign \new_[39347]_  = ~A299 & A298;
  assign \new_[39350]_  = A301 & A300;
  assign \new_[39351]_  = \new_[39350]_  & \new_[39347]_ ;
  assign \new_[39352]_  = \new_[39351]_  & \new_[39344]_ ;
  assign \new_[39356]_  = A199 & A166;
  assign \new_[39357]_  = A167 & \new_[39356]_ ;
  assign \new_[39361]_  = ~A202 & ~A201;
  assign \new_[39362]_  = ~A200 & \new_[39361]_ ;
  assign \new_[39363]_  = \new_[39362]_  & \new_[39357]_ ;
  assign \new_[39367]_  = A269 & ~A267;
  assign \new_[39368]_  = ~A203 & \new_[39367]_ ;
  assign \new_[39371]_  = ~A299 & A298;
  assign \new_[39374]_  = A302 & A300;
  assign \new_[39375]_  = \new_[39374]_  & \new_[39371]_ ;
  assign \new_[39376]_  = \new_[39375]_  & \new_[39368]_ ;
  assign \new_[39380]_  = A199 & A166;
  assign \new_[39381]_  = A167 & \new_[39380]_ ;
  assign \new_[39385]_  = ~A202 & ~A201;
  assign \new_[39386]_  = ~A200 & \new_[39385]_ ;
  assign \new_[39387]_  = \new_[39386]_  & \new_[39381]_ ;
  assign \new_[39391]_  = A269 & ~A267;
  assign \new_[39392]_  = ~A203 & \new_[39391]_ ;
  assign \new_[39395]_  = A299 & ~A298;
  assign \new_[39398]_  = A301 & A300;
  assign \new_[39399]_  = \new_[39398]_  & \new_[39395]_ ;
  assign \new_[39400]_  = \new_[39399]_  & \new_[39392]_ ;
  assign \new_[39404]_  = A199 & A166;
  assign \new_[39405]_  = A167 & \new_[39404]_ ;
  assign \new_[39409]_  = ~A202 & ~A201;
  assign \new_[39410]_  = ~A200 & \new_[39409]_ ;
  assign \new_[39411]_  = \new_[39410]_  & \new_[39405]_ ;
  assign \new_[39415]_  = A269 & ~A267;
  assign \new_[39416]_  = ~A203 & \new_[39415]_ ;
  assign \new_[39419]_  = A299 & ~A298;
  assign \new_[39422]_  = A302 & A300;
  assign \new_[39423]_  = \new_[39422]_  & \new_[39419]_ ;
  assign \new_[39424]_  = \new_[39423]_  & \new_[39416]_ ;
  assign \new_[39428]_  = A199 & A166;
  assign \new_[39429]_  = A167 & \new_[39428]_ ;
  assign \new_[39433]_  = ~A202 & ~A201;
  assign \new_[39434]_  = ~A200 & \new_[39433]_ ;
  assign \new_[39435]_  = \new_[39434]_  & \new_[39429]_ ;
  assign \new_[39439]_  = A266 & A265;
  assign \new_[39440]_  = ~A203 & \new_[39439]_ ;
  assign \new_[39443]_  = ~A299 & A298;
  assign \new_[39446]_  = A301 & A300;
  assign \new_[39447]_  = \new_[39446]_  & \new_[39443]_ ;
  assign \new_[39448]_  = \new_[39447]_  & \new_[39440]_ ;
  assign \new_[39452]_  = A199 & A166;
  assign \new_[39453]_  = A167 & \new_[39452]_ ;
  assign \new_[39457]_  = ~A202 & ~A201;
  assign \new_[39458]_  = ~A200 & \new_[39457]_ ;
  assign \new_[39459]_  = \new_[39458]_  & \new_[39453]_ ;
  assign \new_[39463]_  = A266 & A265;
  assign \new_[39464]_  = ~A203 & \new_[39463]_ ;
  assign \new_[39467]_  = ~A299 & A298;
  assign \new_[39470]_  = A302 & A300;
  assign \new_[39471]_  = \new_[39470]_  & \new_[39467]_ ;
  assign \new_[39472]_  = \new_[39471]_  & \new_[39464]_ ;
  assign \new_[39476]_  = A199 & A166;
  assign \new_[39477]_  = A167 & \new_[39476]_ ;
  assign \new_[39481]_  = ~A202 & ~A201;
  assign \new_[39482]_  = ~A200 & \new_[39481]_ ;
  assign \new_[39483]_  = \new_[39482]_  & \new_[39477]_ ;
  assign \new_[39487]_  = A266 & A265;
  assign \new_[39488]_  = ~A203 & \new_[39487]_ ;
  assign \new_[39491]_  = A299 & ~A298;
  assign \new_[39494]_  = A301 & A300;
  assign \new_[39495]_  = \new_[39494]_  & \new_[39491]_ ;
  assign \new_[39496]_  = \new_[39495]_  & \new_[39488]_ ;
  assign \new_[39500]_  = A199 & A166;
  assign \new_[39501]_  = A167 & \new_[39500]_ ;
  assign \new_[39505]_  = ~A202 & ~A201;
  assign \new_[39506]_  = ~A200 & \new_[39505]_ ;
  assign \new_[39507]_  = \new_[39506]_  & \new_[39501]_ ;
  assign \new_[39511]_  = A266 & A265;
  assign \new_[39512]_  = ~A203 & \new_[39511]_ ;
  assign \new_[39515]_  = A299 & ~A298;
  assign \new_[39518]_  = A302 & A300;
  assign \new_[39519]_  = \new_[39518]_  & \new_[39515]_ ;
  assign \new_[39520]_  = \new_[39519]_  & \new_[39512]_ ;
  assign \new_[39524]_  = A199 & A166;
  assign \new_[39525]_  = A167 & \new_[39524]_ ;
  assign \new_[39529]_  = ~A202 & ~A201;
  assign \new_[39530]_  = ~A200 & \new_[39529]_ ;
  assign \new_[39531]_  = \new_[39530]_  & \new_[39525]_ ;
  assign \new_[39535]_  = ~A266 & ~A265;
  assign \new_[39536]_  = ~A203 & \new_[39535]_ ;
  assign \new_[39539]_  = ~A299 & A298;
  assign \new_[39542]_  = A301 & A300;
  assign \new_[39543]_  = \new_[39542]_  & \new_[39539]_ ;
  assign \new_[39544]_  = \new_[39543]_  & \new_[39536]_ ;
  assign \new_[39548]_  = A199 & A166;
  assign \new_[39549]_  = A167 & \new_[39548]_ ;
  assign \new_[39553]_  = ~A202 & ~A201;
  assign \new_[39554]_  = ~A200 & \new_[39553]_ ;
  assign \new_[39555]_  = \new_[39554]_  & \new_[39549]_ ;
  assign \new_[39559]_  = ~A266 & ~A265;
  assign \new_[39560]_  = ~A203 & \new_[39559]_ ;
  assign \new_[39563]_  = ~A299 & A298;
  assign \new_[39566]_  = A302 & A300;
  assign \new_[39567]_  = \new_[39566]_  & \new_[39563]_ ;
  assign \new_[39568]_  = \new_[39567]_  & \new_[39560]_ ;
  assign \new_[39572]_  = A199 & A166;
  assign \new_[39573]_  = A167 & \new_[39572]_ ;
  assign \new_[39577]_  = ~A202 & ~A201;
  assign \new_[39578]_  = ~A200 & \new_[39577]_ ;
  assign \new_[39579]_  = \new_[39578]_  & \new_[39573]_ ;
  assign \new_[39583]_  = ~A266 & ~A265;
  assign \new_[39584]_  = ~A203 & \new_[39583]_ ;
  assign \new_[39587]_  = A299 & ~A298;
  assign \new_[39590]_  = A301 & A300;
  assign \new_[39591]_  = \new_[39590]_  & \new_[39587]_ ;
  assign \new_[39592]_  = \new_[39591]_  & \new_[39584]_ ;
  assign \new_[39596]_  = A199 & A166;
  assign \new_[39597]_  = A167 & \new_[39596]_ ;
  assign \new_[39601]_  = ~A202 & ~A201;
  assign \new_[39602]_  = ~A200 & \new_[39601]_ ;
  assign \new_[39603]_  = \new_[39602]_  & \new_[39597]_ ;
  assign \new_[39607]_  = ~A266 & ~A265;
  assign \new_[39608]_  = ~A203 & \new_[39607]_ ;
  assign \new_[39611]_  = A299 & ~A298;
  assign \new_[39614]_  = A302 & A300;
  assign \new_[39615]_  = \new_[39614]_  & \new_[39611]_ ;
  assign \new_[39616]_  = \new_[39615]_  & \new_[39608]_ ;
  assign \new_[39620]_  = A201 & ~A166;
  assign \new_[39621]_  = ~A167 & \new_[39620]_ ;
  assign \new_[39625]_  = ~A265 & ~A203;
  assign \new_[39626]_  = ~A202 & \new_[39625]_ ;
  assign \new_[39627]_  = \new_[39626]_  & \new_[39621]_ ;
  assign \new_[39631]_  = ~A268 & ~A267;
  assign \new_[39632]_  = A266 & \new_[39631]_ ;
  assign \new_[39635]_  = A300 & ~A269;
  assign \new_[39638]_  = ~A302 & ~A301;
  assign \new_[39639]_  = \new_[39638]_  & \new_[39635]_ ;
  assign \new_[39640]_  = \new_[39639]_  & \new_[39632]_ ;
  assign \new_[39644]_  = A201 & ~A166;
  assign \new_[39645]_  = ~A167 & \new_[39644]_ ;
  assign \new_[39649]_  = A265 & ~A203;
  assign \new_[39650]_  = ~A202 & \new_[39649]_ ;
  assign \new_[39651]_  = \new_[39650]_  & \new_[39645]_ ;
  assign \new_[39655]_  = ~A268 & ~A267;
  assign \new_[39656]_  = ~A266 & \new_[39655]_ ;
  assign \new_[39659]_  = A300 & ~A269;
  assign \new_[39662]_  = ~A302 & ~A301;
  assign \new_[39663]_  = \new_[39662]_  & \new_[39659]_ ;
  assign \new_[39664]_  = \new_[39663]_  & \new_[39656]_ ;
  assign \new_[39668]_  = ~A199 & ~A166;
  assign \new_[39669]_  = ~A167 & \new_[39668]_ ;
  assign \new_[39673]_  = A202 & A201;
  assign \new_[39674]_  = A200 & \new_[39673]_ ;
  assign \new_[39675]_  = \new_[39674]_  & \new_[39669]_ ;
  assign \new_[39679]_  = ~A269 & ~A268;
  assign \new_[39680]_  = A267 & \new_[39679]_ ;
  assign \new_[39683]_  = ~A299 & A298;
  assign \new_[39686]_  = A301 & A300;
  assign \new_[39687]_  = \new_[39686]_  & \new_[39683]_ ;
  assign \new_[39688]_  = \new_[39687]_  & \new_[39680]_ ;
  assign \new_[39692]_  = ~A199 & ~A166;
  assign \new_[39693]_  = ~A167 & \new_[39692]_ ;
  assign \new_[39697]_  = A202 & A201;
  assign \new_[39698]_  = A200 & \new_[39697]_ ;
  assign \new_[39699]_  = \new_[39698]_  & \new_[39693]_ ;
  assign \new_[39703]_  = ~A269 & ~A268;
  assign \new_[39704]_  = A267 & \new_[39703]_ ;
  assign \new_[39707]_  = ~A299 & A298;
  assign \new_[39710]_  = A302 & A300;
  assign \new_[39711]_  = \new_[39710]_  & \new_[39707]_ ;
  assign \new_[39712]_  = \new_[39711]_  & \new_[39704]_ ;
  assign \new_[39716]_  = ~A199 & ~A166;
  assign \new_[39717]_  = ~A167 & \new_[39716]_ ;
  assign \new_[39721]_  = A202 & A201;
  assign \new_[39722]_  = A200 & \new_[39721]_ ;
  assign \new_[39723]_  = \new_[39722]_  & \new_[39717]_ ;
  assign \new_[39727]_  = ~A269 & ~A268;
  assign \new_[39728]_  = A267 & \new_[39727]_ ;
  assign \new_[39731]_  = A299 & ~A298;
  assign \new_[39734]_  = A301 & A300;
  assign \new_[39735]_  = \new_[39734]_  & \new_[39731]_ ;
  assign \new_[39736]_  = \new_[39735]_  & \new_[39728]_ ;
  assign \new_[39740]_  = ~A199 & ~A166;
  assign \new_[39741]_  = ~A167 & \new_[39740]_ ;
  assign \new_[39745]_  = A202 & A201;
  assign \new_[39746]_  = A200 & \new_[39745]_ ;
  assign \new_[39747]_  = \new_[39746]_  & \new_[39741]_ ;
  assign \new_[39751]_  = ~A269 & ~A268;
  assign \new_[39752]_  = A267 & \new_[39751]_ ;
  assign \new_[39755]_  = A299 & ~A298;
  assign \new_[39758]_  = A302 & A300;
  assign \new_[39759]_  = \new_[39758]_  & \new_[39755]_ ;
  assign \new_[39760]_  = \new_[39759]_  & \new_[39752]_ ;
  assign \new_[39764]_  = ~A199 & ~A166;
  assign \new_[39765]_  = ~A167 & \new_[39764]_ ;
  assign \new_[39769]_  = A202 & A201;
  assign \new_[39770]_  = A200 & \new_[39769]_ ;
  assign \new_[39771]_  = \new_[39770]_  & \new_[39765]_ ;
  assign \new_[39775]_  = A298 & A268;
  assign \new_[39776]_  = ~A267 & \new_[39775]_ ;
  assign \new_[39779]_  = ~A300 & ~A299;
  assign \new_[39782]_  = ~A302 & ~A301;
  assign \new_[39783]_  = \new_[39782]_  & \new_[39779]_ ;
  assign \new_[39784]_  = \new_[39783]_  & \new_[39776]_ ;
  assign \new_[39788]_  = ~A199 & ~A166;
  assign \new_[39789]_  = ~A167 & \new_[39788]_ ;
  assign \new_[39793]_  = A202 & A201;
  assign \new_[39794]_  = A200 & \new_[39793]_ ;
  assign \new_[39795]_  = \new_[39794]_  & \new_[39789]_ ;
  assign \new_[39799]_  = ~A298 & A268;
  assign \new_[39800]_  = ~A267 & \new_[39799]_ ;
  assign \new_[39803]_  = ~A300 & A299;
  assign \new_[39806]_  = ~A302 & ~A301;
  assign \new_[39807]_  = \new_[39806]_  & \new_[39803]_ ;
  assign \new_[39808]_  = \new_[39807]_  & \new_[39800]_ ;
  assign \new_[39812]_  = ~A199 & ~A166;
  assign \new_[39813]_  = ~A167 & \new_[39812]_ ;
  assign \new_[39817]_  = A202 & A201;
  assign \new_[39818]_  = A200 & \new_[39817]_ ;
  assign \new_[39819]_  = \new_[39818]_  & \new_[39813]_ ;
  assign \new_[39823]_  = A298 & A269;
  assign \new_[39824]_  = ~A267 & \new_[39823]_ ;
  assign \new_[39827]_  = ~A300 & ~A299;
  assign \new_[39830]_  = ~A302 & ~A301;
  assign \new_[39831]_  = \new_[39830]_  & \new_[39827]_ ;
  assign \new_[39832]_  = \new_[39831]_  & \new_[39824]_ ;
  assign \new_[39836]_  = ~A199 & ~A166;
  assign \new_[39837]_  = ~A167 & \new_[39836]_ ;
  assign \new_[39841]_  = A202 & A201;
  assign \new_[39842]_  = A200 & \new_[39841]_ ;
  assign \new_[39843]_  = \new_[39842]_  & \new_[39837]_ ;
  assign \new_[39847]_  = ~A298 & A269;
  assign \new_[39848]_  = ~A267 & \new_[39847]_ ;
  assign \new_[39851]_  = ~A300 & A299;
  assign \new_[39854]_  = ~A302 & ~A301;
  assign \new_[39855]_  = \new_[39854]_  & \new_[39851]_ ;
  assign \new_[39856]_  = \new_[39855]_  & \new_[39848]_ ;
  assign \new_[39860]_  = ~A199 & ~A166;
  assign \new_[39861]_  = ~A167 & \new_[39860]_ ;
  assign \new_[39865]_  = A202 & A201;
  assign \new_[39866]_  = A200 & \new_[39865]_ ;
  assign \new_[39867]_  = \new_[39866]_  & \new_[39861]_ ;
  assign \new_[39871]_  = A298 & A266;
  assign \new_[39872]_  = A265 & \new_[39871]_ ;
  assign \new_[39875]_  = ~A300 & ~A299;
  assign \new_[39878]_  = ~A302 & ~A301;
  assign \new_[39879]_  = \new_[39878]_  & \new_[39875]_ ;
  assign \new_[39880]_  = \new_[39879]_  & \new_[39872]_ ;
  assign \new_[39884]_  = ~A199 & ~A166;
  assign \new_[39885]_  = ~A167 & \new_[39884]_ ;
  assign \new_[39889]_  = A202 & A201;
  assign \new_[39890]_  = A200 & \new_[39889]_ ;
  assign \new_[39891]_  = \new_[39890]_  & \new_[39885]_ ;
  assign \new_[39895]_  = ~A298 & A266;
  assign \new_[39896]_  = A265 & \new_[39895]_ ;
  assign \new_[39899]_  = ~A300 & A299;
  assign \new_[39902]_  = ~A302 & ~A301;
  assign \new_[39903]_  = \new_[39902]_  & \new_[39899]_ ;
  assign \new_[39904]_  = \new_[39903]_  & \new_[39896]_ ;
  assign \new_[39908]_  = ~A199 & ~A166;
  assign \new_[39909]_  = ~A167 & \new_[39908]_ ;
  assign \new_[39913]_  = A202 & A201;
  assign \new_[39914]_  = A200 & \new_[39913]_ ;
  assign \new_[39915]_  = \new_[39914]_  & \new_[39909]_ ;
  assign \new_[39919]_  = A298 & ~A266;
  assign \new_[39920]_  = ~A265 & \new_[39919]_ ;
  assign \new_[39923]_  = ~A300 & ~A299;
  assign \new_[39926]_  = ~A302 & ~A301;
  assign \new_[39927]_  = \new_[39926]_  & \new_[39923]_ ;
  assign \new_[39928]_  = \new_[39927]_  & \new_[39920]_ ;
  assign \new_[39932]_  = ~A199 & ~A166;
  assign \new_[39933]_  = ~A167 & \new_[39932]_ ;
  assign \new_[39937]_  = A202 & A201;
  assign \new_[39938]_  = A200 & \new_[39937]_ ;
  assign \new_[39939]_  = \new_[39938]_  & \new_[39933]_ ;
  assign \new_[39943]_  = ~A298 & ~A266;
  assign \new_[39944]_  = ~A265 & \new_[39943]_ ;
  assign \new_[39947]_  = ~A300 & A299;
  assign \new_[39950]_  = ~A302 & ~A301;
  assign \new_[39951]_  = \new_[39950]_  & \new_[39947]_ ;
  assign \new_[39952]_  = \new_[39951]_  & \new_[39944]_ ;
  assign \new_[39956]_  = ~A199 & ~A166;
  assign \new_[39957]_  = ~A167 & \new_[39956]_ ;
  assign \new_[39961]_  = A203 & A201;
  assign \new_[39962]_  = A200 & \new_[39961]_ ;
  assign \new_[39963]_  = \new_[39962]_  & \new_[39957]_ ;
  assign \new_[39967]_  = ~A269 & ~A268;
  assign \new_[39968]_  = A267 & \new_[39967]_ ;
  assign \new_[39971]_  = ~A299 & A298;
  assign \new_[39974]_  = A301 & A300;
  assign \new_[39975]_  = \new_[39974]_  & \new_[39971]_ ;
  assign \new_[39976]_  = \new_[39975]_  & \new_[39968]_ ;
  assign \new_[39980]_  = ~A199 & ~A166;
  assign \new_[39981]_  = ~A167 & \new_[39980]_ ;
  assign \new_[39985]_  = A203 & A201;
  assign \new_[39986]_  = A200 & \new_[39985]_ ;
  assign \new_[39987]_  = \new_[39986]_  & \new_[39981]_ ;
  assign \new_[39991]_  = ~A269 & ~A268;
  assign \new_[39992]_  = A267 & \new_[39991]_ ;
  assign \new_[39995]_  = ~A299 & A298;
  assign \new_[39998]_  = A302 & A300;
  assign \new_[39999]_  = \new_[39998]_  & \new_[39995]_ ;
  assign \new_[40000]_  = \new_[39999]_  & \new_[39992]_ ;
  assign \new_[40004]_  = ~A199 & ~A166;
  assign \new_[40005]_  = ~A167 & \new_[40004]_ ;
  assign \new_[40009]_  = A203 & A201;
  assign \new_[40010]_  = A200 & \new_[40009]_ ;
  assign \new_[40011]_  = \new_[40010]_  & \new_[40005]_ ;
  assign \new_[40015]_  = ~A269 & ~A268;
  assign \new_[40016]_  = A267 & \new_[40015]_ ;
  assign \new_[40019]_  = A299 & ~A298;
  assign \new_[40022]_  = A301 & A300;
  assign \new_[40023]_  = \new_[40022]_  & \new_[40019]_ ;
  assign \new_[40024]_  = \new_[40023]_  & \new_[40016]_ ;
  assign \new_[40028]_  = ~A199 & ~A166;
  assign \new_[40029]_  = ~A167 & \new_[40028]_ ;
  assign \new_[40033]_  = A203 & A201;
  assign \new_[40034]_  = A200 & \new_[40033]_ ;
  assign \new_[40035]_  = \new_[40034]_  & \new_[40029]_ ;
  assign \new_[40039]_  = ~A269 & ~A268;
  assign \new_[40040]_  = A267 & \new_[40039]_ ;
  assign \new_[40043]_  = A299 & ~A298;
  assign \new_[40046]_  = A302 & A300;
  assign \new_[40047]_  = \new_[40046]_  & \new_[40043]_ ;
  assign \new_[40048]_  = \new_[40047]_  & \new_[40040]_ ;
  assign \new_[40052]_  = ~A199 & ~A166;
  assign \new_[40053]_  = ~A167 & \new_[40052]_ ;
  assign \new_[40057]_  = A203 & A201;
  assign \new_[40058]_  = A200 & \new_[40057]_ ;
  assign \new_[40059]_  = \new_[40058]_  & \new_[40053]_ ;
  assign \new_[40063]_  = A298 & A268;
  assign \new_[40064]_  = ~A267 & \new_[40063]_ ;
  assign \new_[40067]_  = ~A300 & ~A299;
  assign \new_[40070]_  = ~A302 & ~A301;
  assign \new_[40071]_  = \new_[40070]_  & \new_[40067]_ ;
  assign \new_[40072]_  = \new_[40071]_  & \new_[40064]_ ;
  assign \new_[40076]_  = ~A199 & ~A166;
  assign \new_[40077]_  = ~A167 & \new_[40076]_ ;
  assign \new_[40081]_  = A203 & A201;
  assign \new_[40082]_  = A200 & \new_[40081]_ ;
  assign \new_[40083]_  = \new_[40082]_  & \new_[40077]_ ;
  assign \new_[40087]_  = ~A298 & A268;
  assign \new_[40088]_  = ~A267 & \new_[40087]_ ;
  assign \new_[40091]_  = ~A300 & A299;
  assign \new_[40094]_  = ~A302 & ~A301;
  assign \new_[40095]_  = \new_[40094]_  & \new_[40091]_ ;
  assign \new_[40096]_  = \new_[40095]_  & \new_[40088]_ ;
  assign \new_[40100]_  = ~A199 & ~A166;
  assign \new_[40101]_  = ~A167 & \new_[40100]_ ;
  assign \new_[40105]_  = A203 & A201;
  assign \new_[40106]_  = A200 & \new_[40105]_ ;
  assign \new_[40107]_  = \new_[40106]_  & \new_[40101]_ ;
  assign \new_[40111]_  = A298 & A269;
  assign \new_[40112]_  = ~A267 & \new_[40111]_ ;
  assign \new_[40115]_  = ~A300 & ~A299;
  assign \new_[40118]_  = ~A302 & ~A301;
  assign \new_[40119]_  = \new_[40118]_  & \new_[40115]_ ;
  assign \new_[40120]_  = \new_[40119]_  & \new_[40112]_ ;
  assign \new_[40124]_  = ~A199 & ~A166;
  assign \new_[40125]_  = ~A167 & \new_[40124]_ ;
  assign \new_[40129]_  = A203 & A201;
  assign \new_[40130]_  = A200 & \new_[40129]_ ;
  assign \new_[40131]_  = \new_[40130]_  & \new_[40125]_ ;
  assign \new_[40135]_  = ~A298 & A269;
  assign \new_[40136]_  = ~A267 & \new_[40135]_ ;
  assign \new_[40139]_  = ~A300 & A299;
  assign \new_[40142]_  = ~A302 & ~A301;
  assign \new_[40143]_  = \new_[40142]_  & \new_[40139]_ ;
  assign \new_[40144]_  = \new_[40143]_  & \new_[40136]_ ;
  assign \new_[40148]_  = ~A199 & ~A166;
  assign \new_[40149]_  = ~A167 & \new_[40148]_ ;
  assign \new_[40153]_  = A203 & A201;
  assign \new_[40154]_  = A200 & \new_[40153]_ ;
  assign \new_[40155]_  = \new_[40154]_  & \new_[40149]_ ;
  assign \new_[40159]_  = A298 & A266;
  assign \new_[40160]_  = A265 & \new_[40159]_ ;
  assign \new_[40163]_  = ~A300 & ~A299;
  assign \new_[40166]_  = ~A302 & ~A301;
  assign \new_[40167]_  = \new_[40166]_  & \new_[40163]_ ;
  assign \new_[40168]_  = \new_[40167]_  & \new_[40160]_ ;
  assign \new_[40172]_  = ~A199 & ~A166;
  assign \new_[40173]_  = ~A167 & \new_[40172]_ ;
  assign \new_[40177]_  = A203 & A201;
  assign \new_[40178]_  = A200 & \new_[40177]_ ;
  assign \new_[40179]_  = \new_[40178]_  & \new_[40173]_ ;
  assign \new_[40183]_  = ~A298 & A266;
  assign \new_[40184]_  = A265 & \new_[40183]_ ;
  assign \new_[40187]_  = ~A300 & A299;
  assign \new_[40190]_  = ~A302 & ~A301;
  assign \new_[40191]_  = \new_[40190]_  & \new_[40187]_ ;
  assign \new_[40192]_  = \new_[40191]_  & \new_[40184]_ ;
  assign \new_[40196]_  = ~A199 & ~A166;
  assign \new_[40197]_  = ~A167 & \new_[40196]_ ;
  assign \new_[40201]_  = A203 & A201;
  assign \new_[40202]_  = A200 & \new_[40201]_ ;
  assign \new_[40203]_  = \new_[40202]_  & \new_[40197]_ ;
  assign \new_[40207]_  = A298 & ~A266;
  assign \new_[40208]_  = ~A265 & \new_[40207]_ ;
  assign \new_[40211]_  = ~A300 & ~A299;
  assign \new_[40214]_  = ~A302 & ~A301;
  assign \new_[40215]_  = \new_[40214]_  & \new_[40211]_ ;
  assign \new_[40216]_  = \new_[40215]_  & \new_[40208]_ ;
  assign \new_[40220]_  = ~A199 & ~A166;
  assign \new_[40221]_  = ~A167 & \new_[40220]_ ;
  assign \new_[40225]_  = A203 & A201;
  assign \new_[40226]_  = A200 & \new_[40225]_ ;
  assign \new_[40227]_  = \new_[40226]_  & \new_[40221]_ ;
  assign \new_[40231]_  = ~A298 & ~A266;
  assign \new_[40232]_  = ~A265 & \new_[40231]_ ;
  assign \new_[40235]_  = ~A300 & A299;
  assign \new_[40238]_  = ~A302 & ~A301;
  assign \new_[40239]_  = \new_[40238]_  & \new_[40235]_ ;
  assign \new_[40240]_  = \new_[40239]_  & \new_[40232]_ ;
  assign \new_[40244]_  = ~A199 & ~A166;
  assign \new_[40245]_  = ~A167 & \new_[40244]_ ;
  assign \new_[40249]_  = ~A202 & ~A201;
  assign \new_[40250]_  = A200 & \new_[40249]_ ;
  assign \new_[40251]_  = \new_[40250]_  & \new_[40245]_ ;
  assign \new_[40255]_  = A268 & ~A267;
  assign \new_[40256]_  = ~A203 & \new_[40255]_ ;
  assign \new_[40259]_  = ~A299 & A298;
  assign \new_[40262]_  = A301 & A300;
  assign \new_[40263]_  = \new_[40262]_  & \new_[40259]_ ;
  assign \new_[40264]_  = \new_[40263]_  & \new_[40256]_ ;
  assign \new_[40268]_  = ~A199 & ~A166;
  assign \new_[40269]_  = ~A167 & \new_[40268]_ ;
  assign \new_[40273]_  = ~A202 & ~A201;
  assign \new_[40274]_  = A200 & \new_[40273]_ ;
  assign \new_[40275]_  = \new_[40274]_  & \new_[40269]_ ;
  assign \new_[40279]_  = A268 & ~A267;
  assign \new_[40280]_  = ~A203 & \new_[40279]_ ;
  assign \new_[40283]_  = ~A299 & A298;
  assign \new_[40286]_  = A302 & A300;
  assign \new_[40287]_  = \new_[40286]_  & \new_[40283]_ ;
  assign \new_[40288]_  = \new_[40287]_  & \new_[40280]_ ;
  assign \new_[40292]_  = ~A199 & ~A166;
  assign \new_[40293]_  = ~A167 & \new_[40292]_ ;
  assign \new_[40297]_  = ~A202 & ~A201;
  assign \new_[40298]_  = A200 & \new_[40297]_ ;
  assign \new_[40299]_  = \new_[40298]_  & \new_[40293]_ ;
  assign \new_[40303]_  = A268 & ~A267;
  assign \new_[40304]_  = ~A203 & \new_[40303]_ ;
  assign \new_[40307]_  = A299 & ~A298;
  assign \new_[40310]_  = A301 & A300;
  assign \new_[40311]_  = \new_[40310]_  & \new_[40307]_ ;
  assign \new_[40312]_  = \new_[40311]_  & \new_[40304]_ ;
  assign \new_[40316]_  = ~A199 & ~A166;
  assign \new_[40317]_  = ~A167 & \new_[40316]_ ;
  assign \new_[40321]_  = ~A202 & ~A201;
  assign \new_[40322]_  = A200 & \new_[40321]_ ;
  assign \new_[40323]_  = \new_[40322]_  & \new_[40317]_ ;
  assign \new_[40327]_  = A268 & ~A267;
  assign \new_[40328]_  = ~A203 & \new_[40327]_ ;
  assign \new_[40331]_  = A299 & ~A298;
  assign \new_[40334]_  = A302 & A300;
  assign \new_[40335]_  = \new_[40334]_  & \new_[40331]_ ;
  assign \new_[40336]_  = \new_[40335]_  & \new_[40328]_ ;
  assign \new_[40340]_  = ~A199 & ~A166;
  assign \new_[40341]_  = ~A167 & \new_[40340]_ ;
  assign \new_[40345]_  = ~A202 & ~A201;
  assign \new_[40346]_  = A200 & \new_[40345]_ ;
  assign \new_[40347]_  = \new_[40346]_  & \new_[40341]_ ;
  assign \new_[40351]_  = A269 & ~A267;
  assign \new_[40352]_  = ~A203 & \new_[40351]_ ;
  assign \new_[40355]_  = ~A299 & A298;
  assign \new_[40358]_  = A301 & A300;
  assign \new_[40359]_  = \new_[40358]_  & \new_[40355]_ ;
  assign \new_[40360]_  = \new_[40359]_  & \new_[40352]_ ;
  assign \new_[40364]_  = ~A199 & ~A166;
  assign \new_[40365]_  = ~A167 & \new_[40364]_ ;
  assign \new_[40369]_  = ~A202 & ~A201;
  assign \new_[40370]_  = A200 & \new_[40369]_ ;
  assign \new_[40371]_  = \new_[40370]_  & \new_[40365]_ ;
  assign \new_[40375]_  = A269 & ~A267;
  assign \new_[40376]_  = ~A203 & \new_[40375]_ ;
  assign \new_[40379]_  = ~A299 & A298;
  assign \new_[40382]_  = A302 & A300;
  assign \new_[40383]_  = \new_[40382]_  & \new_[40379]_ ;
  assign \new_[40384]_  = \new_[40383]_  & \new_[40376]_ ;
  assign \new_[40388]_  = ~A199 & ~A166;
  assign \new_[40389]_  = ~A167 & \new_[40388]_ ;
  assign \new_[40393]_  = ~A202 & ~A201;
  assign \new_[40394]_  = A200 & \new_[40393]_ ;
  assign \new_[40395]_  = \new_[40394]_  & \new_[40389]_ ;
  assign \new_[40399]_  = A269 & ~A267;
  assign \new_[40400]_  = ~A203 & \new_[40399]_ ;
  assign \new_[40403]_  = A299 & ~A298;
  assign \new_[40406]_  = A301 & A300;
  assign \new_[40407]_  = \new_[40406]_  & \new_[40403]_ ;
  assign \new_[40408]_  = \new_[40407]_  & \new_[40400]_ ;
  assign \new_[40412]_  = ~A199 & ~A166;
  assign \new_[40413]_  = ~A167 & \new_[40412]_ ;
  assign \new_[40417]_  = ~A202 & ~A201;
  assign \new_[40418]_  = A200 & \new_[40417]_ ;
  assign \new_[40419]_  = \new_[40418]_  & \new_[40413]_ ;
  assign \new_[40423]_  = A269 & ~A267;
  assign \new_[40424]_  = ~A203 & \new_[40423]_ ;
  assign \new_[40427]_  = A299 & ~A298;
  assign \new_[40430]_  = A302 & A300;
  assign \new_[40431]_  = \new_[40430]_  & \new_[40427]_ ;
  assign \new_[40432]_  = \new_[40431]_  & \new_[40424]_ ;
  assign \new_[40436]_  = ~A199 & ~A166;
  assign \new_[40437]_  = ~A167 & \new_[40436]_ ;
  assign \new_[40441]_  = ~A202 & ~A201;
  assign \new_[40442]_  = A200 & \new_[40441]_ ;
  assign \new_[40443]_  = \new_[40442]_  & \new_[40437]_ ;
  assign \new_[40447]_  = A266 & A265;
  assign \new_[40448]_  = ~A203 & \new_[40447]_ ;
  assign \new_[40451]_  = ~A299 & A298;
  assign \new_[40454]_  = A301 & A300;
  assign \new_[40455]_  = \new_[40454]_  & \new_[40451]_ ;
  assign \new_[40456]_  = \new_[40455]_  & \new_[40448]_ ;
  assign \new_[40460]_  = ~A199 & ~A166;
  assign \new_[40461]_  = ~A167 & \new_[40460]_ ;
  assign \new_[40465]_  = ~A202 & ~A201;
  assign \new_[40466]_  = A200 & \new_[40465]_ ;
  assign \new_[40467]_  = \new_[40466]_  & \new_[40461]_ ;
  assign \new_[40471]_  = A266 & A265;
  assign \new_[40472]_  = ~A203 & \new_[40471]_ ;
  assign \new_[40475]_  = ~A299 & A298;
  assign \new_[40478]_  = A302 & A300;
  assign \new_[40479]_  = \new_[40478]_  & \new_[40475]_ ;
  assign \new_[40480]_  = \new_[40479]_  & \new_[40472]_ ;
  assign \new_[40484]_  = ~A199 & ~A166;
  assign \new_[40485]_  = ~A167 & \new_[40484]_ ;
  assign \new_[40489]_  = ~A202 & ~A201;
  assign \new_[40490]_  = A200 & \new_[40489]_ ;
  assign \new_[40491]_  = \new_[40490]_  & \new_[40485]_ ;
  assign \new_[40495]_  = A266 & A265;
  assign \new_[40496]_  = ~A203 & \new_[40495]_ ;
  assign \new_[40499]_  = A299 & ~A298;
  assign \new_[40502]_  = A301 & A300;
  assign \new_[40503]_  = \new_[40502]_  & \new_[40499]_ ;
  assign \new_[40504]_  = \new_[40503]_  & \new_[40496]_ ;
  assign \new_[40508]_  = ~A199 & ~A166;
  assign \new_[40509]_  = ~A167 & \new_[40508]_ ;
  assign \new_[40513]_  = ~A202 & ~A201;
  assign \new_[40514]_  = A200 & \new_[40513]_ ;
  assign \new_[40515]_  = \new_[40514]_  & \new_[40509]_ ;
  assign \new_[40519]_  = A266 & A265;
  assign \new_[40520]_  = ~A203 & \new_[40519]_ ;
  assign \new_[40523]_  = A299 & ~A298;
  assign \new_[40526]_  = A302 & A300;
  assign \new_[40527]_  = \new_[40526]_  & \new_[40523]_ ;
  assign \new_[40528]_  = \new_[40527]_  & \new_[40520]_ ;
  assign \new_[40532]_  = ~A199 & ~A166;
  assign \new_[40533]_  = ~A167 & \new_[40532]_ ;
  assign \new_[40537]_  = ~A202 & ~A201;
  assign \new_[40538]_  = A200 & \new_[40537]_ ;
  assign \new_[40539]_  = \new_[40538]_  & \new_[40533]_ ;
  assign \new_[40543]_  = ~A266 & ~A265;
  assign \new_[40544]_  = ~A203 & \new_[40543]_ ;
  assign \new_[40547]_  = ~A299 & A298;
  assign \new_[40550]_  = A301 & A300;
  assign \new_[40551]_  = \new_[40550]_  & \new_[40547]_ ;
  assign \new_[40552]_  = \new_[40551]_  & \new_[40544]_ ;
  assign \new_[40556]_  = ~A199 & ~A166;
  assign \new_[40557]_  = ~A167 & \new_[40556]_ ;
  assign \new_[40561]_  = ~A202 & ~A201;
  assign \new_[40562]_  = A200 & \new_[40561]_ ;
  assign \new_[40563]_  = \new_[40562]_  & \new_[40557]_ ;
  assign \new_[40567]_  = ~A266 & ~A265;
  assign \new_[40568]_  = ~A203 & \new_[40567]_ ;
  assign \new_[40571]_  = ~A299 & A298;
  assign \new_[40574]_  = A302 & A300;
  assign \new_[40575]_  = \new_[40574]_  & \new_[40571]_ ;
  assign \new_[40576]_  = \new_[40575]_  & \new_[40568]_ ;
  assign \new_[40580]_  = ~A199 & ~A166;
  assign \new_[40581]_  = ~A167 & \new_[40580]_ ;
  assign \new_[40585]_  = ~A202 & ~A201;
  assign \new_[40586]_  = A200 & \new_[40585]_ ;
  assign \new_[40587]_  = \new_[40586]_  & \new_[40581]_ ;
  assign \new_[40591]_  = ~A266 & ~A265;
  assign \new_[40592]_  = ~A203 & \new_[40591]_ ;
  assign \new_[40595]_  = A299 & ~A298;
  assign \new_[40598]_  = A301 & A300;
  assign \new_[40599]_  = \new_[40598]_  & \new_[40595]_ ;
  assign \new_[40600]_  = \new_[40599]_  & \new_[40592]_ ;
  assign \new_[40604]_  = ~A199 & ~A166;
  assign \new_[40605]_  = ~A167 & \new_[40604]_ ;
  assign \new_[40609]_  = ~A202 & ~A201;
  assign \new_[40610]_  = A200 & \new_[40609]_ ;
  assign \new_[40611]_  = \new_[40610]_  & \new_[40605]_ ;
  assign \new_[40615]_  = ~A266 & ~A265;
  assign \new_[40616]_  = ~A203 & \new_[40615]_ ;
  assign \new_[40619]_  = A299 & ~A298;
  assign \new_[40622]_  = A302 & A300;
  assign \new_[40623]_  = \new_[40622]_  & \new_[40619]_ ;
  assign \new_[40624]_  = \new_[40623]_  & \new_[40616]_ ;
  assign \new_[40628]_  = A199 & ~A166;
  assign \new_[40629]_  = ~A167 & \new_[40628]_ ;
  assign \new_[40633]_  = A202 & A201;
  assign \new_[40634]_  = ~A200 & \new_[40633]_ ;
  assign \new_[40635]_  = \new_[40634]_  & \new_[40629]_ ;
  assign \new_[40639]_  = ~A269 & ~A268;
  assign \new_[40640]_  = A267 & \new_[40639]_ ;
  assign \new_[40643]_  = ~A299 & A298;
  assign \new_[40646]_  = A301 & A300;
  assign \new_[40647]_  = \new_[40646]_  & \new_[40643]_ ;
  assign \new_[40648]_  = \new_[40647]_  & \new_[40640]_ ;
  assign \new_[40652]_  = A199 & ~A166;
  assign \new_[40653]_  = ~A167 & \new_[40652]_ ;
  assign \new_[40657]_  = A202 & A201;
  assign \new_[40658]_  = ~A200 & \new_[40657]_ ;
  assign \new_[40659]_  = \new_[40658]_  & \new_[40653]_ ;
  assign \new_[40663]_  = ~A269 & ~A268;
  assign \new_[40664]_  = A267 & \new_[40663]_ ;
  assign \new_[40667]_  = ~A299 & A298;
  assign \new_[40670]_  = A302 & A300;
  assign \new_[40671]_  = \new_[40670]_  & \new_[40667]_ ;
  assign \new_[40672]_  = \new_[40671]_  & \new_[40664]_ ;
  assign \new_[40676]_  = A199 & ~A166;
  assign \new_[40677]_  = ~A167 & \new_[40676]_ ;
  assign \new_[40681]_  = A202 & A201;
  assign \new_[40682]_  = ~A200 & \new_[40681]_ ;
  assign \new_[40683]_  = \new_[40682]_  & \new_[40677]_ ;
  assign \new_[40687]_  = ~A269 & ~A268;
  assign \new_[40688]_  = A267 & \new_[40687]_ ;
  assign \new_[40691]_  = A299 & ~A298;
  assign \new_[40694]_  = A301 & A300;
  assign \new_[40695]_  = \new_[40694]_  & \new_[40691]_ ;
  assign \new_[40696]_  = \new_[40695]_  & \new_[40688]_ ;
  assign \new_[40700]_  = A199 & ~A166;
  assign \new_[40701]_  = ~A167 & \new_[40700]_ ;
  assign \new_[40705]_  = A202 & A201;
  assign \new_[40706]_  = ~A200 & \new_[40705]_ ;
  assign \new_[40707]_  = \new_[40706]_  & \new_[40701]_ ;
  assign \new_[40711]_  = ~A269 & ~A268;
  assign \new_[40712]_  = A267 & \new_[40711]_ ;
  assign \new_[40715]_  = A299 & ~A298;
  assign \new_[40718]_  = A302 & A300;
  assign \new_[40719]_  = \new_[40718]_  & \new_[40715]_ ;
  assign \new_[40720]_  = \new_[40719]_  & \new_[40712]_ ;
  assign \new_[40724]_  = A199 & ~A166;
  assign \new_[40725]_  = ~A167 & \new_[40724]_ ;
  assign \new_[40729]_  = A202 & A201;
  assign \new_[40730]_  = ~A200 & \new_[40729]_ ;
  assign \new_[40731]_  = \new_[40730]_  & \new_[40725]_ ;
  assign \new_[40735]_  = A298 & A268;
  assign \new_[40736]_  = ~A267 & \new_[40735]_ ;
  assign \new_[40739]_  = ~A300 & ~A299;
  assign \new_[40742]_  = ~A302 & ~A301;
  assign \new_[40743]_  = \new_[40742]_  & \new_[40739]_ ;
  assign \new_[40744]_  = \new_[40743]_  & \new_[40736]_ ;
  assign \new_[40748]_  = A199 & ~A166;
  assign \new_[40749]_  = ~A167 & \new_[40748]_ ;
  assign \new_[40753]_  = A202 & A201;
  assign \new_[40754]_  = ~A200 & \new_[40753]_ ;
  assign \new_[40755]_  = \new_[40754]_  & \new_[40749]_ ;
  assign \new_[40759]_  = ~A298 & A268;
  assign \new_[40760]_  = ~A267 & \new_[40759]_ ;
  assign \new_[40763]_  = ~A300 & A299;
  assign \new_[40766]_  = ~A302 & ~A301;
  assign \new_[40767]_  = \new_[40766]_  & \new_[40763]_ ;
  assign \new_[40768]_  = \new_[40767]_  & \new_[40760]_ ;
  assign \new_[40772]_  = A199 & ~A166;
  assign \new_[40773]_  = ~A167 & \new_[40772]_ ;
  assign \new_[40777]_  = A202 & A201;
  assign \new_[40778]_  = ~A200 & \new_[40777]_ ;
  assign \new_[40779]_  = \new_[40778]_  & \new_[40773]_ ;
  assign \new_[40783]_  = A298 & A269;
  assign \new_[40784]_  = ~A267 & \new_[40783]_ ;
  assign \new_[40787]_  = ~A300 & ~A299;
  assign \new_[40790]_  = ~A302 & ~A301;
  assign \new_[40791]_  = \new_[40790]_  & \new_[40787]_ ;
  assign \new_[40792]_  = \new_[40791]_  & \new_[40784]_ ;
  assign \new_[40796]_  = A199 & ~A166;
  assign \new_[40797]_  = ~A167 & \new_[40796]_ ;
  assign \new_[40801]_  = A202 & A201;
  assign \new_[40802]_  = ~A200 & \new_[40801]_ ;
  assign \new_[40803]_  = \new_[40802]_  & \new_[40797]_ ;
  assign \new_[40807]_  = ~A298 & A269;
  assign \new_[40808]_  = ~A267 & \new_[40807]_ ;
  assign \new_[40811]_  = ~A300 & A299;
  assign \new_[40814]_  = ~A302 & ~A301;
  assign \new_[40815]_  = \new_[40814]_  & \new_[40811]_ ;
  assign \new_[40816]_  = \new_[40815]_  & \new_[40808]_ ;
  assign \new_[40820]_  = A199 & ~A166;
  assign \new_[40821]_  = ~A167 & \new_[40820]_ ;
  assign \new_[40825]_  = A202 & A201;
  assign \new_[40826]_  = ~A200 & \new_[40825]_ ;
  assign \new_[40827]_  = \new_[40826]_  & \new_[40821]_ ;
  assign \new_[40831]_  = A298 & A266;
  assign \new_[40832]_  = A265 & \new_[40831]_ ;
  assign \new_[40835]_  = ~A300 & ~A299;
  assign \new_[40838]_  = ~A302 & ~A301;
  assign \new_[40839]_  = \new_[40838]_  & \new_[40835]_ ;
  assign \new_[40840]_  = \new_[40839]_  & \new_[40832]_ ;
  assign \new_[40844]_  = A199 & ~A166;
  assign \new_[40845]_  = ~A167 & \new_[40844]_ ;
  assign \new_[40849]_  = A202 & A201;
  assign \new_[40850]_  = ~A200 & \new_[40849]_ ;
  assign \new_[40851]_  = \new_[40850]_  & \new_[40845]_ ;
  assign \new_[40855]_  = ~A298 & A266;
  assign \new_[40856]_  = A265 & \new_[40855]_ ;
  assign \new_[40859]_  = ~A300 & A299;
  assign \new_[40862]_  = ~A302 & ~A301;
  assign \new_[40863]_  = \new_[40862]_  & \new_[40859]_ ;
  assign \new_[40864]_  = \new_[40863]_  & \new_[40856]_ ;
  assign \new_[40868]_  = A199 & ~A166;
  assign \new_[40869]_  = ~A167 & \new_[40868]_ ;
  assign \new_[40873]_  = A202 & A201;
  assign \new_[40874]_  = ~A200 & \new_[40873]_ ;
  assign \new_[40875]_  = \new_[40874]_  & \new_[40869]_ ;
  assign \new_[40879]_  = A298 & ~A266;
  assign \new_[40880]_  = ~A265 & \new_[40879]_ ;
  assign \new_[40883]_  = ~A300 & ~A299;
  assign \new_[40886]_  = ~A302 & ~A301;
  assign \new_[40887]_  = \new_[40886]_  & \new_[40883]_ ;
  assign \new_[40888]_  = \new_[40887]_  & \new_[40880]_ ;
  assign \new_[40892]_  = A199 & ~A166;
  assign \new_[40893]_  = ~A167 & \new_[40892]_ ;
  assign \new_[40897]_  = A202 & A201;
  assign \new_[40898]_  = ~A200 & \new_[40897]_ ;
  assign \new_[40899]_  = \new_[40898]_  & \new_[40893]_ ;
  assign \new_[40903]_  = ~A298 & ~A266;
  assign \new_[40904]_  = ~A265 & \new_[40903]_ ;
  assign \new_[40907]_  = ~A300 & A299;
  assign \new_[40910]_  = ~A302 & ~A301;
  assign \new_[40911]_  = \new_[40910]_  & \new_[40907]_ ;
  assign \new_[40912]_  = \new_[40911]_  & \new_[40904]_ ;
  assign \new_[40916]_  = A199 & ~A166;
  assign \new_[40917]_  = ~A167 & \new_[40916]_ ;
  assign \new_[40921]_  = A203 & A201;
  assign \new_[40922]_  = ~A200 & \new_[40921]_ ;
  assign \new_[40923]_  = \new_[40922]_  & \new_[40917]_ ;
  assign \new_[40927]_  = ~A269 & ~A268;
  assign \new_[40928]_  = A267 & \new_[40927]_ ;
  assign \new_[40931]_  = ~A299 & A298;
  assign \new_[40934]_  = A301 & A300;
  assign \new_[40935]_  = \new_[40934]_  & \new_[40931]_ ;
  assign \new_[40936]_  = \new_[40935]_  & \new_[40928]_ ;
  assign \new_[40940]_  = A199 & ~A166;
  assign \new_[40941]_  = ~A167 & \new_[40940]_ ;
  assign \new_[40945]_  = A203 & A201;
  assign \new_[40946]_  = ~A200 & \new_[40945]_ ;
  assign \new_[40947]_  = \new_[40946]_  & \new_[40941]_ ;
  assign \new_[40951]_  = ~A269 & ~A268;
  assign \new_[40952]_  = A267 & \new_[40951]_ ;
  assign \new_[40955]_  = ~A299 & A298;
  assign \new_[40958]_  = A302 & A300;
  assign \new_[40959]_  = \new_[40958]_  & \new_[40955]_ ;
  assign \new_[40960]_  = \new_[40959]_  & \new_[40952]_ ;
  assign \new_[40964]_  = A199 & ~A166;
  assign \new_[40965]_  = ~A167 & \new_[40964]_ ;
  assign \new_[40969]_  = A203 & A201;
  assign \new_[40970]_  = ~A200 & \new_[40969]_ ;
  assign \new_[40971]_  = \new_[40970]_  & \new_[40965]_ ;
  assign \new_[40975]_  = ~A269 & ~A268;
  assign \new_[40976]_  = A267 & \new_[40975]_ ;
  assign \new_[40979]_  = A299 & ~A298;
  assign \new_[40982]_  = A301 & A300;
  assign \new_[40983]_  = \new_[40982]_  & \new_[40979]_ ;
  assign \new_[40984]_  = \new_[40983]_  & \new_[40976]_ ;
  assign \new_[40988]_  = A199 & ~A166;
  assign \new_[40989]_  = ~A167 & \new_[40988]_ ;
  assign \new_[40993]_  = A203 & A201;
  assign \new_[40994]_  = ~A200 & \new_[40993]_ ;
  assign \new_[40995]_  = \new_[40994]_  & \new_[40989]_ ;
  assign \new_[40999]_  = ~A269 & ~A268;
  assign \new_[41000]_  = A267 & \new_[40999]_ ;
  assign \new_[41003]_  = A299 & ~A298;
  assign \new_[41006]_  = A302 & A300;
  assign \new_[41007]_  = \new_[41006]_  & \new_[41003]_ ;
  assign \new_[41008]_  = \new_[41007]_  & \new_[41000]_ ;
  assign \new_[41012]_  = A199 & ~A166;
  assign \new_[41013]_  = ~A167 & \new_[41012]_ ;
  assign \new_[41017]_  = A203 & A201;
  assign \new_[41018]_  = ~A200 & \new_[41017]_ ;
  assign \new_[41019]_  = \new_[41018]_  & \new_[41013]_ ;
  assign \new_[41023]_  = A298 & A268;
  assign \new_[41024]_  = ~A267 & \new_[41023]_ ;
  assign \new_[41027]_  = ~A300 & ~A299;
  assign \new_[41030]_  = ~A302 & ~A301;
  assign \new_[41031]_  = \new_[41030]_  & \new_[41027]_ ;
  assign \new_[41032]_  = \new_[41031]_  & \new_[41024]_ ;
  assign \new_[41036]_  = A199 & ~A166;
  assign \new_[41037]_  = ~A167 & \new_[41036]_ ;
  assign \new_[41041]_  = A203 & A201;
  assign \new_[41042]_  = ~A200 & \new_[41041]_ ;
  assign \new_[41043]_  = \new_[41042]_  & \new_[41037]_ ;
  assign \new_[41047]_  = ~A298 & A268;
  assign \new_[41048]_  = ~A267 & \new_[41047]_ ;
  assign \new_[41051]_  = ~A300 & A299;
  assign \new_[41054]_  = ~A302 & ~A301;
  assign \new_[41055]_  = \new_[41054]_  & \new_[41051]_ ;
  assign \new_[41056]_  = \new_[41055]_  & \new_[41048]_ ;
  assign \new_[41060]_  = A199 & ~A166;
  assign \new_[41061]_  = ~A167 & \new_[41060]_ ;
  assign \new_[41065]_  = A203 & A201;
  assign \new_[41066]_  = ~A200 & \new_[41065]_ ;
  assign \new_[41067]_  = \new_[41066]_  & \new_[41061]_ ;
  assign \new_[41071]_  = A298 & A269;
  assign \new_[41072]_  = ~A267 & \new_[41071]_ ;
  assign \new_[41075]_  = ~A300 & ~A299;
  assign \new_[41078]_  = ~A302 & ~A301;
  assign \new_[41079]_  = \new_[41078]_  & \new_[41075]_ ;
  assign \new_[41080]_  = \new_[41079]_  & \new_[41072]_ ;
  assign \new_[41084]_  = A199 & ~A166;
  assign \new_[41085]_  = ~A167 & \new_[41084]_ ;
  assign \new_[41089]_  = A203 & A201;
  assign \new_[41090]_  = ~A200 & \new_[41089]_ ;
  assign \new_[41091]_  = \new_[41090]_  & \new_[41085]_ ;
  assign \new_[41095]_  = ~A298 & A269;
  assign \new_[41096]_  = ~A267 & \new_[41095]_ ;
  assign \new_[41099]_  = ~A300 & A299;
  assign \new_[41102]_  = ~A302 & ~A301;
  assign \new_[41103]_  = \new_[41102]_  & \new_[41099]_ ;
  assign \new_[41104]_  = \new_[41103]_  & \new_[41096]_ ;
  assign \new_[41108]_  = A199 & ~A166;
  assign \new_[41109]_  = ~A167 & \new_[41108]_ ;
  assign \new_[41113]_  = A203 & A201;
  assign \new_[41114]_  = ~A200 & \new_[41113]_ ;
  assign \new_[41115]_  = \new_[41114]_  & \new_[41109]_ ;
  assign \new_[41119]_  = A298 & A266;
  assign \new_[41120]_  = A265 & \new_[41119]_ ;
  assign \new_[41123]_  = ~A300 & ~A299;
  assign \new_[41126]_  = ~A302 & ~A301;
  assign \new_[41127]_  = \new_[41126]_  & \new_[41123]_ ;
  assign \new_[41128]_  = \new_[41127]_  & \new_[41120]_ ;
  assign \new_[41132]_  = A199 & ~A166;
  assign \new_[41133]_  = ~A167 & \new_[41132]_ ;
  assign \new_[41137]_  = A203 & A201;
  assign \new_[41138]_  = ~A200 & \new_[41137]_ ;
  assign \new_[41139]_  = \new_[41138]_  & \new_[41133]_ ;
  assign \new_[41143]_  = ~A298 & A266;
  assign \new_[41144]_  = A265 & \new_[41143]_ ;
  assign \new_[41147]_  = ~A300 & A299;
  assign \new_[41150]_  = ~A302 & ~A301;
  assign \new_[41151]_  = \new_[41150]_  & \new_[41147]_ ;
  assign \new_[41152]_  = \new_[41151]_  & \new_[41144]_ ;
  assign \new_[41156]_  = A199 & ~A166;
  assign \new_[41157]_  = ~A167 & \new_[41156]_ ;
  assign \new_[41161]_  = A203 & A201;
  assign \new_[41162]_  = ~A200 & \new_[41161]_ ;
  assign \new_[41163]_  = \new_[41162]_  & \new_[41157]_ ;
  assign \new_[41167]_  = A298 & ~A266;
  assign \new_[41168]_  = ~A265 & \new_[41167]_ ;
  assign \new_[41171]_  = ~A300 & ~A299;
  assign \new_[41174]_  = ~A302 & ~A301;
  assign \new_[41175]_  = \new_[41174]_  & \new_[41171]_ ;
  assign \new_[41176]_  = \new_[41175]_  & \new_[41168]_ ;
  assign \new_[41180]_  = A199 & ~A166;
  assign \new_[41181]_  = ~A167 & \new_[41180]_ ;
  assign \new_[41185]_  = A203 & A201;
  assign \new_[41186]_  = ~A200 & \new_[41185]_ ;
  assign \new_[41187]_  = \new_[41186]_  & \new_[41181]_ ;
  assign \new_[41191]_  = ~A298 & ~A266;
  assign \new_[41192]_  = ~A265 & \new_[41191]_ ;
  assign \new_[41195]_  = ~A300 & A299;
  assign \new_[41198]_  = ~A302 & ~A301;
  assign \new_[41199]_  = \new_[41198]_  & \new_[41195]_ ;
  assign \new_[41200]_  = \new_[41199]_  & \new_[41192]_ ;
  assign \new_[41204]_  = A199 & ~A166;
  assign \new_[41205]_  = ~A167 & \new_[41204]_ ;
  assign \new_[41209]_  = ~A202 & ~A201;
  assign \new_[41210]_  = ~A200 & \new_[41209]_ ;
  assign \new_[41211]_  = \new_[41210]_  & \new_[41205]_ ;
  assign \new_[41215]_  = A268 & ~A267;
  assign \new_[41216]_  = ~A203 & \new_[41215]_ ;
  assign \new_[41219]_  = ~A299 & A298;
  assign \new_[41222]_  = A301 & A300;
  assign \new_[41223]_  = \new_[41222]_  & \new_[41219]_ ;
  assign \new_[41224]_  = \new_[41223]_  & \new_[41216]_ ;
  assign \new_[41228]_  = A199 & ~A166;
  assign \new_[41229]_  = ~A167 & \new_[41228]_ ;
  assign \new_[41233]_  = ~A202 & ~A201;
  assign \new_[41234]_  = ~A200 & \new_[41233]_ ;
  assign \new_[41235]_  = \new_[41234]_  & \new_[41229]_ ;
  assign \new_[41239]_  = A268 & ~A267;
  assign \new_[41240]_  = ~A203 & \new_[41239]_ ;
  assign \new_[41243]_  = ~A299 & A298;
  assign \new_[41246]_  = A302 & A300;
  assign \new_[41247]_  = \new_[41246]_  & \new_[41243]_ ;
  assign \new_[41248]_  = \new_[41247]_  & \new_[41240]_ ;
  assign \new_[41252]_  = A199 & ~A166;
  assign \new_[41253]_  = ~A167 & \new_[41252]_ ;
  assign \new_[41257]_  = ~A202 & ~A201;
  assign \new_[41258]_  = ~A200 & \new_[41257]_ ;
  assign \new_[41259]_  = \new_[41258]_  & \new_[41253]_ ;
  assign \new_[41263]_  = A268 & ~A267;
  assign \new_[41264]_  = ~A203 & \new_[41263]_ ;
  assign \new_[41267]_  = A299 & ~A298;
  assign \new_[41270]_  = A301 & A300;
  assign \new_[41271]_  = \new_[41270]_  & \new_[41267]_ ;
  assign \new_[41272]_  = \new_[41271]_  & \new_[41264]_ ;
  assign \new_[41276]_  = A199 & ~A166;
  assign \new_[41277]_  = ~A167 & \new_[41276]_ ;
  assign \new_[41281]_  = ~A202 & ~A201;
  assign \new_[41282]_  = ~A200 & \new_[41281]_ ;
  assign \new_[41283]_  = \new_[41282]_  & \new_[41277]_ ;
  assign \new_[41287]_  = A268 & ~A267;
  assign \new_[41288]_  = ~A203 & \new_[41287]_ ;
  assign \new_[41291]_  = A299 & ~A298;
  assign \new_[41294]_  = A302 & A300;
  assign \new_[41295]_  = \new_[41294]_  & \new_[41291]_ ;
  assign \new_[41296]_  = \new_[41295]_  & \new_[41288]_ ;
  assign \new_[41300]_  = A199 & ~A166;
  assign \new_[41301]_  = ~A167 & \new_[41300]_ ;
  assign \new_[41305]_  = ~A202 & ~A201;
  assign \new_[41306]_  = ~A200 & \new_[41305]_ ;
  assign \new_[41307]_  = \new_[41306]_  & \new_[41301]_ ;
  assign \new_[41311]_  = A269 & ~A267;
  assign \new_[41312]_  = ~A203 & \new_[41311]_ ;
  assign \new_[41315]_  = ~A299 & A298;
  assign \new_[41318]_  = A301 & A300;
  assign \new_[41319]_  = \new_[41318]_  & \new_[41315]_ ;
  assign \new_[41320]_  = \new_[41319]_  & \new_[41312]_ ;
  assign \new_[41324]_  = A199 & ~A166;
  assign \new_[41325]_  = ~A167 & \new_[41324]_ ;
  assign \new_[41329]_  = ~A202 & ~A201;
  assign \new_[41330]_  = ~A200 & \new_[41329]_ ;
  assign \new_[41331]_  = \new_[41330]_  & \new_[41325]_ ;
  assign \new_[41335]_  = A269 & ~A267;
  assign \new_[41336]_  = ~A203 & \new_[41335]_ ;
  assign \new_[41339]_  = ~A299 & A298;
  assign \new_[41342]_  = A302 & A300;
  assign \new_[41343]_  = \new_[41342]_  & \new_[41339]_ ;
  assign \new_[41344]_  = \new_[41343]_  & \new_[41336]_ ;
  assign \new_[41348]_  = A199 & ~A166;
  assign \new_[41349]_  = ~A167 & \new_[41348]_ ;
  assign \new_[41353]_  = ~A202 & ~A201;
  assign \new_[41354]_  = ~A200 & \new_[41353]_ ;
  assign \new_[41355]_  = \new_[41354]_  & \new_[41349]_ ;
  assign \new_[41359]_  = A269 & ~A267;
  assign \new_[41360]_  = ~A203 & \new_[41359]_ ;
  assign \new_[41363]_  = A299 & ~A298;
  assign \new_[41366]_  = A301 & A300;
  assign \new_[41367]_  = \new_[41366]_  & \new_[41363]_ ;
  assign \new_[41368]_  = \new_[41367]_  & \new_[41360]_ ;
  assign \new_[41372]_  = A199 & ~A166;
  assign \new_[41373]_  = ~A167 & \new_[41372]_ ;
  assign \new_[41377]_  = ~A202 & ~A201;
  assign \new_[41378]_  = ~A200 & \new_[41377]_ ;
  assign \new_[41379]_  = \new_[41378]_  & \new_[41373]_ ;
  assign \new_[41383]_  = A269 & ~A267;
  assign \new_[41384]_  = ~A203 & \new_[41383]_ ;
  assign \new_[41387]_  = A299 & ~A298;
  assign \new_[41390]_  = A302 & A300;
  assign \new_[41391]_  = \new_[41390]_  & \new_[41387]_ ;
  assign \new_[41392]_  = \new_[41391]_  & \new_[41384]_ ;
  assign \new_[41396]_  = A199 & ~A166;
  assign \new_[41397]_  = ~A167 & \new_[41396]_ ;
  assign \new_[41401]_  = ~A202 & ~A201;
  assign \new_[41402]_  = ~A200 & \new_[41401]_ ;
  assign \new_[41403]_  = \new_[41402]_  & \new_[41397]_ ;
  assign \new_[41407]_  = A266 & A265;
  assign \new_[41408]_  = ~A203 & \new_[41407]_ ;
  assign \new_[41411]_  = ~A299 & A298;
  assign \new_[41414]_  = A301 & A300;
  assign \new_[41415]_  = \new_[41414]_  & \new_[41411]_ ;
  assign \new_[41416]_  = \new_[41415]_  & \new_[41408]_ ;
  assign \new_[41420]_  = A199 & ~A166;
  assign \new_[41421]_  = ~A167 & \new_[41420]_ ;
  assign \new_[41425]_  = ~A202 & ~A201;
  assign \new_[41426]_  = ~A200 & \new_[41425]_ ;
  assign \new_[41427]_  = \new_[41426]_  & \new_[41421]_ ;
  assign \new_[41431]_  = A266 & A265;
  assign \new_[41432]_  = ~A203 & \new_[41431]_ ;
  assign \new_[41435]_  = ~A299 & A298;
  assign \new_[41438]_  = A302 & A300;
  assign \new_[41439]_  = \new_[41438]_  & \new_[41435]_ ;
  assign \new_[41440]_  = \new_[41439]_  & \new_[41432]_ ;
  assign \new_[41444]_  = A199 & ~A166;
  assign \new_[41445]_  = ~A167 & \new_[41444]_ ;
  assign \new_[41449]_  = ~A202 & ~A201;
  assign \new_[41450]_  = ~A200 & \new_[41449]_ ;
  assign \new_[41451]_  = \new_[41450]_  & \new_[41445]_ ;
  assign \new_[41455]_  = A266 & A265;
  assign \new_[41456]_  = ~A203 & \new_[41455]_ ;
  assign \new_[41459]_  = A299 & ~A298;
  assign \new_[41462]_  = A301 & A300;
  assign \new_[41463]_  = \new_[41462]_  & \new_[41459]_ ;
  assign \new_[41464]_  = \new_[41463]_  & \new_[41456]_ ;
  assign \new_[41468]_  = A199 & ~A166;
  assign \new_[41469]_  = ~A167 & \new_[41468]_ ;
  assign \new_[41473]_  = ~A202 & ~A201;
  assign \new_[41474]_  = ~A200 & \new_[41473]_ ;
  assign \new_[41475]_  = \new_[41474]_  & \new_[41469]_ ;
  assign \new_[41479]_  = A266 & A265;
  assign \new_[41480]_  = ~A203 & \new_[41479]_ ;
  assign \new_[41483]_  = A299 & ~A298;
  assign \new_[41486]_  = A302 & A300;
  assign \new_[41487]_  = \new_[41486]_  & \new_[41483]_ ;
  assign \new_[41488]_  = \new_[41487]_  & \new_[41480]_ ;
  assign \new_[41492]_  = A199 & ~A166;
  assign \new_[41493]_  = ~A167 & \new_[41492]_ ;
  assign \new_[41497]_  = ~A202 & ~A201;
  assign \new_[41498]_  = ~A200 & \new_[41497]_ ;
  assign \new_[41499]_  = \new_[41498]_  & \new_[41493]_ ;
  assign \new_[41503]_  = ~A266 & ~A265;
  assign \new_[41504]_  = ~A203 & \new_[41503]_ ;
  assign \new_[41507]_  = ~A299 & A298;
  assign \new_[41510]_  = A301 & A300;
  assign \new_[41511]_  = \new_[41510]_  & \new_[41507]_ ;
  assign \new_[41512]_  = \new_[41511]_  & \new_[41504]_ ;
  assign \new_[41516]_  = A199 & ~A166;
  assign \new_[41517]_  = ~A167 & \new_[41516]_ ;
  assign \new_[41521]_  = ~A202 & ~A201;
  assign \new_[41522]_  = ~A200 & \new_[41521]_ ;
  assign \new_[41523]_  = \new_[41522]_  & \new_[41517]_ ;
  assign \new_[41527]_  = ~A266 & ~A265;
  assign \new_[41528]_  = ~A203 & \new_[41527]_ ;
  assign \new_[41531]_  = ~A299 & A298;
  assign \new_[41534]_  = A302 & A300;
  assign \new_[41535]_  = \new_[41534]_  & \new_[41531]_ ;
  assign \new_[41536]_  = \new_[41535]_  & \new_[41528]_ ;
  assign \new_[41540]_  = A199 & ~A166;
  assign \new_[41541]_  = ~A167 & \new_[41540]_ ;
  assign \new_[41545]_  = ~A202 & ~A201;
  assign \new_[41546]_  = ~A200 & \new_[41545]_ ;
  assign \new_[41547]_  = \new_[41546]_  & \new_[41541]_ ;
  assign \new_[41551]_  = ~A266 & ~A265;
  assign \new_[41552]_  = ~A203 & \new_[41551]_ ;
  assign \new_[41555]_  = A299 & ~A298;
  assign \new_[41558]_  = A301 & A300;
  assign \new_[41559]_  = \new_[41558]_  & \new_[41555]_ ;
  assign \new_[41560]_  = \new_[41559]_  & \new_[41552]_ ;
  assign \new_[41564]_  = A199 & ~A166;
  assign \new_[41565]_  = ~A167 & \new_[41564]_ ;
  assign \new_[41569]_  = ~A202 & ~A201;
  assign \new_[41570]_  = ~A200 & \new_[41569]_ ;
  assign \new_[41571]_  = \new_[41570]_  & \new_[41565]_ ;
  assign \new_[41575]_  = ~A266 & ~A265;
  assign \new_[41576]_  = ~A203 & \new_[41575]_ ;
  assign \new_[41579]_  = A299 & ~A298;
  assign \new_[41582]_  = A302 & A300;
  assign \new_[41583]_  = \new_[41582]_  & \new_[41579]_ ;
  assign \new_[41584]_  = \new_[41583]_  & \new_[41576]_ ;
  assign \new_[41588]_  = A167 & A168;
  assign \new_[41589]_  = ~A170 & \new_[41588]_ ;
  assign \new_[41593]_  = ~A202 & A201;
  assign \new_[41594]_  = ~A166 & \new_[41593]_ ;
  assign \new_[41595]_  = \new_[41594]_  & \new_[41589]_ ;
  assign \new_[41599]_  = A268 & ~A267;
  assign \new_[41600]_  = ~A203 & \new_[41599]_ ;
  assign \new_[41603]_  = ~A299 & A298;
  assign \new_[41606]_  = A301 & A300;
  assign \new_[41607]_  = \new_[41606]_  & \new_[41603]_ ;
  assign \new_[41608]_  = \new_[41607]_  & \new_[41600]_ ;
  assign \new_[41612]_  = A167 & A168;
  assign \new_[41613]_  = ~A170 & \new_[41612]_ ;
  assign \new_[41617]_  = ~A202 & A201;
  assign \new_[41618]_  = ~A166 & \new_[41617]_ ;
  assign \new_[41619]_  = \new_[41618]_  & \new_[41613]_ ;
  assign \new_[41623]_  = A268 & ~A267;
  assign \new_[41624]_  = ~A203 & \new_[41623]_ ;
  assign \new_[41627]_  = ~A299 & A298;
  assign \new_[41630]_  = A302 & A300;
  assign \new_[41631]_  = \new_[41630]_  & \new_[41627]_ ;
  assign \new_[41632]_  = \new_[41631]_  & \new_[41624]_ ;
  assign \new_[41636]_  = A167 & A168;
  assign \new_[41637]_  = ~A170 & \new_[41636]_ ;
  assign \new_[41641]_  = ~A202 & A201;
  assign \new_[41642]_  = ~A166 & \new_[41641]_ ;
  assign \new_[41643]_  = \new_[41642]_  & \new_[41637]_ ;
  assign \new_[41647]_  = A268 & ~A267;
  assign \new_[41648]_  = ~A203 & \new_[41647]_ ;
  assign \new_[41651]_  = A299 & ~A298;
  assign \new_[41654]_  = A301 & A300;
  assign \new_[41655]_  = \new_[41654]_  & \new_[41651]_ ;
  assign \new_[41656]_  = \new_[41655]_  & \new_[41648]_ ;
  assign \new_[41660]_  = A167 & A168;
  assign \new_[41661]_  = ~A170 & \new_[41660]_ ;
  assign \new_[41665]_  = ~A202 & A201;
  assign \new_[41666]_  = ~A166 & \new_[41665]_ ;
  assign \new_[41667]_  = \new_[41666]_  & \new_[41661]_ ;
  assign \new_[41671]_  = A268 & ~A267;
  assign \new_[41672]_  = ~A203 & \new_[41671]_ ;
  assign \new_[41675]_  = A299 & ~A298;
  assign \new_[41678]_  = A302 & A300;
  assign \new_[41679]_  = \new_[41678]_  & \new_[41675]_ ;
  assign \new_[41680]_  = \new_[41679]_  & \new_[41672]_ ;
  assign \new_[41684]_  = A167 & A168;
  assign \new_[41685]_  = ~A170 & \new_[41684]_ ;
  assign \new_[41689]_  = ~A202 & A201;
  assign \new_[41690]_  = ~A166 & \new_[41689]_ ;
  assign \new_[41691]_  = \new_[41690]_  & \new_[41685]_ ;
  assign \new_[41695]_  = A269 & ~A267;
  assign \new_[41696]_  = ~A203 & \new_[41695]_ ;
  assign \new_[41699]_  = ~A299 & A298;
  assign \new_[41702]_  = A301 & A300;
  assign \new_[41703]_  = \new_[41702]_  & \new_[41699]_ ;
  assign \new_[41704]_  = \new_[41703]_  & \new_[41696]_ ;
  assign \new_[41708]_  = A167 & A168;
  assign \new_[41709]_  = ~A170 & \new_[41708]_ ;
  assign \new_[41713]_  = ~A202 & A201;
  assign \new_[41714]_  = ~A166 & \new_[41713]_ ;
  assign \new_[41715]_  = \new_[41714]_  & \new_[41709]_ ;
  assign \new_[41719]_  = A269 & ~A267;
  assign \new_[41720]_  = ~A203 & \new_[41719]_ ;
  assign \new_[41723]_  = ~A299 & A298;
  assign \new_[41726]_  = A302 & A300;
  assign \new_[41727]_  = \new_[41726]_  & \new_[41723]_ ;
  assign \new_[41728]_  = \new_[41727]_  & \new_[41720]_ ;
  assign \new_[41732]_  = A167 & A168;
  assign \new_[41733]_  = ~A170 & \new_[41732]_ ;
  assign \new_[41737]_  = ~A202 & A201;
  assign \new_[41738]_  = ~A166 & \new_[41737]_ ;
  assign \new_[41739]_  = \new_[41738]_  & \new_[41733]_ ;
  assign \new_[41743]_  = A269 & ~A267;
  assign \new_[41744]_  = ~A203 & \new_[41743]_ ;
  assign \new_[41747]_  = A299 & ~A298;
  assign \new_[41750]_  = A301 & A300;
  assign \new_[41751]_  = \new_[41750]_  & \new_[41747]_ ;
  assign \new_[41752]_  = \new_[41751]_  & \new_[41744]_ ;
  assign \new_[41756]_  = A167 & A168;
  assign \new_[41757]_  = ~A170 & \new_[41756]_ ;
  assign \new_[41761]_  = ~A202 & A201;
  assign \new_[41762]_  = ~A166 & \new_[41761]_ ;
  assign \new_[41763]_  = \new_[41762]_  & \new_[41757]_ ;
  assign \new_[41767]_  = A269 & ~A267;
  assign \new_[41768]_  = ~A203 & \new_[41767]_ ;
  assign \new_[41771]_  = A299 & ~A298;
  assign \new_[41774]_  = A302 & A300;
  assign \new_[41775]_  = \new_[41774]_  & \new_[41771]_ ;
  assign \new_[41776]_  = \new_[41775]_  & \new_[41768]_ ;
  assign \new_[41780]_  = A167 & A168;
  assign \new_[41781]_  = ~A170 & \new_[41780]_ ;
  assign \new_[41785]_  = ~A202 & A201;
  assign \new_[41786]_  = ~A166 & \new_[41785]_ ;
  assign \new_[41787]_  = \new_[41786]_  & \new_[41781]_ ;
  assign \new_[41791]_  = A266 & A265;
  assign \new_[41792]_  = ~A203 & \new_[41791]_ ;
  assign \new_[41795]_  = ~A299 & A298;
  assign \new_[41798]_  = A301 & A300;
  assign \new_[41799]_  = \new_[41798]_  & \new_[41795]_ ;
  assign \new_[41800]_  = \new_[41799]_  & \new_[41792]_ ;
  assign \new_[41804]_  = A167 & A168;
  assign \new_[41805]_  = ~A170 & \new_[41804]_ ;
  assign \new_[41809]_  = ~A202 & A201;
  assign \new_[41810]_  = ~A166 & \new_[41809]_ ;
  assign \new_[41811]_  = \new_[41810]_  & \new_[41805]_ ;
  assign \new_[41815]_  = A266 & A265;
  assign \new_[41816]_  = ~A203 & \new_[41815]_ ;
  assign \new_[41819]_  = ~A299 & A298;
  assign \new_[41822]_  = A302 & A300;
  assign \new_[41823]_  = \new_[41822]_  & \new_[41819]_ ;
  assign \new_[41824]_  = \new_[41823]_  & \new_[41816]_ ;
  assign \new_[41828]_  = A167 & A168;
  assign \new_[41829]_  = ~A170 & \new_[41828]_ ;
  assign \new_[41833]_  = ~A202 & A201;
  assign \new_[41834]_  = ~A166 & \new_[41833]_ ;
  assign \new_[41835]_  = \new_[41834]_  & \new_[41829]_ ;
  assign \new_[41839]_  = A266 & A265;
  assign \new_[41840]_  = ~A203 & \new_[41839]_ ;
  assign \new_[41843]_  = A299 & ~A298;
  assign \new_[41846]_  = A301 & A300;
  assign \new_[41847]_  = \new_[41846]_  & \new_[41843]_ ;
  assign \new_[41848]_  = \new_[41847]_  & \new_[41840]_ ;
  assign \new_[41852]_  = A167 & A168;
  assign \new_[41853]_  = ~A170 & \new_[41852]_ ;
  assign \new_[41857]_  = ~A202 & A201;
  assign \new_[41858]_  = ~A166 & \new_[41857]_ ;
  assign \new_[41859]_  = \new_[41858]_  & \new_[41853]_ ;
  assign \new_[41863]_  = A266 & A265;
  assign \new_[41864]_  = ~A203 & \new_[41863]_ ;
  assign \new_[41867]_  = A299 & ~A298;
  assign \new_[41870]_  = A302 & A300;
  assign \new_[41871]_  = \new_[41870]_  & \new_[41867]_ ;
  assign \new_[41872]_  = \new_[41871]_  & \new_[41864]_ ;
  assign \new_[41876]_  = A167 & A168;
  assign \new_[41877]_  = ~A170 & \new_[41876]_ ;
  assign \new_[41881]_  = ~A202 & A201;
  assign \new_[41882]_  = ~A166 & \new_[41881]_ ;
  assign \new_[41883]_  = \new_[41882]_  & \new_[41877]_ ;
  assign \new_[41887]_  = ~A266 & ~A265;
  assign \new_[41888]_  = ~A203 & \new_[41887]_ ;
  assign \new_[41891]_  = ~A299 & A298;
  assign \new_[41894]_  = A301 & A300;
  assign \new_[41895]_  = \new_[41894]_  & \new_[41891]_ ;
  assign \new_[41896]_  = \new_[41895]_  & \new_[41888]_ ;
  assign \new_[41900]_  = A167 & A168;
  assign \new_[41901]_  = ~A170 & \new_[41900]_ ;
  assign \new_[41905]_  = ~A202 & A201;
  assign \new_[41906]_  = ~A166 & \new_[41905]_ ;
  assign \new_[41907]_  = \new_[41906]_  & \new_[41901]_ ;
  assign \new_[41911]_  = ~A266 & ~A265;
  assign \new_[41912]_  = ~A203 & \new_[41911]_ ;
  assign \new_[41915]_  = ~A299 & A298;
  assign \new_[41918]_  = A302 & A300;
  assign \new_[41919]_  = \new_[41918]_  & \new_[41915]_ ;
  assign \new_[41920]_  = \new_[41919]_  & \new_[41912]_ ;
  assign \new_[41924]_  = A167 & A168;
  assign \new_[41925]_  = ~A170 & \new_[41924]_ ;
  assign \new_[41929]_  = ~A202 & A201;
  assign \new_[41930]_  = ~A166 & \new_[41929]_ ;
  assign \new_[41931]_  = \new_[41930]_  & \new_[41925]_ ;
  assign \new_[41935]_  = ~A266 & ~A265;
  assign \new_[41936]_  = ~A203 & \new_[41935]_ ;
  assign \new_[41939]_  = A299 & ~A298;
  assign \new_[41942]_  = A301 & A300;
  assign \new_[41943]_  = \new_[41942]_  & \new_[41939]_ ;
  assign \new_[41944]_  = \new_[41943]_  & \new_[41936]_ ;
  assign \new_[41948]_  = A167 & A168;
  assign \new_[41949]_  = ~A170 & \new_[41948]_ ;
  assign \new_[41953]_  = ~A202 & A201;
  assign \new_[41954]_  = ~A166 & \new_[41953]_ ;
  assign \new_[41955]_  = \new_[41954]_  & \new_[41949]_ ;
  assign \new_[41959]_  = ~A266 & ~A265;
  assign \new_[41960]_  = ~A203 & \new_[41959]_ ;
  assign \new_[41963]_  = A299 & ~A298;
  assign \new_[41966]_  = A302 & A300;
  assign \new_[41967]_  = \new_[41966]_  & \new_[41963]_ ;
  assign \new_[41968]_  = \new_[41967]_  & \new_[41960]_ ;
  assign \new_[41972]_  = A167 & A168;
  assign \new_[41973]_  = ~A170 & \new_[41972]_ ;
  assign \new_[41977]_  = A202 & ~A201;
  assign \new_[41978]_  = ~A166 & \new_[41977]_ ;
  assign \new_[41979]_  = \new_[41978]_  & \new_[41973]_ ;
  assign \new_[41983]_  = ~A269 & ~A268;
  assign \new_[41984]_  = A267 & \new_[41983]_ ;
  assign \new_[41987]_  = ~A299 & A298;
  assign \new_[41990]_  = A301 & A300;
  assign \new_[41991]_  = \new_[41990]_  & \new_[41987]_ ;
  assign \new_[41992]_  = \new_[41991]_  & \new_[41984]_ ;
  assign \new_[41996]_  = A167 & A168;
  assign \new_[41997]_  = ~A170 & \new_[41996]_ ;
  assign \new_[42001]_  = A202 & ~A201;
  assign \new_[42002]_  = ~A166 & \new_[42001]_ ;
  assign \new_[42003]_  = \new_[42002]_  & \new_[41997]_ ;
  assign \new_[42007]_  = ~A269 & ~A268;
  assign \new_[42008]_  = A267 & \new_[42007]_ ;
  assign \new_[42011]_  = ~A299 & A298;
  assign \new_[42014]_  = A302 & A300;
  assign \new_[42015]_  = \new_[42014]_  & \new_[42011]_ ;
  assign \new_[42016]_  = \new_[42015]_  & \new_[42008]_ ;
  assign \new_[42020]_  = A167 & A168;
  assign \new_[42021]_  = ~A170 & \new_[42020]_ ;
  assign \new_[42025]_  = A202 & ~A201;
  assign \new_[42026]_  = ~A166 & \new_[42025]_ ;
  assign \new_[42027]_  = \new_[42026]_  & \new_[42021]_ ;
  assign \new_[42031]_  = ~A269 & ~A268;
  assign \new_[42032]_  = A267 & \new_[42031]_ ;
  assign \new_[42035]_  = A299 & ~A298;
  assign \new_[42038]_  = A301 & A300;
  assign \new_[42039]_  = \new_[42038]_  & \new_[42035]_ ;
  assign \new_[42040]_  = \new_[42039]_  & \new_[42032]_ ;
  assign \new_[42044]_  = A167 & A168;
  assign \new_[42045]_  = ~A170 & \new_[42044]_ ;
  assign \new_[42049]_  = A202 & ~A201;
  assign \new_[42050]_  = ~A166 & \new_[42049]_ ;
  assign \new_[42051]_  = \new_[42050]_  & \new_[42045]_ ;
  assign \new_[42055]_  = ~A269 & ~A268;
  assign \new_[42056]_  = A267 & \new_[42055]_ ;
  assign \new_[42059]_  = A299 & ~A298;
  assign \new_[42062]_  = A302 & A300;
  assign \new_[42063]_  = \new_[42062]_  & \new_[42059]_ ;
  assign \new_[42064]_  = \new_[42063]_  & \new_[42056]_ ;
  assign \new_[42068]_  = A167 & A168;
  assign \new_[42069]_  = ~A170 & \new_[42068]_ ;
  assign \new_[42073]_  = A202 & ~A201;
  assign \new_[42074]_  = ~A166 & \new_[42073]_ ;
  assign \new_[42075]_  = \new_[42074]_  & \new_[42069]_ ;
  assign \new_[42079]_  = A298 & A268;
  assign \new_[42080]_  = ~A267 & \new_[42079]_ ;
  assign \new_[42083]_  = ~A300 & ~A299;
  assign \new_[42086]_  = ~A302 & ~A301;
  assign \new_[42087]_  = \new_[42086]_  & \new_[42083]_ ;
  assign \new_[42088]_  = \new_[42087]_  & \new_[42080]_ ;
  assign \new_[42092]_  = A167 & A168;
  assign \new_[42093]_  = ~A170 & \new_[42092]_ ;
  assign \new_[42097]_  = A202 & ~A201;
  assign \new_[42098]_  = ~A166 & \new_[42097]_ ;
  assign \new_[42099]_  = \new_[42098]_  & \new_[42093]_ ;
  assign \new_[42103]_  = ~A298 & A268;
  assign \new_[42104]_  = ~A267 & \new_[42103]_ ;
  assign \new_[42107]_  = ~A300 & A299;
  assign \new_[42110]_  = ~A302 & ~A301;
  assign \new_[42111]_  = \new_[42110]_  & \new_[42107]_ ;
  assign \new_[42112]_  = \new_[42111]_  & \new_[42104]_ ;
  assign \new_[42116]_  = A167 & A168;
  assign \new_[42117]_  = ~A170 & \new_[42116]_ ;
  assign \new_[42121]_  = A202 & ~A201;
  assign \new_[42122]_  = ~A166 & \new_[42121]_ ;
  assign \new_[42123]_  = \new_[42122]_  & \new_[42117]_ ;
  assign \new_[42127]_  = A298 & A269;
  assign \new_[42128]_  = ~A267 & \new_[42127]_ ;
  assign \new_[42131]_  = ~A300 & ~A299;
  assign \new_[42134]_  = ~A302 & ~A301;
  assign \new_[42135]_  = \new_[42134]_  & \new_[42131]_ ;
  assign \new_[42136]_  = \new_[42135]_  & \new_[42128]_ ;
  assign \new_[42140]_  = A167 & A168;
  assign \new_[42141]_  = ~A170 & \new_[42140]_ ;
  assign \new_[42145]_  = A202 & ~A201;
  assign \new_[42146]_  = ~A166 & \new_[42145]_ ;
  assign \new_[42147]_  = \new_[42146]_  & \new_[42141]_ ;
  assign \new_[42151]_  = ~A298 & A269;
  assign \new_[42152]_  = ~A267 & \new_[42151]_ ;
  assign \new_[42155]_  = ~A300 & A299;
  assign \new_[42158]_  = ~A302 & ~A301;
  assign \new_[42159]_  = \new_[42158]_  & \new_[42155]_ ;
  assign \new_[42160]_  = \new_[42159]_  & \new_[42152]_ ;
  assign \new_[42164]_  = A167 & A168;
  assign \new_[42165]_  = ~A170 & \new_[42164]_ ;
  assign \new_[42169]_  = A202 & ~A201;
  assign \new_[42170]_  = ~A166 & \new_[42169]_ ;
  assign \new_[42171]_  = \new_[42170]_  & \new_[42165]_ ;
  assign \new_[42175]_  = A298 & A266;
  assign \new_[42176]_  = A265 & \new_[42175]_ ;
  assign \new_[42179]_  = ~A300 & ~A299;
  assign \new_[42182]_  = ~A302 & ~A301;
  assign \new_[42183]_  = \new_[42182]_  & \new_[42179]_ ;
  assign \new_[42184]_  = \new_[42183]_  & \new_[42176]_ ;
  assign \new_[42188]_  = A167 & A168;
  assign \new_[42189]_  = ~A170 & \new_[42188]_ ;
  assign \new_[42193]_  = A202 & ~A201;
  assign \new_[42194]_  = ~A166 & \new_[42193]_ ;
  assign \new_[42195]_  = \new_[42194]_  & \new_[42189]_ ;
  assign \new_[42199]_  = ~A298 & A266;
  assign \new_[42200]_  = A265 & \new_[42199]_ ;
  assign \new_[42203]_  = ~A300 & A299;
  assign \new_[42206]_  = ~A302 & ~A301;
  assign \new_[42207]_  = \new_[42206]_  & \new_[42203]_ ;
  assign \new_[42208]_  = \new_[42207]_  & \new_[42200]_ ;
  assign \new_[42212]_  = A167 & A168;
  assign \new_[42213]_  = ~A170 & \new_[42212]_ ;
  assign \new_[42217]_  = A202 & ~A201;
  assign \new_[42218]_  = ~A166 & \new_[42217]_ ;
  assign \new_[42219]_  = \new_[42218]_  & \new_[42213]_ ;
  assign \new_[42223]_  = A298 & ~A266;
  assign \new_[42224]_  = ~A265 & \new_[42223]_ ;
  assign \new_[42227]_  = ~A300 & ~A299;
  assign \new_[42230]_  = ~A302 & ~A301;
  assign \new_[42231]_  = \new_[42230]_  & \new_[42227]_ ;
  assign \new_[42232]_  = \new_[42231]_  & \new_[42224]_ ;
  assign \new_[42236]_  = A167 & A168;
  assign \new_[42237]_  = ~A170 & \new_[42236]_ ;
  assign \new_[42241]_  = A202 & ~A201;
  assign \new_[42242]_  = ~A166 & \new_[42241]_ ;
  assign \new_[42243]_  = \new_[42242]_  & \new_[42237]_ ;
  assign \new_[42247]_  = ~A298 & ~A266;
  assign \new_[42248]_  = ~A265 & \new_[42247]_ ;
  assign \new_[42251]_  = ~A300 & A299;
  assign \new_[42254]_  = ~A302 & ~A301;
  assign \new_[42255]_  = \new_[42254]_  & \new_[42251]_ ;
  assign \new_[42256]_  = \new_[42255]_  & \new_[42248]_ ;
  assign \new_[42260]_  = A167 & A168;
  assign \new_[42261]_  = ~A170 & \new_[42260]_ ;
  assign \new_[42265]_  = A203 & ~A201;
  assign \new_[42266]_  = ~A166 & \new_[42265]_ ;
  assign \new_[42267]_  = \new_[42266]_  & \new_[42261]_ ;
  assign \new_[42271]_  = ~A269 & ~A268;
  assign \new_[42272]_  = A267 & \new_[42271]_ ;
  assign \new_[42275]_  = ~A299 & A298;
  assign \new_[42278]_  = A301 & A300;
  assign \new_[42279]_  = \new_[42278]_  & \new_[42275]_ ;
  assign \new_[42280]_  = \new_[42279]_  & \new_[42272]_ ;
  assign \new_[42284]_  = A167 & A168;
  assign \new_[42285]_  = ~A170 & \new_[42284]_ ;
  assign \new_[42289]_  = A203 & ~A201;
  assign \new_[42290]_  = ~A166 & \new_[42289]_ ;
  assign \new_[42291]_  = \new_[42290]_  & \new_[42285]_ ;
  assign \new_[42295]_  = ~A269 & ~A268;
  assign \new_[42296]_  = A267 & \new_[42295]_ ;
  assign \new_[42299]_  = ~A299 & A298;
  assign \new_[42302]_  = A302 & A300;
  assign \new_[42303]_  = \new_[42302]_  & \new_[42299]_ ;
  assign \new_[42304]_  = \new_[42303]_  & \new_[42296]_ ;
  assign \new_[42308]_  = A167 & A168;
  assign \new_[42309]_  = ~A170 & \new_[42308]_ ;
  assign \new_[42313]_  = A203 & ~A201;
  assign \new_[42314]_  = ~A166 & \new_[42313]_ ;
  assign \new_[42315]_  = \new_[42314]_  & \new_[42309]_ ;
  assign \new_[42319]_  = ~A269 & ~A268;
  assign \new_[42320]_  = A267 & \new_[42319]_ ;
  assign \new_[42323]_  = A299 & ~A298;
  assign \new_[42326]_  = A301 & A300;
  assign \new_[42327]_  = \new_[42326]_  & \new_[42323]_ ;
  assign \new_[42328]_  = \new_[42327]_  & \new_[42320]_ ;
  assign \new_[42332]_  = A167 & A168;
  assign \new_[42333]_  = ~A170 & \new_[42332]_ ;
  assign \new_[42337]_  = A203 & ~A201;
  assign \new_[42338]_  = ~A166 & \new_[42337]_ ;
  assign \new_[42339]_  = \new_[42338]_  & \new_[42333]_ ;
  assign \new_[42343]_  = ~A269 & ~A268;
  assign \new_[42344]_  = A267 & \new_[42343]_ ;
  assign \new_[42347]_  = A299 & ~A298;
  assign \new_[42350]_  = A302 & A300;
  assign \new_[42351]_  = \new_[42350]_  & \new_[42347]_ ;
  assign \new_[42352]_  = \new_[42351]_  & \new_[42344]_ ;
  assign \new_[42356]_  = A167 & A168;
  assign \new_[42357]_  = ~A170 & \new_[42356]_ ;
  assign \new_[42361]_  = A203 & ~A201;
  assign \new_[42362]_  = ~A166 & \new_[42361]_ ;
  assign \new_[42363]_  = \new_[42362]_  & \new_[42357]_ ;
  assign \new_[42367]_  = A298 & A268;
  assign \new_[42368]_  = ~A267 & \new_[42367]_ ;
  assign \new_[42371]_  = ~A300 & ~A299;
  assign \new_[42374]_  = ~A302 & ~A301;
  assign \new_[42375]_  = \new_[42374]_  & \new_[42371]_ ;
  assign \new_[42376]_  = \new_[42375]_  & \new_[42368]_ ;
  assign \new_[42380]_  = A167 & A168;
  assign \new_[42381]_  = ~A170 & \new_[42380]_ ;
  assign \new_[42385]_  = A203 & ~A201;
  assign \new_[42386]_  = ~A166 & \new_[42385]_ ;
  assign \new_[42387]_  = \new_[42386]_  & \new_[42381]_ ;
  assign \new_[42391]_  = ~A298 & A268;
  assign \new_[42392]_  = ~A267 & \new_[42391]_ ;
  assign \new_[42395]_  = ~A300 & A299;
  assign \new_[42398]_  = ~A302 & ~A301;
  assign \new_[42399]_  = \new_[42398]_  & \new_[42395]_ ;
  assign \new_[42400]_  = \new_[42399]_  & \new_[42392]_ ;
  assign \new_[42404]_  = A167 & A168;
  assign \new_[42405]_  = ~A170 & \new_[42404]_ ;
  assign \new_[42409]_  = A203 & ~A201;
  assign \new_[42410]_  = ~A166 & \new_[42409]_ ;
  assign \new_[42411]_  = \new_[42410]_  & \new_[42405]_ ;
  assign \new_[42415]_  = A298 & A269;
  assign \new_[42416]_  = ~A267 & \new_[42415]_ ;
  assign \new_[42419]_  = ~A300 & ~A299;
  assign \new_[42422]_  = ~A302 & ~A301;
  assign \new_[42423]_  = \new_[42422]_  & \new_[42419]_ ;
  assign \new_[42424]_  = \new_[42423]_  & \new_[42416]_ ;
  assign \new_[42428]_  = A167 & A168;
  assign \new_[42429]_  = ~A170 & \new_[42428]_ ;
  assign \new_[42433]_  = A203 & ~A201;
  assign \new_[42434]_  = ~A166 & \new_[42433]_ ;
  assign \new_[42435]_  = \new_[42434]_  & \new_[42429]_ ;
  assign \new_[42439]_  = ~A298 & A269;
  assign \new_[42440]_  = ~A267 & \new_[42439]_ ;
  assign \new_[42443]_  = ~A300 & A299;
  assign \new_[42446]_  = ~A302 & ~A301;
  assign \new_[42447]_  = \new_[42446]_  & \new_[42443]_ ;
  assign \new_[42448]_  = \new_[42447]_  & \new_[42440]_ ;
  assign \new_[42452]_  = A167 & A168;
  assign \new_[42453]_  = ~A170 & \new_[42452]_ ;
  assign \new_[42457]_  = A203 & ~A201;
  assign \new_[42458]_  = ~A166 & \new_[42457]_ ;
  assign \new_[42459]_  = \new_[42458]_  & \new_[42453]_ ;
  assign \new_[42463]_  = A298 & A266;
  assign \new_[42464]_  = A265 & \new_[42463]_ ;
  assign \new_[42467]_  = ~A300 & ~A299;
  assign \new_[42470]_  = ~A302 & ~A301;
  assign \new_[42471]_  = \new_[42470]_  & \new_[42467]_ ;
  assign \new_[42472]_  = \new_[42471]_  & \new_[42464]_ ;
  assign \new_[42476]_  = A167 & A168;
  assign \new_[42477]_  = ~A170 & \new_[42476]_ ;
  assign \new_[42481]_  = A203 & ~A201;
  assign \new_[42482]_  = ~A166 & \new_[42481]_ ;
  assign \new_[42483]_  = \new_[42482]_  & \new_[42477]_ ;
  assign \new_[42487]_  = ~A298 & A266;
  assign \new_[42488]_  = A265 & \new_[42487]_ ;
  assign \new_[42491]_  = ~A300 & A299;
  assign \new_[42494]_  = ~A302 & ~A301;
  assign \new_[42495]_  = \new_[42494]_  & \new_[42491]_ ;
  assign \new_[42496]_  = \new_[42495]_  & \new_[42488]_ ;
  assign \new_[42500]_  = A167 & A168;
  assign \new_[42501]_  = ~A170 & \new_[42500]_ ;
  assign \new_[42505]_  = A203 & ~A201;
  assign \new_[42506]_  = ~A166 & \new_[42505]_ ;
  assign \new_[42507]_  = \new_[42506]_  & \new_[42501]_ ;
  assign \new_[42511]_  = A298 & ~A266;
  assign \new_[42512]_  = ~A265 & \new_[42511]_ ;
  assign \new_[42515]_  = ~A300 & ~A299;
  assign \new_[42518]_  = ~A302 & ~A301;
  assign \new_[42519]_  = \new_[42518]_  & \new_[42515]_ ;
  assign \new_[42520]_  = \new_[42519]_  & \new_[42512]_ ;
  assign \new_[42524]_  = A167 & A168;
  assign \new_[42525]_  = ~A170 & \new_[42524]_ ;
  assign \new_[42529]_  = A203 & ~A201;
  assign \new_[42530]_  = ~A166 & \new_[42529]_ ;
  assign \new_[42531]_  = \new_[42530]_  & \new_[42525]_ ;
  assign \new_[42535]_  = ~A298 & ~A266;
  assign \new_[42536]_  = ~A265 & \new_[42535]_ ;
  assign \new_[42539]_  = ~A300 & A299;
  assign \new_[42542]_  = ~A302 & ~A301;
  assign \new_[42543]_  = \new_[42542]_  & \new_[42539]_ ;
  assign \new_[42544]_  = \new_[42543]_  & \new_[42536]_ ;
  assign \new_[42548]_  = A167 & A168;
  assign \new_[42549]_  = ~A170 & \new_[42548]_ ;
  assign \new_[42553]_  = A200 & A199;
  assign \new_[42554]_  = ~A166 & \new_[42553]_ ;
  assign \new_[42555]_  = \new_[42554]_  & \new_[42549]_ ;
  assign \new_[42559]_  = ~A269 & ~A268;
  assign \new_[42560]_  = A267 & \new_[42559]_ ;
  assign \new_[42563]_  = ~A299 & A298;
  assign \new_[42566]_  = A301 & A300;
  assign \new_[42567]_  = \new_[42566]_  & \new_[42563]_ ;
  assign \new_[42568]_  = \new_[42567]_  & \new_[42560]_ ;
  assign \new_[42572]_  = A167 & A168;
  assign \new_[42573]_  = ~A170 & \new_[42572]_ ;
  assign \new_[42577]_  = A200 & A199;
  assign \new_[42578]_  = ~A166 & \new_[42577]_ ;
  assign \new_[42579]_  = \new_[42578]_  & \new_[42573]_ ;
  assign \new_[42583]_  = ~A269 & ~A268;
  assign \new_[42584]_  = A267 & \new_[42583]_ ;
  assign \new_[42587]_  = ~A299 & A298;
  assign \new_[42590]_  = A302 & A300;
  assign \new_[42591]_  = \new_[42590]_  & \new_[42587]_ ;
  assign \new_[42592]_  = \new_[42591]_  & \new_[42584]_ ;
  assign \new_[42596]_  = A167 & A168;
  assign \new_[42597]_  = ~A170 & \new_[42596]_ ;
  assign \new_[42601]_  = A200 & A199;
  assign \new_[42602]_  = ~A166 & \new_[42601]_ ;
  assign \new_[42603]_  = \new_[42602]_  & \new_[42597]_ ;
  assign \new_[42607]_  = ~A269 & ~A268;
  assign \new_[42608]_  = A267 & \new_[42607]_ ;
  assign \new_[42611]_  = A299 & ~A298;
  assign \new_[42614]_  = A301 & A300;
  assign \new_[42615]_  = \new_[42614]_  & \new_[42611]_ ;
  assign \new_[42616]_  = \new_[42615]_  & \new_[42608]_ ;
  assign \new_[42620]_  = A167 & A168;
  assign \new_[42621]_  = ~A170 & \new_[42620]_ ;
  assign \new_[42625]_  = A200 & A199;
  assign \new_[42626]_  = ~A166 & \new_[42625]_ ;
  assign \new_[42627]_  = \new_[42626]_  & \new_[42621]_ ;
  assign \new_[42631]_  = ~A269 & ~A268;
  assign \new_[42632]_  = A267 & \new_[42631]_ ;
  assign \new_[42635]_  = A299 & ~A298;
  assign \new_[42638]_  = A302 & A300;
  assign \new_[42639]_  = \new_[42638]_  & \new_[42635]_ ;
  assign \new_[42640]_  = \new_[42639]_  & \new_[42632]_ ;
  assign \new_[42644]_  = A167 & A168;
  assign \new_[42645]_  = ~A170 & \new_[42644]_ ;
  assign \new_[42649]_  = A200 & A199;
  assign \new_[42650]_  = ~A166 & \new_[42649]_ ;
  assign \new_[42651]_  = \new_[42650]_  & \new_[42645]_ ;
  assign \new_[42655]_  = A298 & A268;
  assign \new_[42656]_  = ~A267 & \new_[42655]_ ;
  assign \new_[42659]_  = ~A300 & ~A299;
  assign \new_[42662]_  = ~A302 & ~A301;
  assign \new_[42663]_  = \new_[42662]_  & \new_[42659]_ ;
  assign \new_[42664]_  = \new_[42663]_  & \new_[42656]_ ;
  assign \new_[42668]_  = A167 & A168;
  assign \new_[42669]_  = ~A170 & \new_[42668]_ ;
  assign \new_[42673]_  = A200 & A199;
  assign \new_[42674]_  = ~A166 & \new_[42673]_ ;
  assign \new_[42675]_  = \new_[42674]_  & \new_[42669]_ ;
  assign \new_[42679]_  = ~A298 & A268;
  assign \new_[42680]_  = ~A267 & \new_[42679]_ ;
  assign \new_[42683]_  = ~A300 & A299;
  assign \new_[42686]_  = ~A302 & ~A301;
  assign \new_[42687]_  = \new_[42686]_  & \new_[42683]_ ;
  assign \new_[42688]_  = \new_[42687]_  & \new_[42680]_ ;
  assign \new_[42692]_  = A167 & A168;
  assign \new_[42693]_  = ~A170 & \new_[42692]_ ;
  assign \new_[42697]_  = A200 & A199;
  assign \new_[42698]_  = ~A166 & \new_[42697]_ ;
  assign \new_[42699]_  = \new_[42698]_  & \new_[42693]_ ;
  assign \new_[42703]_  = A298 & A269;
  assign \new_[42704]_  = ~A267 & \new_[42703]_ ;
  assign \new_[42707]_  = ~A300 & ~A299;
  assign \new_[42710]_  = ~A302 & ~A301;
  assign \new_[42711]_  = \new_[42710]_  & \new_[42707]_ ;
  assign \new_[42712]_  = \new_[42711]_  & \new_[42704]_ ;
  assign \new_[42716]_  = A167 & A168;
  assign \new_[42717]_  = ~A170 & \new_[42716]_ ;
  assign \new_[42721]_  = A200 & A199;
  assign \new_[42722]_  = ~A166 & \new_[42721]_ ;
  assign \new_[42723]_  = \new_[42722]_  & \new_[42717]_ ;
  assign \new_[42727]_  = ~A298 & A269;
  assign \new_[42728]_  = ~A267 & \new_[42727]_ ;
  assign \new_[42731]_  = ~A300 & A299;
  assign \new_[42734]_  = ~A302 & ~A301;
  assign \new_[42735]_  = \new_[42734]_  & \new_[42731]_ ;
  assign \new_[42736]_  = \new_[42735]_  & \new_[42728]_ ;
  assign \new_[42740]_  = A167 & A168;
  assign \new_[42741]_  = ~A170 & \new_[42740]_ ;
  assign \new_[42745]_  = A200 & A199;
  assign \new_[42746]_  = ~A166 & \new_[42745]_ ;
  assign \new_[42747]_  = \new_[42746]_  & \new_[42741]_ ;
  assign \new_[42751]_  = A298 & A266;
  assign \new_[42752]_  = A265 & \new_[42751]_ ;
  assign \new_[42755]_  = ~A300 & ~A299;
  assign \new_[42758]_  = ~A302 & ~A301;
  assign \new_[42759]_  = \new_[42758]_  & \new_[42755]_ ;
  assign \new_[42760]_  = \new_[42759]_  & \new_[42752]_ ;
  assign \new_[42764]_  = A167 & A168;
  assign \new_[42765]_  = ~A170 & \new_[42764]_ ;
  assign \new_[42769]_  = A200 & A199;
  assign \new_[42770]_  = ~A166 & \new_[42769]_ ;
  assign \new_[42771]_  = \new_[42770]_  & \new_[42765]_ ;
  assign \new_[42775]_  = ~A298 & A266;
  assign \new_[42776]_  = A265 & \new_[42775]_ ;
  assign \new_[42779]_  = ~A300 & A299;
  assign \new_[42782]_  = ~A302 & ~A301;
  assign \new_[42783]_  = \new_[42782]_  & \new_[42779]_ ;
  assign \new_[42784]_  = \new_[42783]_  & \new_[42776]_ ;
  assign \new_[42788]_  = A167 & A168;
  assign \new_[42789]_  = ~A170 & \new_[42788]_ ;
  assign \new_[42793]_  = A200 & A199;
  assign \new_[42794]_  = ~A166 & \new_[42793]_ ;
  assign \new_[42795]_  = \new_[42794]_  & \new_[42789]_ ;
  assign \new_[42799]_  = A298 & ~A266;
  assign \new_[42800]_  = ~A265 & \new_[42799]_ ;
  assign \new_[42803]_  = ~A300 & ~A299;
  assign \new_[42806]_  = ~A302 & ~A301;
  assign \new_[42807]_  = \new_[42806]_  & \new_[42803]_ ;
  assign \new_[42808]_  = \new_[42807]_  & \new_[42800]_ ;
  assign \new_[42812]_  = A167 & A168;
  assign \new_[42813]_  = ~A170 & \new_[42812]_ ;
  assign \new_[42817]_  = A200 & A199;
  assign \new_[42818]_  = ~A166 & \new_[42817]_ ;
  assign \new_[42819]_  = \new_[42818]_  & \new_[42813]_ ;
  assign \new_[42823]_  = ~A298 & ~A266;
  assign \new_[42824]_  = ~A265 & \new_[42823]_ ;
  assign \new_[42827]_  = ~A300 & A299;
  assign \new_[42830]_  = ~A302 & ~A301;
  assign \new_[42831]_  = \new_[42830]_  & \new_[42827]_ ;
  assign \new_[42832]_  = \new_[42831]_  & \new_[42824]_ ;
  assign \new_[42836]_  = A167 & A168;
  assign \new_[42837]_  = ~A170 & \new_[42836]_ ;
  assign \new_[42841]_  = ~A200 & ~A199;
  assign \new_[42842]_  = ~A166 & \new_[42841]_ ;
  assign \new_[42843]_  = \new_[42842]_  & \new_[42837]_ ;
  assign \new_[42847]_  = ~A269 & ~A268;
  assign \new_[42848]_  = A267 & \new_[42847]_ ;
  assign \new_[42851]_  = ~A299 & A298;
  assign \new_[42854]_  = A301 & A300;
  assign \new_[42855]_  = \new_[42854]_  & \new_[42851]_ ;
  assign \new_[42856]_  = \new_[42855]_  & \new_[42848]_ ;
  assign \new_[42860]_  = A167 & A168;
  assign \new_[42861]_  = ~A170 & \new_[42860]_ ;
  assign \new_[42865]_  = ~A200 & ~A199;
  assign \new_[42866]_  = ~A166 & \new_[42865]_ ;
  assign \new_[42867]_  = \new_[42866]_  & \new_[42861]_ ;
  assign \new_[42871]_  = ~A269 & ~A268;
  assign \new_[42872]_  = A267 & \new_[42871]_ ;
  assign \new_[42875]_  = ~A299 & A298;
  assign \new_[42878]_  = A302 & A300;
  assign \new_[42879]_  = \new_[42878]_  & \new_[42875]_ ;
  assign \new_[42880]_  = \new_[42879]_  & \new_[42872]_ ;
  assign \new_[42884]_  = A167 & A168;
  assign \new_[42885]_  = ~A170 & \new_[42884]_ ;
  assign \new_[42889]_  = ~A200 & ~A199;
  assign \new_[42890]_  = ~A166 & \new_[42889]_ ;
  assign \new_[42891]_  = \new_[42890]_  & \new_[42885]_ ;
  assign \new_[42895]_  = ~A269 & ~A268;
  assign \new_[42896]_  = A267 & \new_[42895]_ ;
  assign \new_[42899]_  = A299 & ~A298;
  assign \new_[42902]_  = A301 & A300;
  assign \new_[42903]_  = \new_[42902]_  & \new_[42899]_ ;
  assign \new_[42904]_  = \new_[42903]_  & \new_[42896]_ ;
  assign \new_[42908]_  = A167 & A168;
  assign \new_[42909]_  = ~A170 & \new_[42908]_ ;
  assign \new_[42913]_  = ~A200 & ~A199;
  assign \new_[42914]_  = ~A166 & \new_[42913]_ ;
  assign \new_[42915]_  = \new_[42914]_  & \new_[42909]_ ;
  assign \new_[42919]_  = ~A269 & ~A268;
  assign \new_[42920]_  = A267 & \new_[42919]_ ;
  assign \new_[42923]_  = A299 & ~A298;
  assign \new_[42926]_  = A302 & A300;
  assign \new_[42927]_  = \new_[42926]_  & \new_[42923]_ ;
  assign \new_[42928]_  = \new_[42927]_  & \new_[42920]_ ;
  assign \new_[42932]_  = A167 & A168;
  assign \new_[42933]_  = ~A170 & \new_[42932]_ ;
  assign \new_[42937]_  = ~A200 & ~A199;
  assign \new_[42938]_  = ~A166 & \new_[42937]_ ;
  assign \new_[42939]_  = \new_[42938]_  & \new_[42933]_ ;
  assign \new_[42943]_  = A298 & A268;
  assign \new_[42944]_  = ~A267 & \new_[42943]_ ;
  assign \new_[42947]_  = ~A300 & ~A299;
  assign \new_[42950]_  = ~A302 & ~A301;
  assign \new_[42951]_  = \new_[42950]_  & \new_[42947]_ ;
  assign \new_[42952]_  = \new_[42951]_  & \new_[42944]_ ;
  assign \new_[42956]_  = A167 & A168;
  assign \new_[42957]_  = ~A170 & \new_[42956]_ ;
  assign \new_[42961]_  = ~A200 & ~A199;
  assign \new_[42962]_  = ~A166 & \new_[42961]_ ;
  assign \new_[42963]_  = \new_[42962]_  & \new_[42957]_ ;
  assign \new_[42967]_  = ~A298 & A268;
  assign \new_[42968]_  = ~A267 & \new_[42967]_ ;
  assign \new_[42971]_  = ~A300 & A299;
  assign \new_[42974]_  = ~A302 & ~A301;
  assign \new_[42975]_  = \new_[42974]_  & \new_[42971]_ ;
  assign \new_[42976]_  = \new_[42975]_  & \new_[42968]_ ;
  assign \new_[42980]_  = A167 & A168;
  assign \new_[42981]_  = ~A170 & \new_[42980]_ ;
  assign \new_[42985]_  = ~A200 & ~A199;
  assign \new_[42986]_  = ~A166 & \new_[42985]_ ;
  assign \new_[42987]_  = \new_[42986]_  & \new_[42981]_ ;
  assign \new_[42991]_  = A298 & A269;
  assign \new_[42992]_  = ~A267 & \new_[42991]_ ;
  assign \new_[42995]_  = ~A300 & ~A299;
  assign \new_[42998]_  = ~A302 & ~A301;
  assign \new_[42999]_  = \new_[42998]_  & \new_[42995]_ ;
  assign \new_[43000]_  = \new_[42999]_  & \new_[42992]_ ;
  assign \new_[43004]_  = A167 & A168;
  assign \new_[43005]_  = ~A170 & \new_[43004]_ ;
  assign \new_[43009]_  = ~A200 & ~A199;
  assign \new_[43010]_  = ~A166 & \new_[43009]_ ;
  assign \new_[43011]_  = \new_[43010]_  & \new_[43005]_ ;
  assign \new_[43015]_  = ~A298 & A269;
  assign \new_[43016]_  = ~A267 & \new_[43015]_ ;
  assign \new_[43019]_  = ~A300 & A299;
  assign \new_[43022]_  = ~A302 & ~A301;
  assign \new_[43023]_  = \new_[43022]_  & \new_[43019]_ ;
  assign \new_[43024]_  = \new_[43023]_  & \new_[43016]_ ;
  assign \new_[43028]_  = A167 & A168;
  assign \new_[43029]_  = ~A170 & \new_[43028]_ ;
  assign \new_[43033]_  = ~A200 & ~A199;
  assign \new_[43034]_  = ~A166 & \new_[43033]_ ;
  assign \new_[43035]_  = \new_[43034]_  & \new_[43029]_ ;
  assign \new_[43039]_  = A298 & A266;
  assign \new_[43040]_  = A265 & \new_[43039]_ ;
  assign \new_[43043]_  = ~A300 & ~A299;
  assign \new_[43046]_  = ~A302 & ~A301;
  assign \new_[43047]_  = \new_[43046]_  & \new_[43043]_ ;
  assign \new_[43048]_  = \new_[43047]_  & \new_[43040]_ ;
  assign \new_[43052]_  = A167 & A168;
  assign \new_[43053]_  = ~A170 & \new_[43052]_ ;
  assign \new_[43057]_  = ~A200 & ~A199;
  assign \new_[43058]_  = ~A166 & \new_[43057]_ ;
  assign \new_[43059]_  = \new_[43058]_  & \new_[43053]_ ;
  assign \new_[43063]_  = ~A298 & A266;
  assign \new_[43064]_  = A265 & \new_[43063]_ ;
  assign \new_[43067]_  = ~A300 & A299;
  assign \new_[43070]_  = ~A302 & ~A301;
  assign \new_[43071]_  = \new_[43070]_  & \new_[43067]_ ;
  assign \new_[43072]_  = \new_[43071]_  & \new_[43064]_ ;
  assign \new_[43076]_  = A167 & A168;
  assign \new_[43077]_  = ~A170 & \new_[43076]_ ;
  assign \new_[43081]_  = ~A200 & ~A199;
  assign \new_[43082]_  = ~A166 & \new_[43081]_ ;
  assign \new_[43083]_  = \new_[43082]_  & \new_[43077]_ ;
  assign \new_[43087]_  = A298 & ~A266;
  assign \new_[43088]_  = ~A265 & \new_[43087]_ ;
  assign \new_[43091]_  = ~A300 & ~A299;
  assign \new_[43094]_  = ~A302 & ~A301;
  assign \new_[43095]_  = \new_[43094]_  & \new_[43091]_ ;
  assign \new_[43096]_  = \new_[43095]_  & \new_[43088]_ ;
  assign \new_[43100]_  = A167 & A168;
  assign \new_[43101]_  = ~A170 & \new_[43100]_ ;
  assign \new_[43105]_  = ~A200 & ~A199;
  assign \new_[43106]_  = ~A166 & \new_[43105]_ ;
  assign \new_[43107]_  = \new_[43106]_  & \new_[43101]_ ;
  assign \new_[43111]_  = ~A298 & ~A266;
  assign \new_[43112]_  = ~A265 & \new_[43111]_ ;
  assign \new_[43115]_  = ~A300 & A299;
  assign \new_[43118]_  = ~A302 & ~A301;
  assign \new_[43119]_  = \new_[43118]_  & \new_[43115]_ ;
  assign \new_[43120]_  = \new_[43119]_  & \new_[43112]_ ;
  assign \new_[43124]_  = ~A167 & A168;
  assign \new_[43125]_  = ~A170 & \new_[43124]_ ;
  assign \new_[43129]_  = ~A202 & A201;
  assign \new_[43130]_  = A166 & \new_[43129]_ ;
  assign \new_[43131]_  = \new_[43130]_  & \new_[43125]_ ;
  assign \new_[43135]_  = A268 & ~A267;
  assign \new_[43136]_  = ~A203 & \new_[43135]_ ;
  assign \new_[43139]_  = ~A299 & A298;
  assign \new_[43142]_  = A301 & A300;
  assign \new_[43143]_  = \new_[43142]_  & \new_[43139]_ ;
  assign \new_[43144]_  = \new_[43143]_  & \new_[43136]_ ;
  assign \new_[43148]_  = ~A167 & A168;
  assign \new_[43149]_  = ~A170 & \new_[43148]_ ;
  assign \new_[43153]_  = ~A202 & A201;
  assign \new_[43154]_  = A166 & \new_[43153]_ ;
  assign \new_[43155]_  = \new_[43154]_  & \new_[43149]_ ;
  assign \new_[43159]_  = A268 & ~A267;
  assign \new_[43160]_  = ~A203 & \new_[43159]_ ;
  assign \new_[43163]_  = ~A299 & A298;
  assign \new_[43166]_  = A302 & A300;
  assign \new_[43167]_  = \new_[43166]_  & \new_[43163]_ ;
  assign \new_[43168]_  = \new_[43167]_  & \new_[43160]_ ;
  assign \new_[43172]_  = ~A167 & A168;
  assign \new_[43173]_  = ~A170 & \new_[43172]_ ;
  assign \new_[43177]_  = ~A202 & A201;
  assign \new_[43178]_  = A166 & \new_[43177]_ ;
  assign \new_[43179]_  = \new_[43178]_  & \new_[43173]_ ;
  assign \new_[43183]_  = A268 & ~A267;
  assign \new_[43184]_  = ~A203 & \new_[43183]_ ;
  assign \new_[43187]_  = A299 & ~A298;
  assign \new_[43190]_  = A301 & A300;
  assign \new_[43191]_  = \new_[43190]_  & \new_[43187]_ ;
  assign \new_[43192]_  = \new_[43191]_  & \new_[43184]_ ;
  assign \new_[43196]_  = ~A167 & A168;
  assign \new_[43197]_  = ~A170 & \new_[43196]_ ;
  assign \new_[43201]_  = ~A202 & A201;
  assign \new_[43202]_  = A166 & \new_[43201]_ ;
  assign \new_[43203]_  = \new_[43202]_  & \new_[43197]_ ;
  assign \new_[43207]_  = A268 & ~A267;
  assign \new_[43208]_  = ~A203 & \new_[43207]_ ;
  assign \new_[43211]_  = A299 & ~A298;
  assign \new_[43214]_  = A302 & A300;
  assign \new_[43215]_  = \new_[43214]_  & \new_[43211]_ ;
  assign \new_[43216]_  = \new_[43215]_  & \new_[43208]_ ;
  assign \new_[43220]_  = ~A167 & A168;
  assign \new_[43221]_  = ~A170 & \new_[43220]_ ;
  assign \new_[43225]_  = ~A202 & A201;
  assign \new_[43226]_  = A166 & \new_[43225]_ ;
  assign \new_[43227]_  = \new_[43226]_  & \new_[43221]_ ;
  assign \new_[43231]_  = A269 & ~A267;
  assign \new_[43232]_  = ~A203 & \new_[43231]_ ;
  assign \new_[43235]_  = ~A299 & A298;
  assign \new_[43238]_  = A301 & A300;
  assign \new_[43239]_  = \new_[43238]_  & \new_[43235]_ ;
  assign \new_[43240]_  = \new_[43239]_  & \new_[43232]_ ;
  assign \new_[43244]_  = ~A167 & A168;
  assign \new_[43245]_  = ~A170 & \new_[43244]_ ;
  assign \new_[43249]_  = ~A202 & A201;
  assign \new_[43250]_  = A166 & \new_[43249]_ ;
  assign \new_[43251]_  = \new_[43250]_  & \new_[43245]_ ;
  assign \new_[43255]_  = A269 & ~A267;
  assign \new_[43256]_  = ~A203 & \new_[43255]_ ;
  assign \new_[43259]_  = ~A299 & A298;
  assign \new_[43262]_  = A302 & A300;
  assign \new_[43263]_  = \new_[43262]_  & \new_[43259]_ ;
  assign \new_[43264]_  = \new_[43263]_  & \new_[43256]_ ;
  assign \new_[43268]_  = ~A167 & A168;
  assign \new_[43269]_  = ~A170 & \new_[43268]_ ;
  assign \new_[43273]_  = ~A202 & A201;
  assign \new_[43274]_  = A166 & \new_[43273]_ ;
  assign \new_[43275]_  = \new_[43274]_  & \new_[43269]_ ;
  assign \new_[43279]_  = A269 & ~A267;
  assign \new_[43280]_  = ~A203 & \new_[43279]_ ;
  assign \new_[43283]_  = A299 & ~A298;
  assign \new_[43286]_  = A301 & A300;
  assign \new_[43287]_  = \new_[43286]_  & \new_[43283]_ ;
  assign \new_[43288]_  = \new_[43287]_  & \new_[43280]_ ;
  assign \new_[43292]_  = ~A167 & A168;
  assign \new_[43293]_  = ~A170 & \new_[43292]_ ;
  assign \new_[43297]_  = ~A202 & A201;
  assign \new_[43298]_  = A166 & \new_[43297]_ ;
  assign \new_[43299]_  = \new_[43298]_  & \new_[43293]_ ;
  assign \new_[43303]_  = A269 & ~A267;
  assign \new_[43304]_  = ~A203 & \new_[43303]_ ;
  assign \new_[43307]_  = A299 & ~A298;
  assign \new_[43310]_  = A302 & A300;
  assign \new_[43311]_  = \new_[43310]_  & \new_[43307]_ ;
  assign \new_[43312]_  = \new_[43311]_  & \new_[43304]_ ;
  assign \new_[43316]_  = ~A167 & A168;
  assign \new_[43317]_  = ~A170 & \new_[43316]_ ;
  assign \new_[43321]_  = ~A202 & A201;
  assign \new_[43322]_  = A166 & \new_[43321]_ ;
  assign \new_[43323]_  = \new_[43322]_  & \new_[43317]_ ;
  assign \new_[43327]_  = A266 & A265;
  assign \new_[43328]_  = ~A203 & \new_[43327]_ ;
  assign \new_[43331]_  = ~A299 & A298;
  assign \new_[43334]_  = A301 & A300;
  assign \new_[43335]_  = \new_[43334]_  & \new_[43331]_ ;
  assign \new_[43336]_  = \new_[43335]_  & \new_[43328]_ ;
  assign \new_[43340]_  = ~A167 & A168;
  assign \new_[43341]_  = ~A170 & \new_[43340]_ ;
  assign \new_[43345]_  = ~A202 & A201;
  assign \new_[43346]_  = A166 & \new_[43345]_ ;
  assign \new_[43347]_  = \new_[43346]_  & \new_[43341]_ ;
  assign \new_[43351]_  = A266 & A265;
  assign \new_[43352]_  = ~A203 & \new_[43351]_ ;
  assign \new_[43355]_  = ~A299 & A298;
  assign \new_[43358]_  = A302 & A300;
  assign \new_[43359]_  = \new_[43358]_  & \new_[43355]_ ;
  assign \new_[43360]_  = \new_[43359]_  & \new_[43352]_ ;
  assign \new_[43364]_  = ~A167 & A168;
  assign \new_[43365]_  = ~A170 & \new_[43364]_ ;
  assign \new_[43369]_  = ~A202 & A201;
  assign \new_[43370]_  = A166 & \new_[43369]_ ;
  assign \new_[43371]_  = \new_[43370]_  & \new_[43365]_ ;
  assign \new_[43375]_  = A266 & A265;
  assign \new_[43376]_  = ~A203 & \new_[43375]_ ;
  assign \new_[43379]_  = A299 & ~A298;
  assign \new_[43382]_  = A301 & A300;
  assign \new_[43383]_  = \new_[43382]_  & \new_[43379]_ ;
  assign \new_[43384]_  = \new_[43383]_  & \new_[43376]_ ;
  assign \new_[43388]_  = ~A167 & A168;
  assign \new_[43389]_  = ~A170 & \new_[43388]_ ;
  assign \new_[43393]_  = ~A202 & A201;
  assign \new_[43394]_  = A166 & \new_[43393]_ ;
  assign \new_[43395]_  = \new_[43394]_  & \new_[43389]_ ;
  assign \new_[43399]_  = A266 & A265;
  assign \new_[43400]_  = ~A203 & \new_[43399]_ ;
  assign \new_[43403]_  = A299 & ~A298;
  assign \new_[43406]_  = A302 & A300;
  assign \new_[43407]_  = \new_[43406]_  & \new_[43403]_ ;
  assign \new_[43408]_  = \new_[43407]_  & \new_[43400]_ ;
  assign \new_[43412]_  = ~A167 & A168;
  assign \new_[43413]_  = ~A170 & \new_[43412]_ ;
  assign \new_[43417]_  = ~A202 & A201;
  assign \new_[43418]_  = A166 & \new_[43417]_ ;
  assign \new_[43419]_  = \new_[43418]_  & \new_[43413]_ ;
  assign \new_[43423]_  = ~A266 & ~A265;
  assign \new_[43424]_  = ~A203 & \new_[43423]_ ;
  assign \new_[43427]_  = ~A299 & A298;
  assign \new_[43430]_  = A301 & A300;
  assign \new_[43431]_  = \new_[43430]_  & \new_[43427]_ ;
  assign \new_[43432]_  = \new_[43431]_  & \new_[43424]_ ;
  assign \new_[43436]_  = ~A167 & A168;
  assign \new_[43437]_  = ~A170 & \new_[43436]_ ;
  assign \new_[43441]_  = ~A202 & A201;
  assign \new_[43442]_  = A166 & \new_[43441]_ ;
  assign \new_[43443]_  = \new_[43442]_  & \new_[43437]_ ;
  assign \new_[43447]_  = ~A266 & ~A265;
  assign \new_[43448]_  = ~A203 & \new_[43447]_ ;
  assign \new_[43451]_  = ~A299 & A298;
  assign \new_[43454]_  = A302 & A300;
  assign \new_[43455]_  = \new_[43454]_  & \new_[43451]_ ;
  assign \new_[43456]_  = \new_[43455]_  & \new_[43448]_ ;
  assign \new_[43460]_  = ~A167 & A168;
  assign \new_[43461]_  = ~A170 & \new_[43460]_ ;
  assign \new_[43465]_  = ~A202 & A201;
  assign \new_[43466]_  = A166 & \new_[43465]_ ;
  assign \new_[43467]_  = \new_[43466]_  & \new_[43461]_ ;
  assign \new_[43471]_  = ~A266 & ~A265;
  assign \new_[43472]_  = ~A203 & \new_[43471]_ ;
  assign \new_[43475]_  = A299 & ~A298;
  assign \new_[43478]_  = A301 & A300;
  assign \new_[43479]_  = \new_[43478]_  & \new_[43475]_ ;
  assign \new_[43480]_  = \new_[43479]_  & \new_[43472]_ ;
  assign \new_[43484]_  = ~A167 & A168;
  assign \new_[43485]_  = ~A170 & \new_[43484]_ ;
  assign \new_[43489]_  = ~A202 & A201;
  assign \new_[43490]_  = A166 & \new_[43489]_ ;
  assign \new_[43491]_  = \new_[43490]_  & \new_[43485]_ ;
  assign \new_[43495]_  = ~A266 & ~A265;
  assign \new_[43496]_  = ~A203 & \new_[43495]_ ;
  assign \new_[43499]_  = A299 & ~A298;
  assign \new_[43502]_  = A302 & A300;
  assign \new_[43503]_  = \new_[43502]_  & \new_[43499]_ ;
  assign \new_[43504]_  = \new_[43503]_  & \new_[43496]_ ;
  assign \new_[43508]_  = ~A167 & A168;
  assign \new_[43509]_  = ~A170 & \new_[43508]_ ;
  assign \new_[43513]_  = A202 & ~A201;
  assign \new_[43514]_  = A166 & \new_[43513]_ ;
  assign \new_[43515]_  = \new_[43514]_  & \new_[43509]_ ;
  assign \new_[43519]_  = ~A269 & ~A268;
  assign \new_[43520]_  = A267 & \new_[43519]_ ;
  assign \new_[43523]_  = ~A299 & A298;
  assign \new_[43526]_  = A301 & A300;
  assign \new_[43527]_  = \new_[43526]_  & \new_[43523]_ ;
  assign \new_[43528]_  = \new_[43527]_  & \new_[43520]_ ;
  assign \new_[43532]_  = ~A167 & A168;
  assign \new_[43533]_  = ~A170 & \new_[43532]_ ;
  assign \new_[43537]_  = A202 & ~A201;
  assign \new_[43538]_  = A166 & \new_[43537]_ ;
  assign \new_[43539]_  = \new_[43538]_  & \new_[43533]_ ;
  assign \new_[43543]_  = ~A269 & ~A268;
  assign \new_[43544]_  = A267 & \new_[43543]_ ;
  assign \new_[43547]_  = ~A299 & A298;
  assign \new_[43550]_  = A302 & A300;
  assign \new_[43551]_  = \new_[43550]_  & \new_[43547]_ ;
  assign \new_[43552]_  = \new_[43551]_  & \new_[43544]_ ;
  assign \new_[43556]_  = ~A167 & A168;
  assign \new_[43557]_  = ~A170 & \new_[43556]_ ;
  assign \new_[43561]_  = A202 & ~A201;
  assign \new_[43562]_  = A166 & \new_[43561]_ ;
  assign \new_[43563]_  = \new_[43562]_  & \new_[43557]_ ;
  assign \new_[43567]_  = ~A269 & ~A268;
  assign \new_[43568]_  = A267 & \new_[43567]_ ;
  assign \new_[43571]_  = A299 & ~A298;
  assign \new_[43574]_  = A301 & A300;
  assign \new_[43575]_  = \new_[43574]_  & \new_[43571]_ ;
  assign \new_[43576]_  = \new_[43575]_  & \new_[43568]_ ;
  assign \new_[43580]_  = ~A167 & A168;
  assign \new_[43581]_  = ~A170 & \new_[43580]_ ;
  assign \new_[43585]_  = A202 & ~A201;
  assign \new_[43586]_  = A166 & \new_[43585]_ ;
  assign \new_[43587]_  = \new_[43586]_  & \new_[43581]_ ;
  assign \new_[43591]_  = ~A269 & ~A268;
  assign \new_[43592]_  = A267 & \new_[43591]_ ;
  assign \new_[43595]_  = A299 & ~A298;
  assign \new_[43598]_  = A302 & A300;
  assign \new_[43599]_  = \new_[43598]_  & \new_[43595]_ ;
  assign \new_[43600]_  = \new_[43599]_  & \new_[43592]_ ;
  assign \new_[43604]_  = ~A167 & A168;
  assign \new_[43605]_  = ~A170 & \new_[43604]_ ;
  assign \new_[43609]_  = A202 & ~A201;
  assign \new_[43610]_  = A166 & \new_[43609]_ ;
  assign \new_[43611]_  = \new_[43610]_  & \new_[43605]_ ;
  assign \new_[43615]_  = A298 & A268;
  assign \new_[43616]_  = ~A267 & \new_[43615]_ ;
  assign \new_[43619]_  = ~A300 & ~A299;
  assign \new_[43622]_  = ~A302 & ~A301;
  assign \new_[43623]_  = \new_[43622]_  & \new_[43619]_ ;
  assign \new_[43624]_  = \new_[43623]_  & \new_[43616]_ ;
  assign \new_[43628]_  = ~A167 & A168;
  assign \new_[43629]_  = ~A170 & \new_[43628]_ ;
  assign \new_[43633]_  = A202 & ~A201;
  assign \new_[43634]_  = A166 & \new_[43633]_ ;
  assign \new_[43635]_  = \new_[43634]_  & \new_[43629]_ ;
  assign \new_[43639]_  = ~A298 & A268;
  assign \new_[43640]_  = ~A267 & \new_[43639]_ ;
  assign \new_[43643]_  = ~A300 & A299;
  assign \new_[43646]_  = ~A302 & ~A301;
  assign \new_[43647]_  = \new_[43646]_  & \new_[43643]_ ;
  assign \new_[43648]_  = \new_[43647]_  & \new_[43640]_ ;
  assign \new_[43652]_  = ~A167 & A168;
  assign \new_[43653]_  = ~A170 & \new_[43652]_ ;
  assign \new_[43657]_  = A202 & ~A201;
  assign \new_[43658]_  = A166 & \new_[43657]_ ;
  assign \new_[43659]_  = \new_[43658]_  & \new_[43653]_ ;
  assign \new_[43663]_  = A298 & A269;
  assign \new_[43664]_  = ~A267 & \new_[43663]_ ;
  assign \new_[43667]_  = ~A300 & ~A299;
  assign \new_[43670]_  = ~A302 & ~A301;
  assign \new_[43671]_  = \new_[43670]_  & \new_[43667]_ ;
  assign \new_[43672]_  = \new_[43671]_  & \new_[43664]_ ;
  assign \new_[43676]_  = ~A167 & A168;
  assign \new_[43677]_  = ~A170 & \new_[43676]_ ;
  assign \new_[43681]_  = A202 & ~A201;
  assign \new_[43682]_  = A166 & \new_[43681]_ ;
  assign \new_[43683]_  = \new_[43682]_  & \new_[43677]_ ;
  assign \new_[43687]_  = ~A298 & A269;
  assign \new_[43688]_  = ~A267 & \new_[43687]_ ;
  assign \new_[43691]_  = ~A300 & A299;
  assign \new_[43694]_  = ~A302 & ~A301;
  assign \new_[43695]_  = \new_[43694]_  & \new_[43691]_ ;
  assign \new_[43696]_  = \new_[43695]_  & \new_[43688]_ ;
  assign \new_[43700]_  = ~A167 & A168;
  assign \new_[43701]_  = ~A170 & \new_[43700]_ ;
  assign \new_[43705]_  = A202 & ~A201;
  assign \new_[43706]_  = A166 & \new_[43705]_ ;
  assign \new_[43707]_  = \new_[43706]_  & \new_[43701]_ ;
  assign \new_[43711]_  = A298 & A266;
  assign \new_[43712]_  = A265 & \new_[43711]_ ;
  assign \new_[43715]_  = ~A300 & ~A299;
  assign \new_[43718]_  = ~A302 & ~A301;
  assign \new_[43719]_  = \new_[43718]_  & \new_[43715]_ ;
  assign \new_[43720]_  = \new_[43719]_  & \new_[43712]_ ;
  assign \new_[43724]_  = ~A167 & A168;
  assign \new_[43725]_  = ~A170 & \new_[43724]_ ;
  assign \new_[43729]_  = A202 & ~A201;
  assign \new_[43730]_  = A166 & \new_[43729]_ ;
  assign \new_[43731]_  = \new_[43730]_  & \new_[43725]_ ;
  assign \new_[43735]_  = ~A298 & A266;
  assign \new_[43736]_  = A265 & \new_[43735]_ ;
  assign \new_[43739]_  = ~A300 & A299;
  assign \new_[43742]_  = ~A302 & ~A301;
  assign \new_[43743]_  = \new_[43742]_  & \new_[43739]_ ;
  assign \new_[43744]_  = \new_[43743]_  & \new_[43736]_ ;
  assign \new_[43748]_  = ~A167 & A168;
  assign \new_[43749]_  = ~A170 & \new_[43748]_ ;
  assign \new_[43753]_  = A202 & ~A201;
  assign \new_[43754]_  = A166 & \new_[43753]_ ;
  assign \new_[43755]_  = \new_[43754]_  & \new_[43749]_ ;
  assign \new_[43759]_  = A298 & ~A266;
  assign \new_[43760]_  = ~A265 & \new_[43759]_ ;
  assign \new_[43763]_  = ~A300 & ~A299;
  assign \new_[43766]_  = ~A302 & ~A301;
  assign \new_[43767]_  = \new_[43766]_  & \new_[43763]_ ;
  assign \new_[43768]_  = \new_[43767]_  & \new_[43760]_ ;
  assign \new_[43772]_  = ~A167 & A168;
  assign \new_[43773]_  = ~A170 & \new_[43772]_ ;
  assign \new_[43777]_  = A202 & ~A201;
  assign \new_[43778]_  = A166 & \new_[43777]_ ;
  assign \new_[43779]_  = \new_[43778]_  & \new_[43773]_ ;
  assign \new_[43783]_  = ~A298 & ~A266;
  assign \new_[43784]_  = ~A265 & \new_[43783]_ ;
  assign \new_[43787]_  = ~A300 & A299;
  assign \new_[43790]_  = ~A302 & ~A301;
  assign \new_[43791]_  = \new_[43790]_  & \new_[43787]_ ;
  assign \new_[43792]_  = \new_[43791]_  & \new_[43784]_ ;
  assign \new_[43796]_  = ~A167 & A168;
  assign \new_[43797]_  = ~A170 & \new_[43796]_ ;
  assign \new_[43801]_  = A203 & ~A201;
  assign \new_[43802]_  = A166 & \new_[43801]_ ;
  assign \new_[43803]_  = \new_[43802]_  & \new_[43797]_ ;
  assign \new_[43807]_  = ~A269 & ~A268;
  assign \new_[43808]_  = A267 & \new_[43807]_ ;
  assign \new_[43811]_  = ~A299 & A298;
  assign \new_[43814]_  = A301 & A300;
  assign \new_[43815]_  = \new_[43814]_  & \new_[43811]_ ;
  assign \new_[43816]_  = \new_[43815]_  & \new_[43808]_ ;
  assign \new_[43820]_  = ~A167 & A168;
  assign \new_[43821]_  = ~A170 & \new_[43820]_ ;
  assign \new_[43825]_  = A203 & ~A201;
  assign \new_[43826]_  = A166 & \new_[43825]_ ;
  assign \new_[43827]_  = \new_[43826]_  & \new_[43821]_ ;
  assign \new_[43831]_  = ~A269 & ~A268;
  assign \new_[43832]_  = A267 & \new_[43831]_ ;
  assign \new_[43835]_  = ~A299 & A298;
  assign \new_[43838]_  = A302 & A300;
  assign \new_[43839]_  = \new_[43838]_  & \new_[43835]_ ;
  assign \new_[43840]_  = \new_[43839]_  & \new_[43832]_ ;
  assign \new_[43844]_  = ~A167 & A168;
  assign \new_[43845]_  = ~A170 & \new_[43844]_ ;
  assign \new_[43849]_  = A203 & ~A201;
  assign \new_[43850]_  = A166 & \new_[43849]_ ;
  assign \new_[43851]_  = \new_[43850]_  & \new_[43845]_ ;
  assign \new_[43855]_  = ~A269 & ~A268;
  assign \new_[43856]_  = A267 & \new_[43855]_ ;
  assign \new_[43859]_  = A299 & ~A298;
  assign \new_[43862]_  = A301 & A300;
  assign \new_[43863]_  = \new_[43862]_  & \new_[43859]_ ;
  assign \new_[43864]_  = \new_[43863]_  & \new_[43856]_ ;
  assign \new_[43868]_  = ~A167 & A168;
  assign \new_[43869]_  = ~A170 & \new_[43868]_ ;
  assign \new_[43873]_  = A203 & ~A201;
  assign \new_[43874]_  = A166 & \new_[43873]_ ;
  assign \new_[43875]_  = \new_[43874]_  & \new_[43869]_ ;
  assign \new_[43879]_  = ~A269 & ~A268;
  assign \new_[43880]_  = A267 & \new_[43879]_ ;
  assign \new_[43883]_  = A299 & ~A298;
  assign \new_[43886]_  = A302 & A300;
  assign \new_[43887]_  = \new_[43886]_  & \new_[43883]_ ;
  assign \new_[43888]_  = \new_[43887]_  & \new_[43880]_ ;
  assign \new_[43892]_  = ~A167 & A168;
  assign \new_[43893]_  = ~A170 & \new_[43892]_ ;
  assign \new_[43897]_  = A203 & ~A201;
  assign \new_[43898]_  = A166 & \new_[43897]_ ;
  assign \new_[43899]_  = \new_[43898]_  & \new_[43893]_ ;
  assign \new_[43903]_  = A298 & A268;
  assign \new_[43904]_  = ~A267 & \new_[43903]_ ;
  assign \new_[43907]_  = ~A300 & ~A299;
  assign \new_[43910]_  = ~A302 & ~A301;
  assign \new_[43911]_  = \new_[43910]_  & \new_[43907]_ ;
  assign \new_[43912]_  = \new_[43911]_  & \new_[43904]_ ;
  assign \new_[43916]_  = ~A167 & A168;
  assign \new_[43917]_  = ~A170 & \new_[43916]_ ;
  assign \new_[43921]_  = A203 & ~A201;
  assign \new_[43922]_  = A166 & \new_[43921]_ ;
  assign \new_[43923]_  = \new_[43922]_  & \new_[43917]_ ;
  assign \new_[43927]_  = ~A298 & A268;
  assign \new_[43928]_  = ~A267 & \new_[43927]_ ;
  assign \new_[43931]_  = ~A300 & A299;
  assign \new_[43934]_  = ~A302 & ~A301;
  assign \new_[43935]_  = \new_[43934]_  & \new_[43931]_ ;
  assign \new_[43936]_  = \new_[43935]_  & \new_[43928]_ ;
  assign \new_[43940]_  = ~A167 & A168;
  assign \new_[43941]_  = ~A170 & \new_[43940]_ ;
  assign \new_[43945]_  = A203 & ~A201;
  assign \new_[43946]_  = A166 & \new_[43945]_ ;
  assign \new_[43947]_  = \new_[43946]_  & \new_[43941]_ ;
  assign \new_[43951]_  = A298 & A269;
  assign \new_[43952]_  = ~A267 & \new_[43951]_ ;
  assign \new_[43955]_  = ~A300 & ~A299;
  assign \new_[43958]_  = ~A302 & ~A301;
  assign \new_[43959]_  = \new_[43958]_  & \new_[43955]_ ;
  assign \new_[43960]_  = \new_[43959]_  & \new_[43952]_ ;
  assign \new_[43964]_  = ~A167 & A168;
  assign \new_[43965]_  = ~A170 & \new_[43964]_ ;
  assign \new_[43969]_  = A203 & ~A201;
  assign \new_[43970]_  = A166 & \new_[43969]_ ;
  assign \new_[43971]_  = \new_[43970]_  & \new_[43965]_ ;
  assign \new_[43975]_  = ~A298 & A269;
  assign \new_[43976]_  = ~A267 & \new_[43975]_ ;
  assign \new_[43979]_  = ~A300 & A299;
  assign \new_[43982]_  = ~A302 & ~A301;
  assign \new_[43983]_  = \new_[43982]_  & \new_[43979]_ ;
  assign \new_[43984]_  = \new_[43983]_  & \new_[43976]_ ;
  assign \new_[43988]_  = ~A167 & A168;
  assign \new_[43989]_  = ~A170 & \new_[43988]_ ;
  assign \new_[43993]_  = A203 & ~A201;
  assign \new_[43994]_  = A166 & \new_[43993]_ ;
  assign \new_[43995]_  = \new_[43994]_  & \new_[43989]_ ;
  assign \new_[43999]_  = A298 & A266;
  assign \new_[44000]_  = A265 & \new_[43999]_ ;
  assign \new_[44003]_  = ~A300 & ~A299;
  assign \new_[44006]_  = ~A302 & ~A301;
  assign \new_[44007]_  = \new_[44006]_  & \new_[44003]_ ;
  assign \new_[44008]_  = \new_[44007]_  & \new_[44000]_ ;
  assign \new_[44012]_  = ~A167 & A168;
  assign \new_[44013]_  = ~A170 & \new_[44012]_ ;
  assign \new_[44017]_  = A203 & ~A201;
  assign \new_[44018]_  = A166 & \new_[44017]_ ;
  assign \new_[44019]_  = \new_[44018]_  & \new_[44013]_ ;
  assign \new_[44023]_  = ~A298 & A266;
  assign \new_[44024]_  = A265 & \new_[44023]_ ;
  assign \new_[44027]_  = ~A300 & A299;
  assign \new_[44030]_  = ~A302 & ~A301;
  assign \new_[44031]_  = \new_[44030]_  & \new_[44027]_ ;
  assign \new_[44032]_  = \new_[44031]_  & \new_[44024]_ ;
  assign \new_[44036]_  = ~A167 & A168;
  assign \new_[44037]_  = ~A170 & \new_[44036]_ ;
  assign \new_[44041]_  = A203 & ~A201;
  assign \new_[44042]_  = A166 & \new_[44041]_ ;
  assign \new_[44043]_  = \new_[44042]_  & \new_[44037]_ ;
  assign \new_[44047]_  = A298 & ~A266;
  assign \new_[44048]_  = ~A265 & \new_[44047]_ ;
  assign \new_[44051]_  = ~A300 & ~A299;
  assign \new_[44054]_  = ~A302 & ~A301;
  assign \new_[44055]_  = \new_[44054]_  & \new_[44051]_ ;
  assign \new_[44056]_  = \new_[44055]_  & \new_[44048]_ ;
  assign \new_[44060]_  = ~A167 & A168;
  assign \new_[44061]_  = ~A170 & \new_[44060]_ ;
  assign \new_[44065]_  = A203 & ~A201;
  assign \new_[44066]_  = A166 & \new_[44065]_ ;
  assign \new_[44067]_  = \new_[44066]_  & \new_[44061]_ ;
  assign \new_[44071]_  = ~A298 & ~A266;
  assign \new_[44072]_  = ~A265 & \new_[44071]_ ;
  assign \new_[44075]_  = ~A300 & A299;
  assign \new_[44078]_  = ~A302 & ~A301;
  assign \new_[44079]_  = \new_[44078]_  & \new_[44075]_ ;
  assign \new_[44080]_  = \new_[44079]_  & \new_[44072]_ ;
  assign \new_[44084]_  = ~A167 & A168;
  assign \new_[44085]_  = ~A170 & \new_[44084]_ ;
  assign \new_[44089]_  = A200 & A199;
  assign \new_[44090]_  = A166 & \new_[44089]_ ;
  assign \new_[44091]_  = \new_[44090]_  & \new_[44085]_ ;
  assign \new_[44095]_  = ~A269 & ~A268;
  assign \new_[44096]_  = A267 & \new_[44095]_ ;
  assign \new_[44099]_  = ~A299 & A298;
  assign \new_[44102]_  = A301 & A300;
  assign \new_[44103]_  = \new_[44102]_  & \new_[44099]_ ;
  assign \new_[44104]_  = \new_[44103]_  & \new_[44096]_ ;
  assign \new_[44108]_  = ~A167 & A168;
  assign \new_[44109]_  = ~A170 & \new_[44108]_ ;
  assign \new_[44113]_  = A200 & A199;
  assign \new_[44114]_  = A166 & \new_[44113]_ ;
  assign \new_[44115]_  = \new_[44114]_  & \new_[44109]_ ;
  assign \new_[44119]_  = ~A269 & ~A268;
  assign \new_[44120]_  = A267 & \new_[44119]_ ;
  assign \new_[44123]_  = ~A299 & A298;
  assign \new_[44126]_  = A302 & A300;
  assign \new_[44127]_  = \new_[44126]_  & \new_[44123]_ ;
  assign \new_[44128]_  = \new_[44127]_  & \new_[44120]_ ;
  assign \new_[44132]_  = ~A167 & A168;
  assign \new_[44133]_  = ~A170 & \new_[44132]_ ;
  assign \new_[44137]_  = A200 & A199;
  assign \new_[44138]_  = A166 & \new_[44137]_ ;
  assign \new_[44139]_  = \new_[44138]_  & \new_[44133]_ ;
  assign \new_[44143]_  = ~A269 & ~A268;
  assign \new_[44144]_  = A267 & \new_[44143]_ ;
  assign \new_[44147]_  = A299 & ~A298;
  assign \new_[44150]_  = A301 & A300;
  assign \new_[44151]_  = \new_[44150]_  & \new_[44147]_ ;
  assign \new_[44152]_  = \new_[44151]_  & \new_[44144]_ ;
  assign \new_[44156]_  = ~A167 & A168;
  assign \new_[44157]_  = ~A170 & \new_[44156]_ ;
  assign \new_[44161]_  = A200 & A199;
  assign \new_[44162]_  = A166 & \new_[44161]_ ;
  assign \new_[44163]_  = \new_[44162]_  & \new_[44157]_ ;
  assign \new_[44167]_  = ~A269 & ~A268;
  assign \new_[44168]_  = A267 & \new_[44167]_ ;
  assign \new_[44171]_  = A299 & ~A298;
  assign \new_[44174]_  = A302 & A300;
  assign \new_[44175]_  = \new_[44174]_  & \new_[44171]_ ;
  assign \new_[44176]_  = \new_[44175]_  & \new_[44168]_ ;
  assign \new_[44180]_  = ~A167 & A168;
  assign \new_[44181]_  = ~A170 & \new_[44180]_ ;
  assign \new_[44185]_  = A200 & A199;
  assign \new_[44186]_  = A166 & \new_[44185]_ ;
  assign \new_[44187]_  = \new_[44186]_  & \new_[44181]_ ;
  assign \new_[44191]_  = A298 & A268;
  assign \new_[44192]_  = ~A267 & \new_[44191]_ ;
  assign \new_[44195]_  = ~A300 & ~A299;
  assign \new_[44198]_  = ~A302 & ~A301;
  assign \new_[44199]_  = \new_[44198]_  & \new_[44195]_ ;
  assign \new_[44200]_  = \new_[44199]_  & \new_[44192]_ ;
  assign \new_[44204]_  = ~A167 & A168;
  assign \new_[44205]_  = ~A170 & \new_[44204]_ ;
  assign \new_[44209]_  = A200 & A199;
  assign \new_[44210]_  = A166 & \new_[44209]_ ;
  assign \new_[44211]_  = \new_[44210]_  & \new_[44205]_ ;
  assign \new_[44215]_  = ~A298 & A268;
  assign \new_[44216]_  = ~A267 & \new_[44215]_ ;
  assign \new_[44219]_  = ~A300 & A299;
  assign \new_[44222]_  = ~A302 & ~A301;
  assign \new_[44223]_  = \new_[44222]_  & \new_[44219]_ ;
  assign \new_[44224]_  = \new_[44223]_  & \new_[44216]_ ;
  assign \new_[44228]_  = ~A167 & A168;
  assign \new_[44229]_  = ~A170 & \new_[44228]_ ;
  assign \new_[44233]_  = A200 & A199;
  assign \new_[44234]_  = A166 & \new_[44233]_ ;
  assign \new_[44235]_  = \new_[44234]_  & \new_[44229]_ ;
  assign \new_[44239]_  = A298 & A269;
  assign \new_[44240]_  = ~A267 & \new_[44239]_ ;
  assign \new_[44243]_  = ~A300 & ~A299;
  assign \new_[44246]_  = ~A302 & ~A301;
  assign \new_[44247]_  = \new_[44246]_  & \new_[44243]_ ;
  assign \new_[44248]_  = \new_[44247]_  & \new_[44240]_ ;
  assign \new_[44252]_  = ~A167 & A168;
  assign \new_[44253]_  = ~A170 & \new_[44252]_ ;
  assign \new_[44257]_  = A200 & A199;
  assign \new_[44258]_  = A166 & \new_[44257]_ ;
  assign \new_[44259]_  = \new_[44258]_  & \new_[44253]_ ;
  assign \new_[44263]_  = ~A298 & A269;
  assign \new_[44264]_  = ~A267 & \new_[44263]_ ;
  assign \new_[44267]_  = ~A300 & A299;
  assign \new_[44270]_  = ~A302 & ~A301;
  assign \new_[44271]_  = \new_[44270]_  & \new_[44267]_ ;
  assign \new_[44272]_  = \new_[44271]_  & \new_[44264]_ ;
  assign \new_[44276]_  = ~A167 & A168;
  assign \new_[44277]_  = ~A170 & \new_[44276]_ ;
  assign \new_[44281]_  = A200 & A199;
  assign \new_[44282]_  = A166 & \new_[44281]_ ;
  assign \new_[44283]_  = \new_[44282]_  & \new_[44277]_ ;
  assign \new_[44287]_  = A298 & A266;
  assign \new_[44288]_  = A265 & \new_[44287]_ ;
  assign \new_[44291]_  = ~A300 & ~A299;
  assign \new_[44294]_  = ~A302 & ~A301;
  assign \new_[44295]_  = \new_[44294]_  & \new_[44291]_ ;
  assign \new_[44296]_  = \new_[44295]_  & \new_[44288]_ ;
  assign \new_[44300]_  = ~A167 & A168;
  assign \new_[44301]_  = ~A170 & \new_[44300]_ ;
  assign \new_[44305]_  = A200 & A199;
  assign \new_[44306]_  = A166 & \new_[44305]_ ;
  assign \new_[44307]_  = \new_[44306]_  & \new_[44301]_ ;
  assign \new_[44311]_  = ~A298 & A266;
  assign \new_[44312]_  = A265 & \new_[44311]_ ;
  assign \new_[44315]_  = ~A300 & A299;
  assign \new_[44318]_  = ~A302 & ~A301;
  assign \new_[44319]_  = \new_[44318]_  & \new_[44315]_ ;
  assign \new_[44320]_  = \new_[44319]_  & \new_[44312]_ ;
  assign \new_[44324]_  = ~A167 & A168;
  assign \new_[44325]_  = ~A170 & \new_[44324]_ ;
  assign \new_[44329]_  = A200 & A199;
  assign \new_[44330]_  = A166 & \new_[44329]_ ;
  assign \new_[44331]_  = \new_[44330]_  & \new_[44325]_ ;
  assign \new_[44335]_  = A298 & ~A266;
  assign \new_[44336]_  = ~A265 & \new_[44335]_ ;
  assign \new_[44339]_  = ~A300 & ~A299;
  assign \new_[44342]_  = ~A302 & ~A301;
  assign \new_[44343]_  = \new_[44342]_  & \new_[44339]_ ;
  assign \new_[44344]_  = \new_[44343]_  & \new_[44336]_ ;
  assign \new_[44348]_  = ~A167 & A168;
  assign \new_[44349]_  = ~A170 & \new_[44348]_ ;
  assign \new_[44353]_  = A200 & A199;
  assign \new_[44354]_  = A166 & \new_[44353]_ ;
  assign \new_[44355]_  = \new_[44354]_  & \new_[44349]_ ;
  assign \new_[44359]_  = ~A298 & ~A266;
  assign \new_[44360]_  = ~A265 & \new_[44359]_ ;
  assign \new_[44363]_  = ~A300 & A299;
  assign \new_[44366]_  = ~A302 & ~A301;
  assign \new_[44367]_  = \new_[44366]_  & \new_[44363]_ ;
  assign \new_[44368]_  = \new_[44367]_  & \new_[44360]_ ;
  assign \new_[44372]_  = ~A167 & A168;
  assign \new_[44373]_  = ~A170 & \new_[44372]_ ;
  assign \new_[44377]_  = ~A200 & ~A199;
  assign \new_[44378]_  = A166 & \new_[44377]_ ;
  assign \new_[44379]_  = \new_[44378]_  & \new_[44373]_ ;
  assign \new_[44383]_  = ~A269 & ~A268;
  assign \new_[44384]_  = A267 & \new_[44383]_ ;
  assign \new_[44387]_  = ~A299 & A298;
  assign \new_[44390]_  = A301 & A300;
  assign \new_[44391]_  = \new_[44390]_  & \new_[44387]_ ;
  assign \new_[44392]_  = \new_[44391]_  & \new_[44384]_ ;
  assign \new_[44396]_  = ~A167 & A168;
  assign \new_[44397]_  = ~A170 & \new_[44396]_ ;
  assign \new_[44401]_  = ~A200 & ~A199;
  assign \new_[44402]_  = A166 & \new_[44401]_ ;
  assign \new_[44403]_  = \new_[44402]_  & \new_[44397]_ ;
  assign \new_[44407]_  = ~A269 & ~A268;
  assign \new_[44408]_  = A267 & \new_[44407]_ ;
  assign \new_[44411]_  = ~A299 & A298;
  assign \new_[44414]_  = A302 & A300;
  assign \new_[44415]_  = \new_[44414]_  & \new_[44411]_ ;
  assign \new_[44416]_  = \new_[44415]_  & \new_[44408]_ ;
  assign \new_[44420]_  = ~A167 & A168;
  assign \new_[44421]_  = ~A170 & \new_[44420]_ ;
  assign \new_[44425]_  = ~A200 & ~A199;
  assign \new_[44426]_  = A166 & \new_[44425]_ ;
  assign \new_[44427]_  = \new_[44426]_  & \new_[44421]_ ;
  assign \new_[44431]_  = ~A269 & ~A268;
  assign \new_[44432]_  = A267 & \new_[44431]_ ;
  assign \new_[44435]_  = A299 & ~A298;
  assign \new_[44438]_  = A301 & A300;
  assign \new_[44439]_  = \new_[44438]_  & \new_[44435]_ ;
  assign \new_[44440]_  = \new_[44439]_  & \new_[44432]_ ;
  assign \new_[44444]_  = ~A167 & A168;
  assign \new_[44445]_  = ~A170 & \new_[44444]_ ;
  assign \new_[44449]_  = ~A200 & ~A199;
  assign \new_[44450]_  = A166 & \new_[44449]_ ;
  assign \new_[44451]_  = \new_[44450]_  & \new_[44445]_ ;
  assign \new_[44455]_  = ~A269 & ~A268;
  assign \new_[44456]_  = A267 & \new_[44455]_ ;
  assign \new_[44459]_  = A299 & ~A298;
  assign \new_[44462]_  = A302 & A300;
  assign \new_[44463]_  = \new_[44462]_  & \new_[44459]_ ;
  assign \new_[44464]_  = \new_[44463]_  & \new_[44456]_ ;
  assign \new_[44468]_  = ~A167 & A168;
  assign \new_[44469]_  = ~A170 & \new_[44468]_ ;
  assign \new_[44473]_  = ~A200 & ~A199;
  assign \new_[44474]_  = A166 & \new_[44473]_ ;
  assign \new_[44475]_  = \new_[44474]_  & \new_[44469]_ ;
  assign \new_[44479]_  = A298 & A268;
  assign \new_[44480]_  = ~A267 & \new_[44479]_ ;
  assign \new_[44483]_  = ~A300 & ~A299;
  assign \new_[44486]_  = ~A302 & ~A301;
  assign \new_[44487]_  = \new_[44486]_  & \new_[44483]_ ;
  assign \new_[44488]_  = \new_[44487]_  & \new_[44480]_ ;
  assign \new_[44492]_  = ~A167 & A168;
  assign \new_[44493]_  = ~A170 & \new_[44492]_ ;
  assign \new_[44497]_  = ~A200 & ~A199;
  assign \new_[44498]_  = A166 & \new_[44497]_ ;
  assign \new_[44499]_  = \new_[44498]_  & \new_[44493]_ ;
  assign \new_[44503]_  = ~A298 & A268;
  assign \new_[44504]_  = ~A267 & \new_[44503]_ ;
  assign \new_[44507]_  = ~A300 & A299;
  assign \new_[44510]_  = ~A302 & ~A301;
  assign \new_[44511]_  = \new_[44510]_  & \new_[44507]_ ;
  assign \new_[44512]_  = \new_[44511]_  & \new_[44504]_ ;
  assign \new_[44516]_  = ~A167 & A168;
  assign \new_[44517]_  = ~A170 & \new_[44516]_ ;
  assign \new_[44521]_  = ~A200 & ~A199;
  assign \new_[44522]_  = A166 & \new_[44521]_ ;
  assign \new_[44523]_  = \new_[44522]_  & \new_[44517]_ ;
  assign \new_[44527]_  = A298 & A269;
  assign \new_[44528]_  = ~A267 & \new_[44527]_ ;
  assign \new_[44531]_  = ~A300 & ~A299;
  assign \new_[44534]_  = ~A302 & ~A301;
  assign \new_[44535]_  = \new_[44534]_  & \new_[44531]_ ;
  assign \new_[44536]_  = \new_[44535]_  & \new_[44528]_ ;
  assign \new_[44540]_  = ~A167 & A168;
  assign \new_[44541]_  = ~A170 & \new_[44540]_ ;
  assign \new_[44545]_  = ~A200 & ~A199;
  assign \new_[44546]_  = A166 & \new_[44545]_ ;
  assign \new_[44547]_  = \new_[44546]_  & \new_[44541]_ ;
  assign \new_[44551]_  = ~A298 & A269;
  assign \new_[44552]_  = ~A267 & \new_[44551]_ ;
  assign \new_[44555]_  = ~A300 & A299;
  assign \new_[44558]_  = ~A302 & ~A301;
  assign \new_[44559]_  = \new_[44558]_  & \new_[44555]_ ;
  assign \new_[44560]_  = \new_[44559]_  & \new_[44552]_ ;
  assign \new_[44564]_  = ~A167 & A168;
  assign \new_[44565]_  = ~A170 & \new_[44564]_ ;
  assign \new_[44569]_  = ~A200 & ~A199;
  assign \new_[44570]_  = A166 & \new_[44569]_ ;
  assign \new_[44571]_  = \new_[44570]_  & \new_[44565]_ ;
  assign \new_[44575]_  = A298 & A266;
  assign \new_[44576]_  = A265 & \new_[44575]_ ;
  assign \new_[44579]_  = ~A300 & ~A299;
  assign \new_[44582]_  = ~A302 & ~A301;
  assign \new_[44583]_  = \new_[44582]_  & \new_[44579]_ ;
  assign \new_[44584]_  = \new_[44583]_  & \new_[44576]_ ;
  assign \new_[44588]_  = ~A167 & A168;
  assign \new_[44589]_  = ~A170 & \new_[44588]_ ;
  assign \new_[44593]_  = ~A200 & ~A199;
  assign \new_[44594]_  = A166 & \new_[44593]_ ;
  assign \new_[44595]_  = \new_[44594]_  & \new_[44589]_ ;
  assign \new_[44599]_  = ~A298 & A266;
  assign \new_[44600]_  = A265 & \new_[44599]_ ;
  assign \new_[44603]_  = ~A300 & A299;
  assign \new_[44606]_  = ~A302 & ~A301;
  assign \new_[44607]_  = \new_[44606]_  & \new_[44603]_ ;
  assign \new_[44608]_  = \new_[44607]_  & \new_[44600]_ ;
  assign \new_[44612]_  = ~A167 & A168;
  assign \new_[44613]_  = ~A170 & \new_[44612]_ ;
  assign \new_[44617]_  = ~A200 & ~A199;
  assign \new_[44618]_  = A166 & \new_[44617]_ ;
  assign \new_[44619]_  = \new_[44618]_  & \new_[44613]_ ;
  assign \new_[44623]_  = A298 & ~A266;
  assign \new_[44624]_  = ~A265 & \new_[44623]_ ;
  assign \new_[44627]_  = ~A300 & ~A299;
  assign \new_[44630]_  = ~A302 & ~A301;
  assign \new_[44631]_  = \new_[44630]_  & \new_[44627]_ ;
  assign \new_[44632]_  = \new_[44631]_  & \new_[44624]_ ;
  assign \new_[44636]_  = ~A167 & A168;
  assign \new_[44637]_  = ~A170 & \new_[44636]_ ;
  assign \new_[44641]_  = ~A200 & ~A199;
  assign \new_[44642]_  = A166 & \new_[44641]_ ;
  assign \new_[44643]_  = \new_[44642]_  & \new_[44637]_ ;
  assign \new_[44647]_  = ~A298 & ~A266;
  assign \new_[44648]_  = ~A265 & \new_[44647]_ ;
  assign \new_[44651]_  = ~A300 & A299;
  assign \new_[44654]_  = ~A302 & ~A301;
  assign \new_[44655]_  = \new_[44654]_  & \new_[44651]_ ;
  assign \new_[44656]_  = \new_[44655]_  & \new_[44648]_ ;
  assign \new_[44660]_  = A201 & ~A168;
  assign \new_[44661]_  = ~A170 & \new_[44660]_ ;
  assign \new_[44665]_  = ~A265 & ~A203;
  assign \new_[44666]_  = ~A202 & \new_[44665]_ ;
  assign \new_[44667]_  = \new_[44666]_  & \new_[44661]_ ;
  assign \new_[44671]_  = ~A268 & ~A267;
  assign \new_[44672]_  = A266 & \new_[44671]_ ;
  assign \new_[44675]_  = A300 & ~A269;
  assign \new_[44678]_  = ~A302 & ~A301;
  assign \new_[44679]_  = \new_[44678]_  & \new_[44675]_ ;
  assign \new_[44680]_  = \new_[44679]_  & \new_[44672]_ ;
  assign \new_[44684]_  = A201 & ~A168;
  assign \new_[44685]_  = ~A170 & \new_[44684]_ ;
  assign \new_[44689]_  = A265 & ~A203;
  assign \new_[44690]_  = ~A202 & \new_[44689]_ ;
  assign \new_[44691]_  = \new_[44690]_  & \new_[44685]_ ;
  assign \new_[44695]_  = ~A268 & ~A267;
  assign \new_[44696]_  = ~A266 & \new_[44695]_ ;
  assign \new_[44699]_  = A300 & ~A269;
  assign \new_[44702]_  = ~A302 & ~A301;
  assign \new_[44703]_  = \new_[44702]_  & \new_[44699]_ ;
  assign \new_[44704]_  = \new_[44703]_  & \new_[44696]_ ;
  assign \new_[44708]_  = ~A199 & ~A168;
  assign \new_[44709]_  = ~A170 & \new_[44708]_ ;
  assign \new_[44713]_  = A202 & A201;
  assign \new_[44714]_  = A200 & \new_[44713]_ ;
  assign \new_[44715]_  = \new_[44714]_  & \new_[44709]_ ;
  assign \new_[44719]_  = ~A269 & ~A268;
  assign \new_[44720]_  = A267 & \new_[44719]_ ;
  assign \new_[44723]_  = ~A299 & A298;
  assign \new_[44726]_  = A301 & A300;
  assign \new_[44727]_  = \new_[44726]_  & \new_[44723]_ ;
  assign \new_[44728]_  = \new_[44727]_  & \new_[44720]_ ;
  assign \new_[44732]_  = ~A199 & ~A168;
  assign \new_[44733]_  = ~A170 & \new_[44732]_ ;
  assign \new_[44737]_  = A202 & A201;
  assign \new_[44738]_  = A200 & \new_[44737]_ ;
  assign \new_[44739]_  = \new_[44738]_  & \new_[44733]_ ;
  assign \new_[44743]_  = ~A269 & ~A268;
  assign \new_[44744]_  = A267 & \new_[44743]_ ;
  assign \new_[44747]_  = ~A299 & A298;
  assign \new_[44750]_  = A302 & A300;
  assign \new_[44751]_  = \new_[44750]_  & \new_[44747]_ ;
  assign \new_[44752]_  = \new_[44751]_  & \new_[44744]_ ;
  assign \new_[44756]_  = ~A199 & ~A168;
  assign \new_[44757]_  = ~A170 & \new_[44756]_ ;
  assign \new_[44761]_  = A202 & A201;
  assign \new_[44762]_  = A200 & \new_[44761]_ ;
  assign \new_[44763]_  = \new_[44762]_  & \new_[44757]_ ;
  assign \new_[44767]_  = ~A269 & ~A268;
  assign \new_[44768]_  = A267 & \new_[44767]_ ;
  assign \new_[44771]_  = A299 & ~A298;
  assign \new_[44774]_  = A301 & A300;
  assign \new_[44775]_  = \new_[44774]_  & \new_[44771]_ ;
  assign \new_[44776]_  = \new_[44775]_  & \new_[44768]_ ;
  assign \new_[44780]_  = ~A199 & ~A168;
  assign \new_[44781]_  = ~A170 & \new_[44780]_ ;
  assign \new_[44785]_  = A202 & A201;
  assign \new_[44786]_  = A200 & \new_[44785]_ ;
  assign \new_[44787]_  = \new_[44786]_  & \new_[44781]_ ;
  assign \new_[44791]_  = ~A269 & ~A268;
  assign \new_[44792]_  = A267 & \new_[44791]_ ;
  assign \new_[44795]_  = A299 & ~A298;
  assign \new_[44798]_  = A302 & A300;
  assign \new_[44799]_  = \new_[44798]_  & \new_[44795]_ ;
  assign \new_[44800]_  = \new_[44799]_  & \new_[44792]_ ;
  assign \new_[44804]_  = ~A199 & ~A168;
  assign \new_[44805]_  = ~A170 & \new_[44804]_ ;
  assign \new_[44809]_  = A202 & A201;
  assign \new_[44810]_  = A200 & \new_[44809]_ ;
  assign \new_[44811]_  = \new_[44810]_  & \new_[44805]_ ;
  assign \new_[44815]_  = A298 & A268;
  assign \new_[44816]_  = ~A267 & \new_[44815]_ ;
  assign \new_[44819]_  = ~A300 & ~A299;
  assign \new_[44822]_  = ~A302 & ~A301;
  assign \new_[44823]_  = \new_[44822]_  & \new_[44819]_ ;
  assign \new_[44824]_  = \new_[44823]_  & \new_[44816]_ ;
  assign \new_[44828]_  = ~A199 & ~A168;
  assign \new_[44829]_  = ~A170 & \new_[44828]_ ;
  assign \new_[44833]_  = A202 & A201;
  assign \new_[44834]_  = A200 & \new_[44833]_ ;
  assign \new_[44835]_  = \new_[44834]_  & \new_[44829]_ ;
  assign \new_[44839]_  = ~A298 & A268;
  assign \new_[44840]_  = ~A267 & \new_[44839]_ ;
  assign \new_[44843]_  = ~A300 & A299;
  assign \new_[44846]_  = ~A302 & ~A301;
  assign \new_[44847]_  = \new_[44846]_  & \new_[44843]_ ;
  assign \new_[44848]_  = \new_[44847]_  & \new_[44840]_ ;
  assign \new_[44852]_  = ~A199 & ~A168;
  assign \new_[44853]_  = ~A170 & \new_[44852]_ ;
  assign \new_[44857]_  = A202 & A201;
  assign \new_[44858]_  = A200 & \new_[44857]_ ;
  assign \new_[44859]_  = \new_[44858]_  & \new_[44853]_ ;
  assign \new_[44863]_  = A298 & A269;
  assign \new_[44864]_  = ~A267 & \new_[44863]_ ;
  assign \new_[44867]_  = ~A300 & ~A299;
  assign \new_[44870]_  = ~A302 & ~A301;
  assign \new_[44871]_  = \new_[44870]_  & \new_[44867]_ ;
  assign \new_[44872]_  = \new_[44871]_  & \new_[44864]_ ;
  assign \new_[44876]_  = ~A199 & ~A168;
  assign \new_[44877]_  = ~A170 & \new_[44876]_ ;
  assign \new_[44881]_  = A202 & A201;
  assign \new_[44882]_  = A200 & \new_[44881]_ ;
  assign \new_[44883]_  = \new_[44882]_  & \new_[44877]_ ;
  assign \new_[44887]_  = ~A298 & A269;
  assign \new_[44888]_  = ~A267 & \new_[44887]_ ;
  assign \new_[44891]_  = ~A300 & A299;
  assign \new_[44894]_  = ~A302 & ~A301;
  assign \new_[44895]_  = \new_[44894]_  & \new_[44891]_ ;
  assign \new_[44896]_  = \new_[44895]_  & \new_[44888]_ ;
  assign \new_[44900]_  = ~A199 & ~A168;
  assign \new_[44901]_  = ~A170 & \new_[44900]_ ;
  assign \new_[44905]_  = A202 & A201;
  assign \new_[44906]_  = A200 & \new_[44905]_ ;
  assign \new_[44907]_  = \new_[44906]_  & \new_[44901]_ ;
  assign \new_[44911]_  = A298 & A266;
  assign \new_[44912]_  = A265 & \new_[44911]_ ;
  assign \new_[44915]_  = ~A300 & ~A299;
  assign \new_[44918]_  = ~A302 & ~A301;
  assign \new_[44919]_  = \new_[44918]_  & \new_[44915]_ ;
  assign \new_[44920]_  = \new_[44919]_  & \new_[44912]_ ;
  assign \new_[44924]_  = ~A199 & ~A168;
  assign \new_[44925]_  = ~A170 & \new_[44924]_ ;
  assign \new_[44929]_  = A202 & A201;
  assign \new_[44930]_  = A200 & \new_[44929]_ ;
  assign \new_[44931]_  = \new_[44930]_  & \new_[44925]_ ;
  assign \new_[44935]_  = ~A298 & A266;
  assign \new_[44936]_  = A265 & \new_[44935]_ ;
  assign \new_[44939]_  = ~A300 & A299;
  assign \new_[44942]_  = ~A302 & ~A301;
  assign \new_[44943]_  = \new_[44942]_  & \new_[44939]_ ;
  assign \new_[44944]_  = \new_[44943]_  & \new_[44936]_ ;
  assign \new_[44948]_  = ~A199 & ~A168;
  assign \new_[44949]_  = ~A170 & \new_[44948]_ ;
  assign \new_[44953]_  = A202 & A201;
  assign \new_[44954]_  = A200 & \new_[44953]_ ;
  assign \new_[44955]_  = \new_[44954]_  & \new_[44949]_ ;
  assign \new_[44959]_  = A298 & ~A266;
  assign \new_[44960]_  = ~A265 & \new_[44959]_ ;
  assign \new_[44963]_  = ~A300 & ~A299;
  assign \new_[44966]_  = ~A302 & ~A301;
  assign \new_[44967]_  = \new_[44966]_  & \new_[44963]_ ;
  assign \new_[44968]_  = \new_[44967]_  & \new_[44960]_ ;
  assign \new_[44972]_  = ~A199 & ~A168;
  assign \new_[44973]_  = ~A170 & \new_[44972]_ ;
  assign \new_[44977]_  = A202 & A201;
  assign \new_[44978]_  = A200 & \new_[44977]_ ;
  assign \new_[44979]_  = \new_[44978]_  & \new_[44973]_ ;
  assign \new_[44983]_  = ~A298 & ~A266;
  assign \new_[44984]_  = ~A265 & \new_[44983]_ ;
  assign \new_[44987]_  = ~A300 & A299;
  assign \new_[44990]_  = ~A302 & ~A301;
  assign \new_[44991]_  = \new_[44990]_  & \new_[44987]_ ;
  assign \new_[44992]_  = \new_[44991]_  & \new_[44984]_ ;
  assign \new_[44996]_  = ~A199 & ~A168;
  assign \new_[44997]_  = ~A170 & \new_[44996]_ ;
  assign \new_[45001]_  = A203 & A201;
  assign \new_[45002]_  = A200 & \new_[45001]_ ;
  assign \new_[45003]_  = \new_[45002]_  & \new_[44997]_ ;
  assign \new_[45007]_  = ~A269 & ~A268;
  assign \new_[45008]_  = A267 & \new_[45007]_ ;
  assign \new_[45011]_  = ~A299 & A298;
  assign \new_[45014]_  = A301 & A300;
  assign \new_[45015]_  = \new_[45014]_  & \new_[45011]_ ;
  assign \new_[45016]_  = \new_[45015]_  & \new_[45008]_ ;
  assign \new_[45020]_  = ~A199 & ~A168;
  assign \new_[45021]_  = ~A170 & \new_[45020]_ ;
  assign \new_[45025]_  = A203 & A201;
  assign \new_[45026]_  = A200 & \new_[45025]_ ;
  assign \new_[45027]_  = \new_[45026]_  & \new_[45021]_ ;
  assign \new_[45031]_  = ~A269 & ~A268;
  assign \new_[45032]_  = A267 & \new_[45031]_ ;
  assign \new_[45035]_  = ~A299 & A298;
  assign \new_[45038]_  = A302 & A300;
  assign \new_[45039]_  = \new_[45038]_  & \new_[45035]_ ;
  assign \new_[45040]_  = \new_[45039]_  & \new_[45032]_ ;
  assign \new_[45044]_  = ~A199 & ~A168;
  assign \new_[45045]_  = ~A170 & \new_[45044]_ ;
  assign \new_[45049]_  = A203 & A201;
  assign \new_[45050]_  = A200 & \new_[45049]_ ;
  assign \new_[45051]_  = \new_[45050]_  & \new_[45045]_ ;
  assign \new_[45055]_  = ~A269 & ~A268;
  assign \new_[45056]_  = A267 & \new_[45055]_ ;
  assign \new_[45059]_  = A299 & ~A298;
  assign \new_[45062]_  = A301 & A300;
  assign \new_[45063]_  = \new_[45062]_  & \new_[45059]_ ;
  assign \new_[45064]_  = \new_[45063]_  & \new_[45056]_ ;
  assign \new_[45068]_  = ~A199 & ~A168;
  assign \new_[45069]_  = ~A170 & \new_[45068]_ ;
  assign \new_[45073]_  = A203 & A201;
  assign \new_[45074]_  = A200 & \new_[45073]_ ;
  assign \new_[45075]_  = \new_[45074]_  & \new_[45069]_ ;
  assign \new_[45079]_  = ~A269 & ~A268;
  assign \new_[45080]_  = A267 & \new_[45079]_ ;
  assign \new_[45083]_  = A299 & ~A298;
  assign \new_[45086]_  = A302 & A300;
  assign \new_[45087]_  = \new_[45086]_  & \new_[45083]_ ;
  assign \new_[45088]_  = \new_[45087]_  & \new_[45080]_ ;
  assign \new_[45092]_  = ~A199 & ~A168;
  assign \new_[45093]_  = ~A170 & \new_[45092]_ ;
  assign \new_[45097]_  = A203 & A201;
  assign \new_[45098]_  = A200 & \new_[45097]_ ;
  assign \new_[45099]_  = \new_[45098]_  & \new_[45093]_ ;
  assign \new_[45103]_  = A298 & A268;
  assign \new_[45104]_  = ~A267 & \new_[45103]_ ;
  assign \new_[45107]_  = ~A300 & ~A299;
  assign \new_[45110]_  = ~A302 & ~A301;
  assign \new_[45111]_  = \new_[45110]_  & \new_[45107]_ ;
  assign \new_[45112]_  = \new_[45111]_  & \new_[45104]_ ;
  assign \new_[45116]_  = ~A199 & ~A168;
  assign \new_[45117]_  = ~A170 & \new_[45116]_ ;
  assign \new_[45121]_  = A203 & A201;
  assign \new_[45122]_  = A200 & \new_[45121]_ ;
  assign \new_[45123]_  = \new_[45122]_  & \new_[45117]_ ;
  assign \new_[45127]_  = ~A298 & A268;
  assign \new_[45128]_  = ~A267 & \new_[45127]_ ;
  assign \new_[45131]_  = ~A300 & A299;
  assign \new_[45134]_  = ~A302 & ~A301;
  assign \new_[45135]_  = \new_[45134]_  & \new_[45131]_ ;
  assign \new_[45136]_  = \new_[45135]_  & \new_[45128]_ ;
  assign \new_[45140]_  = ~A199 & ~A168;
  assign \new_[45141]_  = ~A170 & \new_[45140]_ ;
  assign \new_[45145]_  = A203 & A201;
  assign \new_[45146]_  = A200 & \new_[45145]_ ;
  assign \new_[45147]_  = \new_[45146]_  & \new_[45141]_ ;
  assign \new_[45151]_  = A298 & A269;
  assign \new_[45152]_  = ~A267 & \new_[45151]_ ;
  assign \new_[45155]_  = ~A300 & ~A299;
  assign \new_[45158]_  = ~A302 & ~A301;
  assign \new_[45159]_  = \new_[45158]_  & \new_[45155]_ ;
  assign \new_[45160]_  = \new_[45159]_  & \new_[45152]_ ;
  assign \new_[45164]_  = ~A199 & ~A168;
  assign \new_[45165]_  = ~A170 & \new_[45164]_ ;
  assign \new_[45169]_  = A203 & A201;
  assign \new_[45170]_  = A200 & \new_[45169]_ ;
  assign \new_[45171]_  = \new_[45170]_  & \new_[45165]_ ;
  assign \new_[45175]_  = ~A298 & A269;
  assign \new_[45176]_  = ~A267 & \new_[45175]_ ;
  assign \new_[45179]_  = ~A300 & A299;
  assign \new_[45182]_  = ~A302 & ~A301;
  assign \new_[45183]_  = \new_[45182]_  & \new_[45179]_ ;
  assign \new_[45184]_  = \new_[45183]_  & \new_[45176]_ ;
  assign \new_[45188]_  = ~A199 & ~A168;
  assign \new_[45189]_  = ~A170 & \new_[45188]_ ;
  assign \new_[45193]_  = A203 & A201;
  assign \new_[45194]_  = A200 & \new_[45193]_ ;
  assign \new_[45195]_  = \new_[45194]_  & \new_[45189]_ ;
  assign \new_[45199]_  = A298 & A266;
  assign \new_[45200]_  = A265 & \new_[45199]_ ;
  assign \new_[45203]_  = ~A300 & ~A299;
  assign \new_[45206]_  = ~A302 & ~A301;
  assign \new_[45207]_  = \new_[45206]_  & \new_[45203]_ ;
  assign \new_[45208]_  = \new_[45207]_  & \new_[45200]_ ;
  assign \new_[45212]_  = ~A199 & ~A168;
  assign \new_[45213]_  = ~A170 & \new_[45212]_ ;
  assign \new_[45217]_  = A203 & A201;
  assign \new_[45218]_  = A200 & \new_[45217]_ ;
  assign \new_[45219]_  = \new_[45218]_  & \new_[45213]_ ;
  assign \new_[45223]_  = ~A298 & A266;
  assign \new_[45224]_  = A265 & \new_[45223]_ ;
  assign \new_[45227]_  = ~A300 & A299;
  assign \new_[45230]_  = ~A302 & ~A301;
  assign \new_[45231]_  = \new_[45230]_  & \new_[45227]_ ;
  assign \new_[45232]_  = \new_[45231]_  & \new_[45224]_ ;
  assign \new_[45236]_  = ~A199 & ~A168;
  assign \new_[45237]_  = ~A170 & \new_[45236]_ ;
  assign \new_[45241]_  = A203 & A201;
  assign \new_[45242]_  = A200 & \new_[45241]_ ;
  assign \new_[45243]_  = \new_[45242]_  & \new_[45237]_ ;
  assign \new_[45247]_  = A298 & ~A266;
  assign \new_[45248]_  = ~A265 & \new_[45247]_ ;
  assign \new_[45251]_  = ~A300 & ~A299;
  assign \new_[45254]_  = ~A302 & ~A301;
  assign \new_[45255]_  = \new_[45254]_  & \new_[45251]_ ;
  assign \new_[45256]_  = \new_[45255]_  & \new_[45248]_ ;
  assign \new_[45260]_  = ~A199 & ~A168;
  assign \new_[45261]_  = ~A170 & \new_[45260]_ ;
  assign \new_[45265]_  = A203 & A201;
  assign \new_[45266]_  = A200 & \new_[45265]_ ;
  assign \new_[45267]_  = \new_[45266]_  & \new_[45261]_ ;
  assign \new_[45271]_  = ~A298 & ~A266;
  assign \new_[45272]_  = ~A265 & \new_[45271]_ ;
  assign \new_[45275]_  = ~A300 & A299;
  assign \new_[45278]_  = ~A302 & ~A301;
  assign \new_[45279]_  = \new_[45278]_  & \new_[45275]_ ;
  assign \new_[45280]_  = \new_[45279]_  & \new_[45272]_ ;
  assign \new_[45284]_  = ~A199 & ~A168;
  assign \new_[45285]_  = ~A170 & \new_[45284]_ ;
  assign \new_[45289]_  = ~A202 & ~A201;
  assign \new_[45290]_  = A200 & \new_[45289]_ ;
  assign \new_[45291]_  = \new_[45290]_  & \new_[45285]_ ;
  assign \new_[45295]_  = A268 & ~A267;
  assign \new_[45296]_  = ~A203 & \new_[45295]_ ;
  assign \new_[45299]_  = ~A299 & A298;
  assign \new_[45302]_  = A301 & A300;
  assign \new_[45303]_  = \new_[45302]_  & \new_[45299]_ ;
  assign \new_[45304]_  = \new_[45303]_  & \new_[45296]_ ;
  assign \new_[45308]_  = ~A199 & ~A168;
  assign \new_[45309]_  = ~A170 & \new_[45308]_ ;
  assign \new_[45313]_  = ~A202 & ~A201;
  assign \new_[45314]_  = A200 & \new_[45313]_ ;
  assign \new_[45315]_  = \new_[45314]_  & \new_[45309]_ ;
  assign \new_[45319]_  = A268 & ~A267;
  assign \new_[45320]_  = ~A203 & \new_[45319]_ ;
  assign \new_[45323]_  = ~A299 & A298;
  assign \new_[45326]_  = A302 & A300;
  assign \new_[45327]_  = \new_[45326]_  & \new_[45323]_ ;
  assign \new_[45328]_  = \new_[45327]_  & \new_[45320]_ ;
  assign \new_[45332]_  = ~A199 & ~A168;
  assign \new_[45333]_  = ~A170 & \new_[45332]_ ;
  assign \new_[45337]_  = ~A202 & ~A201;
  assign \new_[45338]_  = A200 & \new_[45337]_ ;
  assign \new_[45339]_  = \new_[45338]_  & \new_[45333]_ ;
  assign \new_[45343]_  = A268 & ~A267;
  assign \new_[45344]_  = ~A203 & \new_[45343]_ ;
  assign \new_[45347]_  = A299 & ~A298;
  assign \new_[45350]_  = A301 & A300;
  assign \new_[45351]_  = \new_[45350]_  & \new_[45347]_ ;
  assign \new_[45352]_  = \new_[45351]_  & \new_[45344]_ ;
  assign \new_[45356]_  = ~A199 & ~A168;
  assign \new_[45357]_  = ~A170 & \new_[45356]_ ;
  assign \new_[45361]_  = ~A202 & ~A201;
  assign \new_[45362]_  = A200 & \new_[45361]_ ;
  assign \new_[45363]_  = \new_[45362]_  & \new_[45357]_ ;
  assign \new_[45367]_  = A268 & ~A267;
  assign \new_[45368]_  = ~A203 & \new_[45367]_ ;
  assign \new_[45371]_  = A299 & ~A298;
  assign \new_[45374]_  = A302 & A300;
  assign \new_[45375]_  = \new_[45374]_  & \new_[45371]_ ;
  assign \new_[45376]_  = \new_[45375]_  & \new_[45368]_ ;
  assign \new_[45380]_  = ~A199 & ~A168;
  assign \new_[45381]_  = ~A170 & \new_[45380]_ ;
  assign \new_[45385]_  = ~A202 & ~A201;
  assign \new_[45386]_  = A200 & \new_[45385]_ ;
  assign \new_[45387]_  = \new_[45386]_  & \new_[45381]_ ;
  assign \new_[45391]_  = A269 & ~A267;
  assign \new_[45392]_  = ~A203 & \new_[45391]_ ;
  assign \new_[45395]_  = ~A299 & A298;
  assign \new_[45398]_  = A301 & A300;
  assign \new_[45399]_  = \new_[45398]_  & \new_[45395]_ ;
  assign \new_[45400]_  = \new_[45399]_  & \new_[45392]_ ;
  assign \new_[45404]_  = ~A199 & ~A168;
  assign \new_[45405]_  = ~A170 & \new_[45404]_ ;
  assign \new_[45409]_  = ~A202 & ~A201;
  assign \new_[45410]_  = A200 & \new_[45409]_ ;
  assign \new_[45411]_  = \new_[45410]_  & \new_[45405]_ ;
  assign \new_[45415]_  = A269 & ~A267;
  assign \new_[45416]_  = ~A203 & \new_[45415]_ ;
  assign \new_[45419]_  = ~A299 & A298;
  assign \new_[45422]_  = A302 & A300;
  assign \new_[45423]_  = \new_[45422]_  & \new_[45419]_ ;
  assign \new_[45424]_  = \new_[45423]_  & \new_[45416]_ ;
  assign \new_[45428]_  = ~A199 & ~A168;
  assign \new_[45429]_  = ~A170 & \new_[45428]_ ;
  assign \new_[45433]_  = ~A202 & ~A201;
  assign \new_[45434]_  = A200 & \new_[45433]_ ;
  assign \new_[45435]_  = \new_[45434]_  & \new_[45429]_ ;
  assign \new_[45439]_  = A269 & ~A267;
  assign \new_[45440]_  = ~A203 & \new_[45439]_ ;
  assign \new_[45443]_  = A299 & ~A298;
  assign \new_[45446]_  = A301 & A300;
  assign \new_[45447]_  = \new_[45446]_  & \new_[45443]_ ;
  assign \new_[45448]_  = \new_[45447]_  & \new_[45440]_ ;
  assign \new_[45452]_  = ~A199 & ~A168;
  assign \new_[45453]_  = ~A170 & \new_[45452]_ ;
  assign \new_[45457]_  = ~A202 & ~A201;
  assign \new_[45458]_  = A200 & \new_[45457]_ ;
  assign \new_[45459]_  = \new_[45458]_  & \new_[45453]_ ;
  assign \new_[45463]_  = A269 & ~A267;
  assign \new_[45464]_  = ~A203 & \new_[45463]_ ;
  assign \new_[45467]_  = A299 & ~A298;
  assign \new_[45470]_  = A302 & A300;
  assign \new_[45471]_  = \new_[45470]_  & \new_[45467]_ ;
  assign \new_[45472]_  = \new_[45471]_  & \new_[45464]_ ;
  assign \new_[45476]_  = ~A199 & ~A168;
  assign \new_[45477]_  = ~A170 & \new_[45476]_ ;
  assign \new_[45481]_  = ~A202 & ~A201;
  assign \new_[45482]_  = A200 & \new_[45481]_ ;
  assign \new_[45483]_  = \new_[45482]_  & \new_[45477]_ ;
  assign \new_[45487]_  = A266 & A265;
  assign \new_[45488]_  = ~A203 & \new_[45487]_ ;
  assign \new_[45491]_  = ~A299 & A298;
  assign \new_[45494]_  = A301 & A300;
  assign \new_[45495]_  = \new_[45494]_  & \new_[45491]_ ;
  assign \new_[45496]_  = \new_[45495]_  & \new_[45488]_ ;
  assign \new_[45500]_  = ~A199 & ~A168;
  assign \new_[45501]_  = ~A170 & \new_[45500]_ ;
  assign \new_[45505]_  = ~A202 & ~A201;
  assign \new_[45506]_  = A200 & \new_[45505]_ ;
  assign \new_[45507]_  = \new_[45506]_  & \new_[45501]_ ;
  assign \new_[45511]_  = A266 & A265;
  assign \new_[45512]_  = ~A203 & \new_[45511]_ ;
  assign \new_[45515]_  = ~A299 & A298;
  assign \new_[45518]_  = A302 & A300;
  assign \new_[45519]_  = \new_[45518]_  & \new_[45515]_ ;
  assign \new_[45520]_  = \new_[45519]_  & \new_[45512]_ ;
  assign \new_[45524]_  = ~A199 & ~A168;
  assign \new_[45525]_  = ~A170 & \new_[45524]_ ;
  assign \new_[45529]_  = ~A202 & ~A201;
  assign \new_[45530]_  = A200 & \new_[45529]_ ;
  assign \new_[45531]_  = \new_[45530]_  & \new_[45525]_ ;
  assign \new_[45535]_  = A266 & A265;
  assign \new_[45536]_  = ~A203 & \new_[45535]_ ;
  assign \new_[45539]_  = A299 & ~A298;
  assign \new_[45542]_  = A301 & A300;
  assign \new_[45543]_  = \new_[45542]_  & \new_[45539]_ ;
  assign \new_[45544]_  = \new_[45543]_  & \new_[45536]_ ;
  assign \new_[45548]_  = ~A199 & ~A168;
  assign \new_[45549]_  = ~A170 & \new_[45548]_ ;
  assign \new_[45553]_  = ~A202 & ~A201;
  assign \new_[45554]_  = A200 & \new_[45553]_ ;
  assign \new_[45555]_  = \new_[45554]_  & \new_[45549]_ ;
  assign \new_[45559]_  = A266 & A265;
  assign \new_[45560]_  = ~A203 & \new_[45559]_ ;
  assign \new_[45563]_  = A299 & ~A298;
  assign \new_[45566]_  = A302 & A300;
  assign \new_[45567]_  = \new_[45566]_  & \new_[45563]_ ;
  assign \new_[45568]_  = \new_[45567]_  & \new_[45560]_ ;
  assign \new_[45572]_  = ~A199 & ~A168;
  assign \new_[45573]_  = ~A170 & \new_[45572]_ ;
  assign \new_[45577]_  = ~A202 & ~A201;
  assign \new_[45578]_  = A200 & \new_[45577]_ ;
  assign \new_[45579]_  = \new_[45578]_  & \new_[45573]_ ;
  assign \new_[45583]_  = ~A266 & ~A265;
  assign \new_[45584]_  = ~A203 & \new_[45583]_ ;
  assign \new_[45587]_  = ~A299 & A298;
  assign \new_[45590]_  = A301 & A300;
  assign \new_[45591]_  = \new_[45590]_  & \new_[45587]_ ;
  assign \new_[45592]_  = \new_[45591]_  & \new_[45584]_ ;
  assign \new_[45596]_  = ~A199 & ~A168;
  assign \new_[45597]_  = ~A170 & \new_[45596]_ ;
  assign \new_[45601]_  = ~A202 & ~A201;
  assign \new_[45602]_  = A200 & \new_[45601]_ ;
  assign \new_[45603]_  = \new_[45602]_  & \new_[45597]_ ;
  assign \new_[45607]_  = ~A266 & ~A265;
  assign \new_[45608]_  = ~A203 & \new_[45607]_ ;
  assign \new_[45611]_  = ~A299 & A298;
  assign \new_[45614]_  = A302 & A300;
  assign \new_[45615]_  = \new_[45614]_  & \new_[45611]_ ;
  assign \new_[45616]_  = \new_[45615]_  & \new_[45608]_ ;
  assign \new_[45620]_  = ~A199 & ~A168;
  assign \new_[45621]_  = ~A170 & \new_[45620]_ ;
  assign \new_[45625]_  = ~A202 & ~A201;
  assign \new_[45626]_  = A200 & \new_[45625]_ ;
  assign \new_[45627]_  = \new_[45626]_  & \new_[45621]_ ;
  assign \new_[45631]_  = ~A266 & ~A265;
  assign \new_[45632]_  = ~A203 & \new_[45631]_ ;
  assign \new_[45635]_  = A299 & ~A298;
  assign \new_[45638]_  = A301 & A300;
  assign \new_[45639]_  = \new_[45638]_  & \new_[45635]_ ;
  assign \new_[45640]_  = \new_[45639]_  & \new_[45632]_ ;
  assign \new_[45644]_  = ~A199 & ~A168;
  assign \new_[45645]_  = ~A170 & \new_[45644]_ ;
  assign \new_[45649]_  = ~A202 & ~A201;
  assign \new_[45650]_  = A200 & \new_[45649]_ ;
  assign \new_[45651]_  = \new_[45650]_  & \new_[45645]_ ;
  assign \new_[45655]_  = ~A266 & ~A265;
  assign \new_[45656]_  = ~A203 & \new_[45655]_ ;
  assign \new_[45659]_  = A299 & ~A298;
  assign \new_[45662]_  = A302 & A300;
  assign \new_[45663]_  = \new_[45662]_  & \new_[45659]_ ;
  assign \new_[45664]_  = \new_[45663]_  & \new_[45656]_ ;
  assign \new_[45668]_  = A199 & ~A168;
  assign \new_[45669]_  = ~A170 & \new_[45668]_ ;
  assign \new_[45673]_  = A202 & A201;
  assign \new_[45674]_  = ~A200 & \new_[45673]_ ;
  assign \new_[45675]_  = \new_[45674]_  & \new_[45669]_ ;
  assign \new_[45679]_  = ~A269 & ~A268;
  assign \new_[45680]_  = A267 & \new_[45679]_ ;
  assign \new_[45683]_  = ~A299 & A298;
  assign \new_[45686]_  = A301 & A300;
  assign \new_[45687]_  = \new_[45686]_  & \new_[45683]_ ;
  assign \new_[45688]_  = \new_[45687]_  & \new_[45680]_ ;
  assign \new_[45692]_  = A199 & ~A168;
  assign \new_[45693]_  = ~A170 & \new_[45692]_ ;
  assign \new_[45697]_  = A202 & A201;
  assign \new_[45698]_  = ~A200 & \new_[45697]_ ;
  assign \new_[45699]_  = \new_[45698]_  & \new_[45693]_ ;
  assign \new_[45703]_  = ~A269 & ~A268;
  assign \new_[45704]_  = A267 & \new_[45703]_ ;
  assign \new_[45707]_  = ~A299 & A298;
  assign \new_[45710]_  = A302 & A300;
  assign \new_[45711]_  = \new_[45710]_  & \new_[45707]_ ;
  assign \new_[45712]_  = \new_[45711]_  & \new_[45704]_ ;
  assign \new_[45716]_  = A199 & ~A168;
  assign \new_[45717]_  = ~A170 & \new_[45716]_ ;
  assign \new_[45721]_  = A202 & A201;
  assign \new_[45722]_  = ~A200 & \new_[45721]_ ;
  assign \new_[45723]_  = \new_[45722]_  & \new_[45717]_ ;
  assign \new_[45727]_  = ~A269 & ~A268;
  assign \new_[45728]_  = A267 & \new_[45727]_ ;
  assign \new_[45731]_  = A299 & ~A298;
  assign \new_[45734]_  = A301 & A300;
  assign \new_[45735]_  = \new_[45734]_  & \new_[45731]_ ;
  assign \new_[45736]_  = \new_[45735]_  & \new_[45728]_ ;
  assign \new_[45740]_  = A199 & ~A168;
  assign \new_[45741]_  = ~A170 & \new_[45740]_ ;
  assign \new_[45745]_  = A202 & A201;
  assign \new_[45746]_  = ~A200 & \new_[45745]_ ;
  assign \new_[45747]_  = \new_[45746]_  & \new_[45741]_ ;
  assign \new_[45751]_  = ~A269 & ~A268;
  assign \new_[45752]_  = A267 & \new_[45751]_ ;
  assign \new_[45755]_  = A299 & ~A298;
  assign \new_[45758]_  = A302 & A300;
  assign \new_[45759]_  = \new_[45758]_  & \new_[45755]_ ;
  assign \new_[45760]_  = \new_[45759]_  & \new_[45752]_ ;
  assign \new_[45764]_  = A199 & ~A168;
  assign \new_[45765]_  = ~A170 & \new_[45764]_ ;
  assign \new_[45769]_  = A202 & A201;
  assign \new_[45770]_  = ~A200 & \new_[45769]_ ;
  assign \new_[45771]_  = \new_[45770]_  & \new_[45765]_ ;
  assign \new_[45775]_  = A298 & A268;
  assign \new_[45776]_  = ~A267 & \new_[45775]_ ;
  assign \new_[45779]_  = ~A300 & ~A299;
  assign \new_[45782]_  = ~A302 & ~A301;
  assign \new_[45783]_  = \new_[45782]_  & \new_[45779]_ ;
  assign \new_[45784]_  = \new_[45783]_  & \new_[45776]_ ;
  assign \new_[45788]_  = A199 & ~A168;
  assign \new_[45789]_  = ~A170 & \new_[45788]_ ;
  assign \new_[45793]_  = A202 & A201;
  assign \new_[45794]_  = ~A200 & \new_[45793]_ ;
  assign \new_[45795]_  = \new_[45794]_  & \new_[45789]_ ;
  assign \new_[45799]_  = ~A298 & A268;
  assign \new_[45800]_  = ~A267 & \new_[45799]_ ;
  assign \new_[45803]_  = ~A300 & A299;
  assign \new_[45806]_  = ~A302 & ~A301;
  assign \new_[45807]_  = \new_[45806]_  & \new_[45803]_ ;
  assign \new_[45808]_  = \new_[45807]_  & \new_[45800]_ ;
  assign \new_[45812]_  = A199 & ~A168;
  assign \new_[45813]_  = ~A170 & \new_[45812]_ ;
  assign \new_[45817]_  = A202 & A201;
  assign \new_[45818]_  = ~A200 & \new_[45817]_ ;
  assign \new_[45819]_  = \new_[45818]_  & \new_[45813]_ ;
  assign \new_[45823]_  = A298 & A269;
  assign \new_[45824]_  = ~A267 & \new_[45823]_ ;
  assign \new_[45827]_  = ~A300 & ~A299;
  assign \new_[45830]_  = ~A302 & ~A301;
  assign \new_[45831]_  = \new_[45830]_  & \new_[45827]_ ;
  assign \new_[45832]_  = \new_[45831]_  & \new_[45824]_ ;
  assign \new_[45836]_  = A199 & ~A168;
  assign \new_[45837]_  = ~A170 & \new_[45836]_ ;
  assign \new_[45841]_  = A202 & A201;
  assign \new_[45842]_  = ~A200 & \new_[45841]_ ;
  assign \new_[45843]_  = \new_[45842]_  & \new_[45837]_ ;
  assign \new_[45847]_  = ~A298 & A269;
  assign \new_[45848]_  = ~A267 & \new_[45847]_ ;
  assign \new_[45851]_  = ~A300 & A299;
  assign \new_[45854]_  = ~A302 & ~A301;
  assign \new_[45855]_  = \new_[45854]_  & \new_[45851]_ ;
  assign \new_[45856]_  = \new_[45855]_  & \new_[45848]_ ;
  assign \new_[45860]_  = A199 & ~A168;
  assign \new_[45861]_  = ~A170 & \new_[45860]_ ;
  assign \new_[45865]_  = A202 & A201;
  assign \new_[45866]_  = ~A200 & \new_[45865]_ ;
  assign \new_[45867]_  = \new_[45866]_  & \new_[45861]_ ;
  assign \new_[45871]_  = A298 & A266;
  assign \new_[45872]_  = A265 & \new_[45871]_ ;
  assign \new_[45875]_  = ~A300 & ~A299;
  assign \new_[45878]_  = ~A302 & ~A301;
  assign \new_[45879]_  = \new_[45878]_  & \new_[45875]_ ;
  assign \new_[45880]_  = \new_[45879]_  & \new_[45872]_ ;
  assign \new_[45884]_  = A199 & ~A168;
  assign \new_[45885]_  = ~A170 & \new_[45884]_ ;
  assign \new_[45889]_  = A202 & A201;
  assign \new_[45890]_  = ~A200 & \new_[45889]_ ;
  assign \new_[45891]_  = \new_[45890]_  & \new_[45885]_ ;
  assign \new_[45895]_  = ~A298 & A266;
  assign \new_[45896]_  = A265 & \new_[45895]_ ;
  assign \new_[45899]_  = ~A300 & A299;
  assign \new_[45902]_  = ~A302 & ~A301;
  assign \new_[45903]_  = \new_[45902]_  & \new_[45899]_ ;
  assign \new_[45904]_  = \new_[45903]_  & \new_[45896]_ ;
  assign \new_[45908]_  = A199 & ~A168;
  assign \new_[45909]_  = ~A170 & \new_[45908]_ ;
  assign \new_[45913]_  = A202 & A201;
  assign \new_[45914]_  = ~A200 & \new_[45913]_ ;
  assign \new_[45915]_  = \new_[45914]_  & \new_[45909]_ ;
  assign \new_[45919]_  = A298 & ~A266;
  assign \new_[45920]_  = ~A265 & \new_[45919]_ ;
  assign \new_[45923]_  = ~A300 & ~A299;
  assign \new_[45926]_  = ~A302 & ~A301;
  assign \new_[45927]_  = \new_[45926]_  & \new_[45923]_ ;
  assign \new_[45928]_  = \new_[45927]_  & \new_[45920]_ ;
  assign \new_[45932]_  = A199 & ~A168;
  assign \new_[45933]_  = ~A170 & \new_[45932]_ ;
  assign \new_[45937]_  = A202 & A201;
  assign \new_[45938]_  = ~A200 & \new_[45937]_ ;
  assign \new_[45939]_  = \new_[45938]_  & \new_[45933]_ ;
  assign \new_[45943]_  = ~A298 & ~A266;
  assign \new_[45944]_  = ~A265 & \new_[45943]_ ;
  assign \new_[45947]_  = ~A300 & A299;
  assign \new_[45950]_  = ~A302 & ~A301;
  assign \new_[45951]_  = \new_[45950]_  & \new_[45947]_ ;
  assign \new_[45952]_  = \new_[45951]_  & \new_[45944]_ ;
  assign \new_[45956]_  = A199 & ~A168;
  assign \new_[45957]_  = ~A170 & \new_[45956]_ ;
  assign \new_[45961]_  = A203 & A201;
  assign \new_[45962]_  = ~A200 & \new_[45961]_ ;
  assign \new_[45963]_  = \new_[45962]_  & \new_[45957]_ ;
  assign \new_[45967]_  = ~A269 & ~A268;
  assign \new_[45968]_  = A267 & \new_[45967]_ ;
  assign \new_[45971]_  = ~A299 & A298;
  assign \new_[45974]_  = A301 & A300;
  assign \new_[45975]_  = \new_[45974]_  & \new_[45971]_ ;
  assign \new_[45976]_  = \new_[45975]_  & \new_[45968]_ ;
  assign \new_[45980]_  = A199 & ~A168;
  assign \new_[45981]_  = ~A170 & \new_[45980]_ ;
  assign \new_[45985]_  = A203 & A201;
  assign \new_[45986]_  = ~A200 & \new_[45985]_ ;
  assign \new_[45987]_  = \new_[45986]_  & \new_[45981]_ ;
  assign \new_[45991]_  = ~A269 & ~A268;
  assign \new_[45992]_  = A267 & \new_[45991]_ ;
  assign \new_[45995]_  = ~A299 & A298;
  assign \new_[45998]_  = A302 & A300;
  assign \new_[45999]_  = \new_[45998]_  & \new_[45995]_ ;
  assign \new_[46000]_  = \new_[45999]_  & \new_[45992]_ ;
  assign \new_[46004]_  = A199 & ~A168;
  assign \new_[46005]_  = ~A170 & \new_[46004]_ ;
  assign \new_[46009]_  = A203 & A201;
  assign \new_[46010]_  = ~A200 & \new_[46009]_ ;
  assign \new_[46011]_  = \new_[46010]_  & \new_[46005]_ ;
  assign \new_[46015]_  = ~A269 & ~A268;
  assign \new_[46016]_  = A267 & \new_[46015]_ ;
  assign \new_[46019]_  = A299 & ~A298;
  assign \new_[46022]_  = A301 & A300;
  assign \new_[46023]_  = \new_[46022]_  & \new_[46019]_ ;
  assign \new_[46024]_  = \new_[46023]_  & \new_[46016]_ ;
  assign \new_[46028]_  = A199 & ~A168;
  assign \new_[46029]_  = ~A170 & \new_[46028]_ ;
  assign \new_[46033]_  = A203 & A201;
  assign \new_[46034]_  = ~A200 & \new_[46033]_ ;
  assign \new_[46035]_  = \new_[46034]_  & \new_[46029]_ ;
  assign \new_[46039]_  = ~A269 & ~A268;
  assign \new_[46040]_  = A267 & \new_[46039]_ ;
  assign \new_[46043]_  = A299 & ~A298;
  assign \new_[46046]_  = A302 & A300;
  assign \new_[46047]_  = \new_[46046]_  & \new_[46043]_ ;
  assign \new_[46048]_  = \new_[46047]_  & \new_[46040]_ ;
  assign \new_[46052]_  = A199 & ~A168;
  assign \new_[46053]_  = ~A170 & \new_[46052]_ ;
  assign \new_[46057]_  = A203 & A201;
  assign \new_[46058]_  = ~A200 & \new_[46057]_ ;
  assign \new_[46059]_  = \new_[46058]_  & \new_[46053]_ ;
  assign \new_[46063]_  = A298 & A268;
  assign \new_[46064]_  = ~A267 & \new_[46063]_ ;
  assign \new_[46067]_  = ~A300 & ~A299;
  assign \new_[46070]_  = ~A302 & ~A301;
  assign \new_[46071]_  = \new_[46070]_  & \new_[46067]_ ;
  assign \new_[46072]_  = \new_[46071]_  & \new_[46064]_ ;
  assign \new_[46076]_  = A199 & ~A168;
  assign \new_[46077]_  = ~A170 & \new_[46076]_ ;
  assign \new_[46081]_  = A203 & A201;
  assign \new_[46082]_  = ~A200 & \new_[46081]_ ;
  assign \new_[46083]_  = \new_[46082]_  & \new_[46077]_ ;
  assign \new_[46087]_  = ~A298 & A268;
  assign \new_[46088]_  = ~A267 & \new_[46087]_ ;
  assign \new_[46091]_  = ~A300 & A299;
  assign \new_[46094]_  = ~A302 & ~A301;
  assign \new_[46095]_  = \new_[46094]_  & \new_[46091]_ ;
  assign \new_[46096]_  = \new_[46095]_  & \new_[46088]_ ;
  assign \new_[46100]_  = A199 & ~A168;
  assign \new_[46101]_  = ~A170 & \new_[46100]_ ;
  assign \new_[46105]_  = A203 & A201;
  assign \new_[46106]_  = ~A200 & \new_[46105]_ ;
  assign \new_[46107]_  = \new_[46106]_  & \new_[46101]_ ;
  assign \new_[46111]_  = A298 & A269;
  assign \new_[46112]_  = ~A267 & \new_[46111]_ ;
  assign \new_[46115]_  = ~A300 & ~A299;
  assign \new_[46118]_  = ~A302 & ~A301;
  assign \new_[46119]_  = \new_[46118]_  & \new_[46115]_ ;
  assign \new_[46120]_  = \new_[46119]_  & \new_[46112]_ ;
  assign \new_[46124]_  = A199 & ~A168;
  assign \new_[46125]_  = ~A170 & \new_[46124]_ ;
  assign \new_[46129]_  = A203 & A201;
  assign \new_[46130]_  = ~A200 & \new_[46129]_ ;
  assign \new_[46131]_  = \new_[46130]_  & \new_[46125]_ ;
  assign \new_[46135]_  = ~A298 & A269;
  assign \new_[46136]_  = ~A267 & \new_[46135]_ ;
  assign \new_[46139]_  = ~A300 & A299;
  assign \new_[46142]_  = ~A302 & ~A301;
  assign \new_[46143]_  = \new_[46142]_  & \new_[46139]_ ;
  assign \new_[46144]_  = \new_[46143]_  & \new_[46136]_ ;
  assign \new_[46148]_  = A199 & ~A168;
  assign \new_[46149]_  = ~A170 & \new_[46148]_ ;
  assign \new_[46153]_  = A203 & A201;
  assign \new_[46154]_  = ~A200 & \new_[46153]_ ;
  assign \new_[46155]_  = \new_[46154]_  & \new_[46149]_ ;
  assign \new_[46159]_  = A298 & A266;
  assign \new_[46160]_  = A265 & \new_[46159]_ ;
  assign \new_[46163]_  = ~A300 & ~A299;
  assign \new_[46166]_  = ~A302 & ~A301;
  assign \new_[46167]_  = \new_[46166]_  & \new_[46163]_ ;
  assign \new_[46168]_  = \new_[46167]_  & \new_[46160]_ ;
  assign \new_[46172]_  = A199 & ~A168;
  assign \new_[46173]_  = ~A170 & \new_[46172]_ ;
  assign \new_[46177]_  = A203 & A201;
  assign \new_[46178]_  = ~A200 & \new_[46177]_ ;
  assign \new_[46179]_  = \new_[46178]_  & \new_[46173]_ ;
  assign \new_[46183]_  = ~A298 & A266;
  assign \new_[46184]_  = A265 & \new_[46183]_ ;
  assign \new_[46187]_  = ~A300 & A299;
  assign \new_[46190]_  = ~A302 & ~A301;
  assign \new_[46191]_  = \new_[46190]_  & \new_[46187]_ ;
  assign \new_[46192]_  = \new_[46191]_  & \new_[46184]_ ;
  assign \new_[46196]_  = A199 & ~A168;
  assign \new_[46197]_  = ~A170 & \new_[46196]_ ;
  assign \new_[46201]_  = A203 & A201;
  assign \new_[46202]_  = ~A200 & \new_[46201]_ ;
  assign \new_[46203]_  = \new_[46202]_  & \new_[46197]_ ;
  assign \new_[46207]_  = A298 & ~A266;
  assign \new_[46208]_  = ~A265 & \new_[46207]_ ;
  assign \new_[46211]_  = ~A300 & ~A299;
  assign \new_[46214]_  = ~A302 & ~A301;
  assign \new_[46215]_  = \new_[46214]_  & \new_[46211]_ ;
  assign \new_[46216]_  = \new_[46215]_  & \new_[46208]_ ;
  assign \new_[46220]_  = A199 & ~A168;
  assign \new_[46221]_  = ~A170 & \new_[46220]_ ;
  assign \new_[46225]_  = A203 & A201;
  assign \new_[46226]_  = ~A200 & \new_[46225]_ ;
  assign \new_[46227]_  = \new_[46226]_  & \new_[46221]_ ;
  assign \new_[46231]_  = ~A298 & ~A266;
  assign \new_[46232]_  = ~A265 & \new_[46231]_ ;
  assign \new_[46235]_  = ~A300 & A299;
  assign \new_[46238]_  = ~A302 & ~A301;
  assign \new_[46239]_  = \new_[46238]_  & \new_[46235]_ ;
  assign \new_[46240]_  = \new_[46239]_  & \new_[46232]_ ;
  assign \new_[46244]_  = A199 & ~A168;
  assign \new_[46245]_  = ~A170 & \new_[46244]_ ;
  assign \new_[46249]_  = ~A202 & ~A201;
  assign \new_[46250]_  = ~A200 & \new_[46249]_ ;
  assign \new_[46251]_  = \new_[46250]_  & \new_[46245]_ ;
  assign \new_[46255]_  = A268 & ~A267;
  assign \new_[46256]_  = ~A203 & \new_[46255]_ ;
  assign \new_[46259]_  = ~A299 & A298;
  assign \new_[46262]_  = A301 & A300;
  assign \new_[46263]_  = \new_[46262]_  & \new_[46259]_ ;
  assign \new_[46264]_  = \new_[46263]_  & \new_[46256]_ ;
  assign \new_[46268]_  = A199 & ~A168;
  assign \new_[46269]_  = ~A170 & \new_[46268]_ ;
  assign \new_[46273]_  = ~A202 & ~A201;
  assign \new_[46274]_  = ~A200 & \new_[46273]_ ;
  assign \new_[46275]_  = \new_[46274]_  & \new_[46269]_ ;
  assign \new_[46279]_  = A268 & ~A267;
  assign \new_[46280]_  = ~A203 & \new_[46279]_ ;
  assign \new_[46283]_  = ~A299 & A298;
  assign \new_[46286]_  = A302 & A300;
  assign \new_[46287]_  = \new_[46286]_  & \new_[46283]_ ;
  assign \new_[46288]_  = \new_[46287]_  & \new_[46280]_ ;
  assign \new_[46292]_  = A199 & ~A168;
  assign \new_[46293]_  = ~A170 & \new_[46292]_ ;
  assign \new_[46297]_  = ~A202 & ~A201;
  assign \new_[46298]_  = ~A200 & \new_[46297]_ ;
  assign \new_[46299]_  = \new_[46298]_  & \new_[46293]_ ;
  assign \new_[46303]_  = A268 & ~A267;
  assign \new_[46304]_  = ~A203 & \new_[46303]_ ;
  assign \new_[46307]_  = A299 & ~A298;
  assign \new_[46310]_  = A301 & A300;
  assign \new_[46311]_  = \new_[46310]_  & \new_[46307]_ ;
  assign \new_[46312]_  = \new_[46311]_  & \new_[46304]_ ;
  assign \new_[46316]_  = A199 & ~A168;
  assign \new_[46317]_  = ~A170 & \new_[46316]_ ;
  assign \new_[46321]_  = ~A202 & ~A201;
  assign \new_[46322]_  = ~A200 & \new_[46321]_ ;
  assign \new_[46323]_  = \new_[46322]_  & \new_[46317]_ ;
  assign \new_[46327]_  = A268 & ~A267;
  assign \new_[46328]_  = ~A203 & \new_[46327]_ ;
  assign \new_[46331]_  = A299 & ~A298;
  assign \new_[46334]_  = A302 & A300;
  assign \new_[46335]_  = \new_[46334]_  & \new_[46331]_ ;
  assign \new_[46336]_  = \new_[46335]_  & \new_[46328]_ ;
  assign \new_[46340]_  = A199 & ~A168;
  assign \new_[46341]_  = ~A170 & \new_[46340]_ ;
  assign \new_[46345]_  = ~A202 & ~A201;
  assign \new_[46346]_  = ~A200 & \new_[46345]_ ;
  assign \new_[46347]_  = \new_[46346]_  & \new_[46341]_ ;
  assign \new_[46351]_  = A269 & ~A267;
  assign \new_[46352]_  = ~A203 & \new_[46351]_ ;
  assign \new_[46355]_  = ~A299 & A298;
  assign \new_[46358]_  = A301 & A300;
  assign \new_[46359]_  = \new_[46358]_  & \new_[46355]_ ;
  assign \new_[46360]_  = \new_[46359]_  & \new_[46352]_ ;
  assign \new_[46364]_  = A199 & ~A168;
  assign \new_[46365]_  = ~A170 & \new_[46364]_ ;
  assign \new_[46369]_  = ~A202 & ~A201;
  assign \new_[46370]_  = ~A200 & \new_[46369]_ ;
  assign \new_[46371]_  = \new_[46370]_  & \new_[46365]_ ;
  assign \new_[46375]_  = A269 & ~A267;
  assign \new_[46376]_  = ~A203 & \new_[46375]_ ;
  assign \new_[46379]_  = ~A299 & A298;
  assign \new_[46382]_  = A302 & A300;
  assign \new_[46383]_  = \new_[46382]_  & \new_[46379]_ ;
  assign \new_[46384]_  = \new_[46383]_  & \new_[46376]_ ;
  assign \new_[46388]_  = A199 & ~A168;
  assign \new_[46389]_  = ~A170 & \new_[46388]_ ;
  assign \new_[46393]_  = ~A202 & ~A201;
  assign \new_[46394]_  = ~A200 & \new_[46393]_ ;
  assign \new_[46395]_  = \new_[46394]_  & \new_[46389]_ ;
  assign \new_[46399]_  = A269 & ~A267;
  assign \new_[46400]_  = ~A203 & \new_[46399]_ ;
  assign \new_[46403]_  = A299 & ~A298;
  assign \new_[46406]_  = A301 & A300;
  assign \new_[46407]_  = \new_[46406]_  & \new_[46403]_ ;
  assign \new_[46408]_  = \new_[46407]_  & \new_[46400]_ ;
  assign \new_[46412]_  = A199 & ~A168;
  assign \new_[46413]_  = ~A170 & \new_[46412]_ ;
  assign \new_[46417]_  = ~A202 & ~A201;
  assign \new_[46418]_  = ~A200 & \new_[46417]_ ;
  assign \new_[46419]_  = \new_[46418]_  & \new_[46413]_ ;
  assign \new_[46423]_  = A269 & ~A267;
  assign \new_[46424]_  = ~A203 & \new_[46423]_ ;
  assign \new_[46427]_  = A299 & ~A298;
  assign \new_[46430]_  = A302 & A300;
  assign \new_[46431]_  = \new_[46430]_  & \new_[46427]_ ;
  assign \new_[46432]_  = \new_[46431]_  & \new_[46424]_ ;
  assign \new_[46436]_  = A199 & ~A168;
  assign \new_[46437]_  = ~A170 & \new_[46436]_ ;
  assign \new_[46441]_  = ~A202 & ~A201;
  assign \new_[46442]_  = ~A200 & \new_[46441]_ ;
  assign \new_[46443]_  = \new_[46442]_  & \new_[46437]_ ;
  assign \new_[46447]_  = A266 & A265;
  assign \new_[46448]_  = ~A203 & \new_[46447]_ ;
  assign \new_[46451]_  = ~A299 & A298;
  assign \new_[46454]_  = A301 & A300;
  assign \new_[46455]_  = \new_[46454]_  & \new_[46451]_ ;
  assign \new_[46456]_  = \new_[46455]_  & \new_[46448]_ ;
  assign \new_[46460]_  = A199 & ~A168;
  assign \new_[46461]_  = ~A170 & \new_[46460]_ ;
  assign \new_[46465]_  = ~A202 & ~A201;
  assign \new_[46466]_  = ~A200 & \new_[46465]_ ;
  assign \new_[46467]_  = \new_[46466]_  & \new_[46461]_ ;
  assign \new_[46471]_  = A266 & A265;
  assign \new_[46472]_  = ~A203 & \new_[46471]_ ;
  assign \new_[46475]_  = ~A299 & A298;
  assign \new_[46478]_  = A302 & A300;
  assign \new_[46479]_  = \new_[46478]_  & \new_[46475]_ ;
  assign \new_[46480]_  = \new_[46479]_  & \new_[46472]_ ;
  assign \new_[46484]_  = A199 & ~A168;
  assign \new_[46485]_  = ~A170 & \new_[46484]_ ;
  assign \new_[46489]_  = ~A202 & ~A201;
  assign \new_[46490]_  = ~A200 & \new_[46489]_ ;
  assign \new_[46491]_  = \new_[46490]_  & \new_[46485]_ ;
  assign \new_[46495]_  = A266 & A265;
  assign \new_[46496]_  = ~A203 & \new_[46495]_ ;
  assign \new_[46499]_  = A299 & ~A298;
  assign \new_[46502]_  = A301 & A300;
  assign \new_[46503]_  = \new_[46502]_  & \new_[46499]_ ;
  assign \new_[46504]_  = \new_[46503]_  & \new_[46496]_ ;
  assign \new_[46508]_  = A199 & ~A168;
  assign \new_[46509]_  = ~A170 & \new_[46508]_ ;
  assign \new_[46513]_  = ~A202 & ~A201;
  assign \new_[46514]_  = ~A200 & \new_[46513]_ ;
  assign \new_[46515]_  = \new_[46514]_  & \new_[46509]_ ;
  assign \new_[46519]_  = A266 & A265;
  assign \new_[46520]_  = ~A203 & \new_[46519]_ ;
  assign \new_[46523]_  = A299 & ~A298;
  assign \new_[46526]_  = A302 & A300;
  assign \new_[46527]_  = \new_[46526]_  & \new_[46523]_ ;
  assign \new_[46528]_  = \new_[46527]_  & \new_[46520]_ ;
  assign \new_[46532]_  = A199 & ~A168;
  assign \new_[46533]_  = ~A170 & \new_[46532]_ ;
  assign \new_[46537]_  = ~A202 & ~A201;
  assign \new_[46538]_  = ~A200 & \new_[46537]_ ;
  assign \new_[46539]_  = \new_[46538]_  & \new_[46533]_ ;
  assign \new_[46543]_  = ~A266 & ~A265;
  assign \new_[46544]_  = ~A203 & \new_[46543]_ ;
  assign \new_[46547]_  = ~A299 & A298;
  assign \new_[46550]_  = A301 & A300;
  assign \new_[46551]_  = \new_[46550]_  & \new_[46547]_ ;
  assign \new_[46552]_  = \new_[46551]_  & \new_[46544]_ ;
  assign \new_[46556]_  = A199 & ~A168;
  assign \new_[46557]_  = ~A170 & \new_[46556]_ ;
  assign \new_[46561]_  = ~A202 & ~A201;
  assign \new_[46562]_  = ~A200 & \new_[46561]_ ;
  assign \new_[46563]_  = \new_[46562]_  & \new_[46557]_ ;
  assign \new_[46567]_  = ~A266 & ~A265;
  assign \new_[46568]_  = ~A203 & \new_[46567]_ ;
  assign \new_[46571]_  = ~A299 & A298;
  assign \new_[46574]_  = A302 & A300;
  assign \new_[46575]_  = \new_[46574]_  & \new_[46571]_ ;
  assign \new_[46576]_  = \new_[46575]_  & \new_[46568]_ ;
  assign \new_[46580]_  = A199 & ~A168;
  assign \new_[46581]_  = ~A170 & \new_[46580]_ ;
  assign \new_[46585]_  = ~A202 & ~A201;
  assign \new_[46586]_  = ~A200 & \new_[46585]_ ;
  assign \new_[46587]_  = \new_[46586]_  & \new_[46581]_ ;
  assign \new_[46591]_  = ~A266 & ~A265;
  assign \new_[46592]_  = ~A203 & \new_[46591]_ ;
  assign \new_[46595]_  = A299 & ~A298;
  assign \new_[46598]_  = A301 & A300;
  assign \new_[46599]_  = \new_[46598]_  & \new_[46595]_ ;
  assign \new_[46600]_  = \new_[46599]_  & \new_[46592]_ ;
  assign \new_[46604]_  = A199 & ~A168;
  assign \new_[46605]_  = ~A170 & \new_[46604]_ ;
  assign \new_[46609]_  = ~A202 & ~A201;
  assign \new_[46610]_  = ~A200 & \new_[46609]_ ;
  assign \new_[46611]_  = \new_[46610]_  & \new_[46605]_ ;
  assign \new_[46615]_  = ~A266 & ~A265;
  assign \new_[46616]_  = ~A203 & \new_[46615]_ ;
  assign \new_[46619]_  = A299 & ~A298;
  assign \new_[46622]_  = A302 & A300;
  assign \new_[46623]_  = \new_[46622]_  & \new_[46619]_ ;
  assign \new_[46624]_  = \new_[46623]_  & \new_[46616]_ ;
  assign \new_[46628]_  = A167 & A168;
  assign \new_[46629]_  = A169 & \new_[46628]_ ;
  assign \new_[46633]_  = ~A202 & A201;
  assign \new_[46634]_  = ~A166 & \new_[46633]_ ;
  assign \new_[46635]_  = \new_[46634]_  & \new_[46629]_ ;
  assign \new_[46639]_  = A268 & ~A267;
  assign \new_[46640]_  = ~A203 & \new_[46639]_ ;
  assign \new_[46643]_  = ~A299 & A298;
  assign \new_[46646]_  = A301 & A300;
  assign \new_[46647]_  = \new_[46646]_  & \new_[46643]_ ;
  assign \new_[46648]_  = \new_[46647]_  & \new_[46640]_ ;
  assign \new_[46652]_  = A167 & A168;
  assign \new_[46653]_  = A169 & \new_[46652]_ ;
  assign \new_[46657]_  = ~A202 & A201;
  assign \new_[46658]_  = ~A166 & \new_[46657]_ ;
  assign \new_[46659]_  = \new_[46658]_  & \new_[46653]_ ;
  assign \new_[46663]_  = A268 & ~A267;
  assign \new_[46664]_  = ~A203 & \new_[46663]_ ;
  assign \new_[46667]_  = ~A299 & A298;
  assign \new_[46670]_  = A302 & A300;
  assign \new_[46671]_  = \new_[46670]_  & \new_[46667]_ ;
  assign \new_[46672]_  = \new_[46671]_  & \new_[46664]_ ;
  assign \new_[46676]_  = A167 & A168;
  assign \new_[46677]_  = A169 & \new_[46676]_ ;
  assign \new_[46681]_  = ~A202 & A201;
  assign \new_[46682]_  = ~A166 & \new_[46681]_ ;
  assign \new_[46683]_  = \new_[46682]_  & \new_[46677]_ ;
  assign \new_[46687]_  = A268 & ~A267;
  assign \new_[46688]_  = ~A203 & \new_[46687]_ ;
  assign \new_[46691]_  = A299 & ~A298;
  assign \new_[46694]_  = A301 & A300;
  assign \new_[46695]_  = \new_[46694]_  & \new_[46691]_ ;
  assign \new_[46696]_  = \new_[46695]_  & \new_[46688]_ ;
  assign \new_[46700]_  = A167 & A168;
  assign \new_[46701]_  = A169 & \new_[46700]_ ;
  assign \new_[46705]_  = ~A202 & A201;
  assign \new_[46706]_  = ~A166 & \new_[46705]_ ;
  assign \new_[46707]_  = \new_[46706]_  & \new_[46701]_ ;
  assign \new_[46711]_  = A268 & ~A267;
  assign \new_[46712]_  = ~A203 & \new_[46711]_ ;
  assign \new_[46715]_  = A299 & ~A298;
  assign \new_[46718]_  = A302 & A300;
  assign \new_[46719]_  = \new_[46718]_  & \new_[46715]_ ;
  assign \new_[46720]_  = \new_[46719]_  & \new_[46712]_ ;
  assign \new_[46724]_  = A167 & A168;
  assign \new_[46725]_  = A169 & \new_[46724]_ ;
  assign \new_[46729]_  = ~A202 & A201;
  assign \new_[46730]_  = ~A166 & \new_[46729]_ ;
  assign \new_[46731]_  = \new_[46730]_  & \new_[46725]_ ;
  assign \new_[46735]_  = A269 & ~A267;
  assign \new_[46736]_  = ~A203 & \new_[46735]_ ;
  assign \new_[46739]_  = ~A299 & A298;
  assign \new_[46742]_  = A301 & A300;
  assign \new_[46743]_  = \new_[46742]_  & \new_[46739]_ ;
  assign \new_[46744]_  = \new_[46743]_  & \new_[46736]_ ;
  assign \new_[46748]_  = A167 & A168;
  assign \new_[46749]_  = A169 & \new_[46748]_ ;
  assign \new_[46753]_  = ~A202 & A201;
  assign \new_[46754]_  = ~A166 & \new_[46753]_ ;
  assign \new_[46755]_  = \new_[46754]_  & \new_[46749]_ ;
  assign \new_[46759]_  = A269 & ~A267;
  assign \new_[46760]_  = ~A203 & \new_[46759]_ ;
  assign \new_[46763]_  = ~A299 & A298;
  assign \new_[46766]_  = A302 & A300;
  assign \new_[46767]_  = \new_[46766]_  & \new_[46763]_ ;
  assign \new_[46768]_  = \new_[46767]_  & \new_[46760]_ ;
  assign \new_[46772]_  = A167 & A168;
  assign \new_[46773]_  = A169 & \new_[46772]_ ;
  assign \new_[46777]_  = ~A202 & A201;
  assign \new_[46778]_  = ~A166 & \new_[46777]_ ;
  assign \new_[46779]_  = \new_[46778]_  & \new_[46773]_ ;
  assign \new_[46783]_  = A269 & ~A267;
  assign \new_[46784]_  = ~A203 & \new_[46783]_ ;
  assign \new_[46787]_  = A299 & ~A298;
  assign \new_[46790]_  = A301 & A300;
  assign \new_[46791]_  = \new_[46790]_  & \new_[46787]_ ;
  assign \new_[46792]_  = \new_[46791]_  & \new_[46784]_ ;
  assign \new_[46796]_  = A167 & A168;
  assign \new_[46797]_  = A169 & \new_[46796]_ ;
  assign \new_[46801]_  = ~A202 & A201;
  assign \new_[46802]_  = ~A166 & \new_[46801]_ ;
  assign \new_[46803]_  = \new_[46802]_  & \new_[46797]_ ;
  assign \new_[46807]_  = A269 & ~A267;
  assign \new_[46808]_  = ~A203 & \new_[46807]_ ;
  assign \new_[46811]_  = A299 & ~A298;
  assign \new_[46814]_  = A302 & A300;
  assign \new_[46815]_  = \new_[46814]_  & \new_[46811]_ ;
  assign \new_[46816]_  = \new_[46815]_  & \new_[46808]_ ;
  assign \new_[46820]_  = A167 & A168;
  assign \new_[46821]_  = A169 & \new_[46820]_ ;
  assign \new_[46825]_  = ~A202 & A201;
  assign \new_[46826]_  = ~A166 & \new_[46825]_ ;
  assign \new_[46827]_  = \new_[46826]_  & \new_[46821]_ ;
  assign \new_[46831]_  = A266 & A265;
  assign \new_[46832]_  = ~A203 & \new_[46831]_ ;
  assign \new_[46835]_  = ~A299 & A298;
  assign \new_[46838]_  = A301 & A300;
  assign \new_[46839]_  = \new_[46838]_  & \new_[46835]_ ;
  assign \new_[46840]_  = \new_[46839]_  & \new_[46832]_ ;
  assign \new_[46844]_  = A167 & A168;
  assign \new_[46845]_  = A169 & \new_[46844]_ ;
  assign \new_[46849]_  = ~A202 & A201;
  assign \new_[46850]_  = ~A166 & \new_[46849]_ ;
  assign \new_[46851]_  = \new_[46850]_  & \new_[46845]_ ;
  assign \new_[46855]_  = A266 & A265;
  assign \new_[46856]_  = ~A203 & \new_[46855]_ ;
  assign \new_[46859]_  = ~A299 & A298;
  assign \new_[46862]_  = A302 & A300;
  assign \new_[46863]_  = \new_[46862]_  & \new_[46859]_ ;
  assign \new_[46864]_  = \new_[46863]_  & \new_[46856]_ ;
  assign \new_[46868]_  = A167 & A168;
  assign \new_[46869]_  = A169 & \new_[46868]_ ;
  assign \new_[46873]_  = ~A202 & A201;
  assign \new_[46874]_  = ~A166 & \new_[46873]_ ;
  assign \new_[46875]_  = \new_[46874]_  & \new_[46869]_ ;
  assign \new_[46879]_  = A266 & A265;
  assign \new_[46880]_  = ~A203 & \new_[46879]_ ;
  assign \new_[46883]_  = A299 & ~A298;
  assign \new_[46886]_  = A301 & A300;
  assign \new_[46887]_  = \new_[46886]_  & \new_[46883]_ ;
  assign \new_[46888]_  = \new_[46887]_  & \new_[46880]_ ;
  assign \new_[46892]_  = A167 & A168;
  assign \new_[46893]_  = A169 & \new_[46892]_ ;
  assign \new_[46897]_  = ~A202 & A201;
  assign \new_[46898]_  = ~A166 & \new_[46897]_ ;
  assign \new_[46899]_  = \new_[46898]_  & \new_[46893]_ ;
  assign \new_[46903]_  = A266 & A265;
  assign \new_[46904]_  = ~A203 & \new_[46903]_ ;
  assign \new_[46907]_  = A299 & ~A298;
  assign \new_[46910]_  = A302 & A300;
  assign \new_[46911]_  = \new_[46910]_  & \new_[46907]_ ;
  assign \new_[46912]_  = \new_[46911]_  & \new_[46904]_ ;
  assign \new_[46916]_  = A167 & A168;
  assign \new_[46917]_  = A169 & \new_[46916]_ ;
  assign \new_[46921]_  = ~A202 & A201;
  assign \new_[46922]_  = ~A166 & \new_[46921]_ ;
  assign \new_[46923]_  = \new_[46922]_  & \new_[46917]_ ;
  assign \new_[46927]_  = ~A266 & ~A265;
  assign \new_[46928]_  = ~A203 & \new_[46927]_ ;
  assign \new_[46931]_  = ~A299 & A298;
  assign \new_[46934]_  = A301 & A300;
  assign \new_[46935]_  = \new_[46934]_  & \new_[46931]_ ;
  assign \new_[46936]_  = \new_[46935]_  & \new_[46928]_ ;
  assign \new_[46940]_  = A167 & A168;
  assign \new_[46941]_  = A169 & \new_[46940]_ ;
  assign \new_[46945]_  = ~A202 & A201;
  assign \new_[46946]_  = ~A166 & \new_[46945]_ ;
  assign \new_[46947]_  = \new_[46946]_  & \new_[46941]_ ;
  assign \new_[46951]_  = ~A266 & ~A265;
  assign \new_[46952]_  = ~A203 & \new_[46951]_ ;
  assign \new_[46955]_  = ~A299 & A298;
  assign \new_[46958]_  = A302 & A300;
  assign \new_[46959]_  = \new_[46958]_  & \new_[46955]_ ;
  assign \new_[46960]_  = \new_[46959]_  & \new_[46952]_ ;
  assign \new_[46964]_  = A167 & A168;
  assign \new_[46965]_  = A169 & \new_[46964]_ ;
  assign \new_[46969]_  = ~A202 & A201;
  assign \new_[46970]_  = ~A166 & \new_[46969]_ ;
  assign \new_[46971]_  = \new_[46970]_  & \new_[46965]_ ;
  assign \new_[46975]_  = ~A266 & ~A265;
  assign \new_[46976]_  = ~A203 & \new_[46975]_ ;
  assign \new_[46979]_  = A299 & ~A298;
  assign \new_[46982]_  = A301 & A300;
  assign \new_[46983]_  = \new_[46982]_  & \new_[46979]_ ;
  assign \new_[46984]_  = \new_[46983]_  & \new_[46976]_ ;
  assign \new_[46988]_  = A167 & A168;
  assign \new_[46989]_  = A169 & \new_[46988]_ ;
  assign \new_[46993]_  = ~A202 & A201;
  assign \new_[46994]_  = ~A166 & \new_[46993]_ ;
  assign \new_[46995]_  = \new_[46994]_  & \new_[46989]_ ;
  assign \new_[46999]_  = ~A266 & ~A265;
  assign \new_[47000]_  = ~A203 & \new_[46999]_ ;
  assign \new_[47003]_  = A299 & ~A298;
  assign \new_[47006]_  = A302 & A300;
  assign \new_[47007]_  = \new_[47006]_  & \new_[47003]_ ;
  assign \new_[47008]_  = \new_[47007]_  & \new_[47000]_ ;
  assign \new_[47012]_  = A167 & A168;
  assign \new_[47013]_  = A169 & \new_[47012]_ ;
  assign \new_[47017]_  = A202 & ~A201;
  assign \new_[47018]_  = ~A166 & \new_[47017]_ ;
  assign \new_[47019]_  = \new_[47018]_  & \new_[47013]_ ;
  assign \new_[47023]_  = ~A269 & ~A268;
  assign \new_[47024]_  = A267 & \new_[47023]_ ;
  assign \new_[47027]_  = ~A299 & A298;
  assign \new_[47030]_  = A301 & A300;
  assign \new_[47031]_  = \new_[47030]_  & \new_[47027]_ ;
  assign \new_[47032]_  = \new_[47031]_  & \new_[47024]_ ;
  assign \new_[47036]_  = A167 & A168;
  assign \new_[47037]_  = A169 & \new_[47036]_ ;
  assign \new_[47041]_  = A202 & ~A201;
  assign \new_[47042]_  = ~A166 & \new_[47041]_ ;
  assign \new_[47043]_  = \new_[47042]_  & \new_[47037]_ ;
  assign \new_[47047]_  = ~A269 & ~A268;
  assign \new_[47048]_  = A267 & \new_[47047]_ ;
  assign \new_[47051]_  = ~A299 & A298;
  assign \new_[47054]_  = A302 & A300;
  assign \new_[47055]_  = \new_[47054]_  & \new_[47051]_ ;
  assign \new_[47056]_  = \new_[47055]_  & \new_[47048]_ ;
  assign \new_[47060]_  = A167 & A168;
  assign \new_[47061]_  = A169 & \new_[47060]_ ;
  assign \new_[47065]_  = A202 & ~A201;
  assign \new_[47066]_  = ~A166 & \new_[47065]_ ;
  assign \new_[47067]_  = \new_[47066]_  & \new_[47061]_ ;
  assign \new_[47071]_  = ~A269 & ~A268;
  assign \new_[47072]_  = A267 & \new_[47071]_ ;
  assign \new_[47075]_  = A299 & ~A298;
  assign \new_[47078]_  = A301 & A300;
  assign \new_[47079]_  = \new_[47078]_  & \new_[47075]_ ;
  assign \new_[47080]_  = \new_[47079]_  & \new_[47072]_ ;
  assign \new_[47084]_  = A167 & A168;
  assign \new_[47085]_  = A169 & \new_[47084]_ ;
  assign \new_[47089]_  = A202 & ~A201;
  assign \new_[47090]_  = ~A166 & \new_[47089]_ ;
  assign \new_[47091]_  = \new_[47090]_  & \new_[47085]_ ;
  assign \new_[47095]_  = ~A269 & ~A268;
  assign \new_[47096]_  = A267 & \new_[47095]_ ;
  assign \new_[47099]_  = A299 & ~A298;
  assign \new_[47102]_  = A302 & A300;
  assign \new_[47103]_  = \new_[47102]_  & \new_[47099]_ ;
  assign \new_[47104]_  = \new_[47103]_  & \new_[47096]_ ;
  assign \new_[47108]_  = A167 & A168;
  assign \new_[47109]_  = A169 & \new_[47108]_ ;
  assign \new_[47113]_  = A202 & ~A201;
  assign \new_[47114]_  = ~A166 & \new_[47113]_ ;
  assign \new_[47115]_  = \new_[47114]_  & \new_[47109]_ ;
  assign \new_[47119]_  = A298 & A268;
  assign \new_[47120]_  = ~A267 & \new_[47119]_ ;
  assign \new_[47123]_  = ~A300 & ~A299;
  assign \new_[47126]_  = ~A302 & ~A301;
  assign \new_[47127]_  = \new_[47126]_  & \new_[47123]_ ;
  assign \new_[47128]_  = \new_[47127]_  & \new_[47120]_ ;
  assign \new_[47132]_  = A167 & A168;
  assign \new_[47133]_  = A169 & \new_[47132]_ ;
  assign \new_[47137]_  = A202 & ~A201;
  assign \new_[47138]_  = ~A166 & \new_[47137]_ ;
  assign \new_[47139]_  = \new_[47138]_  & \new_[47133]_ ;
  assign \new_[47143]_  = ~A298 & A268;
  assign \new_[47144]_  = ~A267 & \new_[47143]_ ;
  assign \new_[47147]_  = ~A300 & A299;
  assign \new_[47150]_  = ~A302 & ~A301;
  assign \new_[47151]_  = \new_[47150]_  & \new_[47147]_ ;
  assign \new_[47152]_  = \new_[47151]_  & \new_[47144]_ ;
  assign \new_[47156]_  = A167 & A168;
  assign \new_[47157]_  = A169 & \new_[47156]_ ;
  assign \new_[47161]_  = A202 & ~A201;
  assign \new_[47162]_  = ~A166 & \new_[47161]_ ;
  assign \new_[47163]_  = \new_[47162]_  & \new_[47157]_ ;
  assign \new_[47167]_  = A298 & A269;
  assign \new_[47168]_  = ~A267 & \new_[47167]_ ;
  assign \new_[47171]_  = ~A300 & ~A299;
  assign \new_[47174]_  = ~A302 & ~A301;
  assign \new_[47175]_  = \new_[47174]_  & \new_[47171]_ ;
  assign \new_[47176]_  = \new_[47175]_  & \new_[47168]_ ;
  assign \new_[47180]_  = A167 & A168;
  assign \new_[47181]_  = A169 & \new_[47180]_ ;
  assign \new_[47185]_  = A202 & ~A201;
  assign \new_[47186]_  = ~A166 & \new_[47185]_ ;
  assign \new_[47187]_  = \new_[47186]_  & \new_[47181]_ ;
  assign \new_[47191]_  = ~A298 & A269;
  assign \new_[47192]_  = ~A267 & \new_[47191]_ ;
  assign \new_[47195]_  = ~A300 & A299;
  assign \new_[47198]_  = ~A302 & ~A301;
  assign \new_[47199]_  = \new_[47198]_  & \new_[47195]_ ;
  assign \new_[47200]_  = \new_[47199]_  & \new_[47192]_ ;
  assign \new_[47204]_  = A167 & A168;
  assign \new_[47205]_  = A169 & \new_[47204]_ ;
  assign \new_[47209]_  = A202 & ~A201;
  assign \new_[47210]_  = ~A166 & \new_[47209]_ ;
  assign \new_[47211]_  = \new_[47210]_  & \new_[47205]_ ;
  assign \new_[47215]_  = A298 & A266;
  assign \new_[47216]_  = A265 & \new_[47215]_ ;
  assign \new_[47219]_  = ~A300 & ~A299;
  assign \new_[47222]_  = ~A302 & ~A301;
  assign \new_[47223]_  = \new_[47222]_  & \new_[47219]_ ;
  assign \new_[47224]_  = \new_[47223]_  & \new_[47216]_ ;
  assign \new_[47228]_  = A167 & A168;
  assign \new_[47229]_  = A169 & \new_[47228]_ ;
  assign \new_[47233]_  = A202 & ~A201;
  assign \new_[47234]_  = ~A166 & \new_[47233]_ ;
  assign \new_[47235]_  = \new_[47234]_  & \new_[47229]_ ;
  assign \new_[47239]_  = ~A298 & A266;
  assign \new_[47240]_  = A265 & \new_[47239]_ ;
  assign \new_[47243]_  = ~A300 & A299;
  assign \new_[47246]_  = ~A302 & ~A301;
  assign \new_[47247]_  = \new_[47246]_  & \new_[47243]_ ;
  assign \new_[47248]_  = \new_[47247]_  & \new_[47240]_ ;
  assign \new_[47252]_  = A167 & A168;
  assign \new_[47253]_  = A169 & \new_[47252]_ ;
  assign \new_[47257]_  = A202 & ~A201;
  assign \new_[47258]_  = ~A166 & \new_[47257]_ ;
  assign \new_[47259]_  = \new_[47258]_  & \new_[47253]_ ;
  assign \new_[47263]_  = A298 & ~A266;
  assign \new_[47264]_  = ~A265 & \new_[47263]_ ;
  assign \new_[47267]_  = ~A300 & ~A299;
  assign \new_[47270]_  = ~A302 & ~A301;
  assign \new_[47271]_  = \new_[47270]_  & \new_[47267]_ ;
  assign \new_[47272]_  = \new_[47271]_  & \new_[47264]_ ;
  assign \new_[47276]_  = A167 & A168;
  assign \new_[47277]_  = A169 & \new_[47276]_ ;
  assign \new_[47281]_  = A202 & ~A201;
  assign \new_[47282]_  = ~A166 & \new_[47281]_ ;
  assign \new_[47283]_  = \new_[47282]_  & \new_[47277]_ ;
  assign \new_[47287]_  = ~A298 & ~A266;
  assign \new_[47288]_  = ~A265 & \new_[47287]_ ;
  assign \new_[47291]_  = ~A300 & A299;
  assign \new_[47294]_  = ~A302 & ~A301;
  assign \new_[47295]_  = \new_[47294]_  & \new_[47291]_ ;
  assign \new_[47296]_  = \new_[47295]_  & \new_[47288]_ ;
  assign \new_[47300]_  = A167 & A168;
  assign \new_[47301]_  = A169 & \new_[47300]_ ;
  assign \new_[47305]_  = A203 & ~A201;
  assign \new_[47306]_  = ~A166 & \new_[47305]_ ;
  assign \new_[47307]_  = \new_[47306]_  & \new_[47301]_ ;
  assign \new_[47311]_  = ~A269 & ~A268;
  assign \new_[47312]_  = A267 & \new_[47311]_ ;
  assign \new_[47315]_  = ~A299 & A298;
  assign \new_[47318]_  = A301 & A300;
  assign \new_[47319]_  = \new_[47318]_  & \new_[47315]_ ;
  assign \new_[47320]_  = \new_[47319]_  & \new_[47312]_ ;
  assign \new_[47324]_  = A167 & A168;
  assign \new_[47325]_  = A169 & \new_[47324]_ ;
  assign \new_[47329]_  = A203 & ~A201;
  assign \new_[47330]_  = ~A166 & \new_[47329]_ ;
  assign \new_[47331]_  = \new_[47330]_  & \new_[47325]_ ;
  assign \new_[47335]_  = ~A269 & ~A268;
  assign \new_[47336]_  = A267 & \new_[47335]_ ;
  assign \new_[47339]_  = ~A299 & A298;
  assign \new_[47342]_  = A302 & A300;
  assign \new_[47343]_  = \new_[47342]_  & \new_[47339]_ ;
  assign \new_[47344]_  = \new_[47343]_  & \new_[47336]_ ;
  assign \new_[47348]_  = A167 & A168;
  assign \new_[47349]_  = A169 & \new_[47348]_ ;
  assign \new_[47353]_  = A203 & ~A201;
  assign \new_[47354]_  = ~A166 & \new_[47353]_ ;
  assign \new_[47355]_  = \new_[47354]_  & \new_[47349]_ ;
  assign \new_[47359]_  = ~A269 & ~A268;
  assign \new_[47360]_  = A267 & \new_[47359]_ ;
  assign \new_[47363]_  = A299 & ~A298;
  assign \new_[47366]_  = A301 & A300;
  assign \new_[47367]_  = \new_[47366]_  & \new_[47363]_ ;
  assign \new_[47368]_  = \new_[47367]_  & \new_[47360]_ ;
  assign \new_[47372]_  = A167 & A168;
  assign \new_[47373]_  = A169 & \new_[47372]_ ;
  assign \new_[47377]_  = A203 & ~A201;
  assign \new_[47378]_  = ~A166 & \new_[47377]_ ;
  assign \new_[47379]_  = \new_[47378]_  & \new_[47373]_ ;
  assign \new_[47383]_  = ~A269 & ~A268;
  assign \new_[47384]_  = A267 & \new_[47383]_ ;
  assign \new_[47387]_  = A299 & ~A298;
  assign \new_[47390]_  = A302 & A300;
  assign \new_[47391]_  = \new_[47390]_  & \new_[47387]_ ;
  assign \new_[47392]_  = \new_[47391]_  & \new_[47384]_ ;
  assign \new_[47396]_  = A167 & A168;
  assign \new_[47397]_  = A169 & \new_[47396]_ ;
  assign \new_[47401]_  = A203 & ~A201;
  assign \new_[47402]_  = ~A166 & \new_[47401]_ ;
  assign \new_[47403]_  = \new_[47402]_  & \new_[47397]_ ;
  assign \new_[47407]_  = A298 & A268;
  assign \new_[47408]_  = ~A267 & \new_[47407]_ ;
  assign \new_[47411]_  = ~A300 & ~A299;
  assign \new_[47414]_  = ~A302 & ~A301;
  assign \new_[47415]_  = \new_[47414]_  & \new_[47411]_ ;
  assign \new_[47416]_  = \new_[47415]_  & \new_[47408]_ ;
  assign \new_[47420]_  = A167 & A168;
  assign \new_[47421]_  = A169 & \new_[47420]_ ;
  assign \new_[47425]_  = A203 & ~A201;
  assign \new_[47426]_  = ~A166 & \new_[47425]_ ;
  assign \new_[47427]_  = \new_[47426]_  & \new_[47421]_ ;
  assign \new_[47431]_  = ~A298 & A268;
  assign \new_[47432]_  = ~A267 & \new_[47431]_ ;
  assign \new_[47435]_  = ~A300 & A299;
  assign \new_[47438]_  = ~A302 & ~A301;
  assign \new_[47439]_  = \new_[47438]_  & \new_[47435]_ ;
  assign \new_[47440]_  = \new_[47439]_  & \new_[47432]_ ;
  assign \new_[47444]_  = A167 & A168;
  assign \new_[47445]_  = A169 & \new_[47444]_ ;
  assign \new_[47449]_  = A203 & ~A201;
  assign \new_[47450]_  = ~A166 & \new_[47449]_ ;
  assign \new_[47451]_  = \new_[47450]_  & \new_[47445]_ ;
  assign \new_[47455]_  = A298 & A269;
  assign \new_[47456]_  = ~A267 & \new_[47455]_ ;
  assign \new_[47459]_  = ~A300 & ~A299;
  assign \new_[47462]_  = ~A302 & ~A301;
  assign \new_[47463]_  = \new_[47462]_  & \new_[47459]_ ;
  assign \new_[47464]_  = \new_[47463]_  & \new_[47456]_ ;
  assign \new_[47468]_  = A167 & A168;
  assign \new_[47469]_  = A169 & \new_[47468]_ ;
  assign \new_[47473]_  = A203 & ~A201;
  assign \new_[47474]_  = ~A166 & \new_[47473]_ ;
  assign \new_[47475]_  = \new_[47474]_  & \new_[47469]_ ;
  assign \new_[47479]_  = ~A298 & A269;
  assign \new_[47480]_  = ~A267 & \new_[47479]_ ;
  assign \new_[47483]_  = ~A300 & A299;
  assign \new_[47486]_  = ~A302 & ~A301;
  assign \new_[47487]_  = \new_[47486]_  & \new_[47483]_ ;
  assign \new_[47488]_  = \new_[47487]_  & \new_[47480]_ ;
  assign \new_[47492]_  = A167 & A168;
  assign \new_[47493]_  = A169 & \new_[47492]_ ;
  assign \new_[47497]_  = A203 & ~A201;
  assign \new_[47498]_  = ~A166 & \new_[47497]_ ;
  assign \new_[47499]_  = \new_[47498]_  & \new_[47493]_ ;
  assign \new_[47503]_  = A298 & A266;
  assign \new_[47504]_  = A265 & \new_[47503]_ ;
  assign \new_[47507]_  = ~A300 & ~A299;
  assign \new_[47510]_  = ~A302 & ~A301;
  assign \new_[47511]_  = \new_[47510]_  & \new_[47507]_ ;
  assign \new_[47512]_  = \new_[47511]_  & \new_[47504]_ ;
  assign \new_[47516]_  = A167 & A168;
  assign \new_[47517]_  = A169 & \new_[47516]_ ;
  assign \new_[47521]_  = A203 & ~A201;
  assign \new_[47522]_  = ~A166 & \new_[47521]_ ;
  assign \new_[47523]_  = \new_[47522]_  & \new_[47517]_ ;
  assign \new_[47527]_  = ~A298 & A266;
  assign \new_[47528]_  = A265 & \new_[47527]_ ;
  assign \new_[47531]_  = ~A300 & A299;
  assign \new_[47534]_  = ~A302 & ~A301;
  assign \new_[47535]_  = \new_[47534]_  & \new_[47531]_ ;
  assign \new_[47536]_  = \new_[47535]_  & \new_[47528]_ ;
  assign \new_[47540]_  = A167 & A168;
  assign \new_[47541]_  = A169 & \new_[47540]_ ;
  assign \new_[47545]_  = A203 & ~A201;
  assign \new_[47546]_  = ~A166 & \new_[47545]_ ;
  assign \new_[47547]_  = \new_[47546]_  & \new_[47541]_ ;
  assign \new_[47551]_  = A298 & ~A266;
  assign \new_[47552]_  = ~A265 & \new_[47551]_ ;
  assign \new_[47555]_  = ~A300 & ~A299;
  assign \new_[47558]_  = ~A302 & ~A301;
  assign \new_[47559]_  = \new_[47558]_  & \new_[47555]_ ;
  assign \new_[47560]_  = \new_[47559]_  & \new_[47552]_ ;
  assign \new_[47564]_  = A167 & A168;
  assign \new_[47565]_  = A169 & \new_[47564]_ ;
  assign \new_[47569]_  = A203 & ~A201;
  assign \new_[47570]_  = ~A166 & \new_[47569]_ ;
  assign \new_[47571]_  = \new_[47570]_  & \new_[47565]_ ;
  assign \new_[47575]_  = ~A298 & ~A266;
  assign \new_[47576]_  = ~A265 & \new_[47575]_ ;
  assign \new_[47579]_  = ~A300 & A299;
  assign \new_[47582]_  = ~A302 & ~A301;
  assign \new_[47583]_  = \new_[47582]_  & \new_[47579]_ ;
  assign \new_[47584]_  = \new_[47583]_  & \new_[47576]_ ;
  assign \new_[47588]_  = A167 & A168;
  assign \new_[47589]_  = A169 & \new_[47588]_ ;
  assign \new_[47593]_  = A200 & A199;
  assign \new_[47594]_  = ~A166 & \new_[47593]_ ;
  assign \new_[47595]_  = \new_[47594]_  & \new_[47589]_ ;
  assign \new_[47599]_  = ~A269 & ~A268;
  assign \new_[47600]_  = A267 & \new_[47599]_ ;
  assign \new_[47603]_  = ~A299 & A298;
  assign \new_[47606]_  = A301 & A300;
  assign \new_[47607]_  = \new_[47606]_  & \new_[47603]_ ;
  assign \new_[47608]_  = \new_[47607]_  & \new_[47600]_ ;
  assign \new_[47612]_  = A167 & A168;
  assign \new_[47613]_  = A169 & \new_[47612]_ ;
  assign \new_[47617]_  = A200 & A199;
  assign \new_[47618]_  = ~A166 & \new_[47617]_ ;
  assign \new_[47619]_  = \new_[47618]_  & \new_[47613]_ ;
  assign \new_[47623]_  = ~A269 & ~A268;
  assign \new_[47624]_  = A267 & \new_[47623]_ ;
  assign \new_[47627]_  = ~A299 & A298;
  assign \new_[47630]_  = A302 & A300;
  assign \new_[47631]_  = \new_[47630]_  & \new_[47627]_ ;
  assign \new_[47632]_  = \new_[47631]_  & \new_[47624]_ ;
  assign \new_[47636]_  = A167 & A168;
  assign \new_[47637]_  = A169 & \new_[47636]_ ;
  assign \new_[47641]_  = A200 & A199;
  assign \new_[47642]_  = ~A166 & \new_[47641]_ ;
  assign \new_[47643]_  = \new_[47642]_  & \new_[47637]_ ;
  assign \new_[47647]_  = ~A269 & ~A268;
  assign \new_[47648]_  = A267 & \new_[47647]_ ;
  assign \new_[47651]_  = A299 & ~A298;
  assign \new_[47654]_  = A301 & A300;
  assign \new_[47655]_  = \new_[47654]_  & \new_[47651]_ ;
  assign \new_[47656]_  = \new_[47655]_  & \new_[47648]_ ;
  assign \new_[47660]_  = A167 & A168;
  assign \new_[47661]_  = A169 & \new_[47660]_ ;
  assign \new_[47665]_  = A200 & A199;
  assign \new_[47666]_  = ~A166 & \new_[47665]_ ;
  assign \new_[47667]_  = \new_[47666]_  & \new_[47661]_ ;
  assign \new_[47671]_  = ~A269 & ~A268;
  assign \new_[47672]_  = A267 & \new_[47671]_ ;
  assign \new_[47675]_  = A299 & ~A298;
  assign \new_[47678]_  = A302 & A300;
  assign \new_[47679]_  = \new_[47678]_  & \new_[47675]_ ;
  assign \new_[47680]_  = \new_[47679]_  & \new_[47672]_ ;
  assign \new_[47684]_  = A167 & A168;
  assign \new_[47685]_  = A169 & \new_[47684]_ ;
  assign \new_[47689]_  = A200 & A199;
  assign \new_[47690]_  = ~A166 & \new_[47689]_ ;
  assign \new_[47691]_  = \new_[47690]_  & \new_[47685]_ ;
  assign \new_[47695]_  = A298 & A268;
  assign \new_[47696]_  = ~A267 & \new_[47695]_ ;
  assign \new_[47699]_  = ~A300 & ~A299;
  assign \new_[47702]_  = ~A302 & ~A301;
  assign \new_[47703]_  = \new_[47702]_  & \new_[47699]_ ;
  assign \new_[47704]_  = \new_[47703]_  & \new_[47696]_ ;
  assign \new_[47708]_  = A167 & A168;
  assign \new_[47709]_  = A169 & \new_[47708]_ ;
  assign \new_[47713]_  = A200 & A199;
  assign \new_[47714]_  = ~A166 & \new_[47713]_ ;
  assign \new_[47715]_  = \new_[47714]_  & \new_[47709]_ ;
  assign \new_[47719]_  = ~A298 & A268;
  assign \new_[47720]_  = ~A267 & \new_[47719]_ ;
  assign \new_[47723]_  = ~A300 & A299;
  assign \new_[47726]_  = ~A302 & ~A301;
  assign \new_[47727]_  = \new_[47726]_  & \new_[47723]_ ;
  assign \new_[47728]_  = \new_[47727]_  & \new_[47720]_ ;
  assign \new_[47732]_  = A167 & A168;
  assign \new_[47733]_  = A169 & \new_[47732]_ ;
  assign \new_[47737]_  = A200 & A199;
  assign \new_[47738]_  = ~A166 & \new_[47737]_ ;
  assign \new_[47739]_  = \new_[47738]_  & \new_[47733]_ ;
  assign \new_[47743]_  = A298 & A269;
  assign \new_[47744]_  = ~A267 & \new_[47743]_ ;
  assign \new_[47747]_  = ~A300 & ~A299;
  assign \new_[47750]_  = ~A302 & ~A301;
  assign \new_[47751]_  = \new_[47750]_  & \new_[47747]_ ;
  assign \new_[47752]_  = \new_[47751]_  & \new_[47744]_ ;
  assign \new_[47756]_  = A167 & A168;
  assign \new_[47757]_  = A169 & \new_[47756]_ ;
  assign \new_[47761]_  = A200 & A199;
  assign \new_[47762]_  = ~A166 & \new_[47761]_ ;
  assign \new_[47763]_  = \new_[47762]_  & \new_[47757]_ ;
  assign \new_[47767]_  = ~A298 & A269;
  assign \new_[47768]_  = ~A267 & \new_[47767]_ ;
  assign \new_[47771]_  = ~A300 & A299;
  assign \new_[47774]_  = ~A302 & ~A301;
  assign \new_[47775]_  = \new_[47774]_  & \new_[47771]_ ;
  assign \new_[47776]_  = \new_[47775]_  & \new_[47768]_ ;
  assign \new_[47780]_  = A167 & A168;
  assign \new_[47781]_  = A169 & \new_[47780]_ ;
  assign \new_[47785]_  = A200 & A199;
  assign \new_[47786]_  = ~A166 & \new_[47785]_ ;
  assign \new_[47787]_  = \new_[47786]_  & \new_[47781]_ ;
  assign \new_[47791]_  = A298 & A266;
  assign \new_[47792]_  = A265 & \new_[47791]_ ;
  assign \new_[47795]_  = ~A300 & ~A299;
  assign \new_[47798]_  = ~A302 & ~A301;
  assign \new_[47799]_  = \new_[47798]_  & \new_[47795]_ ;
  assign \new_[47800]_  = \new_[47799]_  & \new_[47792]_ ;
  assign \new_[47804]_  = A167 & A168;
  assign \new_[47805]_  = A169 & \new_[47804]_ ;
  assign \new_[47809]_  = A200 & A199;
  assign \new_[47810]_  = ~A166 & \new_[47809]_ ;
  assign \new_[47811]_  = \new_[47810]_  & \new_[47805]_ ;
  assign \new_[47815]_  = ~A298 & A266;
  assign \new_[47816]_  = A265 & \new_[47815]_ ;
  assign \new_[47819]_  = ~A300 & A299;
  assign \new_[47822]_  = ~A302 & ~A301;
  assign \new_[47823]_  = \new_[47822]_  & \new_[47819]_ ;
  assign \new_[47824]_  = \new_[47823]_  & \new_[47816]_ ;
  assign \new_[47828]_  = A167 & A168;
  assign \new_[47829]_  = A169 & \new_[47828]_ ;
  assign \new_[47833]_  = A200 & A199;
  assign \new_[47834]_  = ~A166 & \new_[47833]_ ;
  assign \new_[47835]_  = \new_[47834]_  & \new_[47829]_ ;
  assign \new_[47839]_  = A298 & ~A266;
  assign \new_[47840]_  = ~A265 & \new_[47839]_ ;
  assign \new_[47843]_  = ~A300 & ~A299;
  assign \new_[47846]_  = ~A302 & ~A301;
  assign \new_[47847]_  = \new_[47846]_  & \new_[47843]_ ;
  assign \new_[47848]_  = \new_[47847]_  & \new_[47840]_ ;
  assign \new_[47852]_  = A167 & A168;
  assign \new_[47853]_  = A169 & \new_[47852]_ ;
  assign \new_[47857]_  = A200 & A199;
  assign \new_[47858]_  = ~A166 & \new_[47857]_ ;
  assign \new_[47859]_  = \new_[47858]_  & \new_[47853]_ ;
  assign \new_[47863]_  = ~A298 & ~A266;
  assign \new_[47864]_  = ~A265 & \new_[47863]_ ;
  assign \new_[47867]_  = ~A300 & A299;
  assign \new_[47870]_  = ~A302 & ~A301;
  assign \new_[47871]_  = \new_[47870]_  & \new_[47867]_ ;
  assign \new_[47872]_  = \new_[47871]_  & \new_[47864]_ ;
  assign \new_[47876]_  = A167 & A168;
  assign \new_[47877]_  = A169 & \new_[47876]_ ;
  assign \new_[47881]_  = ~A200 & ~A199;
  assign \new_[47882]_  = ~A166 & \new_[47881]_ ;
  assign \new_[47883]_  = \new_[47882]_  & \new_[47877]_ ;
  assign \new_[47887]_  = ~A269 & ~A268;
  assign \new_[47888]_  = A267 & \new_[47887]_ ;
  assign \new_[47891]_  = ~A299 & A298;
  assign \new_[47894]_  = A301 & A300;
  assign \new_[47895]_  = \new_[47894]_  & \new_[47891]_ ;
  assign \new_[47896]_  = \new_[47895]_  & \new_[47888]_ ;
  assign \new_[47900]_  = A167 & A168;
  assign \new_[47901]_  = A169 & \new_[47900]_ ;
  assign \new_[47905]_  = ~A200 & ~A199;
  assign \new_[47906]_  = ~A166 & \new_[47905]_ ;
  assign \new_[47907]_  = \new_[47906]_  & \new_[47901]_ ;
  assign \new_[47911]_  = ~A269 & ~A268;
  assign \new_[47912]_  = A267 & \new_[47911]_ ;
  assign \new_[47915]_  = ~A299 & A298;
  assign \new_[47918]_  = A302 & A300;
  assign \new_[47919]_  = \new_[47918]_  & \new_[47915]_ ;
  assign \new_[47920]_  = \new_[47919]_  & \new_[47912]_ ;
  assign \new_[47924]_  = A167 & A168;
  assign \new_[47925]_  = A169 & \new_[47924]_ ;
  assign \new_[47929]_  = ~A200 & ~A199;
  assign \new_[47930]_  = ~A166 & \new_[47929]_ ;
  assign \new_[47931]_  = \new_[47930]_  & \new_[47925]_ ;
  assign \new_[47935]_  = ~A269 & ~A268;
  assign \new_[47936]_  = A267 & \new_[47935]_ ;
  assign \new_[47939]_  = A299 & ~A298;
  assign \new_[47942]_  = A301 & A300;
  assign \new_[47943]_  = \new_[47942]_  & \new_[47939]_ ;
  assign \new_[47944]_  = \new_[47943]_  & \new_[47936]_ ;
  assign \new_[47948]_  = A167 & A168;
  assign \new_[47949]_  = A169 & \new_[47948]_ ;
  assign \new_[47953]_  = ~A200 & ~A199;
  assign \new_[47954]_  = ~A166 & \new_[47953]_ ;
  assign \new_[47955]_  = \new_[47954]_  & \new_[47949]_ ;
  assign \new_[47959]_  = ~A269 & ~A268;
  assign \new_[47960]_  = A267 & \new_[47959]_ ;
  assign \new_[47963]_  = A299 & ~A298;
  assign \new_[47966]_  = A302 & A300;
  assign \new_[47967]_  = \new_[47966]_  & \new_[47963]_ ;
  assign \new_[47968]_  = \new_[47967]_  & \new_[47960]_ ;
  assign \new_[47972]_  = A167 & A168;
  assign \new_[47973]_  = A169 & \new_[47972]_ ;
  assign \new_[47977]_  = ~A200 & ~A199;
  assign \new_[47978]_  = ~A166 & \new_[47977]_ ;
  assign \new_[47979]_  = \new_[47978]_  & \new_[47973]_ ;
  assign \new_[47983]_  = A298 & A268;
  assign \new_[47984]_  = ~A267 & \new_[47983]_ ;
  assign \new_[47987]_  = ~A300 & ~A299;
  assign \new_[47990]_  = ~A302 & ~A301;
  assign \new_[47991]_  = \new_[47990]_  & \new_[47987]_ ;
  assign \new_[47992]_  = \new_[47991]_  & \new_[47984]_ ;
  assign \new_[47996]_  = A167 & A168;
  assign \new_[47997]_  = A169 & \new_[47996]_ ;
  assign \new_[48001]_  = ~A200 & ~A199;
  assign \new_[48002]_  = ~A166 & \new_[48001]_ ;
  assign \new_[48003]_  = \new_[48002]_  & \new_[47997]_ ;
  assign \new_[48007]_  = ~A298 & A268;
  assign \new_[48008]_  = ~A267 & \new_[48007]_ ;
  assign \new_[48011]_  = ~A300 & A299;
  assign \new_[48014]_  = ~A302 & ~A301;
  assign \new_[48015]_  = \new_[48014]_  & \new_[48011]_ ;
  assign \new_[48016]_  = \new_[48015]_  & \new_[48008]_ ;
  assign \new_[48020]_  = A167 & A168;
  assign \new_[48021]_  = A169 & \new_[48020]_ ;
  assign \new_[48025]_  = ~A200 & ~A199;
  assign \new_[48026]_  = ~A166 & \new_[48025]_ ;
  assign \new_[48027]_  = \new_[48026]_  & \new_[48021]_ ;
  assign \new_[48031]_  = A298 & A269;
  assign \new_[48032]_  = ~A267 & \new_[48031]_ ;
  assign \new_[48035]_  = ~A300 & ~A299;
  assign \new_[48038]_  = ~A302 & ~A301;
  assign \new_[48039]_  = \new_[48038]_  & \new_[48035]_ ;
  assign \new_[48040]_  = \new_[48039]_  & \new_[48032]_ ;
  assign \new_[48044]_  = A167 & A168;
  assign \new_[48045]_  = A169 & \new_[48044]_ ;
  assign \new_[48049]_  = ~A200 & ~A199;
  assign \new_[48050]_  = ~A166 & \new_[48049]_ ;
  assign \new_[48051]_  = \new_[48050]_  & \new_[48045]_ ;
  assign \new_[48055]_  = ~A298 & A269;
  assign \new_[48056]_  = ~A267 & \new_[48055]_ ;
  assign \new_[48059]_  = ~A300 & A299;
  assign \new_[48062]_  = ~A302 & ~A301;
  assign \new_[48063]_  = \new_[48062]_  & \new_[48059]_ ;
  assign \new_[48064]_  = \new_[48063]_  & \new_[48056]_ ;
  assign \new_[48068]_  = A167 & A168;
  assign \new_[48069]_  = A169 & \new_[48068]_ ;
  assign \new_[48073]_  = ~A200 & ~A199;
  assign \new_[48074]_  = ~A166 & \new_[48073]_ ;
  assign \new_[48075]_  = \new_[48074]_  & \new_[48069]_ ;
  assign \new_[48079]_  = A298 & A266;
  assign \new_[48080]_  = A265 & \new_[48079]_ ;
  assign \new_[48083]_  = ~A300 & ~A299;
  assign \new_[48086]_  = ~A302 & ~A301;
  assign \new_[48087]_  = \new_[48086]_  & \new_[48083]_ ;
  assign \new_[48088]_  = \new_[48087]_  & \new_[48080]_ ;
  assign \new_[48092]_  = A167 & A168;
  assign \new_[48093]_  = A169 & \new_[48092]_ ;
  assign \new_[48097]_  = ~A200 & ~A199;
  assign \new_[48098]_  = ~A166 & \new_[48097]_ ;
  assign \new_[48099]_  = \new_[48098]_  & \new_[48093]_ ;
  assign \new_[48103]_  = ~A298 & A266;
  assign \new_[48104]_  = A265 & \new_[48103]_ ;
  assign \new_[48107]_  = ~A300 & A299;
  assign \new_[48110]_  = ~A302 & ~A301;
  assign \new_[48111]_  = \new_[48110]_  & \new_[48107]_ ;
  assign \new_[48112]_  = \new_[48111]_  & \new_[48104]_ ;
  assign \new_[48116]_  = A167 & A168;
  assign \new_[48117]_  = A169 & \new_[48116]_ ;
  assign \new_[48121]_  = ~A200 & ~A199;
  assign \new_[48122]_  = ~A166 & \new_[48121]_ ;
  assign \new_[48123]_  = \new_[48122]_  & \new_[48117]_ ;
  assign \new_[48127]_  = A298 & ~A266;
  assign \new_[48128]_  = ~A265 & \new_[48127]_ ;
  assign \new_[48131]_  = ~A300 & ~A299;
  assign \new_[48134]_  = ~A302 & ~A301;
  assign \new_[48135]_  = \new_[48134]_  & \new_[48131]_ ;
  assign \new_[48136]_  = \new_[48135]_  & \new_[48128]_ ;
  assign \new_[48140]_  = A167 & A168;
  assign \new_[48141]_  = A169 & \new_[48140]_ ;
  assign \new_[48145]_  = ~A200 & ~A199;
  assign \new_[48146]_  = ~A166 & \new_[48145]_ ;
  assign \new_[48147]_  = \new_[48146]_  & \new_[48141]_ ;
  assign \new_[48151]_  = ~A298 & ~A266;
  assign \new_[48152]_  = ~A265 & \new_[48151]_ ;
  assign \new_[48155]_  = ~A300 & A299;
  assign \new_[48158]_  = ~A302 & ~A301;
  assign \new_[48159]_  = \new_[48158]_  & \new_[48155]_ ;
  assign \new_[48160]_  = \new_[48159]_  & \new_[48152]_ ;
  assign \new_[48164]_  = ~A167 & A168;
  assign \new_[48165]_  = A169 & \new_[48164]_ ;
  assign \new_[48169]_  = ~A202 & A201;
  assign \new_[48170]_  = A166 & \new_[48169]_ ;
  assign \new_[48171]_  = \new_[48170]_  & \new_[48165]_ ;
  assign \new_[48175]_  = A268 & ~A267;
  assign \new_[48176]_  = ~A203 & \new_[48175]_ ;
  assign \new_[48179]_  = ~A299 & A298;
  assign \new_[48182]_  = A301 & A300;
  assign \new_[48183]_  = \new_[48182]_  & \new_[48179]_ ;
  assign \new_[48184]_  = \new_[48183]_  & \new_[48176]_ ;
  assign \new_[48188]_  = ~A167 & A168;
  assign \new_[48189]_  = A169 & \new_[48188]_ ;
  assign \new_[48193]_  = ~A202 & A201;
  assign \new_[48194]_  = A166 & \new_[48193]_ ;
  assign \new_[48195]_  = \new_[48194]_  & \new_[48189]_ ;
  assign \new_[48199]_  = A268 & ~A267;
  assign \new_[48200]_  = ~A203 & \new_[48199]_ ;
  assign \new_[48203]_  = ~A299 & A298;
  assign \new_[48206]_  = A302 & A300;
  assign \new_[48207]_  = \new_[48206]_  & \new_[48203]_ ;
  assign \new_[48208]_  = \new_[48207]_  & \new_[48200]_ ;
  assign \new_[48212]_  = ~A167 & A168;
  assign \new_[48213]_  = A169 & \new_[48212]_ ;
  assign \new_[48217]_  = ~A202 & A201;
  assign \new_[48218]_  = A166 & \new_[48217]_ ;
  assign \new_[48219]_  = \new_[48218]_  & \new_[48213]_ ;
  assign \new_[48223]_  = A268 & ~A267;
  assign \new_[48224]_  = ~A203 & \new_[48223]_ ;
  assign \new_[48227]_  = A299 & ~A298;
  assign \new_[48230]_  = A301 & A300;
  assign \new_[48231]_  = \new_[48230]_  & \new_[48227]_ ;
  assign \new_[48232]_  = \new_[48231]_  & \new_[48224]_ ;
  assign \new_[48236]_  = ~A167 & A168;
  assign \new_[48237]_  = A169 & \new_[48236]_ ;
  assign \new_[48241]_  = ~A202 & A201;
  assign \new_[48242]_  = A166 & \new_[48241]_ ;
  assign \new_[48243]_  = \new_[48242]_  & \new_[48237]_ ;
  assign \new_[48247]_  = A268 & ~A267;
  assign \new_[48248]_  = ~A203 & \new_[48247]_ ;
  assign \new_[48251]_  = A299 & ~A298;
  assign \new_[48254]_  = A302 & A300;
  assign \new_[48255]_  = \new_[48254]_  & \new_[48251]_ ;
  assign \new_[48256]_  = \new_[48255]_  & \new_[48248]_ ;
  assign \new_[48260]_  = ~A167 & A168;
  assign \new_[48261]_  = A169 & \new_[48260]_ ;
  assign \new_[48265]_  = ~A202 & A201;
  assign \new_[48266]_  = A166 & \new_[48265]_ ;
  assign \new_[48267]_  = \new_[48266]_  & \new_[48261]_ ;
  assign \new_[48271]_  = A269 & ~A267;
  assign \new_[48272]_  = ~A203 & \new_[48271]_ ;
  assign \new_[48275]_  = ~A299 & A298;
  assign \new_[48278]_  = A301 & A300;
  assign \new_[48279]_  = \new_[48278]_  & \new_[48275]_ ;
  assign \new_[48280]_  = \new_[48279]_  & \new_[48272]_ ;
  assign \new_[48284]_  = ~A167 & A168;
  assign \new_[48285]_  = A169 & \new_[48284]_ ;
  assign \new_[48289]_  = ~A202 & A201;
  assign \new_[48290]_  = A166 & \new_[48289]_ ;
  assign \new_[48291]_  = \new_[48290]_  & \new_[48285]_ ;
  assign \new_[48295]_  = A269 & ~A267;
  assign \new_[48296]_  = ~A203 & \new_[48295]_ ;
  assign \new_[48299]_  = ~A299 & A298;
  assign \new_[48302]_  = A302 & A300;
  assign \new_[48303]_  = \new_[48302]_  & \new_[48299]_ ;
  assign \new_[48304]_  = \new_[48303]_  & \new_[48296]_ ;
  assign \new_[48308]_  = ~A167 & A168;
  assign \new_[48309]_  = A169 & \new_[48308]_ ;
  assign \new_[48313]_  = ~A202 & A201;
  assign \new_[48314]_  = A166 & \new_[48313]_ ;
  assign \new_[48315]_  = \new_[48314]_  & \new_[48309]_ ;
  assign \new_[48319]_  = A269 & ~A267;
  assign \new_[48320]_  = ~A203 & \new_[48319]_ ;
  assign \new_[48323]_  = A299 & ~A298;
  assign \new_[48326]_  = A301 & A300;
  assign \new_[48327]_  = \new_[48326]_  & \new_[48323]_ ;
  assign \new_[48328]_  = \new_[48327]_  & \new_[48320]_ ;
  assign \new_[48332]_  = ~A167 & A168;
  assign \new_[48333]_  = A169 & \new_[48332]_ ;
  assign \new_[48337]_  = ~A202 & A201;
  assign \new_[48338]_  = A166 & \new_[48337]_ ;
  assign \new_[48339]_  = \new_[48338]_  & \new_[48333]_ ;
  assign \new_[48343]_  = A269 & ~A267;
  assign \new_[48344]_  = ~A203 & \new_[48343]_ ;
  assign \new_[48347]_  = A299 & ~A298;
  assign \new_[48350]_  = A302 & A300;
  assign \new_[48351]_  = \new_[48350]_  & \new_[48347]_ ;
  assign \new_[48352]_  = \new_[48351]_  & \new_[48344]_ ;
  assign \new_[48356]_  = ~A167 & A168;
  assign \new_[48357]_  = A169 & \new_[48356]_ ;
  assign \new_[48361]_  = ~A202 & A201;
  assign \new_[48362]_  = A166 & \new_[48361]_ ;
  assign \new_[48363]_  = \new_[48362]_  & \new_[48357]_ ;
  assign \new_[48367]_  = A266 & A265;
  assign \new_[48368]_  = ~A203 & \new_[48367]_ ;
  assign \new_[48371]_  = ~A299 & A298;
  assign \new_[48374]_  = A301 & A300;
  assign \new_[48375]_  = \new_[48374]_  & \new_[48371]_ ;
  assign \new_[48376]_  = \new_[48375]_  & \new_[48368]_ ;
  assign \new_[48380]_  = ~A167 & A168;
  assign \new_[48381]_  = A169 & \new_[48380]_ ;
  assign \new_[48385]_  = ~A202 & A201;
  assign \new_[48386]_  = A166 & \new_[48385]_ ;
  assign \new_[48387]_  = \new_[48386]_  & \new_[48381]_ ;
  assign \new_[48391]_  = A266 & A265;
  assign \new_[48392]_  = ~A203 & \new_[48391]_ ;
  assign \new_[48395]_  = ~A299 & A298;
  assign \new_[48398]_  = A302 & A300;
  assign \new_[48399]_  = \new_[48398]_  & \new_[48395]_ ;
  assign \new_[48400]_  = \new_[48399]_  & \new_[48392]_ ;
  assign \new_[48404]_  = ~A167 & A168;
  assign \new_[48405]_  = A169 & \new_[48404]_ ;
  assign \new_[48409]_  = ~A202 & A201;
  assign \new_[48410]_  = A166 & \new_[48409]_ ;
  assign \new_[48411]_  = \new_[48410]_  & \new_[48405]_ ;
  assign \new_[48415]_  = A266 & A265;
  assign \new_[48416]_  = ~A203 & \new_[48415]_ ;
  assign \new_[48419]_  = A299 & ~A298;
  assign \new_[48422]_  = A301 & A300;
  assign \new_[48423]_  = \new_[48422]_  & \new_[48419]_ ;
  assign \new_[48424]_  = \new_[48423]_  & \new_[48416]_ ;
  assign \new_[48428]_  = ~A167 & A168;
  assign \new_[48429]_  = A169 & \new_[48428]_ ;
  assign \new_[48433]_  = ~A202 & A201;
  assign \new_[48434]_  = A166 & \new_[48433]_ ;
  assign \new_[48435]_  = \new_[48434]_  & \new_[48429]_ ;
  assign \new_[48439]_  = A266 & A265;
  assign \new_[48440]_  = ~A203 & \new_[48439]_ ;
  assign \new_[48443]_  = A299 & ~A298;
  assign \new_[48446]_  = A302 & A300;
  assign \new_[48447]_  = \new_[48446]_  & \new_[48443]_ ;
  assign \new_[48448]_  = \new_[48447]_  & \new_[48440]_ ;
  assign \new_[48452]_  = ~A167 & A168;
  assign \new_[48453]_  = A169 & \new_[48452]_ ;
  assign \new_[48457]_  = ~A202 & A201;
  assign \new_[48458]_  = A166 & \new_[48457]_ ;
  assign \new_[48459]_  = \new_[48458]_  & \new_[48453]_ ;
  assign \new_[48463]_  = ~A266 & ~A265;
  assign \new_[48464]_  = ~A203 & \new_[48463]_ ;
  assign \new_[48467]_  = ~A299 & A298;
  assign \new_[48470]_  = A301 & A300;
  assign \new_[48471]_  = \new_[48470]_  & \new_[48467]_ ;
  assign \new_[48472]_  = \new_[48471]_  & \new_[48464]_ ;
  assign \new_[48476]_  = ~A167 & A168;
  assign \new_[48477]_  = A169 & \new_[48476]_ ;
  assign \new_[48481]_  = ~A202 & A201;
  assign \new_[48482]_  = A166 & \new_[48481]_ ;
  assign \new_[48483]_  = \new_[48482]_  & \new_[48477]_ ;
  assign \new_[48487]_  = ~A266 & ~A265;
  assign \new_[48488]_  = ~A203 & \new_[48487]_ ;
  assign \new_[48491]_  = ~A299 & A298;
  assign \new_[48494]_  = A302 & A300;
  assign \new_[48495]_  = \new_[48494]_  & \new_[48491]_ ;
  assign \new_[48496]_  = \new_[48495]_  & \new_[48488]_ ;
  assign \new_[48500]_  = ~A167 & A168;
  assign \new_[48501]_  = A169 & \new_[48500]_ ;
  assign \new_[48505]_  = ~A202 & A201;
  assign \new_[48506]_  = A166 & \new_[48505]_ ;
  assign \new_[48507]_  = \new_[48506]_  & \new_[48501]_ ;
  assign \new_[48511]_  = ~A266 & ~A265;
  assign \new_[48512]_  = ~A203 & \new_[48511]_ ;
  assign \new_[48515]_  = A299 & ~A298;
  assign \new_[48518]_  = A301 & A300;
  assign \new_[48519]_  = \new_[48518]_  & \new_[48515]_ ;
  assign \new_[48520]_  = \new_[48519]_  & \new_[48512]_ ;
  assign \new_[48524]_  = ~A167 & A168;
  assign \new_[48525]_  = A169 & \new_[48524]_ ;
  assign \new_[48529]_  = ~A202 & A201;
  assign \new_[48530]_  = A166 & \new_[48529]_ ;
  assign \new_[48531]_  = \new_[48530]_  & \new_[48525]_ ;
  assign \new_[48535]_  = ~A266 & ~A265;
  assign \new_[48536]_  = ~A203 & \new_[48535]_ ;
  assign \new_[48539]_  = A299 & ~A298;
  assign \new_[48542]_  = A302 & A300;
  assign \new_[48543]_  = \new_[48542]_  & \new_[48539]_ ;
  assign \new_[48544]_  = \new_[48543]_  & \new_[48536]_ ;
  assign \new_[48548]_  = ~A167 & A168;
  assign \new_[48549]_  = A169 & \new_[48548]_ ;
  assign \new_[48553]_  = A202 & ~A201;
  assign \new_[48554]_  = A166 & \new_[48553]_ ;
  assign \new_[48555]_  = \new_[48554]_  & \new_[48549]_ ;
  assign \new_[48559]_  = ~A269 & ~A268;
  assign \new_[48560]_  = A267 & \new_[48559]_ ;
  assign \new_[48563]_  = ~A299 & A298;
  assign \new_[48566]_  = A301 & A300;
  assign \new_[48567]_  = \new_[48566]_  & \new_[48563]_ ;
  assign \new_[48568]_  = \new_[48567]_  & \new_[48560]_ ;
  assign \new_[48572]_  = ~A167 & A168;
  assign \new_[48573]_  = A169 & \new_[48572]_ ;
  assign \new_[48577]_  = A202 & ~A201;
  assign \new_[48578]_  = A166 & \new_[48577]_ ;
  assign \new_[48579]_  = \new_[48578]_  & \new_[48573]_ ;
  assign \new_[48583]_  = ~A269 & ~A268;
  assign \new_[48584]_  = A267 & \new_[48583]_ ;
  assign \new_[48587]_  = ~A299 & A298;
  assign \new_[48590]_  = A302 & A300;
  assign \new_[48591]_  = \new_[48590]_  & \new_[48587]_ ;
  assign \new_[48592]_  = \new_[48591]_  & \new_[48584]_ ;
  assign \new_[48596]_  = ~A167 & A168;
  assign \new_[48597]_  = A169 & \new_[48596]_ ;
  assign \new_[48601]_  = A202 & ~A201;
  assign \new_[48602]_  = A166 & \new_[48601]_ ;
  assign \new_[48603]_  = \new_[48602]_  & \new_[48597]_ ;
  assign \new_[48607]_  = ~A269 & ~A268;
  assign \new_[48608]_  = A267 & \new_[48607]_ ;
  assign \new_[48611]_  = A299 & ~A298;
  assign \new_[48614]_  = A301 & A300;
  assign \new_[48615]_  = \new_[48614]_  & \new_[48611]_ ;
  assign \new_[48616]_  = \new_[48615]_  & \new_[48608]_ ;
  assign \new_[48620]_  = ~A167 & A168;
  assign \new_[48621]_  = A169 & \new_[48620]_ ;
  assign \new_[48625]_  = A202 & ~A201;
  assign \new_[48626]_  = A166 & \new_[48625]_ ;
  assign \new_[48627]_  = \new_[48626]_  & \new_[48621]_ ;
  assign \new_[48631]_  = ~A269 & ~A268;
  assign \new_[48632]_  = A267 & \new_[48631]_ ;
  assign \new_[48635]_  = A299 & ~A298;
  assign \new_[48638]_  = A302 & A300;
  assign \new_[48639]_  = \new_[48638]_  & \new_[48635]_ ;
  assign \new_[48640]_  = \new_[48639]_  & \new_[48632]_ ;
  assign \new_[48644]_  = ~A167 & A168;
  assign \new_[48645]_  = A169 & \new_[48644]_ ;
  assign \new_[48649]_  = A202 & ~A201;
  assign \new_[48650]_  = A166 & \new_[48649]_ ;
  assign \new_[48651]_  = \new_[48650]_  & \new_[48645]_ ;
  assign \new_[48655]_  = A298 & A268;
  assign \new_[48656]_  = ~A267 & \new_[48655]_ ;
  assign \new_[48659]_  = ~A300 & ~A299;
  assign \new_[48662]_  = ~A302 & ~A301;
  assign \new_[48663]_  = \new_[48662]_  & \new_[48659]_ ;
  assign \new_[48664]_  = \new_[48663]_  & \new_[48656]_ ;
  assign \new_[48668]_  = ~A167 & A168;
  assign \new_[48669]_  = A169 & \new_[48668]_ ;
  assign \new_[48673]_  = A202 & ~A201;
  assign \new_[48674]_  = A166 & \new_[48673]_ ;
  assign \new_[48675]_  = \new_[48674]_  & \new_[48669]_ ;
  assign \new_[48679]_  = ~A298 & A268;
  assign \new_[48680]_  = ~A267 & \new_[48679]_ ;
  assign \new_[48683]_  = ~A300 & A299;
  assign \new_[48686]_  = ~A302 & ~A301;
  assign \new_[48687]_  = \new_[48686]_  & \new_[48683]_ ;
  assign \new_[48688]_  = \new_[48687]_  & \new_[48680]_ ;
  assign \new_[48692]_  = ~A167 & A168;
  assign \new_[48693]_  = A169 & \new_[48692]_ ;
  assign \new_[48697]_  = A202 & ~A201;
  assign \new_[48698]_  = A166 & \new_[48697]_ ;
  assign \new_[48699]_  = \new_[48698]_  & \new_[48693]_ ;
  assign \new_[48703]_  = A298 & A269;
  assign \new_[48704]_  = ~A267 & \new_[48703]_ ;
  assign \new_[48707]_  = ~A300 & ~A299;
  assign \new_[48710]_  = ~A302 & ~A301;
  assign \new_[48711]_  = \new_[48710]_  & \new_[48707]_ ;
  assign \new_[48712]_  = \new_[48711]_  & \new_[48704]_ ;
  assign \new_[48716]_  = ~A167 & A168;
  assign \new_[48717]_  = A169 & \new_[48716]_ ;
  assign \new_[48721]_  = A202 & ~A201;
  assign \new_[48722]_  = A166 & \new_[48721]_ ;
  assign \new_[48723]_  = \new_[48722]_  & \new_[48717]_ ;
  assign \new_[48727]_  = ~A298 & A269;
  assign \new_[48728]_  = ~A267 & \new_[48727]_ ;
  assign \new_[48731]_  = ~A300 & A299;
  assign \new_[48734]_  = ~A302 & ~A301;
  assign \new_[48735]_  = \new_[48734]_  & \new_[48731]_ ;
  assign \new_[48736]_  = \new_[48735]_  & \new_[48728]_ ;
  assign \new_[48740]_  = ~A167 & A168;
  assign \new_[48741]_  = A169 & \new_[48740]_ ;
  assign \new_[48745]_  = A202 & ~A201;
  assign \new_[48746]_  = A166 & \new_[48745]_ ;
  assign \new_[48747]_  = \new_[48746]_  & \new_[48741]_ ;
  assign \new_[48751]_  = A298 & A266;
  assign \new_[48752]_  = A265 & \new_[48751]_ ;
  assign \new_[48755]_  = ~A300 & ~A299;
  assign \new_[48758]_  = ~A302 & ~A301;
  assign \new_[48759]_  = \new_[48758]_  & \new_[48755]_ ;
  assign \new_[48760]_  = \new_[48759]_  & \new_[48752]_ ;
  assign \new_[48764]_  = ~A167 & A168;
  assign \new_[48765]_  = A169 & \new_[48764]_ ;
  assign \new_[48769]_  = A202 & ~A201;
  assign \new_[48770]_  = A166 & \new_[48769]_ ;
  assign \new_[48771]_  = \new_[48770]_  & \new_[48765]_ ;
  assign \new_[48775]_  = ~A298 & A266;
  assign \new_[48776]_  = A265 & \new_[48775]_ ;
  assign \new_[48779]_  = ~A300 & A299;
  assign \new_[48782]_  = ~A302 & ~A301;
  assign \new_[48783]_  = \new_[48782]_  & \new_[48779]_ ;
  assign \new_[48784]_  = \new_[48783]_  & \new_[48776]_ ;
  assign \new_[48788]_  = ~A167 & A168;
  assign \new_[48789]_  = A169 & \new_[48788]_ ;
  assign \new_[48793]_  = A202 & ~A201;
  assign \new_[48794]_  = A166 & \new_[48793]_ ;
  assign \new_[48795]_  = \new_[48794]_  & \new_[48789]_ ;
  assign \new_[48799]_  = A298 & ~A266;
  assign \new_[48800]_  = ~A265 & \new_[48799]_ ;
  assign \new_[48803]_  = ~A300 & ~A299;
  assign \new_[48806]_  = ~A302 & ~A301;
  assign \new_[48807]_  = \new_[48806]_  & \new_[48803]_ ;
  assign \new_[48808]_  = \new_[48807]_  & \new_[48800]_ ;
  assign \new_[48812]_  = ~A167 & A168;
  assign \new_[48813]_  = A169 & \new_[48812]_ ;
  assign \new_[48817]_  = A202 & ~A201;
  assign \new_[48818]_  = A166 & \new_[48817]_ ;
  assign \new_[48819]_  = \new_[48818]_  & \new_[48813]_ ;
  assign \new_[48823]_  = ~A298 & ~A266;
  assign \new_[48824]_  = ~A265 & \new_[48823]_ ;
  assign \new_[48827]_  = ~A300 & A299;
  assign \new_[48830]_  = ~A302 & ~A301;
  assign \new_[48831]_  = \new_[48830]_  & \new_[48827]_ ;
  assign \new_[48832]_  = \new_[48831]_  & \new_[48824]_ ;
  assign \new_[48836]_  = ~A167 & A168;
  assign \new_[48837]_  = A169 & \new_[48836]_ ;
  assign \new_[48841]_  = A203 & ~A201;
  assign \new_[48842]_  = A166 & \new_[48841]_ ;
  assign \new_[48843]_  = \new_[48842]_  & \new_[48837]_ ;
  assign \new_[48847]_  = ~A269 & ~A268;
  assign \new_[48848]_  = A267 & \new_[48847]_ ;
  assign \new_[48851]_  = ~A299 & A298;
  assign \new_[48854]_  = A301 & A300;
  assign \new_[48855]_  = \new_[48854]_  & \new_[48851]_ ;
  assign \new_[48856]_  = \new_[48855]_  & \new_[48848]_ ;
  assign \new_[48860]_  = ~A167 & A168;
  assign \new_[48861]_  = A169 & \new_[48860]_ ;
  assign \new_[48865]_  = A203 & ~A201;
  assign \new_[48866]_  = A166 & \new_[48865]_ ;
  assign \new_[48867]_  = \new_[48866]_  & \new_[48861]_ ;
  assign \new_[48871]_  = ~A269 & ~A268;
  assign \new_[48872]_  = A267 & \new_[48871]_ ;
  assign \new_[48875]_  = ~A299 & A298;
  assign \new_[48878]_  = A302 & A300;
  assign \new_[48879]_  = \new_[48878]_  & \new_[48875]_ ;
  assign \new_[48880]_  = \new_[48879]_  & \new_[48872]_ ;
  assign \new_[48884]_  = ~A167 & A168;
  assign \new_[48885]_  = A169 & \new_[48884]_ ;
  assign \new_[48889]_  = A203 & ~A201;
  assign \new_[48890]_  = A166 & \new_[48889]_ ;
  assign \new_[48891]_  = \new_[48890]_  & \new_[48885]_ ;
  assign \new_[48895]_  = ~A269 & ~A268;
  assign \new_[48896]_  = A267 & \new_[48895]_ ;
  assign \new_[48899]_  = A299 & ~A298;
  assign \new_[48902]_  = A301 & A300;
  assign \new_[48903]_  = \new_[48902]_  & \new_[48899]_ ;
  assign \new_[48904]_  = \new_[48903]_  & \new_[48896]_ ;
  assign \new_[48908]_  = ~A167 & A168;
  assign \new_[48909]_  = A169 & \new_[48908]_ ;
  assign \new_[48913]_  = A203 & ~A201;
  assign \new_[48914]_  = A166 & \new_[48913]_ ;
  assign \new_[48915]_  = \new_[48914]_  & \new_[48909]_ ;
  assign \new_[48919]_  = ~A269 & ~A268;
  assign \new_[48920]_  = A267 & \new_[48919]_ ;
  assign \new_[48923]_  = A299 & ~A298;
  assign \new_[48926]_  = A302 & A300;
  assign \new_[48927]_  = \new_[48926]_  & \new_[48923]_ ;
  assign \new_[48928]_  = \new_[48927]_  & \new_[48920]_ ;
  assign \new_[48932]_  = ~A167 & A168;
  assign \new_[48933]_  = A169 & \new_[48932]_ ;
  assign \new_[48937]_  = A203 & ~A201;
  assign \new_[48938]_  = A166 & \new_[48937]_ ;
  assign \new_[48939]_  = \new_[48938]_  & \new_[48933]_ ;
  assign \new_[48943]_  = A298 & A268;
  assign \new_[48944]_  = ~A267 & \new_[48943]_ ;
  assign \new_[48947]_  = ~A300 & ~A299;
  assign \new_[48950]_  = ~A302 & ~A301;
  assign \new_[48951]_  = \new_[48950]_  & \new_[48947]_ ;
  assign \new_[48952]_  = \new_[48951]_  & \new_[48944]_ ;
  assign \new_[48956]_  = ~A167 & A168;
  assign \new_[48957]_  = A169 & \new_[48956]_ ;
  assign \new_[48961]_  = A203 & ~A201;
  assign \new_[48962]_  = A166 & \new_[48961]_ ;
  assign \new_[48963]_  = \new_[48962]_  & \new_[48957]_ ;
  assign \new_[48967]_  = ~A298 & A268;
  assign \new_[48968]_  = ~A267 & \new_[48967]_ ;
  assign \new_[48971]_  = ~A300 & A299;
  assign \new_[48974]_  = ~A302 & ~A301;
  assign \new_[48975]_  = \new_[48974]_  & \new_[48971]_ ;
  assign \new_[48976]_  = \new_[48975]_  & \new_[48968]_ ;
  assign \new_[48980]_  = ~A167 & A168;
  assign \new_[48981]_  = A169 & \new_[48980]_ ;
  assign \new_[48985]_  = A203 & ~A201;
  assign \new_[48986]_  = A166 & \new_[48985]_ ;
  assign \new_[48987]_  = \new_[48986]_  & \new_[48981]_ ;
  assign \new_[48991]_  = A298 & A269;
  assign \new_[48992]_  = ~A267 & \new_[48991]_ ;
  assign \new_[48995]_  = ~A300 & ~A299;
  assign \new_[48998]_  = ~A302 & ~A301;
  assign \new_[48999]_  = \new_[48998]_  & \new_[48995]_ ;
  assign \new_[49000]_  = \new_[48999]_  & \new_[48992]_ ;
  assign \new_[49004]_  = ~A167 & A168;
  assign \new_[49005]_  = A169 & \new_[49004]_ ;
  assign \new_[49009]_  = A203 & ~A201;
  assign \new_[49010]_  = A166 & \new_[49009]_ ;
  assign \new_[49011]_  = \new_[49010]_  & \new_[49005]_ ;
  assign \new_[49015]_  = ~A298 & A269;
  assign \new_[49016]_  = ~A267 & \new_[49015]_ ;
  assign \new_[49019]_  = ~A300 & A299;
  assign \new_[49022]_  = ~A302 & ~A301;
  assign \new_[49023]_  = \new_[49022]_  & \new_[49019]_ ;
  assign \new_[49024]_  = \new_[49023]_  & \new_[49016]_ ;
  assign \new_[49028]_  = ~A167 & A168;
  assign \new_[49029]_  = A169 & \new_[49028]_ ;
  assign \new_[49033]_  = A203 & ~A201;
  assign \new_[49034]_  = A166 & \new_[49033]_ ;
  assign \new_[49035]_  = \new_[49034]_  & \new_[49029]_ ;
  assign \new_[49039]_  = A298 & A266;
  assign \new_[49040]_  = A265 & \new_[49039]_ ;
  assign \new_[49043]_  = ~A300 & ~A299;
  assign \new_[49046]_  = ~A302 & ~A301;
  assign \new_[49047]_  = \new_[49046]_  & \new_[49043]_ ;
  assign \new_[49048]_  = \new_[49047]_  & \new_[49040]_ ;
  assign \new_[49052]_  = ~A167 & A168;
  assign \new_[49053]_  = A169 & \new_[49052]_ ;
  assign \new_[49057]_  = A203 & ~A201;
  assign \new_[49058]_  = A166 & \new_[49057]_ ;
  assign \new_[49059]_  = \new_[49058]_  & \new_[49053]_ ;
  assign \new_[49063]_  = ~A298 & A266;
  assign \new_[49064]_  = A265 & \new_[49063]_ ;
  assign \new_[49067]_  = ~A300 & A299;
  assign \new_[49070]_  = ~A302 & ~A301;
  assign \new_[49071]_  = \new_[49070]_  & \new_[49067]_ ;
  assign \new_[49072]_  = \new_[49071]_  & \new_[49064]_ ;
  assign \new_[49076]_  = ~A167 & A168;
  assign \new_[49077]_  = A169 & \new_[49076]_ ;
  assign \new_[49081]_  = A203 & ~A201;
  assign \new_[49082]_  = A166 & \new_[49081]_ ;
  assign \new_[49083]_  = \new_[49082]_  & \new_[49077]_ ;
  assign \new_[49087]_  = A298 & ~A266;
  assign \new_[49088]_  = ~A265 & \new_[49087]_ ;
  assign \new_[49091]_  = ~A300 & ~A299;
  assign \new_[49094]_  = ~A302 & ~A301;
  assign \new_[49095]_  = \new_[49094]_  & \new_[49091]_ ;
  assign \new_[49096]_  = \new_[49095]_  & \new_[49088]_ ;
  assign \new_[49100]_  = ~A167 & A168;
  assign \new_[49101]_  = A169 & \new_[49100]_ ;
  assign \new_[49105]_  = A203 & ~A201;
  assign \new_[49106]_  = A166 & \new_[49105]_ ;
  assign \new_[49107]_  = \new_[49106]_  & \new_[49101]_ ;
  assign \new_[49111]_  = ~A298 & ~A266;
  assign \new_[49112]_  = ~A265 & \new_[49111]_ ;
  assign \new_[49115]_  = ~A300 & A299;
  assign \new_[49118]_  = ~A302 & ~A301;
  assign \new_[49119]_  = \new_[49118]_  & \new_[49115]_ ;
  assign \new_[49120]_  = \new_[49119]_  & \new_[49112]_ ;
  assign \new_[49124]_  = ~A167 & A168;
  assign \new_[49125]_  = A169 & \new_[49124]_ ;
  assign \new_[49129]_  = A200 & A199;
  assign \new_[49130]_  = A166 & \new_[49129]_ ;
  assign \new_[49131]_  = \new_[49130]_  & \new_[49125]_ ;
  assign \new_[49135]_  = ~A269 & ~A268;
  assign \new_[49136]_  = A267 & \new_[49135]_ ;
  assign \new_[49139]_  = ~A299 & A298;
  assign \new_[49142]_  = A301 & A300;
  assign \new_[49143]_  = \new_[49142]_  & \new_[49139]_ ;
  assign \new_[49144]_  = \new_[49143]_  & \new_[49136]_ ;
  assign \new_[49148]_  = ~A167 & A168;
  assign \new_[49149]_  = A169 & \new_[49148]_ ;
  assign \new_[49153]_  = A200 & A199;
  assign \new_[49154]_  = A166 & \new_[49153]_ ;
  assign \new_[49155]_  = \new_[49154]_  & \new_[49149]_ ;
  assign \new_[49159]_  = ~A269 & ~A268;
  assign \new_[49160]_  = A267 & \new_[49159]_ ;
  assign \new_[49163]_  = ~A299 & A298;
  assign \new_[49166]_  = A302 & A300;
  assign \new_[49167]_  = \new_[49166]_  & \new_[49163]_ ;
  assign \new_[49168]_  = \new_[49167]_  & \new_[49160]_ ;
  assign \new_[49172]_  = ~A167 & A168;
  assign \new_[49173]_  = A169 & \new_[49172]_ ;
  assign \new_[49177]_  = A200 & A199;
  assign \new_[49178]_  = A166 & \new_[49177]_ ;
  assign \new_[49179]_  = \new_[49178]_  & \new_[49173]_ ;
  assign \new_[49183]_  = ~A269 & ~A268;
  assign \new_[49184]_  = A267 & \new_[49183]_ ;
  assign \new_[49187]_  = A299 & ~A298;
  assign \new_[49190]_  = A301 & A300;
  assign \new_[49191]_  = \new_[49190]_  & \new_[49187]_ ;
  assign \new_[49192]_  = \new_[49191]_  & \new_[49184]_ ;
  assign \new_[49196]_  = ~A167 & A168;
  assign \new_[49197]_  = A169 & \new_[49196]_ ;
  assign \new_[49201]_  = A200 & A199;
  assign \new_[49202]_  = A166 & \new_[49201]_ ;
  assign \new_[49203]_  = \new_[49202]_  & \new_[49197]_ ;
  assign \new_[49207]_  = ~A269 & ~A268;
  assign \new_[49208]_  = A267 & \new_[49207]_ ;
  assign \new_[49211]_  = A299 & ~A298;
  assign \new_[49214]_  = A302 & A300;
  assign \new_[49215]_  = \new_[49214]_  & \new_[49211]_ ;
  assign \new_[49216]_  = \new_[49215]_  & \new_[49208]_ ;
  assign \new_[49220]_  = ~A167 & A168;
  assign \new_[49221]_  = A169 & \new_[49220]_ ;
  assign \new_[49225]_  = A200 & A199;
  assign \new_[49226]_  = A166 & \new_[49225]_ ;
  assign \new_[49227]_  = \new_[49226]_  & \new_[49221]_ ;
  assign \new_[49231]_  = A298 & A268;
  assign \new_[49232]_  = ~A267 & \new_[49231]_ ;
  assign \new_[49235]_  = ~A300 & ~A299;
  assign \new_[49238]_  = ~A302 & ~A301;
  assign \new_[49239]_  = \new_[49238]_  & \new_[49235]_ ;
  assign \new_[49240]_  = \new_[49239]_  & \new_[49232]_ ;
  assign \new_[49244]_  = ~A167 & A168;
  assign \new_[49245]_  = A169 & \new_[49244]_ ;
  assign \new_[49249]_  = A200 & A199;
  assign \new_[49250]_  = A166 & \new_[49249]_ ;
  assign \new_[49251]_  = \new_[49250]_  & \new_[49245]_ ;
  assign \new_[49255]_  = ~A298 & A268;
  assign \new_[49256]_  = ~A267 & \new_[49255]_ ;
  assign \new_[49259]_  = ~A300 & A299;
  assign \new_[49262]_  = ~A302 & ~A301;
  assign \new_[49263]_  = \new_[49262]_  & \new_[49259]_ ;
  assign \new_[49264]_  = \new_[49263]_  & \new_[49256]_ ;
  assign \new_[49268]_  = ~A167 & A168;
  assign \new_[49269]_  = A169 & \new_[49268]_ ;
  assign \new_[49273]_  = A200 & A199;
  assign \new_[49274]_  = A166 & \new_[49273]_ ;
  assign \new_[49275]_  = \new_[49274]_  & \new_[49269]_ ;
  assign \new_[49279]_  = A298 & A269;
  assign \new_[49280]_  = ~A267 & \new_[49279]_ ;
  assign \new_[49283]_  = ~A300 & ~A299;
  assign \new_[49286]_  = ~A302 & ~A301;
  assign \new_[49287]_  = \new_[49286]_  & \new_[49283]_ ;
  assign \new_[49288]_  = \new_[49287]_  & \new_[49280]_ ;
  assign \new_[49292]_  = ~A167 & A168;
  assign \new_[49293]_  = A169 & \new_[49292]_ ;
  assign \new_[49297]_  = A200 & A199;
  assign \new_[49298]_  = A166 & \new_[49297]_ ;
  assign \new_[49299]_  = \new_[49298]_  & \new_[49293]_ ;
  assign \new_[49303]_  = ~A298 & A269;
  assign \new_[49304]_  = ~A267 & \new_[49303]_ ;
  assign \new_[49307]_  = ~A300 & A299;
  assign \new_[49310]_  = ~A302 & ~A301;
  assign \new_[49311]_  = \new_[49310]_  & \new_[49307]_ ;
  assign \new_[49312]_  = \new_[49311]_  & \new_[49304]_ ;
  assign \new_[49316]_  = ~A167 & A168;
  assign \new_[49317]_  = A169 & \new_[49316]_ ;
  assign \new_[49321]_  = A200 & A199;
  assign \new_[49322]_  = A166 & \new_[49321]_ ;
  assign \new_[49323]_  = \new_[49322]_  & \new_[49317]_ ;
  assign \new_[49327]_  = A298 & A266;
  assign \new_[49328]_  = A265 & \new_[49327]_ ;
  assign \new_[49331]_  = ~A300 & ~A299;
  assign \new_[49334]_  = ~A302 & ~A301;
  assign \new_[49335]_  = \new_[49334]_  & \new_[49331]_ ;
  assign \new_[49336]_  = \new_[49335]_  & \new_[49328]_ ;
  assign \new_[49340]_  = ~A167 & A168;
  assign \new_[49341]_  = A169 & \new_[49340]_ ;
  assign \new_[49345]_  = A200 & A199;
  assign \new_[49346]_  = A166 & \new_[49345]_ ;
  assign \new_[49347]_  = \new_[49346]_  & \new_[49341]_ ;
  assign \new_[49351]_  = ~A298 & A266;
  assign \new_[49352]_  = A265 & \new_[49351]_ ;
  assign \new_[49355]_  = ~A300 & A299;
  assign \new_[49358]_  = ~A302 & ~A301;
  assign \new_[49359]_  = \new_[49358]_  & \new_[49355]_ ;
  assign \new_[49360]_  = \new_[49359]_  & \new_[49352]_ ;
  assign \new_[49364]_  = ~A167 & A168;
  assign \new_[49365]_  = A169 & \new_[49364]_ ;
  assign \new_[49369]_  = A200 & A199;
  assign \new_[49370]_  = A166 & \new_[49369]_ ;
  assign \new_[49371]_  = \new_[49370]_  & \new_[49365]_ ;
  assign \new_[49375]_  = A298 & ~A266;
  assign \new_[49376]_  = ~A265 & \new_[49375]_ ;
  assign \new_[49379]_  = ~A300 & ~A299;
  assign \new_[49382]_  = ~A302 & ~A301;
  assign \new_[49383]_  = \new_[49382]_  & \new_[49379]_ ;
  assign \new_[49384]_  = \new_[49383]_  & \new_[49376]_ ;
  assign \new_[49388]_  = ~A167 & A168;
  assign \new_[49389]_  = A169 & \new_[49388]_ ;
  assign \new_[49393]_  = A200 & A199;
  assign \new_[49394]_  = A166 & \new_[49393]_ ;
  assign \new_[49395]_  = \new_[49394]_  & \new_[49389]_ ;
  assign \new_[49399]_  = ~A298 & ~A266;
  assign \new_[49400]_  = ~A265 & \new_[49399]_ ;
  assign \new_[49403]_  = ~A300 & A299;
  assign \new_[49406]_  = ~A302 & ~A301;
  assign \new_[49407]_  = \new_[49406]_  & \new_[49403]_ ;
  assign \new_[49408]_  = \new_[49407]_  & \new_[49400]_ ;
  assign \new_[49412]_  = ~A167 & A168;
  assign \new_[49413]_  = A169 & \new_[49412]_ ;
  assign \new_[49417]_  = ~A200 & ~A199;
  assign \new_[49418]_  = A166 & \new_[49417]_ ;
  assign \new_[49419]_  = \new_[49418]_  & \new_[49413]_ ;
  assign \new_[49423]_  = ~A269 & ~A268;
  assign \new_[49424]_  = A267 & \new_[49423]_ ;
  assign \new_[49427]_  = ~A299 & A298;
  assign \new_[49430]_  = A301 & A300;
  assign \new_[49431]_  = \new_[49430]_  & \new_[49427]_ ;
  assign \new_[49432]_  = \new_[49431]_  & \new_[49424]_ ;
  assign \new_[49436]_  = ~A167 & A168;
  assign \new_[49437]_  = A169 & \new_[49436]_ ;
  assign \new_[49441]_  = ~A200 & ~A199;
  assign \new_[49442]_  = A166 & \new_[49441]_ ;
  assign \new_[49443]_  = \new_[49442]_  & \new_[49437]_ ;
  assign \new_[49447]_  = ~A269 & ~A268;
  assign \new_[49448]_  = A267 & \new_[49447]_ ;
  assign \new_[49451]_  = ~A299 & A298;
  assign \new_[49454]_  = A302 & A300;
  assign \new_[49455]_  = \new_[49454]_  & \new_[49451]_ ;
  assign \new_[49456]_  = \new_[49455]_  & \new_[49448]_ ;
  assign \new_[49460]_  = ~A167 & A168;
  assign \new_[49461]_  = A169 & \new_[49460]_ ;
  assign \new_[49465]_  = ~A200 & ~A199;
  assign \new_[49466]_  = A166 & \new_[49465]_ ;
  assign \new_[49467]_  = \new_[49466]_  & \new_[49461]_ ;
  assign \new_[49471]_  = ~A269 & ~A268;
  assign \new_[49472]_  = A267 & \new_[49471]_ ;
  assign \new_[49475]_  = A299 & ~A298;
  assign \new_[49478]_  = A301 & A300;
  assign \new_[49479]_  = \new_[49478]_  & \new_[49475]_ ;
  assign \new_[49480]_  = \new_[49479]_  & \new_[49472]_ ;
  assign \new_[49484]_  = ~A167 & A168;
  assign \new_[49485]_  = A169 & \new_[49484]_ ;
  assign \new_[49489]_  = ~A200 & ~A199;
  assign \new_[49490]_  = A166 & \new_[49489]_ ;
  assign \new_[49491]_  = \new_[49490]_  & \new_[49485]_ ;
  assign \new_[49495]_  = ~A269 & ~A268;
  assign \new_[49496]_  = A267 & \new_[49495]_ ;
  assign \new_[49499]_  = A299 & ~A298;
  assign \new_[49502]_  = A302 & A300;
  assign \new_[49503]_  = \new_[49502]_  & \new_[49499]_ ;
  assign \new_[49504]_  = \new_[49503]_  & \new_[49496]_ ;
  assign \new_[49508]_  = ~A167 & A168;
  assign \new_[49509]_  = A169 & \new_[49508]_ ;
  assign \new_[49513]_  = ~A200 & ~A199;
  assign \new_[49514]_  = A166 & \new_[49513]_ ;
  assign \new_[49515]_  = \new_[49514]_  & \new_[49509]_ ;
  assign \new_[49519]_  = A298 & A268;
  assign \new_[49520]_  = ~A267 & \new_[49519]_ ;
  assign \new_[49523]_  = ~A300 & ~A299;
  assign \new_[49526]_  = ~A302 & ~A301;
  assign \new_[49527]_  = \new_[49526]_  & \new_[49523]_ ;
  assign \new_[49528]_  = \new_[49527]_  & \new_[49520]_ ;
  assign \new_[49532]_  = ~A167 & A168;
  assign \new_[49533]_  = A169 & \new_[49532]_ ;
  assign \new_[49537]_  = ~A200 & ~A199;
  assign \new_[49538]_  = A166 & \new_[49537]_ ;
  assign \new_[49539]_  = \new_[49538]_  & \new_[49533]_ ;
  assign \new_[49543]_  = ~A298 & A268;
  assign \new_[49544]_  = ~A267 & \new_[49543]_ ;
  assign \new_[49547]_  = ~A300 & A299;
  assign \new_[49550]_  = ~A302 & ~A301;
  assign \new_[49551]_  = \new_[49550]_  & \new_[49547]_ ;
  assign \new_[49552]_  = \new_[49551]_  & \new_[49544]_ ;
  assign \new_[49556]_  = ~A167 & A168;
  assign \new_[49557]_  = A169 & \new_[49556]_ ;
  assign \new_[49561]_  = ~A200 & ~A199;
  assign \new_[49562]_  = A166 & \new_[49561]_ ;
  assign \new_[49563]_  = \new_[49562]_  & \new_[49557]_ ;
  assign \new_[49567]_  = A298 & A269;
  assign \new_[49568]_  = ~A267 & \new_[49567]_ ;
  assign \new_[49571]_  = ~A300 & ~A299;
  assign \new_[49574]_  = ~A302 & ~A301;
  assign \new_[49575]_  = \new_[49574]_  & \new_[49571]_ ;
  assign \new_[49576]_  = \new_[49575]_  & \new_[49568]_ ;
  assign \new_[49580]_  = ~A167 & A168;
  assign \new_[49581]_  = A169 & \new_[49580]_ ;
  assign \new_[49585]_  = ~A200 & ~A199;
  assign \new_[49586]_  = A166 & \new_[49585]_ ;
  assign \new_[49587]_  = \new_[49586]_  & \new_[49581]_ ;
  assign \new_[49591]_  = ~A298 & A269;
  assign \new_[49592]_  = ~A267 & \new_[49591]_ ;
  assign \new_[49595]_  = ~A300 & A299;
  assign \new_[49598]_  = ~A302 & ~A301;
  assign \new_[49599]_  = \new_[49598]_  & \new_[49595]_ ;
  assign \new_[49600]_  = \new_[49599]_  & \new_[49592]_ ;
  assign \new_[49604]_  = ~A167 & A168;
  assign \new_[49605]_  = A169 & \new_[49604]_ ;
  assign \new_[49609]_  = ~A200 & ~A199;
  assign \new_[49610]_  = A166 & \new_[49609]_ ;
  assign \new_[49611]_  = \new_[49610]_  & \new_[49605]_ ;
  assign \new_[49615]_  = A298 & A266;
  assign \new_[49616]_  = A265 & \new_[49615]_ ;
  assign \new_[49619]_  = ~A300 & ~A299;
  assign \new_[49622]_  = ~A302 & ~A301;
  assign \new_[49623]_  = \new_[49622]_  & \new_[49619]_ ;
  assign \new_[49624]_  = \new_[49623]_  & \new_[49616]_ ;
  assign \new_[49628]_  = ~A167 & A168;
  assign \new_[49629]_  = A169 & \new_[49628]_ ;
  assign \new_[49633]_  = ~A200 & ~A199;
  assign \new_[49634]_  = A166 & \new_[49633]_ ;
  assign \new_[49635]_  = \new_[49634]_  & \new_[49629]_ ;
  assign \new_[49639]_  = ~A298 & A266;
  assign \new_[49640]_  = A265 & \new_[49639]_ ;
  assign \new_[49643]_  = ~A300 & A299;
  assign \new_[49646]_  = ~A302 & ~A301;
  assign \new_[49647]_  = \new_[49646]_  & \new_[49643]_ ;
  assign \new_[49648]_  = \new_[49647]_  & \new_[49640]_ ;
  assign \new_[49652]_  = ~A167 & A168;
  assign \new_[49653]_  = A169 & \new_[49652]_ ;
  assign \new_[49657]_  = ~A200 & ~A199;
  assign \new_[49658]_  = A166 & \new_[49657]_ ;
  assign \new_[49659]_  = \new_[49658]_  & \new_[49653]_ ;
  assign \new_[49663]_  = A298 & ~A266;
  assign \new_[49664]_  = ~A265 & \new_[49663]_ ;
  assign \new_[49667]_  = ~A300 & ~A299;
  assign \new_[49670]_  = ~A302 & ~A301;
  assign \new_[49671]_  = \new_[49670]_  & \new_[49667]_ ;
  assign \new_[49672]_  = \new_[49671]_  & \new_[49664]_ ;
  assign \new_[49676]_  = ~A167 & A168;
  assign \new_[49677]_  = A169 & \new_[49676]_ ;
  assign \new_[49681]_  = ~A200 & ~A199;
  assign \new_[49682]_  = A166 & \new_[49681]_ ;
  assign \new_[49683]_  = \new_[49682]_  & \new_[49677]_ ;
  assign \new_[49687]_  = ~A298 & ~A266;
  assign \new_[49688]_  = ~A265 & \new_[49687]_ ;
  assign \new_[49691]_  = ~A300 & A299;
  assign \new_[49694]_  = ~A302 & ~A301;
  assign \new_[49695]_  = \new_[49694]_  & \new_[49691]_ ;
  assign \new_[49696]_  = \new_[49695]_  & \new_[49688]_ ;
  assign \new_[49700]_  = A201 & ~A168;
  assign \new_[49701]_  = A169 & \new_[49700]_ ;
  assign \new_[49705]_  = ~A265 & ~A203;
  assign \new_[49706]_  = ~A202 & \new_[49705]_ ;
  assign \new_[49707]_  = \new_[49706]_  & \new_[49701]_ ;
  assign \new_[49711]_  = ~A268 & ~A267;
  assign \new_[49712]_  = A266 & \new_[49711]_ ;
  assign \new_[49715]_  = A300 & ~A269;
  assign \new_[49718]_  = ~A302 & ~A301;
  assign \new_[49719]_  = \new_[49718]_  & \new_[49715]_ ;
  assign \new_[49720]_  = \new_[49719]_  & \new_[49712]_ ;
  assign \new_[49724]_  = A201 & ~A168;
  assign \new_[49725]_  = A169 & \new_[49724]_ ;
  assign \new_[49729]_  = A265 & ~A203;
  assign \new_[49730]_  = ~A202 & \new_[49729]_ ;
  assign \new_[49731]_  = \new_[49730]_  & \new_[49725]_ ;
  assign \new_[49735]_  = ~A268 & ~A267;
  assign \new_[49736]_  = ~A266 & \new_[49735]_ ;
  assign \new_[49739]_  = A300 & ~A269;
  assign \new_[49742]_  = ~A302 & ~A301;
  assign \new_[49743]_  = \new_[49742]_  & \new_[49739]_ ;
  assign \new_[49744]_  = \new_[49743]_  & \new_[49736]_ ;
  assign \new_[49748]_  = ~A199 & ~A168;
  assign \new_[49749]_  = A169 & \new_[49748]_ ;
  assign \new_[49753]_  = A202 & A201;
  assign \new_[49754]_  = A200 & \new_[49753]_ ;
  assign \new_[49755]_  = \new_[49754]_  & \new_[49749]_ ;
  assign \new_[49759]_  = ~A269 & ~A268;
  assign \new_[49760]_  = A267 & \new_[49759]_ ;
  assign \new_[49763]_  = ~A299 & A298;
  assign \new_[49766]_  = A301 & A300;
  assign \new_[49767]_  = \new_[49766]_  & \new_[49763]_ ;
  assign \new_[49768]_  = \new_[49767]_  & \new_[49760]_ ;
  assign \new_[49772]_  = ~A199 & ~A168;
  assign \new_[49773]_  = A169 & \new_[49772]_ ;
  assign \new_[49777]_  = A202 & A201;
  assign \new_[49778]_  = A200 & \new_[49777]_ ;
  assign \new_[49779]_  = \new_[49778]_  & \new_[49773]_ ;
  assign \new_[49783]_  = ~A269 & ~A268;
  assign \new_[49784]_  = A267 & \new_[49783]_ ;
  assign \new_[49787]_  = ~A299 & A298;
  assign \new_[49790]_  = A302 & A300;
  assign \new_[49791]_  = \new_[49790]_  & \new_[49787]_ ;
  assign \new_[49792]_  = \new_[49791]_  & \new_[49784]_ ;
  assign \new_[49796]_  = ~A199 & ~A168;
  assign \new_[49797]_  = A169 & \new_[49796]_ ;
  assign \new_[49801]_  = A202 & A201;
  assign \new_[49802]_  = A200 & \new_[49801]_ ;
  assign \new_[49803]_  = \new_[49802]_  & \new_[49797]_ ;
  assign \new_[49807]_  = ~A269 & ~A268;
  assign \new_[49808]_  = A267 & \new_[49807]_ ;
  assign \new_[49811]_  = A299 & ~A298;
  assign \new_[49814]_  = A301 & A300;
  assign \new_[49815]_  = \new_[49814]_  & \new_[49811]_ ;
  assign \new_[49816]_  = \new_[49815]_  & \new_[49808]_ ;
  assign \new_[49820]_  = ~A199 & ~A168;
  assign \new_[49821]_  = A169 & \new_[49820]_ ;
  assign \new_[49825]_  = A202 & A201;
  assign \new_[49826]_  = A200 & \new_[49825]_ ;
  assign \new_[49827]_  = \new_[49826]_  & \new_[49821]_ ;
  assign \new_[49831]_  = ~A269 & ~A268;
  assign \new_[49832]_  = A267 & \new_[49831]_ ;
  assign \new_[49835]_  = A299 & ~A298;
  assign \new_[49838]_  = A302 & A300;
  assign \new_[49839]_  = \new_[49838]_  & \new_[49835]_ ;
  assign \new_[49840]_  = \new_[49839]_  & \new_[49832]_ ;
  assign \new_[49844]_  = ~A199 & ~A168;
  assign \new_[49845]_  = A169 & \new_[49844]_ ;
  assign \new_[49849]_  = A202 & A201;
  assign \new_[49850]_  = A200 & \new_[49849]_ ;
  assign \new_[49851]_  = \new_[49850]_  & \new_[49845]_ ;
  assign \new_[49855]_  = A298 & A268;
  assign \new_[49856]_  = ~A267 & \new_[49855]_ ;
  assign \new_[49859]_  = ~A300 & ~A299;
  assign \new_[49862]_  = ~A302 & ~A301;
  assign \new_[49863]_  = \new_[49862]_  & \new_[49859]_ ;
  assign \new_[49864]_  = \new_[49863]_  & \new_[49856]_ ;
  assign \new_[49868]_  = ~A199 & ~A168;
  assign \new_[49869]_  = A169 & \new_[49868]_ ;
  assign \new_[49873]_  = A202 & A201;
  assign \new_[49874]_  = A200 & \new_[49873]_ ;
  assign \new_[49875]_  = \new_[49874]_  & \new_[49869]_ ;
  assign \new_[49879]_  = ~A298 & A268;
  assign \new_[49880]_  = ~A267 & \new_[49879]_ ;
  assign \new_[49883]_  = ~A300 & A299;
  assign \new_[49886]_  = ~A302 & ~A301;
  assign \new_[49887]_  = \new_[49886]_  & \new_[49883]_ ;
  assign \new_[49888]_  = \new_[49887]_  & \new_[49880]_ ;
  assign \new_[49892]_  = ~A199 & ~A168;
  assign \new_[49893]_  = A169 & \new_[49892]_ ;
  assign \new_[49897]_  = A202 & A201;
  assign \new_[49898]_  = A200 & \new_[49897]_ ;
  assign \new_[49899]_  = \new_[49898]_  & \new_[49893]_ ;
  assign \new_[49903]_  = A298 & A269;
  assign \new_[49904]_  = ~A267 & \new_[49903]_ ;
  assign \new_[49907]_  = ~A300 & ~A299;
  assign \new_[49910]_  = ~A302 & ~A301;
  assign \new_[49911]_  = \new_[49910]_  & \new_[49907]_ ;
  assign \new_[49912]_  = \new_[49911]_  & \new_[49904]_ ;
  assign \new_[49916]_  = ~A199 & ~A168;
  assign \new_[49917]_  = A169 & \new_[49916]_ ;
  assign \new_[49921]_  = A202 & A201;
  assign \new_[49922]_  = A200 & \new_[49921]_ ;
  assign \new_[49923]_  = \new_[49922]_  & \new_[49917]_ ;
  assign \new_[49927]_  = ~A298 & A269;
  assign \new_[49928]_  = ~A267 & \new_[49927]_ ;
  assign \new_[49931]_  = ~A300 & A299;
  assign \new_[49934]_  = ~A302 & ~A301;
  assign \new_[49935]_  = \new_[49934]_  & \new_[49931]_ ;
  assign \new_[49936]_  = \new_[49935]_  & \new_[49928]_ ;
  assign \new_[49940]_  = ~A199 & ~A168;
  assign \new_[49941]_  = A169 & \new_[49940]_ ;
  assign \new_[49945]_  = A202 & A201;
  assign \new_[49946]_  = A200 & \new_[49945]_ ;
  assign \new_[49947]_  = \new_[49946]_  & \new_[49941]_ ;
  assign \new_[49951]_  = A298 & A266;
  assign \new_[49952]_  = A265 & \new_[49951]_ ;
  assign \new_[49955]_  = ~A300 & ~A299;
  assign \new_[49958]_  = ~A302 & ~A301;
  assign \new_[49959]_  = \new_[49958]_  & \new_[49955]_ ;
  assign \new_[49960]_  = \new_[49959]_  & \new_[49952]_ ;
  assign \new_[49964]_  = ~A199 & ~A168;
  assign \new_[49965]_  = A169 & \new_[49964]_ ;
  assign \new_[49969]_  = A202 & A201;
  assign \new_[49970]_  = A200 & \new_[49969]_ ;
  assign \new_[49971]_  = \new_[49970]_  & \new_[49965]_ ;
  assign \new_[49975]_  = ~A298 & A266;
  assign \new_[49976]_  = A265 & \new_[49975]_ ;
  assign \new_[49979]_  = ~A300 & A299;
  assign \new_[49982]_  = ~A302 & ~A301;
  assign \new_[49983]_  = \new_[49982]_  & \new_[49979]_ ;
  assign \new_[49984]_  = \new_[49983]_  & \new_[49976]_ ;
  assign \new_[49988]_  = ~A199 & ~A168;
  assign \new_[49989]_  = A169 & \new_[49988]_ ;
  assign \new_[49993]_  = A202 & A201;
  assign \new_[49994]_  = A200 & \new_[49993]_ ;
  assign \new_[49995]_  = \new_[49994]_  & \new_[49989]_ ;
  assign \new_[49999]_  = A298 & ~A266;
  assign \new_[50000]_  = ~A265 & \new_[49999]_ ;
  assign \new_[50003]_  = ~A300 & ~A299;
  assign \new_[50006]_  = ~A302 & ~A301;
  assign \new_[50007]_  = \new_[50006]_  & \new_[50003]_ ;
  assign \new_[50008]_  = \new_[50007]_  & \new_[50000]_ ;
  assign \new_[50012]_  = ~A199 & ~A168;
  assign \new_[50013]_  = A169 & \new_[50012]_ ;
  assign \new_[50017]_  = A202 & A201;
  assign \new_[50018]_  = A200 & \new_[50017]_ ;
  assign \new_[50019]_  = \new_[50018]_  & \new_[50013]_ ;
  assign \new_[50023]_  = ~A298 & ~A266;
  assign \new_[50024]_  = ~A265 & \new_[50023]_ ;
  assign \new_[50027]_  = ~A300 & A299;
  assign \new_[50030]_  = ~A302 & ~A301;
  assign \new_[50031]_  = \new_[50030]_  & \new_[50027]_ ;
  assign \new_[50032]_  = \new_[50031]_  & \new_[50024]_ ;
  assign \new_[50036]_  = ~A199 & ~A168;
  assign \new_[50037]_  = A169 & \new_[50036]_ ;
  assign \new_[50041]_  = A203 & A201;
  assign \new_[50042]_  = A200 & \new_[50041]_ ;
  assign \new_[50043]_  = \new_[50042]_  & \new_[50037]_ ;
  assign \new_[50047]_  = ~A269 & ~A268;
  assign \new_[50048]_  = A267 & \new_[50047]_ ;
  assign \new_[50051]_  = ~A299 & A298;
  assign \new_[50054]_  = A301 & A300;
  assign \new_[50055]_  = \new_[50054]_  & \new_[50051]_ ;
  assign \new_[50056]_  = \new_[50055]_  & \new_[50048]_ ;
  assign \new_[50060]_  = ~A199 & ~A168;
  assign \new_[50061]_  = A169 & \new_[50060]_ ;
  assign \new_[50065]_  = A203 & A201;
  assign \new_[50066]_  = A200 & \new_[50065]_ ;
  assign \new_[50067]_  = \new_[50066]_  & \new_[50061]_ ;
  assign \new_[50071]_  = ~A269 & ~A268;
  assign \new_[50072]_  = A267 & \new_[50071]_ ;
  assign \new_[50075]_  = ~A299 & A298;
  assign \new_[50078]_  = A302 & A300;
  assign \new_[50079]_  = \new_[50078]_  & \new_[50075]_ ;
  assign \new_[50080]_  = \new_[50079]_  & \new_[50072]_ ;
  assign \new_[50084]_  = ~A199 & ~A168;
  assign \new_[50085]_  = A169 & \new_[50084]_ ;
  assign \new_[50089]_  = A203 & A201;
  assign \new_[50090]_  = A200 & \new_[50089]_ ;
  assign \new_[50091]_  = \new_[50090]_  & \new_[50085]_ ;
  assign \new_[50095]_  = ~A269 & ~A268;
  assign \new_[50096]_  = A267 & \new_[50095]_ ;
  assign \new_[50099]_  = A299 & ~A298;
  assign \new_[50102]_  = A301 & A300;
  assign \new_[50103]_  = \new_[50102]_  & \new_[50099]_ ;
  assign \new_[50104]_  = \new_[50103]_  & \new_[50096]_ ;
  assign \new_[50108]_  = ~A199 & ~A168;
  assign \new_[50109]_  = A169 & \new_[50108]_ ;
  assign \new_[50113]_  = A203 & A201;
  assign \new_[50114]_  = A200 & \new_[50113]_ ;
  assign \new_[50115]_  = \new_[50114]_  & \new_[50109]_ ;
  assign \new_[50119]_  = ~A269 & ~A268;
  assign \new_[50120]_  = A267 & \new_[50119]_ ;
  assign \new_[50123]_  = A299 & ~A298;
  assign \new_[50126]_  = A302 & A300;
  assign \new_[50127]_  = \new_[50126]_  & \new_[50123]_ ;
  assign \new_[50128]_  = \new_[50127]_  & \new_[50120]_ ;
  assign \new_[50132]_  = ~A199 & ~A168;
  assign \new_[50133]_  = A169 & \new_[50132]_ ;
  assign \new_[50137]_  = A203 & A201;
  assign \new_[50138]_  = A200 & \new_[50137]_ ;
  assign \new_[50139]_  = \new_[50138]_  & \new_[50133]_ ;
  assign \new_[50143]_  = A298 & A268;
  assign \new_[50144]_  = ~A267 & \new_[50143]_ ;
  assign \new_[50147]_  = ~A300 & ~A299;
  assign \new_[50150]_  = ~A302 & ~A301;
  assign \new_[50151]_  = \new_[50150]_  & \new_[50147]_ ;
  assign \new_[50152]_  = \new_[50151]_  & \new_[50144]_ ;
  assign \new_[50156]_  = ~A199 & ~A168;
  assign \new_[50157]_  = A169 & \new_[50156]_ ;
  assign \new_[50161]_  = A203 & A201;
  assign \new_[50162]_  = A200 & \new_[50161]_ ;
  assign \new_[50163]_  = \new_[50162]_  & \new_[50157]_ ;
  assign \new_[50167]_  = ~A298 & A268;
  assign \new_[50168]_  = ~A267 & \new_[50167]_ ;
  assign \new_[50171]_  = ~A300 & A299;
  assign \new_[50174]_  = ~A302 & ~A301;
  assign \new_[50175]_  = \new_[50174]_  & \new_[50171]_ ;
  assign \new_[50176]_  = \new_[50175]_  & \new_[50168]_ ;
  assign \new_[50180]_  = ~A199 & ~A168;
  assign \new_[50181]_  = A169 & \new_[50180]_ ;
  assign \new_[50185]_  = A203 & A201;
  assign \new_[50186]_  = A200 & \new_[50185]_ ;
  assign \new_[50187]_  = \new_[50186]_  & \new_[50181]_ ;
  assign \new_[50191]_  = A298 & A269;
  assign \new_[50192]_  = ~A267 & \new_[50191]_ ;
  assign \new_[50195]_  = ~A300 & ~A299;
  assign \new_[50198]_  = ~A302 & ~A301;
  assign \new_[50199]_  = \new_[50198]_  & \new_[50195]_ ;
  assign \new_[50200]_  = \new_[50199]_  & \new_[50192]_ ;
  assign \new_[50204]_  = ~A199 & ~A168;
  assign \new_[50205]_  = A169 & \new_[50204]_ ;
  assign \new_[50209]_  = A203 & A201;
  assign \new_[50210]_  = A200 & \new_[50209]_ ;
  assign \new_[50211]_  = \new_[50210]_  & \new_[50205]_ ;
  assign \new_[50215]_  = ~A298 & A269;
  assign \new_[50216]_  = ~A267 & \new_[50215]_ ;
  assign \new_[50219]_  = ~A300 & A299;
  assign \new_[50222]_  = ~A302 & ~A301;
  assign \new_[50223]_  = \new_[50222]_  & \new_[50219]_ ;
  assign \new_[50224]_  = \new_[50223]_  & \new_[50216]_ ;
  assign \new_[50228]_  = ~A199 & ~A168;
  assign \new_[50229]_  = A169 & \new_[50228]_ ;
  assign \new_[50233]_  = A203 & A201;
  assign \new_[50234]_  = A200 & \new_[50233]_ ;
  assign \new_[50235]_  = \new_[50234]_  & \new_[50229]_ ;
  assign \new_[50239]_  = A298 & A266;
  assign \new_[50240]_  = A265 & \new_[50239]_ ;
  assign \new_[50243]_  = ~A300 & ~A299;
  assign \new_[50246]_  = ~A302 & ~A301;
  assign \new_[50247]_  = \new_[50246]_  & \new_[50243]_ ;
  assign \new_[50248]_  = \new_[50247]_  & \new_[50240]_ ;
  assign \new_[50252]_  = ~A199 & ~A168;
  assign \new_[50253]_  = A169 & \new_[50252]_ ;
  assign \new_[50257]_  = A203 & A201;
  assign \new_[50258]_  = A200 & \new_[50257]_ ;
  assign \new_[50259]_  = \new_[50258]_  & \new_[50253]_ ;
  assign \new_[50263]_  = ~A298 & A266;
  assign \new_[50264]_  = A265 & \new_[50263]_ ;
  assign \new_[50267]_  = ~A300 & A299;
  assign \new_[50270]_  = ~A302 & ~A301;
  assign \new_[50271]_  = \new_[50270]_  & \new_[50267]_ ;
  assign \new_[50272]_  = \new_[50271]_  & \new_[50264]_ ;
  assign \new_[50276]_  = ~A199 & ~A168;
  assign \new_[50277]_  = A169 & \new_[50276]_ ;
  assign \new_[50281]_  = A203 & A201;
  assign \new_[50282]_  = A200 & \new_[50281]_ ;
  assign \new_[50283]_  = \new_[50282]_  & \new_[50277]_ ;
  assign \new_[50287]_  = A298 & ~A266;
  assign \new_[50288]_  = ~A265 & \new_[50287]_ ;
  assign \new_[50291]_  = ~A300 & ~A299;
  assign \new_[50294]_  = ~A302 & ~A301;
  assign \new_[50295]_  = \new_[50294]_  & \new_[50291]_ ;
  assign \new_[50296]_  = \new_[50295]_  & \new_[50288]_ ;
  assign \new_[50300]_  = ~A199 & ~A168;
  assign \new_[50301]_  = A169 & \new_[50300]_ ;
  assign \new_[50305]_  = A203 & A201;
  assign \new_[50306]_  = A200 & \new_[50305]_ ;
  assign \new_[50307]_  = \new_[50306]_  & \new_[50301]_ ;
  assign \new_[50311]_  = ~A298 & ~A266;
  assign \new_[50312]_  = ~A265 & \new_[50311]_ ;
  assign \new_[50315]_  = ~A300 & A299;
  assign \new_[50318]_  = ~A302 & ~A301;
  assign \new_[50319]_  = \new_[50318]_  & \new_[50315]_ ;
  assign \new_[50320]_  = \new_[50319]_  & \new_[50312]_ ;
  assign \new_[50324]_  = ~A199 & ~A168;
  assign \new_[50325]_  = A169 & \new_[50324]_ ;
  assign \new_[50329]_  = ~A202 & ~A201;
  assign \new_[50330]_  = A200 & \new_[50329]_ ;
  assign \new_[50331]_  = \new_[50330]_  & \new_[50325]_ ;
  assign \new_[50335]_  = A268 & ~A267;
  assign \new_[50336]_  = ~A203 & \new_[50335]_ ;
  assign \new_[50339]_  = ~A299 & A298;
  assign \new_[50342]_  = A301 & A300;
  assign \new_[50343]_  = \new_[50342]_  & \new_[50339]_ ;
  assign \new_[50344]_  = \new_[50343]_  & \new_[50336]_ ;
  assign \new_[50348]_  = ~A199 & ~A168;
  assign \new_[50349]_  = A169 & \new_[50348]_ ;
  assign \new_[50353]_  = ~A202 & ~A201;
  assign \new_[50354]_  = A200 & \new_[50353]_ ;
  assign \new_[50355]_  = \new_[50354]_  & \new_[50349]_ ;
  assign \new_[50359]_  = A268 & ~A267;
  assign \new_[50360]_  = ~A203 & \new_[50359]_ ;
  assign \new_[50363]_  = ~A299 & A298;
  assign \new_[50366]_  = A302 & A300;
  assign \new_[50367]_  = \new_[50366]_  & \new_[50363]_ ;
  assign \new_[50368]_  = \new_[50367]_  & \new_[50360]_ ;
  assign \new_[50372]_  = ~A199 & ~A168;
  assign \new_[50373]_  = A169 & \new_[50372]_ ;
  assign \new_[50377]_  = ~A202 & ~A201;
  assign \new_[50378]_  = A200 & \new_[50377]_ ;
  assign \new_[50379]_  = \new_[50378]_  & \new_[50373]_ ;
  assign \new_[50383]_  = A268 & ~A267;
  assign \new_[50384]_  = ~A203 & \new_[50383]_ ;
  assign \new_[50387]_  = A299 & ~A298;
  assign \new_[50390]_  = A301 & A300;
  assign \new_[50391]_  = \new_[50390]_  & \new_[50387]_ ;
  assign \new_[50392]_  = \new_[50391]_  & \new_[50384]_ ;
  assign \new_[50396]_  = ~A199 & ~A168;
  assign \new_[50397]_  = A169 & \new_[50396]_ ;
  assign \new_[50401]_  = ~A202 & ~A201;
  assign \new_[50402]_  = A200 & \new_[50401]_ ;
  assign \new_[50403]_  = \new_[50402]_  & \new_[50397]_ ;
  assign \new_[50407]_  = A268 & ~A267;
  assign \new_[50408]_  = ~A203 & \new_[50407]_ ;
  assign \new_[50411]_  = A299 & ~A298;
  assign \new_[50414]_  = A302 & A300;
  assign \new_[50415]_  = \new_[50414]_  & \new_[50411]_ ;
  assign \new_[50416]_  = \new_[50415]_  & \new_[50408]_ ;
  assign \new_[50420]_  = ~A199 & ~A168;
  assign \new_[50421]_  = A169 & \new_[50420]_ ;
  assign \new_[50425]_  = ~A202 & ~A201;
  assign \new_[50426]_  = A200 & \new_[50425]_ ;
  assign \new_[50427]_  = \new_[50426]_  & \new_[50421]_ ;
  assign \new_[50431]_  = A269 & ~A267;
  assign \new_[50432]_  = ~A203 & \new_[50431]_ ;
  assign \new_[50435]_  = ~A299 & A298;
  assign \new_[50438]_  = A301 & A300;
  assign \new_[50439]_  = \new_[50438]_  & \new_[50435]_ ;
  assign \new_[50440]_  = \new_[50439]_  & \new_[50432]_ ;
  assign \new_[50444]_  = ~A199 & ~A168;
  assign \new_[50445]_  = A169 & \new_[50444]_ ;
  assign \new_[50449]_  = ~A202 & ~A201;
  assign \new_[50450]_  = A200 & \new_[50449]_ ;
  assign \new_[50451]_  = \new_[50450]_  & \new_[50445]_ ;
  assign \new_[50455]_  = A269 & ~A267;
  assign \new_[50456]_  = ~A203 & \new_[50455]_ ;
  assign \new_[50459]_  = ~A299 & A298;
  assign \new_[50462]_  = A302 & A300;
  assign \new_[50463]_  = \new_[50462]_  & \new_[50459]_ ;
  assign \new_[50464]_  = \new_[50463]_  & \new_[50456]_ ;
  assign \new_[50468]_  = ~A199 & ~A168;
  assign \new_[50469]_  = A169 & \new_[50468]_ ;
  assign \new_[50473]_  = ~A202 & ~A201;
  assign \new_[50474]_  = A200 & \new_[50473]_ ;
  assign \new_[50475]_  = \new_[50474]_  & \new_[50469]_ ;
  assign \new_[50479]_  = A269 & ~A267;
  assign \new_[50480]_  = ~A203 & \new_[50479]_ ;
  assign \new_[50483]_  = A299 & ~A298;
  assign \new_[50486]_  = A301 & A300;
  assign \new_[50487]_  = \new_[50486]_  & \new_[50483]_ ;
  assign \new_[50488]_  = \new_[50487]_  & \new_[50480]_ ;
  assign \new_[50492]_  = ~A199 & ~A168;
  assign \new_[50493]_  = A169 & \new_[50492]_ ;
  assign \new_[50497]_  = ~A202 & ~A201;
  assign \new_[50498]_  = A200 & \new_[50497]_ ;
  assign \new_[50499]_  = \new_[50498]_  & \new_[50493]_ ;
  assign \new_[50503]_  = A269 & ~A267;
  assign \new_[50504]_  = ~A203 & \new_[50503]_ ;
  assign \new_[50507]_  = A299 & ~A298;
  assign \new_[50510]_  = A302 & A300;
  assign \new_[50511]_  = \new_[50510]_  & \new_[50507]_ ;
  assign \new_[50512]_  = \new_[50511]_  & \new_[50504]_ ;
  assign \new_[50516]_  = ~A199 & ~A168;
  assign \new_[50517]_  = A169 & \new_[50516]_ ;
  assign \new_[50521]_  = ~A202 & ~A201;
  assign \new_[50522]_  = A200 & \new_[50521]_ ;
  assign \new_[50523]_  = \new_[50522]_  & \new_[50517]_ ;
  assign \new_[50527]_  = A266 & A265;
  assign \new_[50528]_  = ~A203 & \new_[50527]_ ;
  assign \new_[50531]_  = ~A299 & A298;
  assign \new_[50534]_  = A301 & A300;
  assign \new_[50535]_  = \new_[50534]_  & \new_[50531]_ ;
  assign \new_[50536]_  = \new_[50535]_  & \new_[50528]_ ;
  assign \new_[50540]_  = ~A199 & ~A168;
  assign \new_[50541]_  = A169 & \new_[50540]_ ;
  assign \new_[50545]_  = ~A202 & ~A201;
  assign \new_[50546]_  = A200 & \new_[50545]_ ;
  assign \new_[50547]_  = \new_[50546]_  & \new_[50541]_ ;
  assign \new_[50551]_  = A266 & A265;
  assign \new_[50552]_  = ~A203 & \new_[50551]_ ;
  assign \new_[50555]_  = ~A299 & A298;
  assign \new_[50558]_  = A302 & A300;
  assign \new_[50559]_  = \new_[50558]_  & \new_[50555]_ ;
  assign \new_[50560]_  = \new_[50559]_  & \new_[50552]_ ;
  assign \new_[50564]_  = ~A199 & ~A168;
  assign \new_[50565]_  = A169 & \new_[50564]_ ;
  assign \new_[50569]_  = ~A202 & ~A201;
  assign \new_[50570]_  = A200 & \new_[50569]_ ;
  assign \new_[50571]_  = \new_[50570]_  & \new_[50565]_ ;
  assign \new_[50575]_  = A266 & A265;
  assign \new_[50576]_  = ~A203 & \new_[50575]_ ;
  assign \new_[50579]_  = A299 & ~A298;
  assign \new_[50582]_  = A301 & A300;
  assign \new_[50583]_  = \new_[50582]_  & \new_[50579]_ ;
  assign \new_[50584]_  = \new_[50583]_  & \new_[50576]_ ;
  assign \new_[50588]_  = ~A199 & ~A168;
  assign \new_[50589]_  = A169 & \new_[50588]_ ;
  assign \new_[50593]_  = ~A202 & ~A201;
  assign \new_[50594]_  = A200 & \new_[50593]_ ;
  assign \new_[50595]_  = \new_[50594]_  & \new_[50589]_ ;
  assign \new_[50599]_  = A266 & A265;
  assign \new_[50600]_  = ~A203 & \new_[50599]_ ;
  assign \new_[50603]_  = A299 & ~A298;
  assign \new_[50606]_  = A302 & A300;
  assign \new_[50607]_  = \new_[50606]_  & \new_[50603]_ ;
  assign \new_[50608]_  = \new_[50607]_  & \new_[50600]_ ;
  assign \new_[50612]_  = ~A199 & ~A168;
  assign \new_[50613]_  = A169 & \new_[50612]_ ;
  assign \new_[50617]_  = ~A202 & ~A201;
  assign \new_[50618]_  = A200 & \new_[50617]_ ;
  assign \new_[50619]_  = \new_[50618]_  & \new_[50613]_ ;
  assign \new_[50623]_  = ~A266 & ~A265;
  assign \new_[50624]_  = ~A203 & \new_[50623]_ ;
  assign \new_[50627]_  = ~A299 & A298;
  assign \new_[50630]_  = A301 & A300;
  assign \new_[50631]_  = \new_[50630]_  & \new_[50627]_ ;
  assign \new_[50632]_  = \new_[50631]_  & \new_[50624]_ ;
  assign \new_[50636]_  = ~A199 & ~A168;
  assign \new_[50637]_  = A169 & \new_[50636]_ ;
  assign \new_[50641]_  = ~A202 & ~A201;
  assign \new_[50642]_  = A200 & \new_[50641]_ ;
  assign \new_[50643]_  = \new_[50642]_  & \new_[50637]_ ;
  assign \new_[50647]_  = ~A266 & ~A265;
  assign \new_[50648]_  = ~A203 & \new_[50647]_ ;
  assign \new_[50651]_  = ~A299 & A298;
  assign \new_[50654]_  = A302 & A300;
  assign \new_[50655]_  = \new_[50654]_  & \new_[50651]_ ;
  assign \new_[50656]_  = \new_[50655]_  & \new_[50648]_ ;
  assign \new_[50660]_  = ~A199 & ~A168;
  assign \new_[50661]_  = A169 & \new_[50660]_ ;
  assign \new_[50665]_  = ~A202 & ~A201;
  assign \new_[50666]_  = A200 & \new_[50665]_ ;
  assign \new_[50667]_  = \new_[50666]_  & \new_[50661]_ ;
  assign \new_[50671]_  = ~A266 & ~A265;
  assign \new_[50672]_  = ~A203 & \new_[50671]_ ;
  assign \new_[50675]_  = A299 & ~A298;
  assign \new_[50678]_  = A301 & A300;
  assign \new_[50679]_  = \new_[50678]_  & \new_[50675]_ ;
  assign \new_[50680]_  = \new_[50679]_  & \new_[50672]_ ;
  assign \new_[50684]_  = ~A199 & ~A168;
  assign \new_[50685]_  = A169 & \new_[50684]_ ;
  assign \new_[50689]_  = ~A202 & ~A201;
  assign \new_[50690]_  = A200 & \new_[50689]_ ;
  assign \new_[50691]_  = \new_[50690]_  & \new_[50685]_ ;
  assign \new_[50695]_  = ~A266 & ~A265;
  assign \new_[50696]_  = ~A203 & \new_[50695]_ ;
  assign \new_[50699]_  = A299 & ~A298;
  assign \new_[50702]_  = A302 & A300;
  assign \new_[50703]_  = \new_[50702]_  & \new_[50699]_ ;
  assign \new_[50704]_  = \new_[50703]_  & \new_[50696]_ ;
  assign \new_[50708]_  = A199 & ~A168;
  assign \new_[50709]_  = A169 & \new_[50708]_ ;
  assign \new_[50713]_  = A202 & A201;
  assign \new_[50714]_  = ~A200 & \new_[50713]_ ;
  assign \new_[50715]_  = \new_[50714]_  & \new_[50709]_ ;
  assign \new_[50719]_  = ~A269 & ~A268;
  assign \new_[50720]_  = A267 & \new_[50719]_ ;
  assign \new_[50723]_  = ~A299 & A298;
  assign \new_[50726]_  = A301 & A300;
  assign \new_[50727]_  = \new_[50726]_  & \new_[50723]_ ;
  assign \new_[50728]_  = \new_[50727]_  & \new_[50720]_ ;
  assign \new_[50732]_  = A199 & ~A168;
  assign \new_[50733]_  = A169 & \new_[50732]_ ;
  assign \new_[50737]_  = A202 & A201;
  assign \new_[50738]_  = ~A200 & \new_[50737]_ ;
  assign \new_[50739]_  = \new_[50738]_  & \new_[50733]_ ;
  assign \new_[50743]_  = ~A269 & ~A268;
  assign \new_[50744]_  = A267 & \new_[50743]_ ;
  assign \new_[50747]_  = ~A299 & A298;
  assign \new_[50750]_  = A302 & A300;
  assign \new_[50751]_  = \new_[50750]_  & \new_[50747]_ ;
  assign \new_[50752]_  = \new_[50751]_  & \new_[50744]_ ;
  assign \new_[50756]_  = A199 & ~A168;
  assign \new_[50757]_  = A169 & \new_[50756]_ ;
  assign \new_[50761]_  = A202 & A201;
  assign \new_[50762]_  = ~A200 & \new_[50761]_ ;
  assign \new_[50763]_  = \new_[50762]_  & \new_[50757]_ ;
  assign \new_[50767]_  = ~A269 & ~A268;
  assign \new_[50768]_  = A267 & \new_[50767]_ ;
  assign \new_[50771]_  = A299 & ~A298;
  assign \new_[50774]_  = A301 & A300;
  assign \new_[50775]_  = \new_[50774]_  & \new_[50771]_ ;
  assign \new_[50776]_  = \new_[50775]_  & \new_[50768]_ ;
  assign \new_[50780]_  = A199 & ~A168;
  assign \new_[50781]_  = A169 & \new_[50780]_ ;
  assign \new_[50785]_  = A202 & A201;
  assign \new_[50786]_  = ~A200 & \new_[50785]_ ;
  assign \new_[50787]_  = \new_[50786]_  & \new_[50781]_ ;
  assign \new_[50791]_  = ~A269 & ~A268;
  assign \new_[50792]_  = A267 & \new_[50791]_ ;
  assign \new_[50795]_  = A299 & ~A298;
  assign \new_[50798]_  = A302 & A300;
  assign \new_[50799]_  = \new_[50798]_  & \new_[50795]_ ;
  assign \new_[50800]_  = \new_[50799]_  & \new_[50792]_ ;
  assign \new_[50804]_  = A199 & ~A168;
  assign \new_[50805]_  = A169 & \new_[50804]_ ;
  assign \new_[50809]_  = A202 & A201;
  assign \new_[50810]_  = ~A200 & \new_[50809]_ ;
  assign \new_[50811]_  = \new_[50810]_  & \new_[50805]_ ;
  assign \new_[50815]_  = A298 & A268;
  assign \new_[50816]_  = ~A267 & \new_[50815]_ ;
  assign \new_[50819]_  = ~A300 & ~A299;
  assign \new_[50822]_  = ~A302 & ~A301;
  assign \new_[50823]_  = \new_[50822]_  & \new_[50819]_ ;
  assign \new_[50824]_  = \new_[50823]_  & \new_[50816]_ ;
  assign \new_[50828]_  = A199 & ~A168;
  assign \new_[50829]_  = A169 & \new_[50828]_ ;
  assign \new_[50833]_  = A202 & A201;
  assign \new_[50834]_  = ~A200 & \new_[50833]_ ;
  assign \new_[50835]_  = \new_[50834]_  & \new_[50829]_ ;
  assign \new_[50839]_  = ~A298 & A268;
  assign \new_[50840]_  = ~A267 & \new_[50839]_ ;
  assign \new_[50843]_  = ~A300 & A299;
  assign \new_[50846]_  = ~A302 & ~A301;
  assign \new_[50847]_  = \new_[50846]_  & \new_[50843]_ ;
  assign \new_[50848]_  = \new_[50847]_  & \new_[50840]_ ;
  assign \new_[50852]_  = A199 & ~A168;
  assign \new_[50853]_  = A169 & \new_[50852]_ ;
  assign \new_[50857]_  = A202 & A201;
  assign \new_[50858]_  = ~A200 & \new_[50857]_ ;
  assign \new_[50859]_  = \new_[50858]_  & \new_[50853]_ ;
  assign \new_[50863]_  = A298 & A269;
  assign \new_[50864]_  = ~A267 & \new_[50863]_ ;
  assign \new_[50867]_  = ~A300 & ~A299;
  assign \new_[50870]_  = ~A302 & ~A301;
  assign \new_[50871]_  = \new_[50870]_  & \new_[50867]_ ;
  assign \new_[50872]_  = \new_[50871]_  & \new_[50864]_ ;
  assign \new_[50876]_  = A199 & ~A168;
  assign \new_[50877]_  = A169 & \new_[50876]_ ;
  assign \new_[50881]_  = A202 & A201;
  assign \new_[50882]_  = ~A200 & \new_[50881]_ ;
  assign \new_[50883]_  = \new_[50882]_  & \new_[50877]_ ;
  assign \new_[50887]_  = ~A298 & A269;
  assign \new_[50888]_  = ~A267 & \new_[50887]_ ;
  assign \new_[50891]_  = ~A300 & A299;
  assign \new_[50894]_  = ~A302 & ~A301;
  assign \new_[50895]_  = \new_[50894]_  & \new_[50891]_ ;
  assign \new_[50896]_  = \new_[50895]_  & \new_[50888]_ ;
  assign \new_[50900]_  = A199 & ~A168;
  assign \new_[50901]_  = A169 & \new_[50900]_ ;
  assign \new_[50905]_  = A202 & A201;
  assign \new_[50906]_  = ~A200 & \new_[50905]_ ;
  assign \new_[50907]_  = \new_[50906]_  & \new_[50901]_ ;
  assign \new_[50911]_  = A298 & A266;
  assign \new_[50912]_  = A265 & \new_[50911]_ ;
  assign \new_[50915]_  = ~A300 & ~A299;
  assign \new_[50918]_  = ~A302 & ~A301;
  assign \new_[50919]_  = \new_[50918]_  & \new_[50915]_ ;
  assign \new_[50920]_  = \new_[50919]_  & \new_[50912]_ ;
  assign \new_[50924]_  = A199 & ~A168;
  assign \new_[50925]_  = A169 & \new_[50924]_ ;
  assign \new_[50929]_  = A202 & A201;
  assign \new_[50930]_  = ~A200 & \new_[50929]_ ;
  assign \new_[50931]_  = \new_[50930]_  & \new_[50925]_ ;
  assign \new_[50935]_  = ~A298 & A266;
  assign \new_[50936]_  = A265 & \new_[50935]_ ;
  assign \new_[50939]_  = ~A300 & A299;
  assign \new_[50942]_  = ~A302 & ~A301;
  assign \new_[50943]_  = \new_[50942]_  & \new_[50939]_ ;
  assign \new_[50944]_  = \new_[50943]_  & \new_[50936]_ ;
  assign \new_[50948]_  = A199 & ~A168;
  assign \new_[50949]_  = A169 & \new_[50948]_ ;
  assign \new_[50953]_  = A202 & A201;
  assign \new_[50954]_  = ~A200 & \new_[50953]_ ;
  assign \new_[50955]_  = \new_[50954]_  & \new_[50949]_ ;
  assign \new_[50959]_  = A298 & ~A266;
  assign \new_[50960]_  = ~A265 & \new_[50959]_ ;
  assign \new_[50963]_  = ~A300 & ~A299;
  assign \new_[50966]_  = ~A302 & ~A301;
  assign \new_[50967]_  = \new_[50966]_  & \new_[50963]_ ;
  assign \new_[50968]_  = \new_[50967]_  & \new_[50960]_ ;
  assign \new_[50972]_  = A199 & ~A168;
  assign \new_[50973]_  = A169 & \new_[50972]_ ;
  assign \new_[50977]_  = A202 & A201;
  assign \new_[50978]_  = ~A200 & \new_[50977]_ ;
  assign \new_[50979]_  = \new_[50978]_  & \new_[50973]_ ;
  assign \new_[50983]_  = ~A298 & ~A266;
  assign \new_[50984]_  = ~A265 & \new_[50983]_ ;
  assign \new_[50987]_  = ~A300 & A299;
  assign \new_[50990]_  = ~A302 & ~A301;
  assign \new_[50991]_  = \new_[50990]_  & \new_[50987]_ ;
  assign \new_[50992]_  = \new_[50991]_  & \new_[50984]_ ;
  assign \new_[50996]_  = A199 & ~A168;
  assign \new_[50997]_  = A169 & \new_[50996]_ ;
  assign \new_[51001]_  = A203 & A201;
  assign \new_[51002]_  = ~A200 & \new_[51001]_ ;
  assign \new_[51003]_  = \new_[51002]_  & \new_[50997]_ ;
  assign \new_[51007]_  = ~A269 & ~A268;
  assign \new_[51008]_  = A267 & \new_[51007]_ ;
  assign \new_[51011]_  = ~A299 & A298;
  assign \new_[51014]_  = A301 & A300;
  assign \new_[51015]_  = \new_[51014]_  & \new_[51011]_ ;
  assign \new_[51016]_  = \new_[51015]_  & \new_[51008]_ ;
  assign \new_[51020]_  = A199 & ~A168;
  assign \new_[51021]_  = A169 & \new_[51020]_ ;
  assign \new_[51025]_  = A203 & A201;
  assign \new_[51026]_  = ~A200 & \new_[51025]_ ;
  assign \new_[51027]_  = \new_[51026]_  & \new_[51021]_ ;
  assign \new_[51031]_  = ~A269 & ~A268;
  assign \new_[51032]_  = A267 & \new_[51031]_ ;
  assign \new_[51035]_  = ~A299 & A298;
  assign \new_[51038]_  = A302 & A300;
  assign \new_[51039]_  = \new_[51038]_  & \new_[51035]_ ;
  assign \new_[51040]_  = \new_[51039]_  & \new_[51032]_ ;
  assign \new_[51044]_  = A199 & ~A168;
  assign \new_[51045]_  = A169 & \new_[51044]_ ;
  assign \new_[51049]_  = A203 & A201;
  assign \new_[51050]_  = ~A200 & \new_[51049]_ ;
  assign \new_[51051]_  = \new_[51050]_  & \new_[51045]_ ;
  assign \new_[51055]_  = ~A269 & ~A268;
  assign \new_[51056]_  = A267 & \new_[51055]_ ;
  assign \new_[51059]_  = A299 & ~A298;
  assign \new_[51062]_  = A301 & A300;
  assign \new_[51063]_  = \new_[51062]_  & \new_[51059]_ ;
  assign \new_[51064]_  = \new_[51063]_  & \new_[51056]_ ;
  assign \new_[51068]_  = A199 & ~A168;
  assign \new_[51069]_  = A169 & \new_[51068]_ ;
  assign \new_[51073]_  = A203 & A201;
  assign \new_[51074]_  = ~A200 & \new_[51073]_ ;
  assign \new_[51075]_  = \new_[51074]_  & \new_[51069]_ ;
  assign \new_[51079]_  = ~A269 & ~A268;
  assign \new_[51080]_  = A267 & \new_[51079]_ ;
  assign \new_[51083]_  = A299 & ~A298;
  assign \new_[51086]_  = A302 & A300;
  assign \new_[51087]_  = \new_[51086]_  & \new_[51083]_ ;
  assign \new_[51088]_  = \new_[51087]_  & \new_[51080]_ ;
  assign \new_[51092]_  = A199 & ~A168;
  assign \new_[51093]_  = A169 & \new_[51092]_ ;
  assign \new_[51097]_  = A203 & A201;
  assign \new_[51098]_  = ~A200 & \new_[51097]_ ;
  assign \new_[51099]_  = \new_[51098]_  & \new_[51093]_ ;
  assign \new_[51103]_  = A298 & A268;
  assign \new_[51104]_  = ~A267 & \new_[51103]_ ;
  assign \new_[51107]_  = ~A300 & ~A299;
  assign \new_[51110]_  = ~A302 & ~A301;
  assign \new_[51111]_  = \new_[51110]_  & \new_[51107]_ ;
  assign \new_[51112]_  = \new_[51111]_  & \new_[51104]_ ;
  assign \new_[51116]_  = A199 & ~A168;
  assign \new_[51117]_  = A169 & \new_[51116]_ ;
  assign \new_[51121]_  = A203 & A201;
  assign \new_[51122]_  = ~A200 & \new_[51121]_ ;
  assign \new_[51123]_  = \new_[51122]_  & \new_[51117]_ ;
  assign \new_[51127]_  = ~A298 & A268;
  assign \new_[51128]_  = ~A267 & \new_[51127]_ ;
  assign \new_[51131]_  = ~A300 & A299;
  assign \new_[51134]_  = ~A302 & ~A301;
  assign \new_[51135]_  = \new_[51134]_  & \new_[51131]_ ;
  assign \new_[51136]_  = \new_[51135]_  & \new_[51128]_ ;
  assign \new_[51140]_  = A199 & ~A168;
  assign \new_[51141]_  = A169 & \new_[51140]_ ;
  assign \new_[51145]_  = A203 & A201;
  assign \new_[51146]_  = ~A200 & \new_[51145]_ ;
  assign \new_[51147]_  = \new_[51146]_  & \new_[51141]_ ;
  assign \new_[51151]_  = A298 & A269;
  assign \new_[51152]_  = ~A267 & \new_[51151]_ ;
  assign \new_[51155]_  = ~A300 & ~A299;
  assign \new_[51158]_  = ~A302 & ~A301;
  assign \new_[51159]_  = \new_[51158]_  & \new_[51155]_ ;
  assign \new_[51160]_  = \new_[51159]_  & \new_[51152]_ ;
  assign \new_[51164]_  = A199 & ~A168;
  assign \new_[51165]_  = A169 & \new_[51164]_ ;
  assign \new_[51169]_  = A203 & A201;
  assign \new_[51170]_  = ~A200 & \new_[51169]_ ;
  assign \new_[51171]_  = \new_[51170]_  & \new_[51165]_ ;
  assign \new_[51175]_  = ~A298 & A269;
  assign \new_[51176]_  = ~A267 & \new_[51175]_ ;
  assign \new_[51179]_  = ~A300 & A299;
  assign \new_[51182]_  = ~A302 & ~A301;
  assign \new_[51183]_  = \new_[51182]_  & \new_[51179]_ ;
  assign \new_[51184]_  = \new_[51183]_  & \new_[51176]_ ;
  assign \new_[51188]_  = A199 & ~A168;
  assign \new_[51189]_  = A169 & \new_[51188]_ ;
  assign \new_[51193]_  = A203 & A201;
  assign \new_[51194]_  = ~A200 & \new_[51193]_ ;
  assign \new_[51195]_  = \new_[51194]_  & \new_[51189]_ ;
  assign \new_[51199]_  = A298 & A266;
  assign \new_[51200]_  = A265 & \new_[51199]_ ;
  assign \new_[51203]_  = ~A300 & ~A299;
  assign \new_[51206]_  = ~A302 & ~A301;
  assign \new_[51207]_  = \new_[51206]_  & \new_[51203]_ ;
  assign \new_[51208]_  = \new_[51207]_  & \new_[51200]_ ;
  assign \new_[51212]_  = A199 & ~A168;
  assign \new_[51213]_  = A169 & \new_[51212]_ ;
  assign \new_[51217]_  = A203 & A201;
  assign \new_[51218]_  = ~A200 & \new_[51217]_ ;
  assign \new_[51219]_  = \new_[51218]_  & \new_[51213]_ ;
  assign \new_[51223]_  = ~A298 & A266;
  assign \new_[51224]_  = A265 & \new_[51223]_ ;
  assign \new_[51227]_  = ~A300 & A299;
  assign \new_[51230]_  = ~A302 & ~A301;
  assign \new_[51231]_  = \new_[51230]_  & \new_[51227]_ ;
  assign \new_[51232]_  = \new_[51231]_  & \new_[51224]_ ;
  assign \new_[51236]_  = A199 & ~A168;
  assign \new_[51237]_  = A169 & \new_[51236]_ ;
  assign \new_[51241]_  = A203 & A201;
  assign \new_[51242]_  = ~A200 & \new_[51241]_ ;
  assign \new_[51243]_  = \new_[51242]_  & \new_[51237]_ ;
  assign \new_[51247]_  = A298 & ~A266;
  assign \new_[51248]_  = ~A265 & \new_[51247]_ ;
  assign \new_[51251]_  = ~A300 & ~A299;
  assign \new_[51254]_  = ~A302 & ~A301;
  assign \new_[51255]_  = \new_[51254]_  & \new_[51251]_ ;
  assign \new_[51256]_  = \new_[51255]_  & \new_[51248]_ ;
  assign \new_[51260]_  = A199 & ~A168;
  assign \new_[51261]_  = A169 & \new_[51260]_ ;
  assign \new_[51265]_  = A203 & A201;
  assign \new_[51266]_  = ~A200 & \new_[51265]_ ;
  assign \new_[51267]_  = \new_[51266]_  & \new_[51261]_ ;
  assign \new_[51271]_  = ~A298 & ~A266;
  assign \new_[51272]_  = ~A265 & \new_[51271]_ ;
  assign \new_[51275]_  = ~A300 & A299;
  assign \new_[51278]_  = ~A302 & ~A301;
  assign \new_[51279]_  = \new_[51278]_  & \new_[51275]_ ;
  assign \new_[51280]_  = \new_[51279]_  & \new_[51272]_ ;
  assign \new_[51284]_  = A199 & ~A168;
  assign \new_[51285]_  = A169 & \new_[51284]_ ;
  assign \new_[51289]_  = ~A202 & ~A201;
  assign \new_[51290]_  = ~A200 & \new_[51289]_ ;
  assign \new_[51291]_  = \new_[51290]_  & \new_[51285]_ ;
  assign \new_[51295]_  = A268 & ~A267;
  assign \new_[51296]_  = ~A203 & \new_[51295]_ ;
  assign \new_[51299]_  = ~A299 & A298;
  assign \new_[51302]_  = A301 & A300;
  assign \new_[51303]_  = \new_[51302]_  & \new_[51299]_ ;
  assign \new_[51304]_  = \new_[51303]_  & \new_[51296]_ ;
  assign \new_[51308]_  = A199 & ~A168;
  assign \new_[51309]_  = A169 & \new_[51308]_ ;
  assign \new_[51313]_  = ~A202 & ~A201;
  assign \new_[51314]_  = ~A200 & \new_[51313]_ ;
  assign \new_[51315]_  = \new_[51314]_  & \new_[51309]_ ;
  assign \new_[51319]_  = A268 & ~A267;
  assign \new_[51320]_  = ~A203 & \new_[51319]_ ;
  assign \new_[51323]_  = ~A299 & A298;
  assign \new_[51326]_  = A302 & A300;
  assign \new_[51327]_  = \new_[51326]_  & \new_[51323]_ ;
  assign \new_[51328]_  = \new_[51327]_  & \new_[51320]_ ;
  assign \new_[51332]_  = A199 & ~A168;
  assign \new_[51333]_  = A169 & \new_[51332]_ ;
  assign \new_[51337]_  = ~A202 & ~A201;
  assign \new_[51338]_  = ~A200 & \new_[51337]_ ;
  assign \new_[51339]_  = \new_[51338]_  & \new_[51333]_ ;
  assign \new_[51343]_  = A268 & ~A267;
  assign \new_[51344]_  = ~A203 & \new_[51343]_ ;
  assign \new_[51347]_  = A299 & ~A298;
  assign \new_[51350]_  = A301 & A300;
  assign \new_[51351]_  = \new_[51350]_  & \new_[51347]_ ;
  assign \new_[51352]_  = \new_[51351]_  & \new_[51344]_ ;
  assign \new_[51356]_  = A199 & ~A168;
  assign \new_[51357]_  = A169 & \new_[51356]_ ;
  assign \new_[51361]_  = ~A202 & ~A201;
  assign \new_[51362]_  = ~A200 & \new_[51361]_ ;
  assign \new_[51363]_  = \new_[51362]_  & \new_[51357]_ ;
  assign \new_[51367]_  = A268 & ~A267;
  assign \new_[51368]_  = ~A203 & \new_[51367]_ ;
  assign \new_[51371]_  = A299 & ~A298;
  assign \new_[51374]_  = A302 & A300;
  assign \new_[51375]_  = \new_[51374]_  & \new_[51371]_ ;
  assign \new_[51376]_  = \new_[51375]_  & \new_[51368]_ ;
  assign \new_[51380]_  = A199 & ~A168;
  assign \new_[51381]_  = A169 & \new_[51380]_ ;
  assign \new_[51385]_  = ~A202 & ~A201;
  assign \new_[51386]_  = ~A200 & \new_[51385]_ ;
  assign \new_[51387]_  = \new_[51386]_  & \new_[51381]_ ;
  assign \new_[51391]_  = A269 & ~A267;
  assign \new_[51392]_  = ~A203 & \new_[51391]_ ;
  assign \new_[51395]_  = ~A299 & A298;
  assign \new_[51398]_  = A301 & A300;
  assign \new_[51399]_  = \new_[51398]_  & \new_[51395]_ ;
  assign \new_[51400]_  = \new_[51399]_  & \new_[51392]_ ;
  assign \new_[51404]_  = A199 & ~A168;
  assign \new_[51405]_  = A169 & \new_[51404]_ ;
  assign \new_[51409]_  = ~A202 & ~A201;
  assign \new_[51410]_  = ~A200 & \new_[51409]_ ;
  assign \new_[51411]_  = \new_[51410]_  & \new_[51405]_ ;
  assign \new_[51415]_  = A269 & ~A267;
  assign \new_[51416]_  = ~A203 & \new_[51415]_ ;
  assign \new_[51419]_  = ~A299 & A298;
  assign \new_[51422]_  = A302 & A300;
  assign \new_[51423]_  = \new_[51422]_  & \new_[51419]_ ;
  assign \new_[51424]_  = \new_[51423]_  & \new_[51416]_ ;
  assign \new_[51428]_  = A199 & ~A168;
  assign \new_[51429]_  = A169 & \new_[51428]_ ;
  assign \new_[51433]_  = ~A202 & ~A201;
  assign \new_[51434]_  = ~A200 & \new_[51433]_ ;
  assign \new_[51435]_  = \new_[51434]_  & \new_[51429]_ ;
  assign \new_[51439]_  = A269 & ~A267;
  assign \new_[51440]_  = ~A203 & \new_[51439]_ ;
  assign \new_[51443]_  = A299 & ~A298;
  assign \new_[51446]_  = A301 & A300;
  assign \new_[51447]_  = \new_[51446]_  & \new_[51443]_ ;
  assign \new_[51448]_  = \new_[51447]_  & \new_[51440]_ ;
  assign \new_[51452]_  = A199 & ~A168;
  assign \new_[51453]_  = A169 & \new_[51452]_ ;
  assign \new_[51457]_  = ~A202 & ~A201;
  assign \new_[51458]_  = ~A200 & \new_[51457]_ ;
  assign \new_[51459]_  = \new_[51458]_  & \new_[51453]_ ;
  assign \new_[51463]_  = A269 & ~A267;
  assign \new_[51464]_  = ~A203 & \new_[51463]_ ;
  assign \new_[51467]_  = A299 & ~A298;
  assign \new_[51470]_  = A302 & A300;
  assign \new_[51471]_  = \new_[51470]_  & \new_[51467]_ ;
  assign \new_[51472]_  = \new_[51471]_  & \new_[51464]_ ;
  assign \new_[51476]_  = A199 & ~A168;
  assign \new_[51477]_  = A169 & \new_[51476]_ ;
  assign \new_[51481]_  = ~A202 & ~A201;
  assign \new_[51482]_  = ~A200 & \new_[51481]_ ;
  assign \new_[51483]_  = \new_[51482]_  & \new_[51477]_ ;
  assign \new_[51487]_  = A266 & A265;
  assign \new_[51488]_  = ~A203 & \new_[51487]_ ;
  assign \new_[51491]_  = ~A299 & A298;
  assign \new_[51494]_  = A301 & A300;
  assign \new_[51495]_  = \new_[51494]_  & \new_[51491]_ ;
  assign \new_[51496]_  = \new_[51495]_  & \new_[51488]_ ;
  assign \new_[51500]_  = A199 & ~A168;
  assign \new_[51501]_  = A169 & \new_[51500]_ ;
  assign \new_[51505]_  = ~A202 & ~A201;
  assign \new_[51506]_  = ~A200 & \new_[51505]_ ;
  assign \new_[51507]_  = \new_[51506]_  & \new_[51501]_ ;
  assign \new_[51511]_  = A266 & A265;
  assign \new_[51512]_  = ~A203 & \new_[51511]_ ;
  assign \new_[51515]_  = ~A299 & A298;
  assign \new_[51518]_  = A302 & A300;
  assign \new_[51519]_  = \new_[51518]_  & \new_[51515]_ ;
  assign \new_[51520]_  = \new_[51519]_  & \new_[51512]_ ;
  assign \new_[51524]_  = A199 & ~A168;
  assign \new_[51525]_  = A169 & \new_[51524]_ ;
  assign \new_[51529]_  = ~A202 & ~A201;
  assign \new_[51530]_  = ~A200 & \new_[51529]_ ;
  assign \new_[51531]_  = \new_[51530]_  & \new_[51525]_ ;
  assign \new_[51535]_  = A266 & A265;
  assign \new_[51536]_  = ~A203 & \new_[51535]_ ;
  assign \new_[51539]_  = A299 & ~A298;
  assign \new_[51542]_  = A301 & A300;
  assign \new_[51543]_  = \new_[51542]_  & \new_[51539]_ ;
  assign \new_[51544]_  = \new_[51543]_  & \new_[51536]_ ;
  assign \new_[51548]_  = A199 & ~A168;
  assign \new_[51549]_  = A169 & \new_[51548]_ ;
  assign \new_[51553]_  = ~A202 & ~A201;
  assign \new_[51554]_  = ~A200 & \new_[51553]_ ;
  assign \new_[51555]_  = \new_[51554]_  & \new_[51549]_ ;
  assign \new_[51559]_  = A266 & A265;
  assign \new_[51560]_  = ~A203 & \new_[51559]_ ;
  assign \new_[51563]_  = A299 & ~A298;
  assign \new_[51566]_  = A302 & A300;
  assign \new_[51567]_  = \new_[51566]_  & \new_[51563]_ ;
  assign \new_[51568]_  = \new_[51567]_  & \new_[51560]_ ;
  assign \new_[51572]_  = A199 & ~A168;
  assign \new_[51573]_  = A169 & \new_[51572]_ ;
  assign \new_[51577]_  = ~A202 & ~A201;
  assign \new_[51578]_  = ~A200 & \new_[51577]_ ;
  assign \new_[51579]_  = \new_[51578]_  & \new_[51573]_ ;
  assign \new_[51583]_  = ~A266 & ~A265;
  assign \new_[51584]_  = ~A203 & \new_[51583]_ ;
  assign \new_[51587]_  = ~A299 & A298;
  assign \new_[51590]_  = A301 & A300;
  assign \new_[51591]_  = \new_[51590]_  & \new_[51587]_ ;
  assign \new_[51592]_  = \new_[51591]_  & \new_[51584]_ ;
  assign \new_[51596]_  = A199 & ~A168;
  assign \new_[51597]_  = A169 & \new_[51596]_ ;
  assign \new_[51601]_  = ~A202 & ~A201;
  assign \new_[51602]_  = ~A200 & \new_[51601]_ ;
  assign \new_[51603]_  = \new_[51602]_  & \new_[51597]_ ;
  assign \new_[51607]_  = ~A266 & ~A265;
  assign \new_[51608]_  = ~A203 & \new_[51607]_ ;
  assign \new_[51611]_  = ~A299 & A298;
  assign \new_[51614]_  = A302 & A300;
  assign \new_[51615]_  = \new_[51614]_  & \new_[51611]_ ;
  assign \new_[51616]_  = \new_[51615]_  & \new_[51608]_ ;
  assign \new_[51620]_  = A199 & ~A168;
  assign \new_[51621]_  = A169 & \new_[51620]_ ;
  assign \new_[51625]_  = ~A202 & ~A201;
  assign \new_[51626]_  = ~A200 & \new_[51625]_ ;
  assign \new_[51627]_  = \new_[51626]_  & \new_[51621]_ ;
  assign \new_[51631]_  = ~A266 & ~A265;
  assign \new_[51632]_  = ~A203 & \new_[51631]_ ;
  assign \new_[51635]_  = A299 & ~A298;
  assign \new_[51638]_  = A301 & A300;
  assign \new_[51639]_  = \new_[51638]_  & \new_[51635]_ ;
  assign \new_[51640]_  = \new_[51639]_  & \new_[51632]_ ;
  assign \new_[51644]_  = A199 & ~A168;
  assign \new_[51645]_  = A169 & \new_[51644]_ ;
  assign \new_[51649]_  = ~A202 & ~A201;
  assign \new_[51650]_  = ~A200 & \new_[51649]_ ;
  assign \new_[51651]_  = \new_[51650]_  & \new_[51645]_ ;
  assign \new_[51655]_  = ~A266 & ~A265;
  assign \new_[51656]_  = ~A203 & \new_[51655]_ ;
  assign \new_[51659]_  = A299 & ~A298;
  assign \new_[51662]_  = A302 & A300;
  assign \new_[51663]_  = \new_[51662]_  & \new_[51659]_ ;
  assign \new_[51664]_  = \new_[51663]_  & \new_[51656]_ ;
  assign \new_[51668]_  = A168 & ~A169;
  assign \new_[51669]_  = A170 & \new_[51668]_ ;
  assign \new_[51673]_  = ~A203 & ~A202;
  assign \new_[51674]_  = A201 & \new_[51673]_ ;
  assign \new_[51675]_  = \new_[51674]_  & \new_[51669]_ ;
  assign \new_[51679]_  = A267 & A266;
  assign \new_[51680]_  = ~A265 & \new_[51679]_ ;
  assign \new_[51683]_  = A300 & A268;
  assign \new_[51686]_  = ~A302 & ~A301;
  assign \new_[51687]_  = \new_[51686]_  & \new_[51683]_ ;
  assign \new_[51688]_  = \new_[51687]_  & \new_[51680]_ ;
  assign \new_[51692]_  = A168 & ~A169;
  assign \new_[51693]_  = A170 & \new_[51692]_ ;
  assign \new_[51697]_  = ~A203 & ~A202;
  assign \new_[51698]_  = A201 & \new_[51697]_ ;
  assign \new_[51699]_  = \new_[51698]_  & \new_[51693]_ ;
  assign \new_[51703]_  = A267 & A266;
  assign \new_[51704]_  = ~A265 & \new_[51703]_ ;
  assign \new_[51707]_  = A300 & A269;
  assign \new_[51710]_  = ~A302 & ~A301;
  assign \new_[51711]_  = \new_[51710]_  & \new_[51707]_ ;
  assign \new_[51712]_  = \new_[51711]_  & \new_[51704]_ ;
  assign \new_[51716]_  = A168 & ~A169;
  assign \new_[51717]_  = A170 & \new_[51716]_ ;
  assign \new_[51721]_  = ~A203 & ~A202;
  assign \new_[51722]_  = A201 & \new_[51721]_ ;
  assign \new_[51723]_  = \new_[51722]_  & \new_[51717]_ ;
  assign \new_[51727]_  = ~A267 & A266;
  assign \new_[51728]_  = ~A265 & \new_[51727]_ ;
  assign \new_[51731]_  = ~A269 & ~A268;
  assign \new_[51734]_  = A301 & ~A300;
  assign \new_[51735]_  = \new_[51734]_  & \new_[51731]_ ;
  assign \new_[51736]_  = \new_[51735]_  & \new_[51728]_ ;
  assign \new_[51740]_  = A168 & ~A169;
  assign \new_[51741]_  = A170 & \new_[51740]_ ;
  assign \new_[51745]_  = ~A203 & ~A202;
  assign \new_[51746]_  = A201 & \new_[51745]_ ;
  assign \new_[51747]_  = \new_[51746]_  & \new_[51741]_ ;
  assign \new_[51751]_  = ~A267 & A266;
  assign \new_[51752]_  = ~A265 & \new_[51751]_ ;
  assign \new_[51755]_  = ~A269 & ~A268;
  assign \new_[51758]_  = A302 & ~A300;
  assign \new_[51759]_  = \new_[51758]_  & \new_[51755]_ ;
  assign \new_[51760]_  = \new_[51759]_  & \new_[51752]_ ;
  assign \new_[51764]_  = A168 & ~A169;
  assign \new_[51765]_  = A170 & \new_[51764]_ ;
  assign \new_[51769]_  = ~A203 & ~A202;
  assign \new_[51770]_  = A201 & \new_[51769]_ ;
  assign \new_[51771]_  = \new_[51770]_  & \new_[51765]_ ;
  assign \new_[51775]_  = ~A267 & A266;
  assign \new_[51776]_  = ~A265 & \new_[51775]_ ;
  assign \new_[51779]_  = ~A269 & ~A268;
  assign \new_[51782]_  = A299 & A298;
  assign \new_[51783]_  = \new_[51782]_  & \new_[51779]_ ;
  assign \new_[51784]_  = \new_[51783]_  & \new_[51776]_ ;
  assign \new_[51788]_  = A168 & ~A169;
  assign \new_[51789]_  = A170 & \new_[51788]_ ;
  assign \new_[51793]_  = ~A203 & ~A202;
  assign \new_[51794]_  = A201 & \new_[51793]_ ;
  assign \new_[51795]_  = \new_[51794]_  & \new_[51789]_ ;
  assign \new_[51799]_  = ~A267 & A266;
  assign \new_[51800]_  = ~A265 & \new_[51799]_ ;
  assign \new_[51803]_  = ~A269 & ~A268;
  assign \new_[51806]_  = ~A299 & ~A298;
  assign \new_[51807]_  = \new_[51806]_  & \new_[51803]_ ;
  assign \new_[51808]_  = \new_[51807]_  & \new_[51800]_ ;
  assign \new_[51812]_  = A168 & ~A169;
  assign \new_[51813]_  = A170 & \new_[51812]_ ;
  assign \new_[51817]_  = ~A203 & ~A202;
  assign \new_[51818]_  = A201 & \new_[51817]_ ;
  assign \new_[51819]_  = \new_[51818]_  & \new_[51813]_ ;
  assign \new_[51823]_  = A267 & ~A266;
  assign \new_[51824]_  = A265 & \new_[51823]_ ;
  assign \new_[51827]_  = A300 & A268;
  assign \new_[51830]_  = ~A302 & ~A301;
  assign \new_[51831]_  = \new_[51830]_  & \new_[51827]_ ;
  assign \new_[51832]_  = \new_[51831]_  & \new_[51824]_ ;
  assign \new_[51836]_  = A168 & ~A169;
  assign \new_[51837]_  = A170 & \new_[51836]_ ;
  assign \new_[51841]_  = ~A203 & ~A202;
  assign \new_[51842]_  = A201 & \new_[51841]_ ;
  assign \new_[51843]_  = \new_[51842]_  & \new_[51837]_ ;
  assign \new_[51847]_  = A267 & ~A266;
  assign \new_[51848]_  = A265 & \new_[51847]_ ;
  assign \new_[51851]_  = A300 & A269;
  assign \new_[51854]_  = ~A302 & ~A301;
  assign \new_[51855]_  = \new_[51854]_  & \new_[51851]_ ;
  assign \new_[51856]_  = \new_[51855]_  & \new_[51848]_ ;
  assign \new_[51860]_  = A168 & ~A169;
  assign \new_[51861]_  = A170 & \new_[51860]_ ;
  assign \new_[51865]_  = ~A203 & ~A202;
  assign \new_[51866]_  = A201 & \new_[51865]_ ;
  assign \new_[51867]_  = \new_[51866]_  & \new_[51861]_ ;
  assign \new_[51871]_  = ~A267 & ~A266;
  assign \new_[51872]_  = A265 & \new_[51871]_ ;
  assign \new_[51875]_  = ~A269 & ~A268;
  assign \new_[51878]_  = A301 & ~A300;
  assign \new_[51879]_  = \new_[51878]_  & \new_[51875]_ ;
  assign \new_[51880]_  = \new_[51879]_  & \new_[51872]_ ;
  assign \new_[51884]_  = A168 & ~A169;
  assign \new_[51885]_  = A170 & \new_[51884]_ ;
  assign \new_[51889]_  = ~A203 & ~A202;
  assign \new_[51890]_  = A201 & \new_[51889]_ ;
  assign \new_[51891]_  = \new_[51890]_  & \new_[51885]_ ;
  assign \new_[51895]_  = ~A267 & ~A266;
  assign \new_[51896]_  = A265 & \new_[51895]_ ;
  assign \new_[51899]_  = ~A269 & ~A268;
  assign \new_[51902]_  = A302 & ~A300;
  assign \new_[51903]_  = \new_[51902]_  & \new_[51899]_ ;
  assign \new_[51904]_  = \new_[51903]_  & \new_[51896]_ ;
  assign \new_[51908]_  = A168 & ~A169;
  assign \new_[51909]_  = A170 & \new_[51908]_ ;
  assign \new_[51913]_  = ~A203 & ~A202;
  assign \new_[51914]_  = A201 & \new_[51913]_ ;
  assign \new_[51915]_  = \new_[51914]_  & \new_[51909]_ ;
  assign \new_[51919]_  = ~A267 & ~A266;
  assign \new_[51920]_  = A265 & \new_[51919]_ ;
  assign \new_[51923]_  = ~A269 & ~A268;
  assign \new_[51926]_  = A299 & A298;
  assign \new_[51927]_  = \new_[51926]_  & \new_[51923]_ ;
  assign \new_[51928]_  = \new_[51927]_  & \new_[51920]_ ;
  assign \new_[51932]_  = A168 & ~A169;
  assign \new_[51933]_  = A170 & \new_[51932]_ ;
  assign \new_[51937]_  = ~A203 & ~A202;
  assign \new_[51938]_  = A201 & \new_[51937]_ ;
  assign \new_[51939]_  = \new_[51938]_  & \new_[51933]_ ;
  assign \new_[51943]_  = ~A267 & ~A266;
  assign \new_[51944]_  = A265 & \new_[51943]_ ;
  assign \new_[51947]_  = ~A269 & ~A268;
  assign \new_[51950]_  = ~A299 & ~A298;
  assign \new_[51951]_  = \new_[51950]_  & \new_[51947]_ ;
  assign \new_[51952]_  = \new_[51951]_  & \new_[51944]_ ;
  assign \new_[51956]_  = A168 & ~A169;
  assign \new_[51957]_  = A170 & \new_[51956]_ ;
  assign \new_[51961]_  = ~A265 & A202;
  assign \new_[51962]_  = ~A201 & \new_[51961]_ ;
  assign \new_[51963]_  = \new_[51962]_  & \new_[51957]_ ;
  assign \new_[51967]_  = ~A268 & ~A267;
  assign \new_[51968]_  = A266 & \new_[51967]_ ;
  assign \new_[51971]_  = A300 & ~A269;
  assign \new_[51974]_  = ~A302 & ~A301;
  assign \new_[51975]_  = \new_[51974]_  & \new_[51971]_ ;
  assign \new_[51976]_  = \new_[51975]_  & \new_[51968]_ ;
  assign \new_[51980]_  = A168 & ~A169;
  assign \new_[51981]_  = A170 & \new_[51980]_ ;
  assign \new_[51985]_  = A265 & A202;
  assign \new_[51986]_  = ~A201 & \new_[51985]_ ;
  assign \new_[51987]_  = \new_[51986]_  & \new_[51981]_ ;
  assign \new_[51991]_  = ~A268 & ~A267;
  assign \new_[51992]_  = ~A266 & \new_[51991]_ ;
  assign \new_[51995]_  = A300 & ~A269;
  assign \new_[51998]_  = ~A302 & ~A301;
  assign \new_[51999]_  = \new_[51998]_  & \new_[51995]_ ;
  assign \new_[52000]_  = \new_[51999]_  & \new_[51992]_ ;
  assign \new_[52004]_  = A168 & ~A169;
  assign \new_[52005]_  = A170 & \new_[52004]_ ;
  assign \new_[52009]_  = ~A265 & A203;
  assign \new_[52010]_  = ~A201 & \new_[52009]_ ;
  assign \new_[52011]_  = \new_[52010]_  & \new_[52005]_ ;
  assign \new_[52015]_  = ~A268 & ~A267;
  assign \new_[52016]_  = A266 & \new_[52015]_ ;
  assign \new_[52019]_  = A300 & ~A269;
  assign \new_[52022]_  = ~A302 & ~A301;
  assign \new_[52023]_  = \new_[52022]_  & \new_[52019]_ ;
  assign \new_[52024]_  = \new_[52023]_  & \new_[52016]_ ;
  assign \new_[52028]_  = A168 & ~A169;
  assign \new_[52029]_  = A170 & \new_[52028]_ ;
  assign \new_[52033]_  = A265 & A203;
  assign \new_[52034]_  = ~A201 & \new_[52033]_ ;
  assign \new_[52035]_  = \new_[52034]_  & \new_[52029]_ ;
  assign \new_[52039]_  = ~A268 & ~A267;
  assign \new_[52040]_  = ~A266 & \new_[52039]_ ;
  assign \new_[52043]_  = A300 & ~A269;
  assign \new_[52046]_  = ~A302 & ~A301;
  assign \new_[52047]_  = \new_[52046]_  & \new_[52043]_ ;
  assign \new_[52048]_  = \new_[52047]_  & \new_[52040]_ ;
  assign \new_[52052]_  = A168 & ~A169;
  assign \new_[52053]_  = A170 & \new_[52052]_ ;
  assign \new_[52057]_  = ~A265 & A200;
  assign \new_[52058]_  = A199 & \new_[52057]_ ;
  assign \new_[52059]_  = \new_[52058]_  & \new_[52053]_ ;
  assign \new_[52063]_  = ~A268 & ~A267;
  assign \new_[52064]_  = A266 & \new_[52063]_ ;
  assign \new_[52067]_  = A300 & ~A269;
  assign \new_[52070]_  = ~A302 & ~A301;
  assign \new_[52071]_  = \new_[52070]_  & \new_[52067]_ ;
  assign \new_[52072]_  = \new_[52071]_  & \new_[52064]_ ;
  assign \new_[52076]_  = A168 & ~A169;
  assign \new_[52077]_  = A170 & \new_[52076]_ ;
  assign \new_[52081]_  = A265 & A200;
  assign \new_[52082]_  = A199 & \new_[52081]_ ;
  assign \new_[52083]_  = \new_[52082]_  & \new_[52077]_ ;
  assign \new_[52087]_  = ~A268 & ~A267;
  assign \new_[52088]_  = ~A266 & \new_[52087]_ ;
  assign \new_[52091]_  = A300 & ~A269;
  assign \new_[52094]_  = ~A302 & ~A301;
  assign \new_[52095]_  = \new_[52094]_  & \new_[52091]_ ;
  assign \new_[52096]_  = \new_[52095]_  & \new_[52088]_ ;
  assign \new_[52100]_  = A168 & ~A169;
  assign \new_[52101]_  = A170 & \new_[52100]_ ;
  assign \new_[52105]_  = A201 & A200;
  assign \new_[52106]_  = ~A199 & \new_[52105]_ ;
  assign \new_[52107]_  = \new_[52106]_  & \new_[52101]_ ;
  assign \new_[52111]_  = A268 & ~A267;
  assign \new_[52112]_  = A202 & \new_[52111]_ ;
  assign \new_[52115]_  = ~A299 & A298;
  assign \new_[52118]_  = A301 & A300;
  assign \new_[52119]_  = \new_[52118]_  & \new_[52115]_ ;
  assign \new_[52120]_  = \new_[52119]_  & \new_[52112]_ ;
  assign \new_[52124]_  = A168 & ~A169;
  assign \new_[52125]_  = A170 & \new_[52124]_ ;
  assign \new_[52129]_  = A201 & A200;
  assign \new_[52130]_  = ~A199 & \new_[52129]_ ;
  assign \new_[52131]_  = \new_[52130]_  & \new_[52125]_ ;
  assign \new_[52135]_  = A268 & ~A267;
  assign \new_[52136]_  = A202 & \new_[52135]_ ;
  assign \new_[52139]_  = ~A299 & A298;
  assign \new_[52142]_  = A302 & A300;
  assign \new_[52143]_  = \new_[52142]_  & \new_[52139]_ ;
  assign \new_[52144]_  = \new_[52143]_  & \new_[52136]_ ;
  assign \new_[52148]_  = A168 & ~A169;
  assign \new_[52149]_  = A170 & \new_[52148]_ ;
  assign \new_[52153]_  = A201 & A200;
  assign \new_[52154]_  = ~A199 & \new_[52153]_ ;
  assign \new_[52155]_  = \new_[52154]_  & \new_[52149]_ ;
  assign \new_[52159]_  = A268 & ~A267;
  assign \new_[52160]_  = A202 & \new_[52159]_ ;
  assign \new_[52163]_  = A299 & ~A298;
  assign \new_[52166]_  = A301 & A300;
  assign \new_[52167]_  = \new_[52166]_  & \new_[52163]_ ;
  assign \new_[52168]_  = \new_[52167]_  & \new_[52160]_ ;
  assign \new_[52172]_  = A168 & ~A169;
  assign \new_[52173]_  = A170 & \new_[52172]_ ;
  assign \new_[52177]_  = A201 & A200;
  assign \new_[52178]_  = ~A199 & \new_[52177]_ ;
  assign \new_[52179]_  = \new_[52178]_  & \new_[52173]_ ;
  assign \new_[52183]_  = A268 & ~A267;
  assign \new_[52184]_  = A202 & \new_[52183]_ ;
  assign \new_[52187]_  = A299 & ~A298;
  assign \new_[52190]_  = A302 & A300;
  assign \new_[52191]_  = \new_[52190]_  & \new_[52187]_ ;
  assign \new_[52192]_  = \new_[52191]_  & \new_[52184]_ ;
  assign \new_[52196]_  = A168 & ~A169;
  assign \new_[52197]_  = A170 & \new_[52196]_ ;
  assign \new_[52201]_  = A201 & A200;
  assign \new_[52202]_  = ~A199 & \new_[52201]_ ;
  assign \new_[52203]_  = \new_[52202]_  & \new_[52197]_ ;
  assign \new_[52207]_  = A269 & ~A267;
  assign \new_[52208]_  = A202 & \new_[52207]_ ;
  assign \new_[52211]_  = ~A299 & A298;
  assign \new_[52214]_  = A301 & A300;
  assign \new_[52215]_  = \new_[52214]_  & \new_[52211]_ ;
  assign \new_[52216]_  = \new_[52215]_  & \new_[52208]_ ;
  assign \new_[52220]_  = A168 & ~A169;
  assign \new_[52221]_  = A170 & \new_[52220]_ ;
  assign \new_[52225]_  = A201 & A200;
  assign \new_[52226]_  = ~A199 & \new_[52225]_ ;
  assign \new_[52227]_  = \new_[52226]_  & \new_[52221]_ ;
  assign \new_[52231]_  = A269 & ~A267;
  assign \new_[52232]_  = A202 & \new_[52231]_ ;
  assign \new_[52235]_  = ~A299 & A298;
  assign \new_[52238]_  = A302 & A300;
  assign \new_[52239]_  = \new_[52238]_  & \new_[52235]_ ;
  assign \new_[52240]_  = \new_[52239]_  & \new_[52232]_ ;
  assign \new_[52244]_  = A168 & ~A169;
  assign \new_[52245]_  = A170 & \new_[52244]_ ;
  assign \new_[52249]_  = A201 & A200;
  assign \new_[52250]_  = ~A199 & \new_[52249]_ ;
  assign \new_[52251]_  = \new_[52250]_  & \new_[52245]_ ;
  assign \new_[52255]_  = A269 & ~A267;
  assign \new_[52256]_  = A202 & \new_[52255]_ ;
  assign \new_[52259]_  = A299 & ~A298;
  assign \new_[52262]_  = A301 & A300;
  assign \new_[52263]_  = \new_[52262]_  & \new_[52259]_ ;
  assign \new_[52264]_  = \new_[52263]_  & \new_[52256]_ ;
  assign \new_[52268]_  = A168 & ~A169;
  assign \new_[52269]_  = A170 & \new_[52268]_ ;
  assign \new_[52273]_  = A201 & A200;
  assign \new_[52274]_  = ~A199 & \new_[52273]_ ;
  assign \new_[52275]_  = \new_[52274]_  & \new_[52269]_ ;
  assign \new_[52279]_  = A269 & ~A267;
  assign \new_[52280]_  = A202 & \new_[52279]_ ;
  assign \new_[52283]_  = A299 & ~A298;
  assign \new_[52286]_  = A302 & A300;
  assign \new_[52287]_  = \new_[52286]_  & \new_[52283]_ ;
  assign \new_[52288]_  = \new_[52287]_  & \new_[52280]_ ;
  assign \new_[52292]_  = A168 & ~A169;
  assign \new_[52293]_  = A170 & \new_[52292]_ ;
  assign \new_[52297]_  = A201 & A200;
  assign \new_[52298]_  = ~A199 & \new_[52297]_ ;
  assign \new_[52299]_  = \new_[52298]_  & \new_[52293]_ ;
  assign \new_[52303]_  = A266 & A265;
  assign \new_[52304]_  = A202 & \new_[52303]_ ;
  assign \new_[52307]_  = ~A299 & A298;
  assign \new_[52310]_  = A301 & A300;
  assign \new_[52311]_  = \new_[52310]_  & \new_[52307]_ ;
  assign \new_[52312]_  = \new_[52311]_  & \new_[52304]_ ;
  assign \new_[52316]_  = A168 & ~A169;
  assign \new_[52317]_  = A170 & \new_[52316]_ ;
  assign \new_[52321]_  = A201 & A200;
  assign \new_[52322]_  = ~A199 & \new_[52321]_ ;
  assign \new_[52323]_  = \new_[52322]_  & \new_[52317]_ ;
  assign \new_[52327]_  = A266 & A265;
  assign \new_[52328]_  = A202 & \new_[52327]_ ;
  assign \new_[52331]_  = ~A299 & A298;
  assign \new_[52334]_  = A302 & A300;
  assign \new_[52335]_  = \new_[52334]_  & \new_[52331]_ ;
  assign \new_[52336]_  = \new_[52335]_  & \new_[52328]_ ;
  assign \new_[52340]_  = A168 & ~A169;
  assign \new_[52341]_  = A170 & \new_[52340]_ ;
  assign \new_[52345]_  = A201 & A200;
  assign \new_[52346]_  = ~A199 & \new_[52345]_ ;
  assign \new_[52347]_  = \new_[52346]_  & \new_[52341]_ ;
  assign \new_[52351]_  = A266 & A265;
  assign \new_[52352]_  = A202 & \new_[52351]_ ;
  assign \new_[52355]_  = A299 & ~A298;
  assign \new_[52358]_  = A301 & A300;
  assign \new_[52359]_  = \new_[52358]_  & \new_[52355]_ ;
  assign \new_[52360]_  = \new_[52359]_  & \new_[52352]_ ;
  assign \new_[52364]_  = A168 & ~A169;
  assign \new_[52365]_  = A170 & \new_[52364]_ ;
  assign \new_[52369]_  = A201 & A200;
  assign \new_[52370]_  = ~A199 & \new_[52369]_ ;
  assign \new_[52371]_  = \new_[52370]_  & \new_[52365]_ ;
  assign \new_[52375]_  = A266 & A265;
  assign \new_[52376]_  = A202 & \new_[52375]_ ;
  assign \new_[52379]_  = A299 & ~A298;
  assign \new_[52382]_  = A302 & A300;
  assign \new_[52383]_  = \new_[52382]_  & \new_[52379]_ ;
  assign \new_[52384]_  = \new_[52383]_  & \new_[52376]_ ;
  assign \new_[52388]_  = A168 & ~A169;
  assign \new_[52389]_  = A170 & \new_[52388]_ ;
  assign \new_[52393]_  = A201 & A200;
  assign \new_[52394]_  = ~A199 & \new_[52393]_ ;
  assign \new_[52395]_  = \new_[52394]_  & \new_[52389]_ ;
  assign \new_[52399]_  = ~A266 & ~A265;
  assign \new_[52400]_  = A202 & \new_[52399]_ ;
  assign \new_[52403]_  = ~A299 & A298;
  assign \new_[52406]_  = A301 & A300;
  assign \new_[52407]_  = \new_[52406]_  & \new_[52403]_ ;
  assign \new_[52408]_  = \new_[52407]_  & \new_[52400]_ ;
  assign \new_[52412]_  = A168 & ~A169;
  assign \new_[52413]_  = A170 & \new_[52412]_ ;
  assign \new_[52417]_  = A201 & A200;
  assign \new_[52418]_  = ~A199 & \new_[52417]_ ;
  assign \new_[52419]_  = \new_[52418]_  & \new_[52413]_ ;
  assign \new_[52423]_  = ~A266 & ~A265;
  assign \new_[52424]_  = A202 & \new_[52423]_ ;
  assign \new_[52427]_  = ~A299 & A298;
  assign \new_[52430]_  = A302 & A300;
  assign \new_[52431]_  = \new_[52430]_  & \new_[52427]_ ;
  assign \new_[52432]_  = \new_[52431]_  & \new_[52424]_ ;
  assign \new_[52436]_  = A168 & ~A169;
  assign \new_[52437]_  = A170 & \new_[52436]_ ;
  assign \new_[52441]_  = A201 & A200;
  assign \new_[52442]_  = ~A199 & \new_[52441]_ ;
  assign \new_[52443]_  = \new_[52442]_  & \new_[52437]_ ;
  assign \new_[52447]_  = ~A266 & ~A265;
  assign \new_[52448]_  = A202 & \new_[52447]_ ;
  assign \new_[52451]_  = A299 & ~A298;
  assign \new_[52454]_  = A301 & A300;
  assign \new_[52455]_  = \new_[52454]_  & \new_[52451]_ ;
  assign \new_[52456]_  = \new_[52455]_  & \new_[52448]_ ;
  assign \new_[52460]_  = A168 & ~A169;
  assign \new_[52461]_  = A170 & \new_[52460]_ ;
  assign \new_[52465]_  = A201 & A200;
  assign \new_[52466]_  = ~A199 & \new_[52465]_ ;
  assign \new_[52467]_  = \new_[52466]_  & \new_[52461]_ ;
  assign \new_[52471]_  = ~A266 & ~A265;
  assign \new_[52472]_  = A202 & \new_[52471]_ ;
  assign \new_[52475]_  = A299 & ~A298;
  assign \new_[52478]_  = A302 & A300;
  assign \new_[52479]_  = \new_[52478]_  & \new_[52475]_ ;
  assign \new_[52480]_  = \new_[52479]_  & \new_[52472]_ ;
  assign \new_[52484]_  = A168 & ~A169;
  assign \new_[52485]_  = A170 & \new_[52484]_ ;
  assign \new_[52489]_  = A201 & A200;
  assign \new_[52490]_  = ~A199 & \new_[52489]_ ;
  assign \new_[52491]_  = \new_[52490]_  & \new_[52485]_ ;
  assign \new_[52495]_  = A268 & ~A267;
  assign \new_[52496]_  = A203 & \new_[52495]_ ;
  assign \new_[52499]_  = ~A299 & A298;
  assign \new_[52502]_  = A301 & A300;
  assign \new_[52503]_  = \new_[52502]_  & \new_[52499]_ ;
  assign \new_[52504]_  = \new_[52503]_  & \new_[52496]_ ;
  assign \new_[52508]_  = A168 & ~A169;
  assign \new_[52509]_  = A170 & \new_[52508]_ ;
  assign \new_[52513]_  = A201 & A200;
  assign \new_[52514]_  = ~A199 & \new_[52513]_ ;
  assign \new_[52515]_  = \new_[52514]_  & \new_[52509]_ ;
  assign \new_[52519]_  = A268 & ~A267;
  assign \new_[52520]_  = A203 & \new_[52519]_ ;
  assign \new_[52523]_  = ~A299 & A298;
  assign \new_[52526]_  = A302 & A300;
  assign \new_[52527]_  = \new_[52526]_  & \new_[52523]_ ;
  assign \new_[52528]_  = \new_[52527]_  & \new_[52520]_ ;
  assign \new_[52532]_  = A168 & ~A169;
  assign \new_[52533]_  = A170 & \new_[52532]_ ;
  assign \new_[52537]_  = A201 & A200;
  assign \new_[52538]_  = ~A199 & \new_[52537]_ ;
  assign \new_[52539]_  = \new_[52538]_  & \new_[52533]_ ;
  assign \new_[52543]_  = A268 & ~A267;
  assign \new_[52544]_  = A203 & \new_[52543]_ ;
  assign \new_[52547]_  = A299 & ~A298;
  assign \new_[52550]_  = A301 & A300;
  assign \new_[52551]_  = \new_[52550]_  & \new_[52547]_ ;
  assign \new_[52552]_  = \new_[52551]_  & \new_[52544]_ ;
  assign \new_[52556]_  = A168 & ~A169;
  assign \new_[52557]_  = A170 & \new_[52556]_ ;
  assign \new_[52561]_  = A201 & A200;
  assign \new_[52562]_  = ~A199 & \new_[52561]_ ;
  assign \new_[52563]_  = \new_[52562]_  & \new_[52557]_ ;
  assign \new_[52567]_  = A268 & ~A267;
  assign \new_[52568]_  = A203 & \new_[52567]_ ;
  assign \new_[52571]_  = A299 & ~A298;
  assign \new_[52574]_  = A302 & A300;
  assign \new_[52575]_  = \new_[52574]_  & \new_[52571]_ ;
  assign \new_[52576]_  = \new_[52575]_  & \new_[52568]_ ;
  assign \new_[52580]_  = A168 & ~A169;
  assign \new_[52581]_  = A170 & \new_[52580]_ ;
  assign \new_[52585]_  = A201 & A200;
  assign \new_[52586]_  = ~A199 & \new_[52585]_ ;
  assign \new_[52587]_  = \new_[52586]_  & \new_[52581]_ ;
  assign \new_[52591]_  = A269 & ~A267;
  assign \new_[52592]_  = A203 & \new_[52591]_ ;
  assign \new_[52595]_  = ~A299 & A298;
  assign \new_[52598]_  = A301 & A300;
  assign \new_[52599]_  = \new_[52598]_  & \new_[52595]_ ;
  assign \new_[52600]_  = \new_[52599]_  & \new_[52592]_ ;
  assign \new_[52604]_  = A168 & ~A169;
  assign \new_[52605]_  = A170 & \new_[52604]_ ;
  assign \new_[52609]_  = A201 & A200;
  assign \new_[52610]_  = ~A199 & \new_[52609]_ ;
  assign \new_[52611]_  = \new_[52610]_  & \new_[52605]_ ;
  assign \new_[52615]_  = A269 & ~A267;
  assign \new_[52616]_  = A203 & \new_[52615]_ ;
  assign \new_[52619]_  = ~A299 & A298;
  assign \new_[52622]_  = A302 & A300;
  assign \new_[52623]_  = \new_[52622]_  & \new_[52619]_ ;
  assign \new_[52624]_  = \new_[52623]_  & \new_[52616]_ ;
  assign \new_[52628]_  = A168 & ~A169;
  assign \new_[52629]_  = A170 & \new_[52628]_ ;
  assign \new_[52633]_  = A201 & A200;
  assign \new_[52634]_  = ~A199 & \new_[52633]_ ;
  assign \new_[52635]_  = \new_[52634]_  & \new_[52629]_ ;
  assign \new_[52639]_  = A269 & ~A267;
  assign \new_[52640]_  = A203 & \new_[52639]_ ;
  assign \new_[52643]_  = A299 & ~A298;
  assign \new_[52646]_  = A301 & A300;
  assign \new_[52647]_  = \new_[52646]_  & \new_[52643]_ ;
  assign \new_[52648]_  = \new_[52647]_  & \new_[52640]_ ;
  assign \new_[52652]_  = A168 & ~A169;
  assign \new_[52653]_  = A170 & \new_[52652]_ ;
  assign \new_[52657]_  = A201 & A200;
  assign \new_[52658]_  = ~A199 & \new_[52657]_ ;
  assign \new_[52659]_  = \new_[52658]_  & \new_[52653]_ ;
  assign \new_[52663]_  = A269 & ~A267;
  assign \new_[52664]_  = A203 & \new_[52663]_ ;
  assign \new_[52667]_  = A299 & ~A298;
  assign \new_[52670]_  = A302 & A300;
  assign \new_[52671]_  = \new_[52670]_  & \new_[52667]_ ;
  assign \new_[52672]_  = \new_[52671]_  & \new_[52664]_ ;
  assign \new_[52676]_  = A168 & ~A169;
  assign \new_[52677]_  = A170 & \new_[52676]_ ;
  assign \new_[52681]_  = A201 & A200;
  assign \new_[52682]_  = ~A199 & \new_[52681]_ ;
  assign \new_[52683]_  = \new_[52682]_  & \new_[52677]_ ;
  assign \new_[52687]_  = A266 & A265;
  assign \new_[52688]_  = A203 & \new_[52687]_ ;
  assign \new_[52691]_  = ~A299 & A298;
  assign \new_[52694]_  = A301 & A300;
  assign \new_[52695]_  = \new_[52694]_  & \new_[52691]_ ;
  assign \new_[52696]_  = \new_[52695]_  & \new_[52688]_ ;
  assign \new_[52700]_  = A168 & ~A169;
  assign \new_[52701]_  = A170 & \new_[52700]_ ;
  assign \new_[52705]_  = A201 & A200;
  assign \new_[52706]_  = ~A199 & \new_[52705]_ ;
  assign \new_[52707]_  = \new_[52706]_  & \new_[52701]_ ;
  assign \new_[52711]_  = A266 & A265;
  assign \new_[52712]_  = A203 & \new_[52711]_ ;
  assign \new_[52715]_  = ~A299 & A298;
  assign \new_[52718]_  = A302 & A300;
  assign \new_[52719]_  = \new_[52718]_  & \new_[52715]_ ;
  assign \new_[52720]_  = \new_[52719]_  & \new_[52712]_ ;
  assign \new_[52724]_  = A168 & ~A169;
  assign \new_[52725]_  = A170 & \new_[52724]_ ;
  assign \new_[52729]_  = A201 & A200;
  assign \new_[52730]_  = ~A199 & \new_[52729]_ ;
  assign \new_[52731]_  = \new_[52730]_  & \new_[52725]_ ;
  assign \new_[52735]_  = A266 & A265;
  assign \new_[52736]_  = A203 & \new_[52735]_ ;
  assign \new_[52739]_  = A299 & ~A298;
  assign \new_[52742]_  = A301 & A300;
  assign \new_[52743]_  = \new_[52742]_  & \new_[52739]_ ;
  assign \new_[52744]_  = \new_[52743]_  & \new_[52736]_ ;
  assign \new_[52748]_  = A168 & ~A169;
  assign \new_[52749]_  = A170 & \new_[52748]_ ;
  assign \new_[52753]_  = A201 & A200;
  assign \new_[52754]_  = ~A199 & \new_[52753]_ ;
  assign \new_[52755]_  = \new_[52754]_  & \new_[52749]_ ;
  assign \new_[52759]_  = A266 & A265;
  assign \new_[52760]_  = A203 & \new_[52759]_ ;
  assign \new_[52763]_  = A299 & ~A298;
  assign \new_[52766]_  = A302 & A300;
  assign \new_[52767]_  = \new_[52766]_  & \new_[52763]_ ;
  assign \new_[52768]_  = \new_[52767]_  & \new_[52760]_ ;
  assign \new_[52772]_  = A168 & ~A169;
  assign \new_[52773]_  = A170 & \new_[52772]_ ;
  assign \new_[52777]_  = A201 & A200;
  assign \new_[52778]_  = ~A199 & \new_[52777]_ ;
  assign \new_[52779]_  = \new_[52778]_  & \new_[52773]_ ;
  assign \new_[52783]_  = ~A266 & ~A265;
  assign \new_[52784]_  = A203 & \new_[52783]_ ;
  assign \new_[52787]_  = ~A299 & A298;
  assign \new_[52790]_  = A301 & A300;
  assign \new_[52791]_  = \new_[52790]_  & \new_[52787]_ ;
  assign \new_[52792]_  = \new_[52791]_  & \new_[52784]_ ;
  assign \new_[52796]_  = A168 & ~A169;
  assign \new_[52797]_  = A170 & \new_[52796]_ ;
  assign \new_[52801]_  = A201 & A200;
  assign \new_[52802]_  = ~A199 & \new_[52801]_ ;
  assign \new_[52803]_  = \new_[52802]_  & \new_[52797]_ ;
  assign \new_[52807]_  = ~A266 & ~A265;
  assign \new_[52808]_  = A203 & \new_[52807]_ ;
  assign \new_[52811]_  = ~A299 & A298;
  assign \new_[52814]_  = A302 & A300;
  assign \new_[52815]_  = \new_[52814]_  & \new_[52811]_ ;
  assign \new_[52816]_  = \new_[52815]_  & \new_[52808]_ ;
  assign \new_[52820]_  = A168 & ~A169;
  assign \new_[52821]_  = A170 & \new_[52820]_ ;
  assign \new_[52825]_  = A201 & A200;
  assign \new_[52826]_  = ~A199 & \new_[52825]_ ;
  assign \new_[52827]_  = \new_[52826]_  & \new_[52821]_ ;
  assign \new_[52831]_  = ~A266 & ~A265;
  assign \new_[52832]_  = A203 & \new_[52831]_ ;
  assign \new_[52835]_  = A299 & ~A298;
  assign \new_[52838]_  = A301 & A300;
  assign \new_[52839]_  = \new_[52838]_  & \new_[52835]_ ;
  assign \new_[52840]_  = \new_[52839]_  & \new_[52832]_ ;
  assign \new_[52844]_  = A168 & ~A169;
  assign \new_[52845]_  = A170 & \new_[52844]_ ;
  assign \new_[52849]_  = A201 & A200;
  assign \new_[52850]_  = ~A199 & \new_[52849]_ ;
  assign \new_[52851]_  = \new_[52850]_  & \new_[52845]_ ;
  assign \new_[52855]_  = ~A266 & ~A265;
  assign \new_[52856]_  = A203 & \new_[52855]_ ;
  assign \new_[52859]_  = A299 & ~A298;
  assign \new_[52862]_  = A302 & A300;
  assign \new_[52863]_  = \new_[52862]_  & \new_[52859]_ ;
  assign \new_[52864]_  = \new_[52863]_  & \new_[52856]_ ;
  assign \new_[52868]_  = A168 & ~A169;
  assign \new_[52869]_  = A170 & \new_[52868]_ ;
  assign \new_[52873]_  = A201 & ~A200;
  assign \new_[52874]_  = A199 & \new_[52873]_ ;
  assign \new_[52875]_  = \new_[52874]_  & \new_[52869]_ ;
  assign \new_[52879]_  = A268 & ~A267;
  assign \new_[52880]_  = A202 & \new_[52879]_ ;
  assign \new_[52883]_  = ~A299 & A298;
  assign \new_[52886]_  = A301 & A300;
  assign \new_[52887]_  = \new_[52886]_  & \new_[52883]_ ;
  assign \new_[52888]_  = \new_[52887]_  & \new_[52880]_ ;
  assign \new_[52892]_  = A168 & ~A169;
  assign \new_[52893]_  = A170 & \new_[52892]_ ;
  assign \new_[52897]_  = A201 & ~A200;
  assign \new_[52898]_  = A199 & \new_[52897]_ ;
  assign \new_[52899]_  = \new_[52898]_  & \new_[52893]_ ;
  assign \new_[52903]_  = A268 & ~A267;
  assign \new_[52904]_  = A202 & \new_[52903]_ ;
  assign \new_[52907]_  = ~A299 & A298;
  assign \new_[52910]_  = A302 & A300;
  assign \new_[52911]_  = \new_[52910]_  & \new_[52907]_ ;
  assign \new_[52912]_  = \new_[52911]_  & \new_[52904]_ ;
  assign \new_[52916]_  = A168 & ~A169;
  assign \new_[52917]_  = A170 & \new_[52916]_ ;
  assign \new_[52921]_  = A201 & ~A200;
  assign \new_[52922]_  = A199 & \new_[52921]_ ;
  assign \new_[52923]_  = \new_[52922]_  & \new_[52917]_ ;
  assign \new_[52927]_  = A268 & ~A267;
  assign \new_[52928]_  = A202 & \new_[52927]_ ;
  assign \new_[52931]_  = A299 & ~A298;
  assign \new_[52934]_  = A301 & A300;
  assign \new_[52935]_  = \new_[52934]_  & \new_[52931]_ ;
  assign \new_[52936]_  = \new_[52935]_  & \new_[52928]_ ;
  assign \new_[52940]_  = A168 & ~A169;
  assign \new_[52941]_  = A170 & \new_[52940]_ ;
  assign \new_[52945]_  = A201 & ~A200;
  assign \new_[52946]_  = A199 & \new_[52945]_ ;
  assign \new_[52947]_  = \new_[52946]_  & \new_[52941]_ ;
  assign \new_[52951]_  = A268 & ~A267;
  assign \new_[52952]_  = A202 & \new_[52951]_ ;
  assign \new_[52955]_  = A299 & ~A298;
  assign \new_[52958]_  = A302 & A300;
  assign \new_[52959]_  = \new_[52958]_  & \new_[52955]_ ;
  assign \new_[52960]_  = \new_[52959]_  & \new_[52952]_ ;
  assign \new_[52964]_  = A168 & ~A169;
  assign \new_[52965]_  = A170 & \new_[52964]_ ;
  assign \new_[52969]_  = A201 & ~A200;
  assign \new_[52970]_  = A199 & \new_[52969]_ ;
  assign \new_[52971]_  = \new_[52970]_  & \new_[52965]_ ;
  assign \new_[52975]_  = A269 & ~A267;
  assign \new_[52976]_  = A202 & \new_[52975]_ ;
  assign \new_[52979]_  = ~A299 & A298;
  assign \new_[52982]_  = A301 & A300;
  assign \new_[52983]_  = \new_[52982]_  & \new_[52979]_ ;
  assign \new_[52984]_  = \new_[52983]_  & \new_[52976]_ ;
  assign \new_[52988]_  = A168 & ~A169;
  assign \new_[52989]_  = A170 & \new_[52988]_ ;
  assign \new_[52993]_  = A201 & ~A200;
  assign \new_[52994]_  = A199 & \new_[52993]_ ;
  assign \new_[52995]_  = \new_[52994]_  & \new_[52989]_ ;
  assign \new_[52999]_  = A269 & ~A267;
  assign \new_[53000]_  = A202 & \new_[52999]_ ;
  assign \new_[53003]_  = ~A299 & A298;
  assign \new_[53006]_  = A302 & A300;
  assign \new_[53007]_  = \new_[53006]_  & \new_[53003]_ ;
  assign \new_[53008]_  = \new_[53007]_  & \new_[53000]_ ;
  assign \new_[53012]_  = A168 & ~A169;
  assign \new_[53013]_  = A170 & \new_[53012]_ ;
  assign \new_[53017]_  = A201 & ~A200;
  assign \new_[53018]_  = A199 & \new_[53017]_ ;
  assign \new_[53019]_  = \new_[53018]_  & \new_[53013]_ ;
  assign \new_[53023]_  = A269 & ~A267;
  assign \new_[53024]_  = A202 & \new_[53023]_ ;
  assign \new_[53027]_  = A299 & ~A298;
  assign \new_[53030]_  = A301 & A300;
  assign \new_[53031]_  = \new_[53030]_  & \new_[53027]_ ;
  assign \new_[53032]_  = \new_[53031]_  & \new_[53024]_ ;
  assign \new_[53036]_  = A168 & ~A169;
  assign \new_[53037]_  = A170 & \new_[53036]_ ;
  assign \new_[53041]_  = A201 & ~A200;
  assign \new_[53042]_  = A199 & \new_[53041]_ ;
  assign \new_[53043]_  = \new_[53042]_  & \new_[53037]_ ;
  assign \new_[53047]_  = A269 & ~A267;
  assign \new_[53048]_  = A202 & \new_[53047]_ ;
  assign \new_[53051]_  = A299 & ~A298;
  assign \new_[53054]_  = A302 & A300;
  assign \new_[53055]_  = \new_[53054]_  & \new_[53051]_ ;
  assign \new_[53056]_  = \new_[53055]_  & \new_[53048]_ ;
  assign \new_[53060]_  = A168 & ~A169;
  assign \new_[53061]_  = A170 & \new_[53060]_ ;
  assign \new_[53065]_  = A201 & ~A200;
  assign \new_[53066]_  = A199 & \new_[53065]_ ;
  assign \new_[53067]_  = \new_[53066]_  & \new_[53061]_ ;
  assign \new_[53071]_  = A266 & A265;
  assign \new_[53072]_  = A202 & \new_[53071]_ ;
  assign \new_[53075]_  = ~A299 & A298;
  assign \new_[53078]_  = A301 & A300;
  assign \new_[53079]_  = \new_[53078]_  & \new_[53075]_ ;
  assign \new_[53080]_  = \new_[53079]_  & \new_[53072]_ ;
  assign \new_[53084]_  = A168 & ~A169;
  assign \new_[53085]_  = A170 & \new_[53084]_ ;
  assign \new_[53089]_  = A201 & ~A200;
  assign \new_[53090]_  = A199 & \new_[53089]_ ;
  assign \new_[53091]_  = \new_[53090]_  & \new_[53085]_ ;
  assign \new_[53095]_  = A266 & A265;
  assign \new_[53096]_  = A202 & \new_[53095]_ ;
  assign \new_[53099]_  = ~A299 & A298;
  assign \new_[53102]_  = A302 & A300;
  assign \new_[53103]_  = \new_[53102]_  & \new_[53099]_ ;
  assign \new_[53104]_  = \new_[53103]_  & \new_[53096]_ ;
  assign \new_[53108]_  = A168 & ~A169;
  assign \new_[53109]_  = A170 & \new_[53108]_ ;
  assign \new_[53113]_  = A201 & ~A200;
  assign \new_[53114]_  = A199 & \new_[53113]_ ;
  assign \new_[53115]_  = \new_[53114]_  & \new_[53109]_ ;
  assign \new_[53119]_  = A266 & A265;
  assign \new_[53120]_  = A202 & \new_[53119]_ ;
  assign \new_[53123]_  = A299 & ~A298;
  assign \new_[53126]_  = A301 & A300;
  assign \new_[53127]_  = \new_[53126]_  & \new_[53123]_ ;
  assign \new_[53128]_  = \new_[53127]_  & \new_[53120]_ ;
  assign \new_[53132]_  = A168 & ~A169;
  assign \new_[53133]_  = A170 & \new_[53132]_ ;
  assign \new_[53137]_  = A201 & ~A200;
  assign \new_[53138]_  = A199 & \new_[53137]_ ;
  assign \new_[53139]_  = \new_[53138]_  & \new_[53133]_ ;
  assign \new_[53143]_  = A266 & A265;
  assign \new_[53144]_  = A202 & \new_[53143]_ ;
  assign \new_[53147]_  = A299 & ~A298;
  assign \new_[53150]_  = A302 & A300;
  assign \new_[53151]_  = \new_[53150]_  & \new_[53147]_ ;
  assign \new_[53152]_  = \new_[53151]_  & \new_[53144]_ ;
  assign \new_[53156]_  = A168 & ~A169;
  assign \new_[53157]_  = A170 & \new_[53156]_ ;
  assign \new_[53161]_  = A201 & ~A200;
  assign \new_[53162]_  = A199 & \new_[53161]_ ;
  assign \new_[53163]_  = \new_[53162]_  & \new_[53157]_ ;
  assign \new_[53167]_  = ~A266 & ~A265;
  assign \new_[53168]_  = A202 & \new_[53167]_ ;
  assign \new_[53171]_  = ~A299 & A298;
  assign \new_[53174]_  = A301 & A300;
  assign \new_[53175]_  = \new_[53174]_  & \new_[53171]_ ;
  assign \new_[53176]_  = \new_[53175]_  & \new_[53168]_ ;
  assign \new_[53180]_  = A168 & ~A169;
  assign \new_[53181]_  = A170 & \new_[53180]_ ;
  assign \new_[53185]_  = A201 & ~A200;
  assign \new_[53186]_  = A199 & \new_[53185]_ ;
  assign \new_[53187]_  = \new_[53186]_  & \new_[53181]_ ;
  assign \new_[53191]_  = ~A266 & ~A265;
  assign \new_[53192]_  = A202 & \new_[53191]_ ;
  assign \new_[53195]_  = ~A299 & A298;
  assign \new_[53198]_  = A302 & A300;
  assign \new_[53199]_  = \new_[53198]_  & \new_[53195]_ ;
  assign \new_[53200]_  = \new_[53199]_  & \new_[53192]_ ;
  assign \new_[53204]_  = A168 & ~A169;
  assign \new_[53205]_  = A170 & \new_[53204]_ ;
  assign \new_[53209]_  = A201 & ~A200;
  assign \new_[53210]_  = A199 & \new_[53209]_ ;
  assign \new_[53211]_  = \new_[53210]_  & \new_[53205]_ ;
  assign \new_[53215]_  = ~A266 & ~A265;
  assign \new_[53216]_  = A202 & \new_[53215]_ ;
  assign \new_[53219]_  = A299 & ~A298;
  assign \new_[53222]_  = A301 & A300;
  assign \new_[53223]_  = \new_[53222]_  & \new_[53219]_ ;
  assign \new_[53224]_  = \new_[53223]_  & \new_[53216]_ ;
  assign \new_[53228]_  = A168 & ~A169;
  assign \new_[53229]_  = A170 & \new_[53228]_ ;
  assign \new_[53233]_  = A201 & ~A200;
  assign \new_[53234]_  = A199 & \new_[53233]_ ;
  assign \new_[53235]_  = \new_[53234]_  & \new_[53229]_ ;
  assign \new_[53239]_  = ~A266 & ~A265;
  assign \new_[53240]_  = A202 & \new_[53239]_ ;
  assign \new_[53243]_  = A299 & ~A298;
  assign \new_[53246]_  = A302 & A300;
  assign \new_[53247]_  = \new_[53246]_  & \new_[53243]_ ;
  assign \new_[53248]_  = \new_[53247]_  & \new_[53240]_ ;
  assign \new_[53252]_  = A168 & ~A169;
  assign \new_[53253]_  = A170 & \new_[53252]_ ;
  assign \new_[53257]_  = A201 & ~A200;
  assign \new_[53258]_  = A199 & \new_[53257]_ ;
  assign \new_[53259]_  = \new_[53258]_  & \new_[53253]_ ;
  assign \new_[53263]_  = A268 & ~A267;
  assign \new_[53264]_  = A203 & \new_[53263]_ ;
  assign \new_[53267]_  = ~A299 & A298;
  assign \new_[53270]_  = A301 & A300;
  assign \new_[53271]_  = \new_[53270]_  & \new_[53267]_ ;
  assign \new_[53272]_  = \new_[53271]_  & \new_[53264]_ ;
  assign \new_[53276]_  = A168 & ~A169;
  assign \new_[53277]_  = A170 & \new_[53276]_ ;
  assign \new_[53281]_  = A201 & ~A200;
  assign \new_[53282]_  = A199 & \new_[53281]_ ;
  assign \new_[53283]_  = \new_[53282]_  & \new_[53277]_ ;
  assign \new_[53287]_  = A268 & ~A267;
  assign \new_[53288]_  = A203 & \new_[53287]_ ;
  assign \new_[53291]_  = ~A299 & A298;
  assign \new_[53294]_  = A302 & A300;
  assign \new_[53295]_  = \new_[53294]_  & \new_[53291]_ ;
  assign \new_[53296]_  = \new_[53295]_  & \new_[53288]_ ;
  assign \new_[53300]_  = A168 & ~A169;
  assign \new_[53301]_  = A170 & \new_[53300]_ ;
  assign \new_[53305]_  = A201 & ~A200;
  assign \new_[53306]_  = A199 & \new_[53305]_ ;
  assign \new_[53307]_  = \new_[53306]_  & \new_[53301]_ ;
  assign \new_[53311]_  = A268 & ~A267;
  assign \new_[53312]_  = A203 & \new_[53311]_ ;
  assign \new_[53315]_  = A299 & ~A298;
  assign \new_[53318]_  = A301 & A300;
  assign \new_[53319]_  = \new_[53318]_  & \new_[53315]_ ;
  assign \new_[53320]_  = \new_[53319]_  & \new_[53312]_ ;
  assign \new_[53324]_  = A168 & ~A169;
  assign \new_[53325]_  = A170 & \new_[53324]_ ;
  assign \new_[53329]_  = A201 & ~A200;
  assign \new_[53330]_  = A199 & \new_[53329]_ ;
  assign \new_[53331]_  = \new_[53330]_  & \new_[53325]_ ;
  assign \new_[53335]_  = A268 & ~A267;
  assign \new_[53336]_  = A203 & \new_[53335]_ ;
  assign \new_[53339]_  = A299 & ~A298;
  assign \new_[53342]_  = A302 & A300;
  assign \new_[53343]_  = \new_[53342]_  & \new_[53339]_ ;
  assign \new_[53344]_  = \new_[53343]_  & \new_[53336]_ ;
  assign \new_[53348]_  = A168 & ~A169;
  assign \new_[53349]_  = A170 & \new_[53348]_ ;
  assign \new_[53353]_  = A201 & ~A200;
  assign \new_[53354]_  = A199 & \new_[53353]_ ;
  assign \new_[53355]_  = \new_[53354]_  & \new_[53349]_ ;
  assign \new_[53359]_  = A269 & ~A267;
  assign \new_[53360]_  = A203 & \new_[53359]_ ;
  assign \new_[53363]_  = ~A299 & A298;
  assign \new_[53366]_  = A301 & A300;
  assign \new_[53367]_  = \new_[53366]_  & \new_[53363]_ ;
  assign \new_[53368]_  = \new_[53367]_  & \new_[53360]_ ;
  assign \new_[53372]_  = A168 & ~A169;
  assign \new_[53373]_  = A170 & \new_[53372]_ ;
  assign \new_[53377]_  = A201 & ~A200;
  assign \new_[53378]_  = A199 & \new_[53377]_ ;
  assign \new_[53379]_  = \new_[53378]_  & \new_[53373]_ ;
  assign \new_[53383]_  = A269 & ~A267;
  assign \new_[53384]_  = A203 & \new_[53383]_ ;
  assign \new_[53387]_  = ~A299 & A298;
  assign \new_[53390]_  = A302 & A300;
  assign \new_[53391]_  = \new_[53390]_  & \new_[53387]_ ;
  assign \new_[53392]_  = \new_[53391]_  & \new_[53384]_ ;
  assign \new_[53396]_  = A168 & ~A169;
  assign \new_[53397]_  = A170 & \new_[53396]_ ;
  assign \new_[53401]_  = A201 & ~A200;
  assign \new_[53402]_  = A199 & \new_[53401]_ ;
  assign \new_[53403]_  = \new_[53402]_  & \new_[53397]_ ;
  assign \new_[53407]_  = A269 & ~A267;
  assign \new_[53408]_  = A203 & \new_[53407]_ ;
  assign \new_[53411]_  = A299 & ~A298;
  assign \new_[53414]_  = A301 & A300;
  assign \new_[53415]_  = \new_[53414]_  & \new_[53411]_ ;
  assign \new_[53416]_  = \new_[53415]_  & \new_[53408]_ ;
  assign \new_[53420]_  = A168 & ~A169;
  assign \new_[53421]_  = A170 & \new_[53420]_ ;
  assign \new_[53425]_  = A201 & ~A200;
  assign \new_[53426]_  = A199 & \new_[53425]_ ;
  assign \new_[53427]_  = \new_[53426]_  & \new_[53421]_ ;
  assign \new_[53431]_  = A269 & ~A267;
  assign \new_[53432]_  = A203 & \new_[53431]_ ;
  assign \new_[53435]_  = A299 & ~A298;
  assign \new_[53438]_  = A302 & A300;
  assign \new_[53439]_  = \new_[53438]_  & \new_[53435]_ ;
  assign \new_[53440]_  = \new_[53439]_  & \new_[53432]_ ;
  assign \new_[53444]_  = A168 & ~A169;
  assign \new_[53445]_  = A170 & \new_[53444]_ ;
  assign \new_[53449]_  = A201 & ~A200;
  assign \new_[53450]_  = A199 & \new_[53449]_ ;
  assign \new_[53451]_  = \new_[53450]_  & \new_[53445]_ ;
  assign \new_[53455]_  = A266 & A265;
  assign \new_[53456]_  = A203 & \new_[53455]_ ;
  assign \new_[53459]_  = ~A299 & A298;
  assign \new_[53462]_  = A301 & A300;
  assign \new_[53463]_  = \new_[53462]_  & \new_[53459]_ ;
  assign \new_[53464]_  = \new_[53463]_  & \new_[53456]_ ;
  assign \new_[53468]_  = A168 & ~A169;
  assign \new_[53469]_  = A170 & \new_[53468]_ ;
  assign \new_[53473]_  = A201 & ~A200;
  assign \new_[53474]_  = A199 & \new_[53473]_ ;
  assign \new_[53475]_  = \new_[53474]_  & \new_[53469]_ ;
  assign \new_[53479]_  = A266 & A265;
  assign \new_[53480]_  = A203 & \new_[53479]_ ;
  assign \new_[53483]_  = ~A299 & A298;
  assign \new_[53486]_  = A302 & A300;
  assign \new_[53487]_  = \new_[53486]_  & \new_[53483]_ ;
  assign \new_[53488]_  = \new_[53487]_  & \new_[53480]_ ;
  assign \new_[53492]_  = A168 & ~A169;
  assign \new_[53493]_  = A170 & \new_[53492]_ ;
  assign \new_[53497]_  = A201 & ~A200;
  assign \new_[53498]_  = A199 & \new_[53497]_ ;
  assign \new_[53499]_  = \new_[53498]_  & \new_[53493]_ ;
  assign \new_[53503]_  = A266 & A265;
  assign \new_[53504]_  = A203 & \new_[53503]_ ;
  assign \new_[53507]_  = A299 & ~A298;
  assign \new_[53510]_  = A301 & A300;
  assign \new_[53511]_  = \new_[53510]_  & \new_[53507]_ ;
  assign \new_[53512]_  = \new_[53511]_  & \new_[53504]_ ;
  assign \new_[53516]_  = A168 & ~A169;
  assign \new_[53517]_  = A170 & \new_[53516]_ ;
  assign \new_[53521]_  = A201 & ~A200;
  assign \new_[53522]_  = A199 & \new_[53521]_ ;
  assign \new_[53523]_  = \new_[53522]_  & \new_[53517]_ ;
  assign \new_[53527]_  = A266 & A265;
  assign \new_[53528]_  = A203 & \new_[53527]_ ;
  assign \new_[53531]_  = A299 & ~A298;
  assign \new_[53534]_  = A302 & A300;
  assign \new_[53535]_  = \new_[53534]_  & \new_[53531]_ ;
  assign \new_[53536]_  = \new_[53535]_  & \new_[53528]_ ;
  assign \new_[53540]_  = A168 & ~A169;
  assign \new_[53541]_  = A170 & \new_[53540]_ ;
  assign \new_[53545]_  = A201 & ~A200;
  assign \new_[53546]_  = A199 & \new_[53545]_ ;
  assign \new_[53547]_  = \new_[53546]_  & \new_[53541]_ ;
  assign \new_[53551]_  = ~A266 & ~A265;
  assign \new_[53552]_  = A203 & \new_[53551]_ ;
  assign \new_[53555]_  = ~A299 & A298;
  assign \new_[53558]_  = A301 & A300;
  assign \new_[53559]_  = \new_[53558]_  & \new_[53555]_ ;
  assign \new_[53560]_  = \new_[53559]_  & \new_[53552]_ ;
  assign \new_[53564]_  = A168 & ~A169;
  assign \new_[53565]_  = A170 & \new_[53564]_ ;
  assign \new_[53569]_  = A201 & ~A200;
  assign \new_[53570]_  = A199 & \new_[53569]_ ;
  assign \new_[53571]_  = \new_[53570]_  & \new_[53565]_ ;
  assign \new_[53575]_  = ~A266 & ~A265;
  assign \new_[53576]_  = A203 & \new_[53575]_ ;
  assign \new_[53579]_  = ~A299 & A298;
  assign \new_[53582]_  = A302 & A300;
  assign \new_[53583]_  = \new_[53582]_  & \new_[53579]_ ;
  assign \new_[53584]_  = \new_[53583]_  & \new_[53576]_ ;
  assign \new_[53588]_  = A168 & ~A169;
  assign \new_[53589]_  = A170 & \new_[53588]_ ;
  assign \new_[53593]_  = A201 & ~A200;
  assign \new_[53594]_  = A199 & \new_[53593]_ ;
  assign \new_[53595]_  = \new_[53594]_  & \new_[53589]_ ;
  assign \new_[53599]_  = ~A266 & ~A265;
  assign \new_[53600]_  = A203 & \new_[53599]_ ;
  assign \new_[53603]_  = A299 & ~A298;
  assign \new_[53606]_  = A301 & A300;
  assign \new_[53607]_  = \new_[53606]_  & \new_[53603]_ ;
  assign \new_[53608]_  = \new_[53607]_  & \new_[53600]_ ;
  assign \new_[53612]_  = A168 & ~A169;
  assign \new_[53613]_  = A170 & \new_[53612]_ ;
  assign \new_[53617]_  = A201 & ~A200;
  assign \new_[53618]_  = A199 & \new_[53617]_ ;
  assign \new_[53619]_  = \new_[53618]_  & \new_[53613]_ ;
  assign \new_[53623]_  = ~A266 & ~A265;
  assign \new_[53624]_  = A203 & \new_[53623]_ ;
  assign \new_[53627]_  = A299 & ~A298;
  assign \new_[53630]_  = A302 & A300;
  assign \new_[53631]_  = \new_[53630]_  & \new_[53627]_ ;
  assign \new_[53632]_  = \new_[53631]_  & \new_[53624]_ ;
  assign \new_[53636]_  = A168 & ~A169;
  assign \new_[53637]_  = A170 & \new_[53636]_ ;
  assign \new_[53641]_  = ~A265 & ~A200;
  assign \new_[53642]_  = ~A199 & \new_[53641]_ ;
  assign \new_[53643]_  = \new_[53642]_  & \new_[53637]_ ;
  assign \new_[53647]_  = ~A268 & ~A267;
  assign \new_[53648]_  = A266 & \new_[53647]_ ;
  assign \new_[53651]_  = A300 & ~A269;
  assign \new_[53654]_  = ~A302 & ~A301;
  assign \new_[53655]_  = \new_[53654]_  & \new_[53651]_ ;
  assign \new_[53656]_  = \new_[53655]_  & \new_[53648]_ ;
  assign \new_[53660]_  = A168 & ~A169;
  assign \new_[53661]_  = A170 & \new_[53660]_ ;
  assign \new_[53665]_  = A265 & ~A200;
  assign \new_[53666]_  = ~A199 & \new_[53665]_ ;
  assign \new_[53667]_  = \new_[53666]_  & \new_[53661]_ ;
  assign \new_[53671]_  = ~A268 & ~A267;
  assign \new_[53672]_  = ~A266 & \new_[53671]_ ;
  assign \new_[53675]_  = A300 & ~A269;
  assign \new_[53678]_  = ~A302 & ~A301;
  assign \new_[53679]_  = \new_[53678]_  & \new_[53675]_ ;
  assign \new_[53680]_  = \new_[53679]_  & \new_[53672]_ ;
  assign \new_[53684]_  = ~A168 & ~A169;
  assign \new_[53685]_  = A170 & \new_[53684]_ ;
  assign \new_[53689]_  = ~A201 & ~A166;
  assign \new_[53690]_  = A167 & \new_[53689]_ ;
  assign \new_[53691]_  = \new_[53690]_  & \new_[53685]_ ;
  assign \new_[53695]_  = A268 & ~A267;
  assign \new_[53696]_  = A202 & \new_[53695]_ ;
  assign \new_[53699]_  = ~A299 & A298;
  assign \new_[53702]_  = A301 & A300;
  assign \new_[53703]_  = \new_[53702]_  & \new_[53699]_ ;
  assign \new_[53704]_  = \new_[53703]_  & \new_[53696]_ ;
  assign \new_[53708]_  = ~A168 & ~A169;
  assign \new_[53709]_  = A170 & \new_[53708]_ ;
  assign \new_[53713]_  = ~A201 & ~A166;
  assign \new_[53714]_  = A167 & \new_[53713]_ ;
  assign \new_[53715]_  = \new_[53714]_  & \new_[53709]_ ;
  assign \new_[53719]_  = A268 & ~A267;
  assign \new_[53720]_  = A202 & \new_[53719]_ ;
  assign \new_[53723]_  = ~A299 & A298;
  assign \new_[53726]_  = A302 & A300;
  assign \new_[53727]_  = \new_[53726]_  & \new_[53723]_ ;
  assign \new_[53728]_  = \new_[53727]_  & \new_[53720]_ ;
  assign \new_[53732]_  = ~A168 & ~A169;
  assign \new_[53733]_  = A170 & \new_[53732]_ ;
  assign \new_[53737]_  = ~A201 & ~A166;
  assign \new_[53738]_  = A167 & \new_[53737]_ ;
  assign \new_[53739]_  = \new_[53738]_  & \new_[53733]_ ;
  assign \new_[53743]_  = A268 & ~A267;
  assign \new_[53744]_  = A202 & \new_[53743]_ ;
  assign \new_[53747]_  = A299 & ~A298;
  assign \new_[53750]_  = A301 & A300;
  assign \new_[53751]_  = \new_[53750]_  & \new_[53747]_ ;
  assign \new_[53752]_  = \new_[53751]_  & \new_[53744]_ ;
  assign \new_[53756]_  = ~A168 & ~A169;
  assign \new_[53757]_  = A170 & \new_[53756]_ ;
  assign \new_[53761]_  = ~A201 & ~A166;
  assign \new_[53762]_  = A167 & \new_[53761]_ ;
  assign \new_[53763]_  = \new_[53762]_  & \new_[53757]_ ;
  assign \new_[53767]_  = A268 & ~A267;
  assign \new_[53768]_  = A202 & \new_[53767]_ ;
  assign \new_[53771]_  = A299 & ~A298;
  assign \new_[53774]_  = A302 & A300;
  assign \new_[53775]_  = \new_[53774]_  & \new_[53771]_ ;
  assign \new_[53776]_  = \new_[53775]_  & \new_[53768]_ ;
  assign \new_[53780]_  = ~A168 & ~A169;
  assign \new_[53781]_  = A170 & \new_[53780]_ ;
  assign \new_[53785]_  = ~A201 & ~A166;
  assign \new_[53786]_  = A167 & \new_[53785]_ ;
  assign \new_[53787]_  = \new_[53786]_  & \new_[53781]_ ;
  assign \new_[53791]_  = A269 & ~A267;
  assign \new_[53792]_  = A202 & \new_[53791]_ ;
  assign \new_[53795]_  = ~A299 & A298;
  assign \new_[53798]_  = A301 & A300;
  assign \new_[53799]_  = \new_[53798]_  & \new_[53795]_ ;
  assign \new_[53800]_  = \new_[53799]_  & \new_[53792]_ ;
  assign \new_[53804]_  = ~A168 & ~A169;
  assign \new_[53805]_  = A170 & \new_[53804]_ ;
  assign \new_[53809]_  = ~A201 & ~A166;
  assign \new_[53810]_  = A167 & \new_[53809]_ ;
  assign \new_[53811]_  = \new_[53810]_  & \new_[53805]_ ;
  assign \new_[53815]_  = A269 & ~A267;
  assign \new_[53816]_  = A202 & \new_[53815]_ ;
  assign \new_[53819]_  = ~A299 & A298;
  assign \new_[53822]_  = A302 & A300;
  assign \new_[53823]_  = \new_[53822]_  & \new_[53819]_ ;
  assign \new_[53824]_  = \new_[53823]_  & \new_[53816]_ ;
  assign \new_[53828]_  = ~A168 & ~A169;
  assign \new_[53829]_  = A170 & \new_[53828]_ ;
  assign \new_[53833]_  = ~A201 & ~A166;
  assign \new_[53834]_  = A167 & \new_[53833]_ ;
  assign \new_[53835]_  = \new_[53834]_  & \new_[53829]_ ;
  assign \new_[53839]_  = A269 & ~A267;
  assign \new_[53840]_  = A202 & \new_[53839]_ ;
  assign \new_[53843]_  = A299 & ~A298;
  assign \new_[53846]_  = A301 & A300;
  assign \new_[53847]_  = \new_[53846]_  & \new_[53843]_ ;
  assign \new_[53848]_  = \new_[53847]_  & \new_[53840]_ ;
  assign \new_[53852]_  = ~A168 & ~A169;
  assign \new_[53853]_  = A170 & \new_[53852]_ ;
  assign \new_[53857]_  = ~A201 & ~A166;
  assign \new_[53858]_  = A167 & \new_[53857]_ ;
  assign \new_[53859]_  = \new_[53858]_  & \new_[53853]_ ;
  assign \new_[53863]_  = A269 & ~A267;
  assign \new_[53864]_  = A202 & \new_[53863]_ ;
  assign \new_[53867]_  = A299 & ~A298;
  assign \new_[53870]_  = A302 & A300;
  assign \new_[53871]_  = \new_[53870]_  & \new_[53867]_ ;
  assign \new_[53872]_  = \new_[53871]_  & \new_[53864]_ ;
  assign \new_[53876]_  = ~A168 & ~A169;
  assign \new_[53877]_  = A170 & \new_[53876]_ ;
  assign \new_[53881]_  = ~A201 & ~A166;
  assign \new_[53882]_  = A167 & \new_[53881]_ ;
  assign \new_[53883]_  = \new_[53882]_  & \new_[53877]_ ;
  assign \new_[53887]_  = A266 & A265;
  assign \new_[53888]_  = A202 & \new_[53887]_ ;
  assign \new_[53891]_  = ~A299 & A298;
  assign \new_[53894]_  = A301 & A300;
  assign \new_[53895]_  = \new_[53894]_  & \new_[53891]_ ;
  assign \new_[53896]_  = \new_[53895]_  & \new_[53888]_ ;
  assign \new_[53900]_  = ~A168 & ~A169;
  assign \new_[53901]_  = A170 & \new_[53900]_ ;
  assign \new_[53905]_  = ~A201 & ~A166;
  assign \new_[53906]_  = A167 & \new_[53905]_ ;
  assign \new_[53907]_  = \new_[53906]_  & \new_[53901]_ ;
  assign \new_[53911]_  = A266 & A265;
  assign \new_[53912]_  = A202 & \new_[53911]_ ;
  assign \new_[53915]_  = ~A299 & A298;
  assign \new_[53918]_  = A302 & A300;
  assign \new_[53919]_  = \new_[53918]_  & \new_[53915]_ ;
  assign \new_[53920]_  = \new_[53919]_  & \new_[53912]_ ;
  assign \new_[53924]_  = ~A168 & ~A169;
  assign \new_[53925]_  = A170 & \new_[53924]_ ;
  assign \new_[53929]_  = ~A201 & ~A166;
  assign \new_[53930]_  = A167 & \new_[53929]_ ;
  assign \new_[53931]_  = \new_[53930]_  & \new_[53925]_ ;
  assign \new_[53935]_  = A266 & A265;
  assign \new_[53936]_  = A202 & \new_[53935]_ ;
  assign \new_[53939]_  = A299 & ~A298;
  assign \new_[53942]_  = A301 & A300;
  assign \new_[53943]_  = \new_[53942]_  & \new_[53939]_ ;
  assign \new_[53944]_  = \new_[53943]_  & \new_[53936]_ ;
  assign \new_[53948]_  = ~A168 & ~A169;
  assign \new_[53949]_  = A170 & \new_[53948]_ ;
  assign \new_[53953]_  = ~A201 & ~A166;
  assign \new_[53954]_  = A167 & \new_[53953]_ ;
  assign \new_[53955]_  = \new_[53954]_  & \new_[53949]_ ;
  assign \new_[53959]_  = A266 & A265;
  assign \new_[53960]_  = A202 & \new_[53959]_ ;
  assign \new_[53963]_  = A299 & ~A298;
  assign \new_[53966]_  = A302 & A300;
  assign \new_[53967]_  = \new_[53966]_  & \new_[53963]_ ;
  assign \new_[53968]_  = \new_[53967]_  & \new_[53960]_ ;
  assign \new_[53972]_  = ~A168 & ~A169;
  assign \new_[53973]_  = A170 & \new_[53972]_ ;
  assign \new_[53977]_  = ~A201 & ~A166;
  assign \new_[53978]_  = A167 & \new_[53977]_ ;
  assign \new_[53979]_  = \new_[53978]_  & \new_[53973]_ ;
  assign \new_[53983]_  = ~A266 & ~A265;
  assign \new_[53984]_  = A202 & \new_[53983]_ ;
  assign \new_[53987]_  = ~A299 & A298;
  assign \new_[53990]_  = A301 & A300;
  assign \new_[53991]_  = \new_[53990]_  & \new_[53987]_ ;
  assign \new_[53992]_  = \new_[53991]_  & \new_[53984]_ ;
  assign \new_[53996]_  = ~A168 & ~A169;
  assign \new_[53997]_  = A170 & \new_[53996]_ ;
  assign \new_[54001]_  = ~A201 & ~A166;
  assign \new_[54002]_  = A167 & \new_[54001]_ ;
  assign \new_[54003]_  = \new_[54002]_  & \new_[53997]_ ;
  assign \new_[54007]_  = ~A266 & ~A265;
  assign \new_[54008]_  = A202 & \new_[54007]_ ;
  assign \new_[54011]_  = ~A299 & A298;
  assign \new_[54014]_  = A302 & A300;
  assign \new_[54015]_  = \new_[54014]_  & \new_[54011]_ ;
  assign \new_[54016]_  = \new_[54015]_  & \new_[54008]_ ;
  assign \new_[54020]_  = ~A168 & ~A169;
  assign \new_[54021]_  = A170 & \new_[54020]_ ;
  assign \new_[54025]_  = ~A201 & ~A166;
  assign \new_[54026]_  = A167 & \new_[54025]_ ;
  assign \new_[54027]_  = \new_[54026]_  & \new_[54021]_ ;
  assign \new_[54031]_  = ~A266 & ~A265;
  assign \new_[54032]_  = A202 & \new_[54031]_ ;
  assign \new_[54035]_  = A299 & ~A298;
  assign \new_[54038]_  = A301 & A300;
  assign \new_[54039]_  = \new_[54038]_  & \new_[54035]_ ;
  assign \new_[54040]_  = \new_[54039]_  & \new_[54032]_ ;
  assign \new_[54044]_  = ~A168 & ~A169;
  assign \new_[54045]_  = A170 & \new_[54044]_ ;
  assign \new_[54049]_  = ~A201 & ~A166;
  assign \new_[54050]_  = A167 & \new_[54049]_ ;
  assign \new_[54051]_  = \new_[54050]_  & \new_[54045]_ ;
  assign \new_[54055]_  = ~A266 & ~A265;
  assign \new_[54056]_  = A202 & \new_[54055]_ ;
  assign \new_[54059]_  = A299 & ~A298;
  assign \new_[54062]_  = A302 & A300;
  assign \new_[54063]_  = \new_[54062]_  & \new_[54059]_ ;
  assign \new_[54064]_  = \new_[54063]_  & \new_[54056]_ ;
  assign \new_[54068]_  = ~A168 & ~A169;
  assign \new_[54069]_  = A170 & \new_[54068]_ ;
  assign \new_[54073]_  = ~A201 & ~A166;
  assign \new_[54074]_  = A167 & \new_[54073]_ ;
  assign \new_[54075]_  = \new_[54074]_  & \new_[54069]_ ;
  assign \new_[54079]_  = A268 & ~A267;
  assign \new_[54080]_  = A203 & \new_[54079]_ ;
  assign \new_[54083]_  = ~A299 & A298;
  assign \new_[54086]_  = A301 & A300;
  assign \new_[54087]_  = \new_[54086]_  & \new_[54083]_ ;
  assign \new_[54088]_  = \new_[54087]_  & \new_[54080]_ ;
  assign \new_[54092]_  = ~A168 & ~A169;
  assign \new_[54093]_  = A170 & \new_[54092]_ ;
  assign \new_[54097]_  = ~A201 & ~A166;
  assign \new_[54098]_  = A167 & \new_[54097]_ ;
  assign \new_[54099]_  = \new_[54098]_  & \new_[54093]_ ;
  assign \new_[54103]_  = A268 & ~A267;
  assign \new_[54104]_  = A203 & \new_[54103]_ ;
  assign \new_[54107]_  = ~A299 & A298;
  assign \new_[54110]_  = A302 & A300;
  assign \new_[54111]_  = \new_[54110]_  & \new_[54107]_ ;
  assign \new_[54112]_  = \new_[54111]_  & \new_[54104]_ ;
  assign \new_[54116]_  = ~A168 & ~A169;
  assign \new_[54117]_  = A170 & \new_[54116]_ ;
  assign \new_[54121]_  = ~A201 & ~A166;
  assign \new_[54122]_  = A167 & \new_[54121]_ ;
  assign \new_[54123]_  = \new_[54122]_  & \new_[54117]_ ;
  assign \new_[54127]_  = A268 & ~A267;
  assign \new_[54128]_  = A203 & \new_[54127]_ ;
  assign \new_[54131]_  = A299 & ~A298;
  assign \new_[54134]_  = A301 & A300;
  assign \new_[54135]_  = \new_[54134]_  & \new_[54131]_ ;
  assign \new_[54136]_  = \new_[54135]_  & \new_[54128]_ ;
  assign \new_[54140]_  = ~A168 & ~A169;
  assign \new_[54141]_  = A170 & \new_[54140]_ ;
  assign \new_[54145]_  = ~A201 & ~A166;
  assign \new_[54146]_  = A167 & \new_[54145]_ ;
  assign \new_[54147]_  = \new_[54146]_  & \new_[54141]_ ;
  assign \new_[54151]_  = A268 & ~A267;
  assign \new_[54152]_  = A203 & \new_[54151]_ ;
  assign \new_[54155]_  = A299 & ~A298;
  assign \new_[54158]_  = A302 & A300;
  assign \new_[54159]_  = \new_[54158]_  & \new_[54155]_ ;
  assign \new_[54160]_  = \new_[54159]_  & \new_[54152]_ ;
  assign \new_[54164]_  = ~A168 & ~A169;
  assign \new_[54165]_  = A170 & \new_[54164]_ ;
  assign \new_[54169]_  = ~A201 & ~A166;
  assign \new_[54170]_  = A167 & \new_[54169]_ ;
  assign \new_[54171]_  = \new_[54170]_  & \new_[54165]_ ;
  assign \new_[54175]_  = A269 & ~A267;
  assign \new_[54176]_  = A203 & \new_[54175]_ ;
  assign \new_[54179]_  = ~A299 & A298;
  assign \new_[54182]_  = A301 & A300;
  assign \new_[54183]_  = \new_[54182]_  & \new_[54179]_ ;
  assign \new_[54184]_  = \new_[54183]_  & \new_[54176]_ ;
  assign \new_[54188]_  = ~A168 & ~A169;
  assign \new_[54189]_  = A170 & \new_[54188]_ ;
  assign \new_[54193]_  = ~A201 & ~A166;
  assign \new_[54194]_  = A167 & \new_[54193]_ ;
  assign \new_[54195]_  = \new_[54194]_  & \new_[54189]_ ;
  assign \new_[54199]_  = A269 & ~A267;
  assign \new_[54200]_  = A203 & \new_[54199]_ ;
  assign \new_[54203]_  = ~A299 & A298;
  assign \new_[54206]_  = A302 & A300;
  assign \new_[54207]_  = \new_[54206]_  & \new_[54203]_ ;
  assign \new_[54208]_  = \new_[54207]_  & \new_[54200]_ ;
  assign \new_[54212]_  = ~A168 & ~A169;
  assign \new_[54213]_  = A170 & \new_[54212]_ ;
  assign \new_[54217]_  = ~A201 & ~A166;
  assign \new_[54218]_  = A167 & \new_[54217]_ ;
  assign \new_[54219]_  = \new_[54218]_  & \new_[54213]_ ;
  assign \new_[54223]_  = A269 & ~A267;
  assign \new_[54224]_  = A203 & \new_[54223]_ ;
  assign \new_[54227]_  = A299 & ~A298;
  assign \new_[54230]_  = A301 & A300;
  assign \new_[54231]_  = \new_[54230]_  & \new_[54227]_ ;
  assign \new_[54232]_  = \new_[54231]_  & \new_[54224]_ ;
  assign \new_[54236]_  = ~A168 & ~A169;
  assign \new_[54237]_  = A170 & \new_[54236]_ ;
  assign \new_[54241]_  = ~A201 & ~A166;
  assign \new_[54242]_  = A167 & \new_[54241]_ ;
  assign \new_[54243]_  = \new_[54242]_  & \new_[54237]_ ;
  assign \new_[54247]_  = A269 & ~A267;
  assign \new_[54248]_  = A203 & \new_[54247]_ ;
  assign \new_[54251]_  = A299 & ~A298;
  assign \new_[54254]_  = A302 & A300;
  assign \new_[54255]_  = \new_[54254]_  & \new_[54251]_ ;
  assign \new_[54256]_  = \new_[54255]_  & \new_[54248]_ ;
  assign \new_[54260]_  = ~A168 & ~A169;
  assign \new_[54261]_  = A170 & \new_[54260]_ ;
  assign \new_[54265]_  = ~A201 & ~A166;
  assign \new_[54266]_  = A167 & \new_[54265]_ ;
  assign \new_[54267]_  = \new_[54266]_  & \new_[54261]_ ;
  assign \new_[54271]_  = A266 & A265;
  assign \new_[54272]_  = A203 & \new_[54271]_ ;
  assign \new_[54275]_  = ~A299 & A298;
  assign \new_[54278]_  = A301 & A300;
  assign \new_[54279]_  = \new_[54278]_  & \new_[54275]_ ;
  assign \new_[54280]_  = \new_[54279]_  & \new_[54272]_ ;
  assign \new_[54284]_  = ~A168 & ~A169;
  assign \new_[54285]_  = A170 & \new_[54284]_ ;
  assign \new_[54289]_  = ~A201 & ~A166;
  assign \new_[54290]_  = A167 & \new_[54289]_ ;
  assign \new_[54291]_  = \new_[54290]_  & \new_[54285]_ ;
  assign \new_[54295]_  = A266 & A265;
  assign \new_[54296]_  = A203 & \new_[54295]_ ;
  assign \new_[54299]_  = ~A299 & A298;
  assign \new_[54302]_  = A302 & A300;
  assign \new_[54303]_  = \new_[54302]_  & \new_[54299]_ ;
  assign \new_[54304]_  = \new_[54303]_  & \new_[54296]_ ;
  assign \new_[54308]_  = ~A168 & ~A169;
  assign \new_[54309]_  = A170 & \new_[54308]_ ;
  assign \new_[54313]_  = ~A201 & ~A166;
  assign \new_[54314]_  = A167 & \new_[54313]_ ;
  assign \new_[54315]_  = \new_[54314]_  & \new_[54309]_ ;
  assign \new_[54319]_  = A266 & A265;
  assign \new_[54320]_  = A203 & \new_[54319]_ ;
  assign \new_[54323]_  = A299 & ~A298;
  assign \new_[54326]_  = A301 & A300;
  assign \new_[54327]_  = \new_[54326]_  & \new_[54323]_ ;
  assign \new_[54328]_  = \new_[54327]_  & \new_[54320]_ ;
  assign \new_[54332]_  = ~A168 & ~A169;
  assign \new_[54333]_  = A170 & \new_[54332]_ ;
  assign \new_[54337]_  = ~A201 & ~A166;
  assign \new_[54338]_  = A167 & \new_[54337]_ ;
  assign \new_[54339]_  = \new_[54338]_  & \new_[54333]_ ;
  assign \new_[54343]_  = A266 & A265;
  assign \new_[54344]_  = A203 & \new_[54343]_ ;
  assign \new_[54347]_  = A299 & ~A298;
  assign \new_[54350]_  = A302 & A300;
  assign \new_[54351]_  = \new_[54350]_  & \new_[54347]_ ;
  assign \new_[54352]_  = \new_[54351]_  & \new_[54344]_ ;
  assign \new_[54356]_  = ~A168 & ~A169;
  assign \new_[54357]_  = A170 & \new_[54356]_ ;
  assign \new_[54361]_  = ~A201 & ~A166;
  assign \new_[54362]_  = A167 & \new_[54361]_ ;
  assign \new_[54363]_  = \new_[54362]_  & \new_[54357]_ ;
  assign \new_[54367]_  = ~A266 & ~A265;
  assign \new_[54368]_  = A203 & \new_[54367]_ ;
  assign \new_[54371]_  = ~A299 & A298;
  assign \new_[54374]_  = A301 & A300;
  assign \new_[54375]_  = \new_[54374]_  & \new_[54371]_ ;
  assign \new_[54376]_  = \new_[54375]_  & \new_[54368]_ ;
  assign \new_[54380]_  = ~A168 & ~A169;
  assign \new_[54381]_  = A170 & \new_[54380]_ ;
  assign \new_[54385]_  = ~A201 & ~A166;
  assign \new_[54386]_  = A167 & \new_[54385]_ ;
  assign \new_[54387]_  = \new_[54386]_  & \new_[54381]_ ;
  assign \new_[54391]_  = ~A266 & ~A265;
  assign \new_[54392]_  = A203 & \new_[54391]_ ;
  assign \new_[54395]_  = ~A299 & A298;
  assign \new_[54398]_  = A302 & A300;
  assign \new_[54399]_  = \new_[54398]_  & \new_[54395]_ ;
  assign \new_[54400]_  = \new_[54399]_  & \new_[54392]_ ;
  assign \new_[54404]_  = ~A168 & ~A169;
  assign \new_[54405]_  = A170 & \new_[54404]_ ;
  assign \new_[54409]_  = ~A201 & ~A166;
  assign \new_[54410]_  = A167 & \new_[54409]_ ;
  assign \new_[54411]_  = \new_[54410]_  & \new_[54405]_ ;
  assign \new_[54415]_  = ~A266 & ~A265;
  assign \new_[54416]_  = A203 & \new_[54415]_ ;
  assign \new_[54419]_  = A299 & ~A298;
  assign \new_[54422]_  = A301 & A300;
  assign \new_[54423]_  = \new_[54422]_  & \new_[54419]_ ;
  assign \new_[54424]_  = \new_[54423]_  & \new_[54416]_ ;
  assign \new_[54428]_  = ~A168 & ~A169;
  assign \new_[54429]_  = A170 & \new_[54428]_ ;
  assign \new_[54433]_  = ~A201 & ~A166;
  assign \new_[54434]_  = A167 & \new_[54433]_ ;
  assign \new_[54435]_  = \new_[54434]_  & \new_[54429]_ ;
  assign \new_[54439]_  = ~A266 & ~A265;
  assign \new_[54440]_  = A203 & \new_[54439]_ ;
  assign \new_[54443]_  = A299 & ~A298;
  assign \new_[54446]_  = A302 & A300;
  assign \new_[54447]_  = \new_[54446]_  & \new_[54443]_ ;
  assign \new_[54448]_  = \new_[54447]_  & \new_[54440]_ ;
  assign \new_[54452]_  = ~A168 & ~A169;
  assign \new_[54453]_  = A170 & \new_[54452]_ ;
  assign \new_[54457]_  = A199 & ~A166;
  assign \new_[54458]_  = A167 & \new_[54457]_ ;
  assign \new_[54459]_  = \new_[54458]_  & \new_[54453]_ ;
  assign \new_[54463]_  = A268 & ~A267;
  assign \new_[54464]_  = A200 & \new_[54463]_ ;
  assign \new_[54467]_  = ~A299 & A298;
  assign \new_[54470]_  = A301 & A300;
  assign \new_[54471]_  = \new_[54470]_  & \new_[54467]_ ;
  assign \new_[54472]_  = \new_[54471]_  & \new_[54464]_ ;
  assign \new_[54476]_  = ~A168 & ~A169;
  assign \new_[54477]_  = A170 & \new_[54476]_ ;
  assign \new_[54481]_  = A199 & ~A166;
  assign \new_[54482]_  = A167 & \new_[54481]_ ;
  assign \new_[54483]_  = \new_[54482]_  & \new_[54477]_ ;
  assign \new_[54487]_  = A268 & ~A267;
  assign \new_[54488]_  = A200 & \new_[54487]_ ;
  assign \new_[54491]_  = ~A299 & A298;
  assign \new_[54494]_  = A302 & A300;
  assign \new_[54495]_  = \new_[54494]_  & \new_[54491]_ ;
  assign \new_[54496]_  = \new_[54495]_  & \new_[54488]_ ;
  assign \new_[54500]_  = ~A168 & ~A169;
  assign \new_[54501]_  = A170 & \new_[54500]_ ;
  assign \new_[54505]_  = A199 & ~A166;
  assign \new_[54506]_  = A167 & \new_[54505]_ ;
  assign \new_[54507]_  = \new_[54506]_  & \new_[54501]_ ;
  assign \new_[54511]_  = A268 & ~A267;
  assign \new_[54512]_  = A200 & \new_[54511]_ ;
  assign \new_[54515]_  = A299 & ~A298;
  assign \new_[54518]_  = A301 & A300;
  assign \new_[54519]_  = \new_[54518]_  & \new_[54515]_ ;
  assign \new_[54520]_  = \new_[54519]_  & \new_[54512]_ ;
  assign \new_[54524]_  = ~A168 & ~A169;
  assign \new_[54525]_  = A170 & \new_[54524]_ ;
  assign \new_[54529]_  = A199 & ~A166;
  assign \new_[54530]_  = A167 & \new_[54529]_ ;
  assign \new_[54531]_  = \new_[54530]_  & \new_[54525]_ ;
  assign \new_[54535]_  = A268 & ~A267;
  assign \new_[54536]_  = A200 & \new_[54535]_ ;
  assign \new_[54539]_  = A299 & ~A298;
  assign \new_[54542]_  = A302 & A300;
  assign \new_[54543]_  = \new_[54542]_  & \new_[54539]_ ;
  assign \new_[54544]_  = \new_[54543]_  & \new_[54536]_ ;
  assign \new_[54548]_  = ~A168 & ~A169;
  assign \new_[54549]_  = A170 & \new_[54548]_ ;
  assign \new_[54553]_  = A199 & ~A166;
  assign \new_[54554]_  = A167 & \new_[54553]_ ;
  assign \new_[54555]_  = \new_[54554]_  & \new_[54549]_ ;
  assign \new_[54559]_  = A269 & ~A267;
  assign \new_[54560]_  = A200 & \new_[54559]_ ;
  assign \new_[54563]_  = ~A299 & A298;
  assign \new_[54566]_  = A301 & A300;
  assign \new_[54567]_  = \new_[54566]_  & \new_[54563]_ ;
  assign \new_[54568]_  = \new_[54567]_  & \new_[54560]_ ;
  assign \new_[54572]_  = ~A168 & ~A169;
  assign \new_[54573]_  = A170 & \new_[54572]_ ;
  assign \new_[54577]_  = A199 & ~A166;
  assign \new_[54578]_  = A167 & \new_[54577]_ ;
  assign \new_[54579]_  = \new_[54578]_  & \new_[54573]_ ;
  assign \new_[54583]_  = A269 & ~A267;
  assign \new_[54584]_  = A200 & \new_[54583]_ ;
  assign \new_[54587]_  = ~A299 & A298;
  assign \new_[54590]_  = A302 & A300;
  assign \new_[54591]_  = \new_[54590]_  & \new_[54587]_ ;
  assign \new_[54592]_  = \new_[54591]_  & \new_[54584]_ ;
  assign \new_[54596]_  = ~A168 & ~A169;
  assign \new_[54597]_  = A170 & \new_[54596]_ ;
  assign \new_[54601]_  = A199 & ~A166;
  assign \new_[54602]_  = A167 & \new_[54601]_ ;
  assign \new_[54603]_  = \new_[54602]_  & \new_[54597]_ ;
  assign \new_[54607]_  = A269 & ~A267;
  assign \new_[54608]_  = A200 & \new_[54607]_ ;
  assign \new_[54611]_  = A299 & ~A298;
  assign \new_[54614]_  = A301 & A300;
  assign \new_[54615]_  = \new_[54614]_  & \new_[54611]_ ;
  assign \new_[54616]_  = \new_[54615]_  & \new_[54608]_ ;
  assign \new_[54620]_  = ~A168 & ~A169;
  assign \new_[54621]_  = A170 & \new_[54620]_ ;
  assign \new_[54625]_  = A199 & ~A166;
  assign \new_[54626]_  = A167 & \new_[54625]_ ;
  assign \new_[54627]_  = \new_[54626]_  & \new_[54621]_ ;
  assign \new_[54631]_  = A269 & ~A267;
  assign \new_[54632]_  = A200 & \new_[54631]_ ;
  assign \new_[54635]_  = A299 & ~A298;
  assign \new_[54638]_  = A302 & A300;
  assign \new_[54639]_  = \new_[54638]_  & \new_[54635]_ ;
  assign \new_[54640]_  = \new_[54639]_  & \new_[54632]_ ;
  assign \new_[54644]_  = ~A168 & ~A169;
  assign \new_[54645]_  = A170 & \new_[54644]_ ;
  assign \new_[54649]_  = A199 & ~A166;
  assign \new_[54650]_  = A167 & \new_[54649]_ ;
  assign \new_[54651]_  = \new_[54650]_  & \new_[54645]_ ;
  assign \new_[54655]_  = A266 & A265;
  assign \new_[54656]_  = A200 & \new_[54655]_ ;
  assign \new_[54659]_  = ~A299 & A298;
  assign \new_[54662]_  = A301 & A300;
  assign \new_[54663]_  = \new_[54662]_  & \new_[54659]_ ;
  assign \new_[54664]_  = \new_[54663]_  & \new_[54656]_ ;
  assign \new_[54668]_  = ~A168 & ~A169;
  assign \new_[54669]_  = A170 & \new_[54668]_ ;
  assign \new_[54673]_  = A199 & ~A166;
  assign \new_[54674]_  = A167 & \new_[54673]_ ;
  assign \new_[54675]_  = \new_[54674]_  & \new_[54669]_ ;
  assign \new_[54679]_  = A266 & A265;
  assign \new_[54680]_  = A200 & \new_[54679]_ ;
  assign \new_[54683]_  = ~A299 & A298;
  assign \new_[54686]_  = A302 & A300;
  assign \new_[54687]_  = \new_[54686]_  & \new_[54683]_ ;
  assign \new_[54688]_  = \new_[54687]_  & \new_[54680]_ ;
  assign \new_[54692]_  = ~A168 & ~A169;
  assign \new_[54693]_  = A170 & \new_[54692]_ ;
  assign \new_[54697]_  = A199 & ~A166;
  assign \new_[54698]_  = A167 & \new_[54697]_ ;
  assign \new_[54699]_  = \new_[54698]_  & \new_[54693]_ ;
  assign \new_[54703]_  = A266 & A265;
  assign \new_[54704]_  = A200 & \new_[54703]_ ;
  assign \new_[54707]_  = A299 & ~A298;
  assign \new_[54710]_  = A301 & A300;
  assign \new_[54711]_  = \new_[54710]_  & \new_[54707]_ ;
  assign \new_[54712]_  = \new_[54711]_  & \new_[54704]_ ;
  assign \new_[54716]_  = ~A168 & ~A169;
  assign \new_[54717]_  = A170 & \new_[54716]_ ;
  assign \new_[54721]_  = A199 & ~A166;
  assign \new_[54722]_  = A167 & \new_[54721]_ ;
  assign \new_[54723]_  = \new_[54722]_  & \new_[54717]_ ;
  assign \new_[54727]_  = A266 & A265;
  assign \new_[54728]_  = A200 & \new_[54727]_ ;
  assign \new_[54731]_  = A299 & ~A298;
  assign \new_[54734]_  = A302 & A300;
  assign \new_[54735]_  = \new_[54734]_  & \new_[54731]_ ;
  assign \new_[54736]_  = \new_[54735]_  & \new_[54728]_ ;
  assign \new_[54740]_  = ~A168 & ~A169;
  assign \new_[54741]_  = A170 & \new_[54740]_ ;
  assign \new_[54745]_  = A199 & ~A166;
  assign \new_[54746]_  = A167 & \new_[54745]_ ;
  assign \new_[54747]_  = \new_[54746]_  & \new_[54741]_ ;
  assign \new_[54751]_  = ~A266 & ~A265;
  assign \new_[54752]_  = A200 & \new_[54751]_ ;
  assign \new_[54755]_  = ~A299 & A298;
  assign \new_[54758]_  = A301 & A300;
  assign \new_[54759]_  = \new_[54758]_  & \new_[54755]_ ;
  assign \new_[54760]_  = \new_[54759]_  & \new_[54752]_ ;
  assign \new_[54764]_  = ~A168 & ~A169;
  assign \new_[54765]_  = A170 & \new_[54764]_ ;
  assign \new_[54769]_  = A199 & ~A166;
  assign \new_[54770]_  = A167 & \new_[54769]_ ;
  assign \new_[54771]_  = \new_[54770]_  & \new_[54765]_ ;
  assign \new_[54775]_  = ~A266 & ~A265;
  assign \new_[54776]_  = A200 & \new_[54775]_ ;
  assign \new_[54779]_  = ~A299 & A298;
  assign \new_[54782]_  = A302 & A300;
  assign \new_[54783]_  = \new_[54782]_  & \new_[54779]_ ;
  assign \new_[54784]_  = \new_[54783]_  & \new_[54776]_ ;
  assign \new_[54788]_  = ~A168 & ~A169;
  assign \new_[54789]_  = A170 & \new_[54788]_ ;
  assign \new_[54793]_  = A199 & ~A166;
  assign \new_[54794]_  = A167 & \new_[54793]_ ;
  assign \new_[54795]_  = \new_[54794]_  & \new_[54789]_ ;
  assign \new_[54799]_  = ~A266 & ~A265;
  assign \new_[54800]_  = A200 & \new_[54799]_ ;
  assign \new_[54803]_  = A299 & ~A298;
  assign \new_[54806]_  = A301 & A300;
  assign \new_[54807]_  = \new_[54806]_  & \new_[54803]_ ;
  assign \new_[54808]_  = \new_[54807]_  & \new_[54800]_ ;
  assign \new_[54812]_  = ~A168 & ~A169;
  assign \new_[54813]_  = A170 & \new_[54812]_ ;
  assign \new_[54817]_  = A199 & ~A166;
  assign \new_[54818]_  = A167 & \new_[54817]_ ;
  assign \new_[54819]_  = \new_[54818]_  & \new_[54813]_ ;
  assign \new_[54823]_  = ~A266 & ~A265;
  assign \new_[54824]_  = A200 & \new_[54823]_ ;
  assign \new_[54827]_  = A299 & ~A298;
  assign \new_[54830]_  = A302 & A300;
  assign \new_[54831]_  = \new_[54830]_  & \new_[54827]_ ;
  assign \new_[54832]_  = \new_[54831]_  & \new_[54824]_ ;
  assign \new_[54836]_  = ~A168 & ~A169;
  assign \new_[54837]_  = A170 & \new_[54836]_ ;
  assign \new_[54841]_  = ~A199 & ~A166;
  assign \new_[54842]_  = A167 & \new_[54841]_ ;
  assign \new_[54843]_  = \new_[54842]_  & \new_[54837]_ ;
  assign \new_[54847]_  = A268 & ~A267;
  assign \new_[54848]_  = ~A200 & \new_[54847]_ ;
  assign \new_[54851]_  = ~A299 & A298;
  assign \new_[54854]_  = A301 & A300;
  assign \new_[54855]_  = \new_[54854]_  & \new_[54851]_ ;
  assign \new_[54856]_  = \new_[54855]_  & \new_[54848]_ ;
  assign \new_[54860]_  = ~A168 & ~A169;
  assign \new_[54861]_  = A170 & \new_[54860]_ ;
  assign \new_[54865]_  = ~A199 & ~A166;
  assign \new_[54866]_  = A167 & \new_[54865]_ ;
  assign \new_[54867]_  = \new_[54866]_  & \new_[54861]_ ;
  assign \new_[54871]_  = A268 & ~A267;
  assign \new_[54872]_  = ~A200 & \new_[54871]_ ;
  assign \new_[54875]_  = ~A299 & A298;
  assign \new_[54878]_  = A302 & A300;
  assign \new_[54879]_  = \new_[54878]_  & \new_[54875]_ ;
  assign \new_[54880]_  = \new_[54879]_  & \new_[54872]_ ;
  assign \new_[54884]_  = ~A168 & ~A169;
  assign \new_[54885]_  = A170 & \new_[54884]_ ;
  assign \new_[54889]_  = ~A199 & ~A166;
  assign \new_[54890]_  = A167 & \new_[54889]_ ;
  assign \new_[54891]_  = \new_[54890]_  & \new_[54885]_ ;
  assign \new_[54895]_  = A268 & ~A267;
  assign \new_[54896]_  = ~A200 & \new_[54895]_ ;
  assign \new_[54899]_  = A299 & ~A298;
  assign \new_[54902]_  = A301 & A300;
  assign \new_[54903]_  = \new_[54902]_  & \new_[54899]_ ;
  assign \new_[54904]_  = \new_[54903]_  & \new_[54896]_ ;
  assign \new_[54908]_  = ~A168 & ~A169;
  assign \new_[54909]_  = A170 & \new_[54908]_ ;
  assign \new_[54913]_  = ~A199 & ~A166;
  assign \new_[54914]_  = A167 & \new_[54913]_ ;
  assign \new_[54915]_  = \new_[54914]_  & \new_[54909]_ ;
  assign \new_[54919]_  = A268 & ~A267;
  assign \new_[54920]_  = ~A200 & \new_[54919]_ ;
  assign \new_[54923]_  = A299 & ~A298;
  assign \new_[54926]_  = A302 & A300;
  assign \new_[54927]_  = \new_[54926]_  & \new_[54923]_ ;
  assign \new_[54928]_  = \new_[54927]_  & \new_[54920]_ ;
  assign \new_[54932]_  = ~A168 & ~A169;
  assign \new_[54933]_  = A170 & \new_[54932]_ ;
  assign \new_[54937]_  = ~A199 & ~A166;
  assign \new_[54938]_  = A167 & \new_[54937]_ ;
  assign \new_[54939]_  = \new_[54938]_  & \new_[54933]_ ;
  assign \new_[54943]_  = A269 & ~A267;
  assign \new_[54944]_  = ~A200 & \new_[54943]_ ;
  assign \new_[54947]_  = ~A299 & A298;
  assign \new_[54950]_  = A301 & A300;
  assign \new_[54951]_  = \new_[54950]_  & \new_[54947]_ ;
  assign \new_[54952]_  = \new_[54951]_  & \new_[54944]_ ;
  assign \new_[54956]_  = ~A168 & ~A169;
  assign \new_[54957]_  = A170 & \new_[54956]_ ;
  assign \new_[54961]_  = ~A199 & ~A166;
  assign \new_[54962]_  = A167 & \new_[54961]_ ;
  assign \new_[54963]_  = \new_[54962]_  & \new_[54957]_ ;
  assign \new_[54967]_  = A269 & ~A267;
  assign \new_[54968]_  = ~A200 & \new_[54967]_ ;
  assign \new_[54971]_  = ~A299 & A298;
  assign \new_[54974]_  = A302 & A300;
  assign \new_[54975]_  = \new_[54974]_  & \new_[54971]_ ;
  assign \new_[54976]_  = \new_[54975]_  & \new_[54968]_ ;
  assign \new_[54980]_  = ~A168 & ~A169;
  assign \new_[54981]_  = A170 & \new_[54980]_ ;
  assign \new_[54985]_  = ~A199 & ~A166;
  assign \new_[54986]_  = A167 & \new_[54985]_ ;
  assign \new_[54987]_  = \new_[54986]_  & \new_[54981]_ ;
  assign \new_[54991]_  = A269 & ~A267;
  assign \new_[54992]_  = ~A200 & \new_[54991]_ ;
  assign \new_[54995]_  = A299 & ~A298;
  assign \new_[54998]_  = A301 & A300;
  assign \new_[54999]_  = \new_[54998]_  & \new_[54995]_ ;
  assign \new_[55000]_  = \new_[54999]_  & \new_[54992]_ ;
  assign \new_[55004]_  = ~A168 & ~A169;
  assign \new_[55005]_  = A170 & \new_[55004]_ ;
  assign \new_[55009]_  = ~A199 & ~A166;
  assign \new_[55010]_  = A167 & \new_[55009]_ ;
  assign \new_[55011]_  = \new_[55010]_  & \new_[55005]_ ;
  assign \new_[55015]_  = A269 & ~A267;
  assign \new_[55016]_  = ~A200 & \new_[55015]_ ;
  assign \new_[55019]_  = A299 & ~A298;
  assign \new_[55022]_  = A302 & A300;
  assign \new_[55023]_  = \new_[55022]_  & \new_[55019]_ ;
  assign \new_[55024]_  = \new_[55023]_  & \new_[55016]_ ;
  assign \new_[55028]_  = ~A168 & ~A169;
  assign \new_[55029]_  = A170 & \new_[55028]_ ;
  assign \new_[55033]_  = ~A199 & ~A166;
  assign \new_[55034]_  = A167 & \new_[55033]_ ;
  assign \new_[55035]_  = \new_[55034]_  & \new_[55029]_ ;
  assign \new_[55039]_  = A266 & A265;
  assign \new_[55040]_  = ~A200 & \new_[55039]_ ;
  assign \new_[55043]_  = ~A299 & A298;
  assign \new_[55046]_  = A301 & A300;
  assign \new_[55047]_  = \new_[55046]_  & \new_[55043]_ ;
  assign \new_[55048]_  = \new_[55047]_  & \new_[55040]_ ;
  assign \new_[55052]_  = ~A168 & ~A169;
  assign \new_[55053]_  = A170 & \new_[55052]_ ;
  assign \new_[55057]_  = ~A199 & ~A166;
  assign \new_[55058]_  = A167 & \new_[55057]_ ;
  assign \new_[55059]_  = \new_[55058]_  & \new_[55053]_ ;
  assign \new_[55063]_  = A266 & A265;
  assign \new_[55064]_  = ~A200 & \new_[55063]_ ;
  assign \new_[55067]_  = ~A299 & A298;
  assign \new_[55070]_  = A302 & A300;
  assign \new_[55071]_  = \new_[55070]_  & \new_[55067]_ ;
  assign \new_[55072]_  = \new_[55071]_  & \new_[55064]_ ;
  assign \new_[55076]_  = ~A168 & ~A169;
  assign \new_[55077]_  = A170 & \new_[55076]_ ;
  assign \new_[55081]_  = ~A199 & ~A166;
  assign \new_[55082]_  = A167 & \new_[55081]_ ;
  assign \new_[55083]_  = \new_[55082]_  & \new_[55077]_ ;
  assign \new_[55087]_  = A266 & A265;
  assign \new_[55088]_  = ~A200 & \new_[55087]_ ;
  assign \new_[55091]_  = A299 & ~A298;
  assign \new_[55094]_  = A301 & A300;
  assign \new_[55095]_  = \new_[55094]_  & \new_[55091]_ ;
  assign \new_[55096]_  = \new_[55095]_  & \new_[55088]_ ;
  assign \new_[55100]_  = ~A168 & ~A169;
  assign \new_[55101]_  = A170 & \new_[55100]_ ;
  assign \new_[55105]_  = ~A199 & ~A166;
  assign \new_[55106]_  = A167 & \new_[55105]_ ;
  assign \new_[55107]_  = \new_[55106]_  & \new_[55101]_ ;
  assign \new_[55111]_  = A266 & A265;
  assign \new_[55112]_  = ~A200 & \new_[55111]_ ;
  assign \new_[55115]_  = A299 & ~A298;
  assign \new_[55118]_  = A302 & A300;
  assign \new_[55119]_  = \new_[55118]_  & \new_[55115]_ ;
  assign \new_[55120]_  = \new_[55119]_  & \new_[55112]_ ;
  assign \new_[55124]_  = ~A168 & ~A169;
  assign \new_[55125]_  = A170 & \new_[55124]_ ;
  assign \new_[55129]_  = ~A199 & ~A166;
  assign \new_[55130]_  = A167 & \new_[55129]_ ;
  assign \new_[55131]_  = \new_[55130]_  & \new_[55125]_ ;
  assign \new_[55135]_  = ~A266 & ~A265;
  assign \new_[55136]_  = ~A200 & \new_[55135]_ ;
  assign \new_[55139]_  = ~A299 & A298;
  assign \new_[55142]_  = A301 & A300;
  assign \new_[55143]_  = \new_[55142]_  & \new_[55139]_ ;
  assign \new_[55144]_  = \new_[55143]_  & \new_[55136]_ ;
  assign \new_[55148]_  = ~A168 & ~A169;
  assign \new_[55149]_  = A170 & \new_[55148]_ ;
  assign \new_[55153]_  = ~A199 & ~A166;
  assign \new_[55154]_  = A167 & \new_[55153]_ ;
  assign \new_[55155]_  = \new_[55154]_  & \new_[55149]_ ;
  assign \new_[55159]_  = ~A266 & ~A265;
  assign \new_[55160]_  = ~A200 & \new_[55159]_ ;
  assign \new_[55163]_  = ~A299 & A298;
  assign \new_[55166]_  = A302 & A300;
  assign \new_[55167]_  = \new_[55166]_  & \new_[55163]_ ;
  assign \new_[55168]_  = \new_[55167]_  & \new_[55160]_ ;
  assign \new_[55172]_  = ~A168 & ~A169;
  assign \new_[55173]_  = A170 & \new_[55172]_ ;
  assign \new_[55177]_  = ~A199 & ~A166;
  assign \new_[55178]_  = A167 & \new_[55177]_ ;
  assign \new_[55179]_  = \new_[55178]_  & \new_[55173]_ ;
  assign \new_[55183]_  = ~A266 & ~A265;
  assign \new_[55184]_  = ~A200 & \new_[55183]_ ;
  assign \new_[55187]_  = A299 & ~A298;
  assign \new_[55190]_  = A301 & A300;
  assign \new_[55191]_  = \new_[55190]_  & \new_[55187]_ ;
  assign \new_[55192]_  = \new_[55191]_  & \new_[55184]_ ;
  assign \new_[55196]_  = ~A168 & ~A169;
  assign \new_[55197]_  = A170 & \new_[55196]_ ;
  assign \new_[55201]_  = ~A199 & ~A166;
  assign \new_[55202]_  = A167 & \new_[55201]_ ;
  assign \new_[55203]_  = \new_[55202]_  & \new_[55197]_ ;
  assign \new_[55207]_  = ~A266 & ~A265;
  assign \new_[55208]_  = ~A200 & \new_[55207]_ ;
  assign \new_[55211]_  = A299 & ~A298;
  assign \new_[55214]_  = A302 & A300;
  assign \new_[55215]_  = \new_[55214]_  & \new_[55211]_ ;
  assign \new_[55216]_  = \new_[55215]_  & \new_[55208]_ ;
  assign \new_[55220]_  = ~A168 & ~A169;
  assign \new_[55221]_  = A170 & \new_[55220]_ ;
  assign \new_[55225]_  = ~A201 & A166;
  assign \new_[55226]_  = ~A167 & \new_[55225]_ ;
  assign \new_[55227]_  = \new_[55226]_  & \new_[55221]_ ;
  assign \new_[55231]_  = A268 & ~A267;
  assign \new_[55232]_  = A202 & \new_[55231]_ ;
  assign \new_[55235]_  = ~A299 & A298;
  assign \new_[55238]_  = A301 & A300;
  assign \new_[55239]_  = \new_[55238]_  & \new_[55235]_ ;
  assign \new_[55240]_  = \new_[55239]_  & \new_[55232]_ ;
  assign \new_[55244]_  = ~A168 & ~A169;
  assign \new_[55245]_  = A170 & \new_[55244]_ ;
  assign \new_[55249]_  = ~A201 & A166;
  assign \new_[55250]_  = ~A167 & \new_[55249]_ ;
  assign \new_[55251]_  = \new_[55250]_  & \new_[55245]_ ;
  assign \new_[55255]_  = A268 & ~A267;
  assign \new_[55256]_  = A202 & \new_[55255]_ ;
  assign \new_[55259]_  = ~A299 & A298;
  assign \new_[55262]_  = A302 & A300;
  assign \new_[55263]_  = \new_[55262]_  & \new_[55259]_ ;
  assign \new_[55264]_  = \new_[55263]_  & \new_[55256]_ ;
  assign \new_[55268]_  = ~A168 & ~A169;
  assign \new_[55269]_  = A170 & \new_[55268]_ ;
  assign \new_[55273]_  = ~A201 & A166;
  assign \new_[55274]_  = ~A167 & \new_[55273]_ ;
  assign \new_[55275]_  = \new_[55274]_  & \new_[55269]_ ;
  assign \new_[55279]_  = A268 & ~A267;
  assign \new_[55280]_  = A202 & \new_[55279]_ ;
  assign \new_[55283]_  = A299 & ~A298;
  assign \new_[55286]_  = A301 & A300;
  assign \new_[55287]_  = \new_[55286]_  & \new_[55283]_ ;
  assign \new_[55288]_  = \new_[55287]_  & \new_[55280]_ ;
  assign \new_[55292]_  = ~A168 & ~A169;
  assign \new_[55293]_  = A170 & \new_[55292]_ ;
  assign \new_[55297]_  = ~A201 & A166;
  assign \new_[55298]_  = ~A167 & \new_[55297]_ ;
  assign \new_[55299]_  = \new_[55298]_  & \new_[55293]_ ;
  assign \new_[55303]_  = A268 & ~A267;
  assign \new_[55304]_  = A202 & \new_[55303]_ ;
  assign \new_[55307]_  = A299 & ~A298;
  assign \new_[55310]_  = A302 & A300;
  assign \new_[55311]_  = \new_[55310]_  & \new_[55307]_ ;
  assign \new_[55312]_  = \new_[55311]_  & \new_[55304]_ ;
  assign \new_[55316]_  = ~A168 & ~A169;
  assign \new_[55317]_  = A170 & \new_[55316]_ ;
  assign \new_[55321]_  = ~A201 & A166;
  assign \new_[55322]_  = ~A167 & \new_[55321]_ ;
  assign \new_[55323]_  = \new_[55322]_  & \new_[55317]_ ;
  assign \new_[55327]_  = A269 & ~A267;
  assign \new_[55328]_  = A202 & \new_[55327]_ ;
  assign \new_[55331]_  = ~A299 & A298;
  assign \new_[55334]_  = A301 & A300;
  assign \new_[55335]_  = \new_[55334]_  & \new_[55331]_ ;
  assign \new_[55336]_  = \new_[55335]_  & \new_[55328]_ ;
  assign \new_[55340]_  = ~A168 & ~A169;
  assign \new_[55341]_  = A170 & \new_[55340]_ ;
  assign \new_[55345]_  = ~A201 & A166;
  assign \new_[55346]_  = ~A167 & \new_[55345]_ ;
  assign \new_[55347]_  = \new_[55346]_  & \new_[55341]_ ;
  assign \new_[55351]_  = A269 & ~A267;
  assign \new_[55352]_  = A202 & \new_[55351]_ ;
  assign \new_[55355]_  = ~A299 & A298;
  assign \new_[55358]_  = A302 & A300;
  assign \new_[55359]_  = \new_[55358]_  & \new_[55355]_ ;
  assign \new_[55360]_  = \new_[55359]_  & \new_[55352]_ ;
  assign \new_[55364]_  = ~A168 & ~A169;
  assign \new_[55365]_  = A170 & \new_[55364]_ ;
  assign \new_[55369]_  = ~A201 & A166;
  assign \new_[55370]_  = ~A167 & \new_[55369]_ ;
  assign \new_[55371]_  = \new_[55370]_  & \new_[55365]_ ;
  assign \new_[55375]_  = A269 & ~A267;
  assign \new_[55376]_  = A202 & \new_[55375]_ ;
  assign \new_[55379]_  = A299 & ~A298;
  assign \new_[55382]_  = A301 & A300;
  assign \new_[55383]_  = \new_[55382]_  & \new_[55379]_ ;
  assign \new_[55384]_  = \new_[55383]_  & \new_[55376]_ ;
  assign \new_[55388]_  = ~A168 & ~A169;
  assign \new_[55389]_  = A170 & \new_[55388]_ ;
  assign \new_[55393]_  = ~A201 & A166;
  assign \new_[55394]_  = ~A167 & \new_[55393]_ ;
  assign \new_[55395]_  = \new_[55394]_  & \new_[55389]_ ;
  assign \new_[55399]_  = A269 & ~A267;
  assign \new_[55400]_  = A202 & \new_[55399]_ ;
  assign \new_[55403]_  = A299 & ~A298;
  assign \new_[55406]_  = A302 & A300;
  assign \new_[55407]_  = \new_[55406]_  & \new_[55403]_ ;
  assign \new_[55408]_  = \new_[55407]_  & \new_[55400]_ ;
  assign \new_[55412]_  = ~A168 & ~A169;
  assign \new_[55413]_  = A170 & \new_[55412]_ ;
  assign \new_[55417]_  = ~A201 & A166;
  assign \new_[55418]_  = ~A167 & \new_[55417]_ ;
  assign \new_[55419]_  = \new_[55418]_  & \new_[55413]_ ;
  assign \new_[55423]_  = A266 & A265;
  assign \new_[55424]_  = A202 & \new_[55423]_ ;
  assign \new_[55427]_  = ~A299 & A298;
  assign \new_[55430]_  = A301 & A300;
  assign \new_[55431]_  = \new_[55430]_  & \new_[55427]_ ;
  assign \new_[55432]_  = \new_[55431]_  & \new_[55424]_ ;
  assign \new_[55436]_  = ~A168 & ~A169;
  assign \new_[55437]_  = A170 & \new_[55436]_ ;
  assign \new_[55441]_  = ~A201 & A166;
  assign \new_[55442]_  = ~A167 & \new_[55441]_ ;
  assign \new_[55443]_  = \new_[55442]_  & \new_[55437]_ ;
  assign \new_[55447]_  = A266 & A265;
  assign \new_[55448]_  = A202 & \new_[55447]_ ;
  assign \new_[55451]_  = ~A299 & A298;
  assign \new_[55454]_  = A302 & A300;
  assign \new_[55455]_  = \new_[55454]_  & \new_[55451]_ ;
  assign \new_[55456]_  = \new_[55455]_  & \new_[55448]_ ;
  assign \new_[55460]_  = ~A168 & ~A169;
  assign \new_[55461]_  = A170 & \new_[55460]_ ;
  assign \new_[55465]_  = ~A201 & A166;
  assign \new_[55466]_  = ~A167 & \new_[55465]_ ;
  assign \new_[55467]_  = \new_[55466]_  & \new_[55461]_ ;
  assign \new_[55471]_  = A266 & A265;
  assign \new_[55472]_  = A202 & \new_[55471]_ ;
  assign \new_[55475]_  = A299 & ~A298;
  assign \new_[55478]_  = A301 & A300;
  assign \new_[55479]_  = \new_[55478]_  & \new_[55475]_ ;
  assign \new_[55480]_  = \new_[55479]_  & \new_[55472]_ ;
  assign \new_[55484]_  = ~A168 & ~A169;
  assign \new_[55485]_  = A170 & \new_[55484]_ ;
  assign \new_[55489]_  = ~A201 & A166;
  assign \new_[55490]_  = ~A167 & \new_[55489]_ ;
  assign \new_[55491]_  = \new_[55490]_  & \new_[55485]_ ;
  assign \new_[55495]_  = A266 & A265;
  assign \new_[55496]_  = A202 & \new_[55495]_ ;
  assign \new_[55499]_  = A299 & ~A298;
  assign \new_[55502]_  = A302 & A300;
  assign \new_[55503]_  = \new_[55502]_  & \new_[55499]_ ;
  assign \new_[55504]_  = \new_[55503]_  & \new_[55496]_ ;
  assign \new_[55508]_  = ~A168 & ~A169;
  assign \new_[55509]_  = A170 & \new_[55508]_ ;
  assign \new_[55513]_  = ~A201 & A166;
  assign \new_[55514]_  = ~A167 & \new_[55513]_ ;
  assign \new_[55515]_  = \new_[55514]_  & \new_[55509]_ ;
  assign \new_[55519]_  = ~A266 & ~A265;
  assign \new_[55520]_  = A202 & \new_[55519]_ ;
  assign \new_[55523]_  = ~A299 & A298;
  assign \new_[55526]_  = A301 & A300;
  assign \new_[55527]_  = \new_[55526]_  & \new_[55523]_ ;
  assign \new_[55528]_  = \new_[55527]_  & \new_[55520]_ ;
  assign \new_[55532]_  = ~A168 & ~A169;
  assign \new_[55533]_  = A170 & \new_[55532]_ ;
  assign \new_[55537]_  = ~A201 & A166;
  assign \new_[55538]_  = ~A167 & \new_[55537]_ ;
  assign \new_[55539]_  = \new_[55538]_  & \new_[55533]_ ;
  assign \new_[55543]_  = ~A266 & ~A265;
  assign \new_[55544]_  = A202 & \new_[55543]_ ;
  assign \new_[55547]_  = ~A299 & A298;
  assign \new_[55550]_  = A302 & A300;
  assign \new_[55551]_  = \new_[55550]_  & \new_[55547]_ ;
  assign \new_[55552]_  = \new_[55551]_  & \new_[55544]_ ;
  assign \new_[55556]_  = ~A168 & ~A169;
  assign \new_[55557]_  = A170 & \new_[55556]_ ;
  assign \new_[55561]_  = ~A201 & A166;
  assign \new_[55562]_  = ~A167 & \new_[55561]_ ;
  assign \new_[55563]_  = \new_[55562]_  & \new_[55557]_ ;
  assign \new_[55567]_  = ~A266 & ~A265;
  assign \new_[55568]_  = A202 & \new_[55567]_ ;
  assign \new_[55571]_  = A299 & ~A298;
  assign \new_[55574]_  = A301 & A300;
  assign \new_[55575]_  = \new_[55574]_  & \new_[55571]_ ;
  assign \new_[55576]_  = \new_[55575]_  & \new_[55568]_ ;
  assign \new_[55580]_  = ~A168 & ~A169;
  assign \new_[55581]_  = A170 & \new_[55580]_ ;
  assign \new_[55585]_  = ~A201 & A166;
  assign \new_[55586]_  = ~A167 & \new_[55585]_ ;
  assign \new_[55587]_  = \new_[55586]_  & \new_[55581]_ ;
  assign \new_[55591]_  = ~A266 & ~A265;
  assign \new_[55592]_  = A202 & \new_[55591]_ ;
  assign \new_[55595]_  = A299 & ~A298;
  assign \new_[55598]_  = A302 & A300;
  assign \new_[55599]_  = \new_[55598]_  & \new_[55595]_ ;
  assign \new_[55600]_  = \new_[55599]_  & \new_[55592]_ ;
  assign \new_[55604]_  = ~A168 & ~A169;
  assign \new_[55605]_  = A170 & \new_[55604]_ ;
  assign \new_[55609]_  = ~A201 & A166;
  assign \new_[55610]_  = ~A167 & \new_[55609]_ ;
  assign \new_[55611]_  = \new_[55610]_  & \new_[55605]_ ;
  assign \new_[55615]_  = A268 & ~A267;
  assign \new_[55616]_  = A203 & \new_[55615]_ ;
  assign \new_[55619]_  = ~A299 & A298;
  assign \new_[55622]_  = A301 & A300;
  assign \new_[55623]_  = \new_[55622]_  & \new_[55619]_ ;
  assign \new_[55624]_  = \new_[55623]_  & \new_[55616]_ ;
  assign \new_[55628]_  = ~A168 & ~A169;
  assign \new_[55629]_  = A170 & \new_[55628]_ ;
  assign \new_[55633]_  = ~A201 & A166;
  assign \new_[55634]_  = ~A167 & \new_[55633]_ ;
  assign \new_[55635]_  = \new_[55634]_  & \new_[55629]_ ;
  assign \new_[55639]_  = A268 & ~A267;
  assign \new_[55640]_  = A203 & \new_[55639]_ ;
  assign \new_[55643]_  = ~A299 & A298;
  assign \new_[55646]_  = A302 & A300;
  assign \new_[55647]_  = \new_[55646]_  & \new_[55643]_ ;
  assign \new_[55648]_  = \new_[55647]_  & \new_[55640]_ ;
  assign \new_[55652]_  = ~A168 & ~A169;
  assign \new_[55653]_  = A170 & \new_[55652]_ ;
  assign \new_[55657]_  = ~A201 & A166;
  assign \new_[55658]_  = ~A167 & \new_[55657]_ ;
  assign \new_[55659]_  = \new_[55658]_  & \new_[55653]_ ;
  assign \new_[55663]_  = A268 & ~A267;
  assign \new_[55664]_  = A203 & \new_[55663]_ ;
  assign \new_[55667]_  = A299 & ~A298;
  assign \new_[55670]_  = A301 & A300;
  assign \new_[55671]_  = \new_[55670]_  & \new_[55667]_ ;
  assign \new_[55672]_  = \new_[55671]_  & \new_[55664]_ ;
  assign \new_[55676]_  = ~A168 & ~A169;
  assign \new_[55677]_  = A170 & \new_[55676]_ ;
  assign \new_[55681]_  = ~A201 & A166;
  assign \new_[55682]_  = ~A167 & \new_[55681]_ ;
  assign \new_[55683]_  = \new_[55682]_  & \new_[55677]_ ;
  assign \new_[55687]_  = A268 & ~A267;
  assign \new_[55688]_  = A203 & \new_[55687]_ ;
  assign \new_[55691]_  = A299 & ~A298;
  assign \new_[55694]_  = A302 & A300;
  assign \new_[55695]_  = \new_[55694]_  & \new_[55691]_ ;
  assign \new_[55696]_  = \new_[55695]_  & \new_[55688]_ ;
  assign \new_[55700]_  = ~A168 & ~A169;
  assign \new_[55701]_  = A170 & \new_[55700]_ ;
  assign \new_[55705]_  = ~A201 & A166;
  assign \new_[55706]_  = ~A167 & \new_[55705]_ ;
  assign \new_[55707]_  = \new_[55706]_  & \new_[55701]_ ;
  assign \new_[55711]_  = A269 & ~A267;
  assign \new_[55712]_  = A203 & \new_[55711]_ ;
  assign \new_[55715]_  = ~A299 & A298;
  assign \new_[55718]_  = A301 & A300;
  assign \new_[55719]_  = \new_[55718]_  & \new_[55715]_ ;
  assign \new_[55720]_  = \new_[55719]_  & \new_[55712]_ ;
  assign \new_[55724]_  = ~A168 & ~A169;
  assign \new_[55725]_  = A170 & \new_[55724]_ ;
  assign \new_[55729]_  = ~A201 & A166;
  assign \new_[55730]_  = ~A167 & \new_[55729]_ ;
  assign \new_[55731]_  = \new_[55730]_  & \new_[55725]_ ;
  assign \new_[55735]_  = A269 & ~A267;
  assign \new_[55736]_  = A203 & \new_[55735]_ ;
  assign \new_[55739]_  = ~A299 & A298;
  assign \new_[55742]_  = A302 & A300;
  assign \new_[55743]_  = \new_[55742]_  & \new_[55739]_ ;
  assign \new_[55744]_  = \new_[55743]_  & \new_[55736]_ ;
  assign \new_[55748]_  = ~A168 & ~A169;
  assign \new_[55749]_  = A170 & \new_[55748]_ ;
  assign \new_[55753]_  = ~A201 & A166;
  assign \new_[55754]_  = ~A167 & \new_[55753]_ ;
  assign \new_[55755]_  = \new_[55754]_  & \new_[55749]_ ;
  assign \new_[55759]_  = A269 & ~A267;
  assign \new_[55760]_  = A203 & \new_[55759]_ ;
  assign \new_[55763]_  = A299 & ~A298;
  assign \new_[55766]_  = A301 & A300;
  assign \new_[55767]_  = \new_[55766]_  & \new_[55763]_ ;
  assign \new_[55768]_  = \new_[55767]_  & \new_[55760]_ ;
  assign \new_[55772]_  = ~A168 & ~A169;
  assign \new_[55773]_  = A170 & \new_[55772]_ ;
  assign \new_[55777]_  = ~A201 & A166;
  assign \new_[55778]_  = ~A167 & \new_[55777]_ ;
  assign \new_[55779]_  = \new_[55778]_  & \new_[55773]_ ;
  assign \new_[55783]_  = A269 & ~A267;
  assign \new_[55784]_  = A203 & \new_[55783]_ ;
  assign \new_[55787]_  = A299 & ~A298;
  assign \new_[55790]_  = A302 & A300;
  assign \new_[55791]_  = \new_[55790]_  & \new_[55787]_ ;
  assign \new_[55792]_  = \new_[55791]_  & \new_[55784]_ ;
  assign \new_[55796]_  = ~A168 & ~A169;
  assign \new_[55797]_  = A170 & \new_[55796]_ ;
  assign \new_[55801]_  = ~A201 & A166;
  assign \new_[55802]_  = ~A167 & \new_[55801]_ ;
  assign \new_[55803]_  = \new_[55802]_  & \new_[55797]_ ;
  assign \new_[55807]_  = A266 & A265;
  assign \new_[55808]_  = A203 & \new_[55807]_ ;
  assign \new_[55811]_  = ~A299 & A298;
  assign \new_[55814]_  = A301 & A300;
  assign \new_[55815]_  = \new_[55814]_  & \new_[55811]_ ;
  assign \new_[55816]_  = \new_[55815]_  & \new_[55808]_ ;
  assign \new_[55820]_  = ~A168 & ~A169;
  assign \new_[55821]_  = A170 & \new_[55820]_ ;
  assign \new_[55825]_  = ~A201 & A166;
  assign \new_[55826]_  = ~A167 & \new_[55825]_ ;
  assign \new_[55827]_  = \new_[55826]_  & \new_[55821]_ ;
  assign \new_[55831]_  = A266 & A265;
  assign \new_[55832]_  = A203 & \new_[55831]_ ;
  assign \new_[55835]_  = ~A299 & A298;
  assign \new_[55838]_  = A302 & A300;
  assign \new_[55839]_  = \new_[55838]_  & \new_[55835]_ ;
  assign \new_[55840]_  = \new_[55839]_  & \new_[55832]_ ;
  assign \new_[55844]_  = ~A168 & ~A169;
  assign \new_[55845]_  = A170 & \new_[55844]_ ;
  assign \new_[55849]_  = ~A201 & A166;
  assign \new_[55850]_  = ~A167 & \new_[55849]_ ;
  assign \new_[55851]_  = \new_[55850]_  & \new_[55845]_ ;
  assign \new_[55855]_  = A266 & A265;
  assign \new_[55856]_  = A203 & \new_[55855]_ ;
  assign \new_[55859]_  = A299 & ~A298;
  assign \new_[55862]_  = A301 & A300;
  assign \new_[55863]_  = \new_[55862]_  & \new_[55859]_ ;
  assign \new_[55864]_  = \new_[55863]_  & \new_[55856]_ ;
  assign \new_[55868]_  = ~A168 & ~A169;
  assign \new_[55869]_  = A170 & \new_[55868]_ ;
  assign \new_[55873]_  = ~A201 & A166;
  assign \new_[55874]_  = ~A167 & \new_[55873]_ ;
  assign \new_[55875]_  = \new_[55874]_  & \new_[55869]_ ;
  assign \new_[55879]_  = A266 & A265;
  assign \new_[55880]_  = A203 & \new_[55879]_ ;
  assign \new_[55883]_  = A299 & ~A298;
  assign \new_[55886]_  = A302 & A300;
  assign \new_[55887]_  = \new_[55886]_  & \new_[55883]_ ;
  assign \new_[55888]_  = \new_[55887]_  & \new_[55880]_ ;
  assign \new_[55892]_  = ~A168 & ~A169;
  assign \new_[55893]_  = A170 & \new_[55892]_ ;
  assign \new_[55897]_  = ~A201 & A166;
  assign \new_[55898]_  = ~A167 & \new_[55897]_ ;
  assign \new_[55899]_  = \new_[55898]_  & \new_[55893]_ ;
  assign \new_[55903]_  = ~A266 & ~A265;
  assign \new_[55904]_  = A203 & \new_[55903]_ ;
  assign \new_[55907]_  = ~A299 & A298;
  assign \new_[55910]_  = A301 & A300;
  assign \new_[55911]_  = \new_[55910]_  & \new_[55907]_ ;
  assign \new_[55912]_  = \new_[55911]_  & \new_[55904]_ ;
  assign \new_[55916]_  = ~A168 & ~A169;
  assign \new_[55917]_  = A170 & \new_[55916]_ ;
  assign \new_[55921]_  = ~A201 & A166;
  assign \new_[55922]_  = ~A167 & \new_[55921]_ ;
  assign \new_[55923]_  = \new_[55922]_  & \new_[55917]_ ;
  assign \new_[55927]_  = ~A266 & ~A265;
  assign \new_[55928]_  = A203 & \new_[55927]_ ;
  assign \new_[55931]_  = ~A299 & A298;
  assign \new_[55934]_  = A302 & A300;
  assign \new_[55935]_  = \new_[55934]_  & \new_[55931]_ ;
  assign \new_[55936]_  = \new_[55935]_  & \new_[55928]_ ;
  assign \new_[55940]_  = ~A168 & ~A169;
  assign \new_[55941]_  = A170 & \new_[55940]_ ;
  assign \new_[55945]_  = ~A201 & A166;
  assign \new_[55946]_  = ~A167 & \new_[55945]_ ;
  assign \new_[55947]_  = \new_[55946]_  & \new_[55941]_ ;
  assign \new_[55951]_  = ~A266 & ~A265;
  assign \new_[55952]_  = A203 & \new_[55951]_ ;
  assign \new_[55955]_  = A299 & ~A298;
  assign \new_[55958]_  = A301 & A300;
  assign \new_[55959]_  = \new_[55958]_  & \new_[55955]_ ;
  assign \new_[55960]_  = \new_[55959]_  & \new_[55952]_ ;
  assign \new_[55964]_  = ~A168 & ~A169;
  assign \new_[55965]_  = A170 & \new_[55964]_ ;
  assign \new_[55969]_  = ~A201 & A166;
  assign \new_[55970]_  = ~A167 & \new_[55969]_ ;
  assign \new_[55971]_  = \new_[55970]_  & \new_[55965]_ ;
  assign \new_[55975]_  = ~A266 & ~A265;
  assign \new_[55976]_  = A203 & \new_[55975]_ ;
  assign \new_[55979]_  = A299 & ~A298;
  assign \new_[55982]_  = A302 & A300;
  assign \new_[55983]_  = \new_[55982]_  & \new_[55979]_ ;
  assign \new_[55984]_  = \new_[55983]_  & \new_[55976]_ ;
  assign \new_[55988]_  = ~A168 & ~A169;
  assign \new_[55989]_  = A170 & \new_[55988]_ ;
  assign \new_[55993]_  = A199 & A166;
  assign \new_[55994]_  = ~A167 & \new_[55993]_ ;
  assign \new_[55995]_  = \new_[55994]_  & \new_[55989]_ ;
  assign \new_[55999]_  = A268 & ~A267;
  assign \new_[56000]_  = A200 & \new_[55999]_ ;
  assign \new_[56003]_  = ~A299 & A298;
  assign \new_[56006]_  = A301 & A300;
  assign \new_[56007]_  = \new_[56006]_  & \new_[56003]_ ;
  assign \new_[56008]_  = \new_[56007]_  & \new_[56000]_ ;
  assign \new_[56012]_  = ~A168 & ~A169;
  assign \new_[56013]_  = A170 & \new_[56012]_ ;
  assign \new_[56017]_  = A199 & A166;
  assign \new_[56018]_  = ~A167 & \new_[56017]_ ;
  assign \new_[56019]_  = \new_[56018]_  & \new_[56013]_ ;
  assign \new_[56023]_  = A268 & ~A267;
  assign \new_[56024]_  = A200 & \new_[56023]_ ;
  assign \new_[56027]_  = ~A299 & A298;
  assign \new_[56030]_  = A302 & A300;
  assign \new_[56031]_  = \new_[56030]_  & \new_[56027]_ ;
  assign \new_[56032]_  = \new_[56031]_  & \new_[56024]_ ;
  assign \new_[56036]_  = ~A168 & ~A169;
  assign \new_[56037]_  = A170 & \new_[56036]_ ;
  assign \new_[56041]_  = A199 & A166;
  assign \new_[56042]_  = ~A167 & \new_[56041]_ ;
  assign \new_[56043]_  = \new_[56042]_  & \new_[56037]_ ;
  assign \new_[56047]_  = A268 & ~A267;
  assign \new_[56048]_  = A200 & \new_[56047]_ ;
  assign \new_[56051]_  = A299 & ~A298;
  assign \new_[56054]_  = A301 & A300;
  assign \new_[56055]_  = \new_[56054]_  & \new_[56051]_ ;
  assign \new_[56056]_  = \new_[56055]_  & \new_[56048]_ ;
  assign \new_[56060]_  = ~A168 & ~A169;
  assign \new_[56061]_  = A170 & \new_[56060]_ ;
  assign \new_[56065]_  = A199 & A166;
  assign \new_[56066]_  = ~A167 & \new_[56065]_ ;
  assign \new_[56067]_  = \new_[56066]_  & \new_[56061]_ ;
  assign \new_[56071]_  = A268 & ~A267;
  assign \new_[56072]_  = A200 & \new_[56071]_ ;
  assign \new_[56075]_  = A299 & ~A298;
  assign \new_[56078]_  = A302 & A300;
  assign \new_[56079]_  = \new_[56078]_  & \new_[56075]_ ;
  assign \new_[56080]_  = \new_[56079]_  & \new_[56072]_ ;
  assign \new_[56084]_  = ~A168 & ~A169;
  assign \new_[56085]_  = A170 & \new_[56084]_ ;
  assign \new_[56089]_  = A199 & A166;
  assign \new_[56090]_  = ~A167 & \new_[56089]_ ;
  assign \new_[56091]_  = \new_[56090]_  & \new_[56085]_ ;
  assign \new_[56095]_  = A269 & ~A267;
  assign \new_[56096]_  = A200 & \new_[56095]_ ;
  assign \new_[56099]_  = ~A299 & A298;
  assign \new_[56102]_  = A301 & A300;
  assign \new_[56103]_  = \new_[56102]_  & \new_[56099]_ ;
  assign \new_[56104]_  = \new_[56103]_  & \new_[56096]_ ;
  assign \new_[56108]_  = ~A168 & ~A169;
  assign \new_[56109]_  = A170 & \new_[56108]_ ;
  assign \new_[56113]_  = A199 & A166;
  assign \new_[56114]_  = ~A167 & \new_[56113]_ ;
  assign \new_[56115]_  = \new_[56114]_  & \new_[56109]_ ;
  assign \new_[56119]_  = A269 & ~A267;
  assign \new_[56120]_  = A200 & \new_[56119]_ ;
  assign \new_[56123]_  = ~A299 & A298;
  assign \new_[56126]_  = A302 & A300;
  assign \new_[56127]_  = \new_[56126]_  & \new_[56123]_ ;
  assign \new_[56128]_  = \new_[56127]_  & \new_[56120]_ ;
  assign \new_[56132]_  = ~A168 & ~A169;
  assign \new_[56133]_  = A170 & \new_[56132]_ ;
  assign \new_[56137]_  = A199 & A166;
  assign \new_[56138]_  = ~A167 & \new_[56137]_ ;
  assign \new_[56139]_  = \new_[56138]_  & \new_[56133]_ ;
  assign \new_[56143]_  = A269 & ~A267;
  assign \new_[56144]_  = A200 & \new_[56143]_ ;
  assign \new_[56147]_  = A299 & ~A298;
  assign \new_[56150]_  = A301 & A300;
  assign \new_[56151]_  = \new_[56150]_  & \new_[56147]_ ;
  assign \new_[56152]_  = \new_[56151]_  & \new_[56144]_ ;
  assign \new_[56156]_  = ~A168 & ~A169;
  assign \new_[56157]_  = A170 & \new_[56156]_ ;
  assign \new_[56161]_  = A199 & A166;
  assign \new_[56162]_  = ~A167 & \new_[56161]_ ;
  assign \new_[56163]_  = \new_[56162]_  & \new_[56157]_ ;
  assign \new_[56167]_  = A269 & ~A267;
  assign \new_[56168]_  = A200 & \new_[56167]_ ;
  assign \new_[56171]_  = A299 & ~A298;
  assign \new_[56174]_  = A302 & A300;
  assign \new_[56175]_  = \new_[56174]_  & \new_[56171]_ ;
  assign \new_[56176]_  = \new_[56175]_  & \new_[56168]_ ;
  assign \new_[56180]_  = ~A168 & ~A169;
  assign \new_[56181]_  = A170 & \new_[56180]_ ;
  assign \new_[56185]_  = A199 & A166;
  assign \new_[56186]_  = ~A167 & \new_[56185]_ ;
  assign \new_[56187]_  = \new_[56186]_  & \new_[56181]_ ;
  assign \new_[56191]_  = A266 & A265;
  assign \new_[56192]_  = A200 & \new_[56191]_ ;
  assign \new_[56195]_  = ~A299 & A298;
  assign \new_[56198]_  = A301 & A300;
  assign \new_[56199]_  = \new_[56198]_  & \new_[56195]_ ;
  assign \new_[56200]_  = \new_[56199]_  & \new_[56192]_ ;
  assign \new_[56204]_  = ~A168 & ~A169;
  assign \new_[56205]_  = A170 & \new_[56204]_ ;
  assign \new_[56209]_  = A199 & A166;
  assign \new_[56210]_  = ~A167 & \new_[56209]_ ;
  assign \new_[56211]_  = \new_[56210]_  & \new_[56205]_ ;
  assign \new_[56215]_  = A266 & A265;
  assign \new_[56216]_  = A200 & \new_[56215]_ ;
  assign \new_[56219]_  = ~A299 & A298;
  assign \new_[56222]_  = A302 & A300;
  assign \new_[56223]_  = \new_[56222]_  & \new_[56219]_ ;
  assign \new_[56224]_  = \new_[56223]_  & \new_[56216]_ ;
  assign \new_[56228]_  = ~A168 & ~A169;
  assign \new_[56229]_  = A170 & \new_[56228]_ ;
  assign \new_[56233]_  = A199 & A166;
  assign \new_[56234]_  = ~A167 & \new_[56233]_ ;
  assign \new_[56235]_  = \new_[56234]_  & \new_[56229]_ ;
  assign \new_[56239]_  = A266 & A265;
  assign \new_[56240]_  = A200 & \new_[56239]_ ;
  assign \new_[56243]_  = A299 & ~A298;
  assign \new_[56246]_  = A301 & A300;
  assign \new_[56247]_  = \new_[56246]_  & \new_[56243]_ ;
  assign \new_[56248]_  = \new_[56247]_  & \new_[56240]_ ;
  assign \new_[56252]_  = ~A168 & ~A169;
  assign \new_[56253]_  = A170 & \new_[56252]_ ;
  assign \new_[56257]_  = A199 & A166;
  assign \new_[56258]_  = ~A167 & \new_[56257]_ ;
  assign \new_[56259]_  = \new_[56258]_  & \new_[56253]_ ;
  assign \new_[56263]_  = A266 & A265;
  assign \new_[56264]_  = A200 & \new_[56263]_ ;
  assign \new_[56267]_  = A299 & ~A298;
  assign \new_[56270]_  = A302 & A300;
  assign \new_[56271]_  = \new_[56270]_  & \new_[56267]_ ;
  assign \new_[56272]_  = \new_[56271]_  & \new_[56264]_ ;
  assign \new_[56276]_  = ~A168 & ~A169;
  assign \new_[56277]_  = A170 & \new_[56276]_ ;
  assign \new_[56281]_  = A199 & A166;
  assign \new_[56282]_  = ~A167 & \new_[56281]_ ;
  assign \new_[56283]_  = \new_[56282]_  & \new_[56277]_ ;
  assign \new_[56287]_  = ~A266 & ~A265;
  assign \new_[56288]_  = A200 & \new_[56287]_ ;
  assign \new_[56291]_  = ~A299 & A298;
  assign \new_[56294]_  = A301 & A300;
  assign \new_[56295]_  = \new_[56294]_  & \new_[56291]_ ;
  assign \new_[56296]_  = \new_[56295]_  & \new_[56288]_ ;
  assign \new_[56300]_  = ~A168 & ~A169;
  assign \new_[56301]_  = A170 & \new_[56300]_ ;
  assign \new_[56305]_  = A199 & A166;
  assign \new_[56306]_  = ~A167 & \new_[56305]_ ;
  assign \new_[56307]_  = \new_[56306]_  & \new_[56301]_ ;
  assign \new_[56311]_  = ~A266 & ~A265;
  assign \new_[56312]_  = A200 & \new_[56311]_ ;
  assign \new_[56315]_  = ~A299 & A298;
  assign \new_[56318]_  = A302 & A300;
  assign \new_[56319]_  = \new_[56318]_  & \new_[56315]_ ;
  assign \new_[56320]_  = \new_[56319]_  & \new_[56312]_ ;
  assign \new_[56324]_  = ~A168 & ~A169;
  assign \new_[56325]_  = A170 & \new_[56324]_ ;
  assign \new_[56329]_  = A199 & A166;
  assign \new_[56330]_  = ~A167 & \new_[56329]_ ;
  assign \new_[56331]_  = \new_[56330]_  & \new_[56325]_ ;
  assign \new_[56335]_  = ~A266 & ~A265;
  assign \new_[56336]_  = A200 & \new_[56335]_ ;
  assign \new_[56339]_  = A299 & ~A298;
  assign \new_[56342]_  = A301 & A300;
  assign \new_[56343]_  = \new_[56342]_  & \new_[56339]_ ;
  assign \new_[56344]_  = \new_[56343]_  & \new_[56336]_ ;
  assign \new_[56348]_  = ~A168 & ~A169;
  assign \new_[56349]_  = A170 & \new_[56348]_ ;
  assign \new_[56353]_  = A199 & A166;
  assign \new_[56354]_  = ~A167 & \new_[56353]_ ;
  assign \new_[56355]_  = \new_[56354]_  & \new_[56349]_ ;
  assign \new_[56359]_  = ~A266 & ~A265;
  assign \new_[56360]_  = A200 & \new_[56359]_ ;
  assign \new_[56363]_  = A299 & ~A298;
  assign \new_[56366]_  = A302 & A300;
  assign \new_[56367]_  = \new_[56366]_  & \new_[56363]_ ;
  assign \new_[56368]_  = \new_[56367]_  & \new_[56360]_ ;
  assign \new_[56372]_  = ~A168 & ~A169;
  assign \new_[56373]_  = A170 & \new_[56372]_ ;
  assign \new_[56377]_  = ~A199 & A166;
  assign \new_[56378]_  = ~A167 & \new_[56377]_ ;
  assign \new_[56379]_  = \new_[56378]_  & \new_[56373]_ ;
  assign \new_[56383]_  = A268 & ~A267;
  assign \new_[56384]_  = ~A200 & \new_[56383]_ ;
  assign \new_[56387]_  = ~A299 & A298;
  assign \new_[56390]_  = A301 & A300;
  assign \new_[56391]_  = \new_[56390]_  & \new_[56387]_ ;
  assign \new_[56392]_  = \new_[56391]_  & \new_[56384]_ ;
  assign \new_[56396]_  = ~A168 & ~A169;
  assign \new_[56397]_  = A170 & \new_[56396]_ ;
  assign \new_[56401]_  = ~A199 & A166;
  assign \new_[56402]_  = ~A167 & \new_[56401]_ ;
  assign \new_[56403]_  = \new_[56402]_  & \new_[56397]_ ;
  assign \new_[56407]_  = A268 & ~A267;
  assign \new_[56408]_  = ~A200 & \new_[56407]_ ;
  assign \new_[56411]_  = ~A299 & A298;
  assign \new_[56414]_  = A302 & A300;
  assign \new_[56415]_  = \new_[56414]_  & \new_[56411]_ ;
  assign \new_[56416]_  = \new_[56415]_  & \new_[56408]_ ;
  assign \new_[56420]_  = ~A168 & ~A169;
  assign \new_[56421]_  = A170 & \new_[56420]_ ;
  assign \new_[56425]_  = ~A199 & A166;
  assign \new_[56426]_  = ~A167 & \new_[56425]_ ;
  assign \new_[56427]_  = \new_[56426]_  & \new_[56421]_ ;
  assign \new_[56431]_  = A268 & ~A267;
  assign \new_[56432]_  = ~A200 & \new_[56431]_ ;
  assign \new_[56435]_  = A299 & ~A298;
  assign \new_[56438]_  = A301 & A300;
  assign \new_[56439]_  = \new_[56438]_  & \new_[56435]_ ;
  assign \new_[56440]_  = \new_[56439]_  & \new_[56432]_ ;
  assign \new_[56444]_  = ~A168 & ~A169;
  assign \new_[56445]_  = A170 & \new_[56444]_ ;
  assign \new_[56449]_  = ~A199 & A166;
  assign \new_[56450]_  = ~A167 & \new_[56449]_ ;
  assign \new_[56451]_  = \new_[56450]_  & \new_[56445]_ ;
  assign \new_[56455]_  = A268 & ~A267;
  assign \new_[56456]_  = ~A200 & \new_[56455]_ ;
  assign \new_[56459]_  = A299 & ~A298;
  assign \new_[56462]_  = A302 & A300;
  assign \new_[56463]_  = \new_[56462]_  & \new_[56459]_ ;
  assign \new_[56464]_  = \new_[56463]_  & \new_[56456]_ ;
  assign \new_[56468]_  = ~A168 & ~A169;
  assign \new_[56469]_  = A170 & \new_[56468]_ ;
  assign \new_[56473]_  = ~A199 & A166;
  assign \new_[56474]_  = ~A167 & \new_[56473]_ ;
  assign \new_[56475]_  = \new_[56474]_  & \new_[56469]_ ;
  assign \new_[56479]_  = A269 & ~A267;
  assign \new_[56480]_  = ~A200 & \new_[56479]_ ;
  assign \new_[56483]_  = ~A299 & A298;
  assign \new_[56486]_  = A301 & A300;
  assign \new_[56487]_  = \new_[56486]_  & \new_[56483]_ ;
  assign \new_[56488]_  = \new_[56487]_  & \new_[56480]_ ;
  assign \new_[56492]_  = ~A168 & ~A169;
  assign \new_[56493]_  = A170 & \new_[56492]_ ;
  assign \new_[56497]_  = ~A199 & A166;
  assign \new_[56498]_  = ~A167 & \new_[56497]_ ;
  assign \new_[56499]_  = \new_[56498]_  & \new_[56493]_ ;
  assign \new_[56503]_  = A269 & ~A267;
  assign \new_[56504]_  = ~A200 & \new_[56503]_ ;
  assign \new_[56507]_  = ~A299 & A298;
  assign \new_[56510]_  = A302 & A300;
  assign \new_[56511]_  = \new_[56510]_  & \new_[56507]_ ;
  assign \new_[56512]_  = \new_[56511]_  & \new_[56504]_ ;
  assign \new_[56516]_  = ~A168 & ~A169;
  assign \new_[56517]_  = A170 & \new_[56516]_ ;
  assign \new_[56521]_  = ~A199 & A166;
  assign \new_[56522]_  = ~A167 & \new_[56521]_ ;
  assign \new_[56523]_  = \new_[56522]_  & \new_[56517]_ ;
  assign \new_[56527]_  = A269 & ~A267;
  assign \new_[56528]_  = ~A200 & \new_[56527]_ ;
  assign \new_[56531]_  = A299 & ~A298;
  assign \new_[56534]_  = A301 & A300;
  assign \new_[56535]_  = \new_[56534]_  & \new_[56531]_ ;
  assign \new_[56536]_  = \new_[56535]_  & \new_[56528]_ ;
  assign \new_[56540]_  = ~A168 & ~A169;
  assign \new_[56541]_  = A170 & \new_[56540]_ ;
  assign \new_[56545]_  = ~A199 & A166;
  assign \new_[56546]_  = ~A167 & \new_[56545]_ ;
  assign \new_[56547]_  = \new_[56546]_  & \new_[56541]_ ;
  assign \new_[56551]_  = A269 & ~A267;
  assign \new_[56552]_  = ~A200 & \new_[56551]_ ;
  assign \new_[56555]_  = A299 & ~A298;
  assign \new_[56558]_  = A302 & A300;
  assign \new_[56559]_  = \new_[56558]_  & \new_[56555]_ ;
  assign \new_[56560]_  = \new_[56559]_  & \new_[56552]_ ;
  assign \new_[56564]_  = ~A168 & ~A169;
  assign \new_[56565]_  = A170 & \new_[56564]_ ;
  assign \new_[56569]_  = ~A199 & A166;
  assign \new_[56570]_  = ~A167 & \new_[56569]_ ;
  assign \new_[56571]_  = \new_[56570]_  & \new_[56565]_ ;
  assign \new_[56575]_  = A266 & A265;
  assign \new_[56576]_  = ~A200 & \new_[56575]_ ;
  assign \new_[56579]_  = ~A299 & A298;
  assign \new_[56582]_  = A301 & A300;
  assign \new_[56583]_  = \new_[56582]_  & \new_[56579]_ ;
  assign \new_[56584]_  = \new_[56583]_  & \new_[56576]_ ;
  assign \new_[56588]_  = ~A168 & ~A169;
  assign \new_[56589]_  = A170 & \new_[56588]_ ;
  assign \new_[56593]_  = ~A199 & A166;
  assign \new_[56594]_  = ~A167 & \new_[56593]_ ;
  assign \new_[56595]_  = \new_[56594]_  & \new_[56589]_ ;
  assign \new_[56599]_  = A266 & A265;
  assign \new_[56600]_  = ~A200 & \new_[56599]_ ;
  assign \new_[56603]_  = ~A299 & A298;
  assign \new_[56606]_  = A302 & A300;
  assign \new_[56607]_  = \new_[56606]_  & \new_[56603]_ ;
  assign \new_[56608]_  = \new_[56607]_  & \new_[56600]_ ;
  assign \new_[56612]_  = ~A168 & ~A169;
  assign \new_[56613]_  = A170 & \new_[56612]_ ;
  assign \new_[56617]_  = ~A199 & A166;
  assign \new_[56618]_  = ~A167 & \new_[56617]_ ;
  assign \new_[56619]_  = \new_[56618]_  & \new_[56613]_ ;
  assign \new_[56623]_  = A266 & A265;
  assign \new_[56624]_  = ~A200 & \new_[56623]_ ;
  assign \new_[56627]_  = A299 & ~A298;
  assign \new_[56630]_  = A301 & A300;
  assign \new_[56631]_  = \new_[56630]_  & \new_[56627]_ ;
  assign \new_[56632]_  = \new_[56631]_  & \new_[56624]_ ;
  assign \new_[56636]_  = ~A168 & ~A169;
  assign \new_[56637]_  = A170 & \new_[56636]_ ;
  assign \new_[56641]_  = ~A199 & A166;
  assign \new_[56642]_  = ~A167 & \new_[56641]_ ;
  assign \new_[56643]_  = \new_[56642]_  & \new_[56637]_ ;
  assign \new_[56647]_  = A266 & A265;
  assign \new_[56648]_  = ~A200 & \new_[56647]_ ;
  assign \new_[56651]_  = A299 & ~A298;
  assign \new_[56654]_  = A302 & A300;
  assign \new_[56655]_  = \new_[56654]_  & \new_[56651]_ ;
  assign \new_[56656]_  = \new_[56655]_  & \new_[56648]_ ;
  assign \new_[56660]_  = ~A168 & ~A169;
  assign \new_[56661]_  = A170 & \new_[56660]_ ;
  assign \new_[56665]_  = ~A199 & A166;
  assign \new_[56666]_  = ~A167 & \new_[56665]_ ;
  assign \new_[56667]_  = \new_[56666]_  & \new_[56661]_ ;
  assign \new_[56671]_  = ~A266 & ~A265;
  assign \new_[56672]_  = ~A200 & \new_[56671]_ ;
  assign \new_[56675]_  = ~A299 & A298;
  assign \new_[56678]_  = A301 & A300;
  assign \new_[56679]_  = \new_[56678]_  & \new_[56675]_ ;
  assign \new_[56680]_  = \new_[56679]_  & \new_[56672]_ ;
  assign \new_[56684]_  = ~A168 & ~A169;
  assign \new_[56685]_  = A170 & \new_[56684]_ ;
  assign \new_[56689]_  = ~A199 & A166;
  assign \new_[56690]_  = ~A167 & \new_[56689]_ ;
  assign \new_[56691]_  = \new_[56690]_  & \new_[56685]_ ;
  assign \new_[56695]_  = ~A266 & ~A265;
  assign \new_[56696]_  = ~A200 & \new_[56695]_ ;
  assign \new_[56699]_  = ~A299 & A298;
  assign \new_[56702]_  = A302 & A300;
  assign \new_[56703]_  = \new_[56702]_  & \new_[56699]_ ;
  assign \new_[56704]_  = \new_[56703]_  & \new_[56696]_ ;
  assign \new_[56708]_  = ~A168 & ~A169;
  assign \new_[56709]_  = A170 & \new_[56708]_ ;
  assign \new_[56713]_  = ~A199 & A166;
  assign \new_[56714]_  = ~A167 & \new_[56713]_ ;
  assign \new_[56715]_  = \new_[56714]_  & \new_[56709]_ ;
  assign \new_[56719]_  = ~A266 & ~A265;
  assign \new_[56720]_  = ~A200 & \new_[56719]_ ;
  assign \new_[56723]_  = A299 & ~A298;
  assign \new_[56726]_  = A301 & A300;
  assign \new_[56727]_  = \new_[56726]_  & \new_[56723]_ ;
  assign \new_[56728]_  = \new_[56727]_  & \new_[56720]_ ;
  assign \new_[56732]_  = ~A168 & ~A169;
  assign \new_[56733]_  = A170 & \new_[56732]_ ;
  assign \new_[56737]_  = ~A199 & A166;
  assign \new_[56738]_  = ~A167 & \new_[56737]_ ;
  assign \new_[56739]_  = \new_[56738]_  & \new_[56733]_ ;
  assign \new_[56743]_  = ~A266 & ~A265;
  assign \new_[56744]_  = ~A200 & \new_[56743]_ ;
  assign \new_[56747]_  = A299 & ~A298;
  assign \new_[56750]_  = A302 & A300;
  assign \new_[56751]_  = \new_[56750]_  & \new_[56747]_ ;
  assign \new_[56752]_  = \new_[56751]_  & \new_[56744]_ ;
  assign \new_[56756]_  = ~A199 & A166;
  assign \new_[56757]_  = A167 & \new_[56756]_ ;
  assign \new_[56760]_  = A201 & A200;
  assign \new_[56763]_  = A267 & A202;
  assign \new_[56764]_  = \new_[56763]_  & \new_[56760]_ ;
  assign \new_[56765]_  = \new_[56764]_  & \new_[56757]_ ;
  assign \new_[56769]_  = A298 & ~A269;
  assign \new_[56770]_  = ~A268 & \new_[56769]_ ;
  assign \new_[56773]_  = ~A300 & ~A299;
  assign \new_[56776]_  = ~A302 & ~A301;
  assign \new_[56777]_  = \new_[56776]_  & \new_[56773]_ ;
  assign \new_[56778]_  = \new_[56777]_  & \new_[56770]_ ;
  assign \new_[56782]_  = ~A199 & A166;
  assign \new_[56783]_  = A167 & \new_[56782]_ ;
  assign \new_[56786]_  = A201 & A200;
  assign \new_[56789]_  = A267 & A202;
  assign \new_[56790]_  = \new_[56789]_  & \new_[56786]_ ;
  assign \new_[56791]_  = \new_[56790]_  & \new_[56783]_ ;
  assign \new_[56795]_  = ~A298 & ~A269;
  assign \new_[56796]_  = ~A268 & \new_[56795]_ ;
  assign \new_[56799]_  = ~A300 & A299;
  assign \new_[56802]_  = ~A302 & ~A301;
  assign \new_[56803]_  = \new_[56802]_  & \new_[56799]_ ;
  assign \new_[56804]_  = \new_[56803]_  & \new_[56796]_ ;
  assign \new_[56808]_  = ~A199 & A166;
  assign \new_[56809]_  = A167 & \new_[56808]_ ;
  assign \new_[56812]_  = A201 & A200;
  assign \new_[56815]_  = A267 & A203;
  assign \new_[56816]_  = \new_[56815]_  & \new_[56812]_ ;
  assign \new_[56817]_  = \new_[56816]_  & \new_[56809]_ ;
  assign \new_[56821]_  = A298 & ~A269;
  assign \new_[56822]_  = ~A268 & \new_[56821]_ ;
  assign \new_[56825]_  = ~A300 & ~A299;
  assign \new_[56828]_  = ~A302 & ~A301;
  assign \new_[56829]_  = \new_[56828]_  & \new_[56825]_ ;
  assign \new_[56830]_  = \new_[56829]_  & \new_[56822]_ ;
  assign \new_[56834]_  = ~A199 & A166;
  assign \new_[56835]_  = A167 & \new_[56834]_ ;
  assign \new_[56838]_  = A201 & A200;
  assign \new_[56841]_  = A267 & A203;
  assign \new_[56842]_  = \new_[56841]_  & \new_[56838]_ ;
  assign \new_[56843]_  = \new_[56842]_  & \new_[56835]_ ;
  assign \new_[56847]_  = ~A298 & ~A269;
  assign \new_[56848]_  = ~A268 & \new_[56847]_ ;
  assign \new_[56851]_  = ~A300 & A299;
  assign \new_[56854]_  = ~A302 & ~A301;
  assign \new_[56855]_  = \new_[56854]_  & \new_[56851]_ ;
  assign \new_[56856]_  = \new_[56855]_  & \new_[56848]_ ;
  assign \new_[56860]_  = ~A199 & A166;
  assign \new_[56861]_  = A167 & \new_[56860]_ ;
  assign \new_[56864]_  = ~A201 & A200;
  assign \new_[56867]_  = ~A203 & ~A202;
  assign \new_[56868]_  = \new_[56867]_  & \new_[56864]_ ;
  assign \new_[56869]_  = \new_[56868]_  & \new_[56861]_ ;
  assign \new_[56873]_  = ~A269 & ~A268;
  assign \new_[56874]_  = A267 & \new_[56873]_ ;
  assign \new_[56877]_  = ~A299 & A298;
  assign \new_[56880]_  = A301 & A300;
  assign \new_[56881]_  = \new_[56880]_  & \new_[56877]_ ;
  assign \new_[56882]_  = \new_[56881]_  & \new_[56874]_ ;
  assign \new_[56886]_  = ~A199 & A166;
  assign \new_[56887]_  = A167 & \new_[56886]_ ;
  assign \new_[56890]_  = ~A201 & A200;
  assign \new_[56893]_  = ~A203 & ~A202;
  assign \new_[56894]_  = \new_[56893]_  & \new_[56890]_ ;
  assign \new_[56895]_  = \new_[56894]_  & \new_[56887]_ ;
  assign \new_[56899]_  = ~A269 & ~A268;
  assign \new_[56900]_  = A267 & \new_[56899]_ ;
  assign \new_[56903]_  = ~A299 & A298;
  assign \new_[56906]_  = A302 & A300;
  assign \new_[56907]_  = \new_[56906]_  & \new_[56903]_ ;
  assign \new_[56908]_  = \new_[56907]_  & \new_[56900]_ ;
  assign \new_[56912]_  = ~A199 & A166;
  assign \new_[56913]_  = A167 & \new_[56912]_ ;
  assign \new_[56916]_  = ~A201 & A200;
  assign \new_[56919]_  = ~A203 & ~A202;
  assign \new_[56920]_  = \new_[56919]_  & \new_[56916]_ ;
  assign \new_[56921]_  = \new_[56920]_  & \new_[56913]_ ;
  assign \new_[56925]_  = ~A269 & ~A268;
  assign \new_[56926]_  = A267 & \new_[56925]_ ;
  assign \new_[56929]_  = A299 & ~A298;
  assign \new_[56932]_  = A301 & A300;
  assign \new_[56933]_  = \new_[56932]_  & \new_[56929]_ ;
  assign \new_[56934]_  = \new_[56933]_  & \new_[56926]_ ;
  assign \new_[56938]_  = ~A199 & A166;
  assign \new_[56939]_  = A167 & \new_[56938]_ ;
  assign \new_[56942]_  = ~A201 & A200;
  assign \new_[56945]_  = ~A203 & ~A202;
  assign \new_[56946]_  = \new_[56945]_  & \new_[56942]_ ;
  assign \new_[56947]_  = \new_[56946]_  & \new_[56939]_ ;
  assign \new_[56951]_  = ~A269 & ~A268;
  assign \new_[56952]_  = A267 & \new_[56951]_ ;
  assign \new_[56955]_  = A299 & ~A298;
  assign \new_[56958]_  = A302 & A300;
  assign \new_[56959]_  = \new_[56958]_  & \new_[56955]_ ;
  assign \new_[56960]_  = \new_[56959]_  & \new_[56952]_ ;
  assign \new_[56964]_  = ~A199 & A166;
  assign \new_[56965]_  = A167 & \new_[56964]_ ;
  assign \new_[56968]_  = ~A201 & A200;
  assign \new_[56971]_  = ~A203 & ~A202;
  assign \new_[56972]_  = \new_[56971]_  & \new_[56968]_ ;
  assign \new_[56973]_  = \new_[56972]_  & \new_[56965]_ ;
  assign \new_[56977]_  = A298 & A268;
  assign \new_[56978]_  = ~A267 & \new_[56977]_ ;
  assign \new_[56981]_  = ~A300 & ~A299;
  assign \new_[56984]_  = ~A302 & ~A301;
  assign \new_[56985]_  = \new_[56984]_  & \new_[56981]_ ;
  assign \new_[56986]_  = \new_[56985]_  & \new_[56978]_ ;
  assign \new_[56990]_  = ~A199 & A166;
  assign \new_[56991]_  = A167 & \new_[56990]_ ;
  assign \new_[56994]_  = ~A201 & A200;
  assign \new_[56997]_  = ~A203 & ~A202;
  assign \new_[56998]_  = \new_[56997]_  & \new_[56994]_ ;
  assign \new_[56999]_  = \new_[56998]_  & \new_[56991]_ ;
  assign \new_[57003]_  = ~A298 & A268;
  assign \new_[57004]_  = ~A267 & \new_[57003]_ ;
  assign \new_[57007]_  = ~A300 & A299;
  assign \new_[57010]_  = ~A302 & ~A301;
  assign \new_[57011]_  = \new_[57010]_  & \new_[57007]_ ;
  assign \new_[57012]_  = \new_[57011]_  & \new_[57004]_ ;
  assign \new_[57016]_  = ~A199 & A166;
  assign \new_[57017]_  = A167 & \new_[57016]_ ;
  assign \new_[57020]_  = ~A201 & A200;
  assign \new_[57023]_  = ~A203 & ~A202;
  assign \new_[57024]_  = \new_[57023]_  & \new_[57020]_ ;
  assign \new_[57025]_  = \new_[57024]_  & \new_[57017]_ ;
  assign \new_[57029]_  = A298 & A269;
  assign \new_[57030]_  = ~A267 & \new_[57029]_ ;
  assign \new_[57033]_  = ~A300 & ~A299;
  assign \new_[57036]_  = ~A302 & ~A301;
  assign \new_[57037]_  = \new_[57036]_  & \new_[57033]_ ;
  assign \new_[57038]_  = \new_[57037]_  & \new_[57030]_ ;
  assign \new_[57042]_  = ~A199 & A166;
  assign \new_[57043]_  = A167 & \new_[57042]_ ;
  assign \new_[57046]_  = ~A201 & A200;
  assign \new_[57049]_  = ~A203 & ~A202;
  assign \new_[57050]_  = \new_[57049]_  & \new_[57046]_ ;
  assign \new_[57051]_  = \new_[57050]_  & \new_[57043]_ ;
  assign \new_[57055]_  = ~A298 & A269;
  assign \new_[57056]_  = ~A267 & \new_[57055]_ ;
  assign \new_[57059]_  = ~A300 & A299;
  assign \new_[57062]_  = ~A302 & ~A301;
  assign \new_[57063]_  = \new_[57062]_  & \new_[57059]_ ;
  assign \new_[57064]_  = \new_[57063]_  & \new_[57056]_ ;
  assign \new_[57068]_  = ~A199 & A166;
  assign \new_[57069]_  = A167 & \new_[57068]_ ;
  assign \new_[57072]_  = ~A201 & A200;
  assign \new_[57075]_  = ~A203 & ~A202;
  assign \new_[57076]_  = \new_[57075]_  & \new_[57072]_ ;
  assign \new_[57077]_  = \new_[57076]_  & \new_[57069]_ ;
  assign \new_[57081]_  = A298 & A266;
  assign \new_[57082]_  = A265 & \new_[57081]_ ;
  assign \new_[57085]_  = ~A300 & ~A299;
  assign \new_[57088]_  = ~A302 & ~A301;
  assign \new_[57089]_  = \new_[57088]_  & \new_[57085]_ ;
  assign \new_[57090]_  = \new_[57089]_  & \new_[57082]_ ;
  assign \new_[57094]_  = ~A199 & A166;
  assign \new_[57095]_  = A167 & \new_[57094]_ ;
  assign \new_[57098]_  = ~A201 & A200;
  assign \new_[57101]_  = ~A203 & ~A202;
  assign \new_[57102]_  = \new_[57101]_  & \new_[57098]_ ;
  assign \new_[57103]_  = \new_[57102]_  & \new_[57095]_ ;
  assign \new_[57107]_  = ~A298 & A266;
  assign \new_[57108]_  = A265 & \new_[57107]_ ;
  assign \new_[57111]_  = ~A300 & A299;
  assign \new_[57114]_  = ~A302 & ~A301;
  assign \new_[57115]_  = \new_[57114]_  & \new_[57111]_ ;
  assign \new_[57116]_  = \new_[57115]_  & \new_[57108]_ ;
  assign \new_[57120]_  = ~A199 & A166;
  assign \new_[57121]_  = A167 & \new_[57120]_ ;
  assign \new_[57124]_  = ~A201 & A200;
  assign \new_[57127]_  = ~A203 & ~A202;
  assign \new_[57128]_  = \new_[57127]_  & \new_[57124]_ ;
  assign \new_[57129]_  = \new_[57128]_  & \new_[57121]_ ;
  assign \new_[57133]_  = A298 & ~A266;
  assign \new_[57134]_  = ~A265 & \new_[57133]_ ;
  assign \new_[57137]_  = ~A300 & ~A299;
  assign \new_[57140]_  = ~A302 & ~A301;
  assign \new_[57141]_  = \new_[57140]_  & \new_[57137]_ ;
  assign \new_[57142]_  = \new_[57141]_  & \new_[57134]_ ;
  assign \new_[57146]_  = ~A199 & A166;
  assign \new_[57147]_  = A167 & \new_[57146]_ ;
  assign \new_[57150]_  = ~A201 & A200;
  assign \new_[57153]_  = ~A203 & ~A202;
  assign \new_[57154]_  = \new_[57153]_  & \new_[57150]_ ;
  assign \new_[57155]_  = \new_[57154]_  & \new_[57147]_ ;
  assign \new_[57159]_  = ~A298 & ~A266;
  assign \new_[57160]_  = ~A265 & \new_[57159]_ ;
  assign \new_[57163]_  = ~A300 & A299;
  assign \new_[57166]_  = ~A302 & ~A301;
  assign \new_[57167]_  = \new_[57166]_  & \new_[57163]_ ;
  assign \new_[57168]_  = \new_[57167]_  & \new_[57160]_ ;
  assign \new_[57172]_  = A199 & A166;
  assign \new_[57173]_  = A167 & \new_[57172]_ ;
  assign \new_[57176]_  = A201 & ~A200;
  assign \new_[57179]_  = A267 & A202;
  assign \new_[57180]_  = \new_[57179]_  & \new_[57176]_ ;
  assign \new_[57181]_  = \new_[57180]_  & \new_[57173]_ ;
  assign \new_[57185]_  = A298 & ~A269;
  assign \new_[57186]_  = ~A268 & \new_[57185]_ ;
  assign \new_[57189]_  = ~A300 & ~A299;
  assign \new_[57192]_  = ~A302 & ~A301;
  assign \new_[57193]_  = \new_[57192]_  & \new_[57189]_ ;
  assign \new_[57194]_  = \new_[57193]_  & \new_[57186]_ ;
  assign \new_[57198]_  = A199 & A166;
  assign \new_[57199]_  = A167 & \new_[57198]_ ;
  assign \new_[57202]_  = A201 & ~A200;
  assign \new_[57205]_  = A267 & A202;
  assign \new_[57206]_  = \new_[57205]_  & \new_[57202]_ ;
  assign \new_[57207]_  = \new_[57206]_  & \new_[57199]_ ;
  assign \new_[57211]_  = ~A298 & ~A269;
  assign \new_[57212]_  = ~A268 & \new_[57211]_ ;
  assign \new_[57215]_  = ~A300 & A299;
  assign \new_[57218]_  = ~A302 & ~A301;
  assign \new_[57219]_  = \new_[57218]_  & \new_[57215]_ ;
  assign \new_[57220]_  = \new_[57219]_  & \new_[57212]_ ;
  assign \new_[57224]_  = A199 & A166;
  assign \new_[57225]_  = A167 & \new_[57224]_ ;
  assign \new_[57228]_  = A201 & ~A200;
  assign \new_[57231]_  = A267 & A203;
  assign \new_[57232]_  = \new_[57231]_  & \new_[57228]_ ;
  assign \new_[57233]_  = \new_[57232]_  & \new_[57225]_ ;
  assign \new_[57237]_  = A298 & ~A269;
  assign \new_[57238]_  = ~A268 & \new_[57237]_ ;
  assign \new_[57241]_  = ~A300 & ~A299;
  assign \new_[57244]_  = ~A302 & ~A301;
  assign \new_[57245]_  = \new_[57244]_  & \new_[57241]_ ;
  assign \new_[57246]_  = \new_[57245]_  & \new_[57238]_ ;
  assign \new_[57250]_  = A199 & A166;
  assign \new_[57251]_  = A167 & \new_[57250]_ ;
  assign \new_[57254]_  = A201 & ~A200;
  assign \new_[57257]_  = A267 & A203;
  assign \new_[57258]_  = \new_[57257]_  & \new_[57254]_ ;
  assign \new_[57259]_  = \new_[57258]_  & \new_[57251]_ ;
  assign \new_[57263]_  = ~A298 & ~A269;
  assign \new_[57264]_  = ~A268 & \new_[57263]_ ;
  assign \new_[57267]_  = ~A300 & A299;
  assign \new_[57270]_  = ~A302 & ~A301;
  assign \new_[57271]_  = \new_[57270]_  & \new_[57267]_ ;
  assign \new_[57272]_  = \new_[57271]_  & \new_[57264]_ ;
  assign \new_[57276]_  = A199 & A166;
  assign \new_[57277]_  = A167 & \new_[57276]_ ;
  assign \new_[57280]_  = ~A201 & ~A200;
  assign \new_[57283]_  = ~A203 & ~A202;
  assign \new_[57284]_  = \new_[57283]_  & \new_[57280]_ ;
  assign \new_[57285]_  = \new_[57284]_  & \new_[57277]_ ;
  assign \new_[57289]_  = ~A269 & ~A268;
  assign \new_[57290]_  = A267 & \new_[57289]_ ;
  assign \new_[57293]_  = ~A299 & A298;
  assign \new_[57296]_  = A301 & A300;
  assign \new_[57297]_  = \new_[57296]_  & \new_[57293]_ ;
  assign \new_[57298]_  = \new_[57297]_  & \new_[57290]_ ;
  assign \new_[57302]_  = A199 & A166;
  assign \new_[57303]_  = A167 & \new_[57302]_ ;
  assign \new_[57306]_  = ~A201 & ~A200;
  assign \new_[57309]_  = ~A203 & ~A202;
  assign \new_[57310]_  = \new_[57309]_  & \new_[57306]_ ;
  assign \new_[57311]_  = \new_[57310]_  & \new_[57303]_ ;
  assign \new_[57315]_  = ~A269 & ~A268;
  assign \new_[57316]_  = A267 & \new_[57315]_ ;
  assign \new_[57319]_  = ~A299 & A298;
  assign \new_[57322]_  = A302 & A300;
  assign \new_[57323]_  = \new_[57322]_  & \new_[57319]_ ;
  assign \new_[57324]_  = \new_[57323]_  & \new_[57316]_ ;
  assign \new_[57328]_  = A199 & A166;
  assign \new_[57329]_  = A167 & \new_[57328]_ ;
  assign \new_[57332]_  = ~A201 & ~A200;
  assign \new_[57335]_  = ~A203 & ~A202;
  assign \new_[57336]_  = \new_[57335]_  & \new_[57332]_ ;
  assign \new_[57337]_  = \new_[57336]_  & \new_[57329]_ ;
  assign \new_[57341]_  = ~A269 & ~A268;
  assign \new_[57342]_  = A267 & \new_[57341]_ ;
  assign \new_[57345]_  = A299 & ~A298;
  assign \new_[57348]_  = A301 & A300;
  assign \new_[57349]_  = \new_[57348]_  & \new_[57345]_ ;
  assign \new_[57350]_  = \new_[57349]_  & \new_[57342]_ ;
  assign \new_[57354]_  = A199 & A166;
  assign \new_[57355]_  = A167 & \new_[57354]_ ;
  assign \new_[57358]_  = ~A201 & ~A200;
  assign \new_[57361]_  = ~A203 & ~A202;
  assign \new_[57362]_  = \new_[57361]_  & \new_[57358]_ ;
  assign \new_[57363]_  = \new_[57362]_  & \new_[57355]_ ;
  assign \new_[57367]_  = ~A269 & ~A268;
  assign \new_[57368]_  = A267 & \new_[57367]_ ;
  assign \new_[57371]_  = A299 & ~A298;
  assign \new_[57374]_  = A302 & A300;
  assign \new_[57375]_  = \new_[57374]_  & \new_[57371]_ ;
  assign \new_[57376]_  = \new_[57375]_  & \new_[57368]_ ;
  assign \new_[57380]_  = A199 & A166;
  assign \new_[57381]_  = A167 & \new_[57380]_ ;
  assign \new_[57384]_  = ~A201 & ~A200;
  assign \new_[57387]_  = ~A203 & ~A202;
  assign \new_[57388]_  = \new_[57387]_  & \new_[57384]_ ;
  assign \new_[57389]_  = \new_[57388]_  & \new_[57381]_ ;
  assign \new_[57393]_  = A298 & A268;
  assign \new_[57394]_  = ~A267 & \new_[57393]_ ;
  assign \new_[57397]_  = ~A300 & ~A299;
  assign \new_[57400]_  = ~A302 & ~A301;
  assign \new_[57401]_  = \new_[57400]_  & \new_[57397]_ ;
  assign \new_[57402]_  = \new_[57401]_  & \new_[57394]_ ;
  assign \new_[57406]_  = A199 & A166;
  assign \new_[57407]_  = A167 & \new_[57406]_ ;
  assign \new_[57410]_  = ~A201 & ~A200;
  assign \new_[57413]_  = ~A203 & ~A202;
  assign \new_[57414]_  = \new_[57413]_  & \new_[57410]_ ;
  assign \new_[57415]_  = \new_[57414]_  & \new_[57407]_ ;
  assign \new_[57419]_  = ~A298 & A268;
  assign \new_[57420]_  = ~A267 & \new_[57419]_ ;
  assign \new_[57423]_  = ~A300 & A299;
  assign \new_[57426]_  = ~A302 & ~A301;
  assign \new_[57427]_  = \new_[57426]_  & \new_[57423]_ ;
  assign \new_[57428]_  = \new_[57427]_  & \new_[57420]_ ;
  assign \new_[57432]_  = A199 & A166;
  assign \new_[57433]_  = A167 & \new_[57432]_ ;
  assign \new_[57436]_  = ~A201 & ~A200;
  assign \new_[57439]_  = ~A203 & ~A202;
  assign \new_[57440]_  = \new_[57439]_  & \new_[57436]_ ;
  assign \new_[57441]_  = \new_[57440]_  & \new_[57433]_ ;
  assign \new_[57445]_  = A298 & A269;
  assign \new_[57446]_  = ~A267 & \new_[57445]_ ;
  assign \new_[57449]_  = ~A300 & ~A299;
  assign \new_[57452]_  = ~A302 & ~A301;
  assign \new_[57453]_  = \new_[57452]_  & \new_[57449]_ ;
  assign \new_[57454]_  = \new_[57453]_  & \new_[57446]_ ;
  assign \new_[57458]_  = A199 & A166;
  assign \new_[57459]_  = A167 & \new_[57458]_ ;
  assign \new_[57462]_  = ~A201 & ~A200;
  assign \new_[57465]_  = ~A203 & ~A202;
  assign \new_[57466]_  = \new_[57465]_  & \new_[57462]_ ;
  assign \new_[57467]_  = \new_[57466]_  & \new_[57459]_ ;
  assign \new_[57471]_  = ~A298 & A269;
  assign \new_[57472]_  = ~A267 & \new_[57471]_ ;
  assign \new_[57475]_  = ~A300 & A299;
  assign \new_[57478]_  = ~A302 & ~A301;
  assign \new_[57479]_  = \new_[57478]_  & \new_[57475]_ ;
  assign \new_[57480]_  = \new_[57479]_  & \new_[57472]_ ;
  assign \new_[57484]_  = A199 & A166;
  assign \new_[57485]_  = A167 & \new_[57484]_ ;
  assign \new_[57488]_  = ~A201 & ~A200;
  assign \new_[57491]_  = ~A203 & ~A202;
  assign \new_[57492]_  = \new_[57491]_  & \new_[57488]_ ;
  assign \new_[57493]_  = \new_[57492]_  & \new_[57485]_ ;
  assign \new_[57497]_  = A298 & A266;
  assign \new_[57498]_  = A265 & \new_[57497]_ ;
  assign \new_[57501]_  = ~A300 & ~A299;
  assign \new_[57504]_  = ~A302 & ~A301;
  assign \new_[57505]_  = \new_[57504]_  & \new_[57501]_ ;
  assign \new_[57506]_  = \new_[57505]_  & \new_[57498]_ ;
  assign \new_[57510]_  = A199 & A166;
  assign \new_[57511]_  = A167 & \new_[57510]_ ;
  assign \new_[57514]_  = ~A201 & ~A200;
  assign \new_[57517]_  = ~A203 & ~A202;
  assign \new_[57518]_  = \new_[57517]_  & \new_[57514]_ ;
  assign \new_[57519]_  = \new_[57518]_  & \new_[57511]_ ;
  assign \new_[57523]_  = ~A298 & A266;
  assign \new_[57524]_  = A265 & \new_[57523]_ ;
  assign \new_[57527]_  = ~A300 & A299;
  assign \new_[57530]_  = ~A302 & ~A301;
  assign \new_[57531]_  = \new_[57530]_  & \new_[57527]_ ;
  assign \new_[57532]_  = \new_[57531]_  & \new_[57524]_ ;
  assign \new_[57536]_  = A199 & A166;
  assign \new_[57537]_  = A167 & \new_[57536]_ ;
  assign \new_[57540]_  = ~A201 & ~A200;
  assign \new_[57543]_  = ~A203 & ~A202;
  assign \new_[57544]_  = \new_[57543]_  & \new_[57540]_ ;
  assign \new_[57545]_  = \new_[57544]_  & \new_[57537]_ ;
  assign \new_[57549]_  = A298 & ~A266;
  assign \new_[57550]_  = ~A265 & \new_[57549]_ ;
  assign \new_[57553]_  = ~A300 & ~A299;
  assign \new_[57556]_  = ~A302 & ~A301;
  assign \new_[57557]_  = \new_[57556]_  & \new_[57553]_ ;
  assign \new_[57558]_  = \new_[57557]_  & \new_[57550]_ ;
  assign \new_[57562]_  = A199 & A166;
  assign \new_[57563]_  = A167 & \new_[57562]_ ;
  assign \new_[57566]_  = ~A201 & ~A200;
  assign \new_[57569]_  = ~A203 & ~A202;
  assign \new_[57570]_  = \new_[57569]_  & \new_[57566]_ ;
  assign \new_[57571]_  = \new_[57570]_  & \new_[57563]_ ;
  assign \new_[57575]_  = ~A298 & ~A266;
  assign \new_[57576]_  = ~A265 & \new_[57575]_ ;
  assign \new_[57579]_  = ~A300 & A299;
  assign \new_[57582]_  = ~A302 & ~A301;
  assign \new_[57583]_  = \new_[57582]_  & \new_[57579]_ ;
  assign \new_[57584]_  = \new_[57583]_  & \new_[57576]_ ;
  assign \new_[57588]_  = ~A199 & ~A166;
  assign \new_[57589]_  = ~A167 & \new_[57588]_ ;
  assign \new_[57592]_  = A201 & A200;
  assign \new_[57595]_  = A267 & A202;
  assign \new_[57596]_  = \new_[57595]_  & \new_[57592]_ ;
  assign \new_[57597]_  = \new_[57596]_  & \new_[57589]_ ;
  assign \new_[57601]_  = A298 & ~A269;
  assign \new_[57602]_  = ~A268 & \new_[57601]_ ;
  assign \new_[57605]_  = ~A300 & ~A299;
  assign \new_[57608]_  = ~A302 & ~A301;
  assign \new_[57609]_  = \new_[57608]_  & \new_[57605]_ ;
  assign \new_[57610]_  = \new_[57609]_  & \new_[57602]_ ;
  assign \new_[57614]_  = ~A199 & ~A166;
  assign \new_[57615]_  = ~A167 & \new_[57614]_ ;
  assign \new_[57618]_  = A201 & A200;
  assign \new_[57621]_  = A267 & A202;
  assign \new_[57622]_  = \new_[57621]_  & \new_[57618]_ ;
  assign \new_[57623]_  = \new_[57622]_  & \new_[57615]_ ;
  assign \new_[57627]_  = ~A298 & ~A269;
  assign \new_[57628]_  = ~A268 & \new_[57627]_ ;
  assign \new_[57631]_  = ~A300 & A299;
  assign \new_[57634]_  = ~A302 & ~A301;
  assign \new_[57635]_  = \new_[57634]_  & \new_[57631]_ ;
  assign \new_[57636]_  = \new_[57635]_  & \new_[57628]_ ;
  assign \new_[57640]_  = ~A199 & ~A166;
  assign \new_[57641]_  = ~A167 & \new_[57640]_ ;
  assign \new_[57644]_  = A201 & A200;
  assign \new_[57647]_  = A267 & A203;
  assign \new_[57648]_  = \new_[57647]_  & \new_[57644]_ ;
  assign \new_[57649]_  = \new_[57648]_  & \new_[57641]_ ;
  assign \new_[57653]_  = A298 & ~A269;
  assign \new_[57654]_  = ~A268 & \new_[57653]_ ;
  assign \new_[57657]_  = ~A300 & ~A299;
  assign \new_[57660]_  = ~A302 & ~A301;
  assign \new_[57661]_  = \new_[57660]_  & \new_[57657]_ ;
  assign \new_[57662]_  = \new_[57661]_  & \new_[57654]_ ;
  assign \new_[57666]_  = ~A199 & ~A166;
  assign \new_[57667]_  = ~A167 & \new_[57666]_ ;
  assign \new_[57670]_  = A201 & A200;
  assign \new_[57673]_  = A267 & A203;
  assign \new_[57674]_  = \new_[57673]_  & \new_[57670]_ ;
  assign \new_[57675]_  = \new_[57674]_  & \new_[57667]_ ;
  assign \new_[57679]_  = ~A298 & ~A269;
  assign \new_[57680]_  = ~A268 & \new_[57679]_ ;
  assign \new_[57683]_  = ~A300 & A299;
  assign \new_[57686]_  = ~A302 & ~A301;
  assign \new_[57687]_  = \new_[57686]_  & \new_[57683]_ ;
  assign \new_[57688]_  = \new_[57687]_  & \new_[57680]_ ;
  assign \new_[57692]_  = ~A199 & ~A166;
  assign \new_[57693]_  = ~A167 & \new_[57692]_ ;
  assign \new_[57696]_  = ~A201 & A200;
  assign \new_[57699]_  = ~A203 & ~A202;
  assign \new_[57700]_  = \new_[57699]_  & \new_[57696]_ ;
  assign \new_[57701]_  = \new_[57700]_  & \new_[57693]_ ;
  assign \new_[57705]_  = ~A269 & ~A268;
  assign \new_[57706]_  = A267 & \new_[57705]_ ;
  assign \new_[57709]_  = ~A299 & A298;
  assign \new_[57712]_  = A301 & A300;
  assign \new_[57713]_  = \new_[57712]_  & \new_[57709]_ ;
  assign \new_[57714]_  = \new_[57713]_  & \new_[57706]_ ;
  assign \new_[57718]_  = ~A199 & ~A166;
  assign \new_[57719]_  = ~A167 & \new_[57718]_ ;
  assign \new_[57722]_  = ~A201 & A200;
  assign \new_[57725]_  = ~A203 & ~A202;
  assign \new_[57726]_  = \new_[57725]_  & \new_[57722]_ ;
  assign \new_[57727]_  = \new_[57726]_  & \new_[57719]_ ;
  assign \new_[57731]_  = ~A269 & ~A268;
  assign \new_[57732]_  = A267 & \new_[57731]_ ;
  assign \new_[57735]_  = ~A299 & A298;
  assign \new_[57738]_  = A302 & A300;
  assign \new_[57739]_  = \new_[57738]_  & \new_[57735]_ ;
  assign \new_[57740]_  = \new_[57739]_  & \new_[57732]_ ;
  assign \new_[57744]_  = ~A199 & ~A166;
  assign \new_[57745]_  = ~A167 & \new_[57744]_ ;
  assign \new_[57748]_  = ~A201 & A200;
  assign \new_[57751]_  = ~A203 & ~A202;
  assign \new_[57752]_  = \new_[57751]_  & \new_[57748]_ ;
  assign \new_[57753]_  = \new_[57752]_  & \new_[57745]_ ;
  assign \new_[57757]_  = ~A269 & ~A268;
  assign \new_[57758]_  = A267 & \new_[57757]_ ;
  assign \new_[57761]_  = A299 & ~A298;
  assign \new_[57764]_  = A301 & A300;
  assign \new_[57765]_  = \new_[57764]_  & \new_[57761]_ ;
  assign \new_[57766]_  = \new_[57765]_  & \new_[57758]_ ;
  assign \new_[57770]_  = ~A199 & ~A166;
  assign \new_[57771]_  = ~A167 & \new_[57770]_ ;
  assign \new_[57774]_  = ~A201 & A200;
  assign \new_[57777]_  = ~A203 & ~A202;
  assign \new_[57778]_  = \new_[57777]_  & \new_[57774]_ ;
  assign \new_[57779]_  = \new_[57778]_  & \new_[57771]_ ;
  assign \new_[57783]_  = ~A269 & ~A268;
  assign \new_[57784]_  = A267 & \new_[57783]_ ;
  assign \new_[57787]_  = A299 & ~A298;
  assign \new_[57790]_  = A302 & A300;
  assign \new_[57791]_  = \new_[57790]_  & \new_[57787]_ ;
  assign \new_[57792]_  = \new_[57791]_  & \new_[57784]_ ;
  assign \new_[57796]_  = ~A199 & ~A166;
  assign \new_[57797]_  = ~A167 & \new_[57796]_ ;
  assign \new_[57800]_  = ~A201 & A200;
  assign \new_[57803]_  = ~A203 & ~A202;
  assign \new_[57804]_  = \new_[57803]_  & \new_[57800]_ ;
  assign \new_[57805]_  = \new_[57804]_  & \new_[57797]_ ;
  assign \new_[57809]_  = A298 & A268;
  assign \new_[57810]_  = ~A267 & \new_[57809]_ ;
  assign \new_[57813]_  = ~A300 & ~A299;
  assign \new_[57816]_  = ~A302 & ~A301;
  assign \new_[57817]_  = \new_[57816]_  & \new_[57813]_ ;
  assign \new_[57818]_  = \new_[57817]_  & \new_[57810]_ ;
  assign \new_[57822]_  = ~A199 & ~A166;
  assign \new_[57823]_  = ~A167 & \new_[57822]_ ;
  assign \new_[57826]_  = ~A201 & A200;
  assign \new_[57829]_  = ~A203 & ~A202;
  assign \new_[57830]_  = \new_[57829]_  & \new_[57826]_ ;
  assign \new_[57831]_  = \new_[57830]_  & \new_[57823]_ ;
  assign \new_[57835]_  = ~A298 & A268;
  assign \new_[57836]_  = ~A267 & \new_[57835]_ ;
  assign \new_[57839]_  = ~A300 & A299;
  assign \new_[57842]_  = ~A302 & ~A301;
  assign \new_[57843]_  = \new_[57842]_  & \new_[57839]_ ;
  assign \new_[57844]_  = \new_[57843]_  & \new_[57836]_ ;
  assign \new_[57848]_  = ~A199 & ~A166;
  assign \new_[57849]_  = ~A167 & \new_[57848]_ ;
  assign \new_[57852]_  = ~A201 & A200;
  assign \new_[57855]_  = ~A203 & ~A202;
  assign \new_[57856]_  = \new_[57855]_  & \new_[57852]_ ;
  assign \new_[57857]_  = \new_[57856]_  & \new_[57849]_ ;
  assign \new_[57861]_  = A298 & A269;
  assign \new_[57862]_  = ~A267 & \new_[57861]_ ;
  assign \new_[57865]_  = ~A300 & ~A299;
  assign \new_[57868]_  = ~A302 & ~A301;
  assign \new_[57869]_  = \new_[57868]_  & \new_[57865]_ ;
  assign \new_[57870]_  = \new_[57869]_  & \new_[57862]_ ;
  assign \new_[57874]_  = ~A199 & ~A166;
  assign \new_[57875]_  = ~A167 & \new_[57874]_ ;
  assign \new_[57878]_  = ~A201 & A200;
  assign \new_[57881]_  = ~A203 & ~A202;
  assign \new_[57882]_  = \new_[57881]_  & \new_[57878]_ ;
  assign \new_[57883]_  = \new_[57882]_  & \new_[57875]_ ;
  assign \new_[57887]_  = ~A298 & A269;
  assign \new_[57888]_  = ~A267 & \new_[57887]_ ;
  assign \new_[57891]_  = ~A300 & A299;
  assign \new_[57894]_  = ~A302 & ~A301;
  assign \new_[57895]_  = \new_[57894]_  & \new_[57891]_ ;
  assign \new_[57896]_  = \new_[57895]_  & \new_[57888]_ ;
  assign \new_[57900]_  = ~A199 & ~A166;
  assign \new_[57901]_  = ~A167 & \new_[57900]_ ;
  assign \new_[57904]_  = ~A201 & A200;
  assign \new_[57907]_  = ~A203 & ~A202;
  assign \new_[57908]_  = \new_[57907]_  & \new_[57904]_ ;
  assign \new_[57909]_  = \new_[57908]_  & \new_[57901]_ ;
  assign \new_[57913]_  = A298 & A266;
  assign \new_[57914]_  = A265 & \new_[57913]_ ;
  assign \new_[57917]_  = ~A300 & ~A299;
  assign \new_[57920]_  = ~A302 & ~A301;
  assign \new_[57921]_  = \new_[57920]_  & \new_[57917]_ ;
  assign \new_[57922]_  = \new_[57921]_  & \new_[57914]_ ;
  assign \new_[57926]_  = ~A199 & ~A166;
  assign \new_[57927]_  = ~A167 & \new_[57926]_ ;
  assign \new_[57930]_  = ~A201 & A200;
  assign \new_[57933]_  = ~A203 & ~A202;
  assign \new_[57934]_  = \new_[57933]_  & \new_[57930]_ ;
  assign \new_[57935]_  = \new_[57934]_  & \new_[57927]_ ;
  assign \new_[57939]_  = ~A298 & A266;
  assign \new_[57940]_  = A265 & \new_[57939]_ ;
  assign \new_[57943]_  = ~A300 & A299;
  assign \new_[57946]_  = ~A302 & ~A301;
  assign \new_[57947]_  = \new_[57946]_  & \new_[57943]_ ;
  assign \new_[57948]_  = \new_[57947]_  & \new_[57940]_ ;
  assign \new_[57952]_  = ~A199 & ~A166;
  assign \new_[57953]_  = ~A167 & \new_[57952]_ ;
  assign \new_[57956]_  = ~A201 & A200;
  assign \new_[57959]_  = ~A203 & ~A202;
  assign \new_[57960]_  = \new_[57959]_  & \new_[57956]_ ;
  assign \new_[57961]_  = \new_[57960]_  & \new_[57953]_ ;
  assign \new_[57965]_  = A298 & ~A266;
  assign \new_[57966]_  = ~A265 & \new_[57965]_ ;
  assign \new_[57969]_  = ~A300 & ~A299;
  assign \new_[57972]_  = ~A302 & ~A301;
  assign \new_[57973]_  = \new_[57972]_  & \new_[57969]_ ;
  assign \new_[57974]_  = \new_[57973]_  & \new_[57966]_ ;
  assign \new_[57978]_  = ~A199 & ~A166;
  assign \new_[57979]_  = ~A167 & \new_[57978]_ ;
  assign \new_[57982]_  = ~A201 & A200;
  assign \new_[57985]_  = ~A203 & ~A202;
  assign \new_[57986]_  = \new_[57985]_  & \new_[57982]_ ;
  assign \new_[57987]_  = \new_[57986]_  & \new_[57979]_ ;
  assign \new_[57991]_  = ~A298 & ~A266;
  assign \new_[57992]_  = ~A265 & \new_[57991]_ ;
  assign \new_[57995]_  = ~A300 & A299;
  assign \new_[57998]_  = ~A302 & ~A301;
  assign \new_[57999]_  = \new_[57998]_  & \new_[57995]_ ;
  assign \new_[58000]_  = \new_[57999]_  & \new_[57992]_ ;
  assign \new_[58004]_  = A199 & ~A166;
  assign \new_[58005]_  = ~A167 & \new_[58004]_ ;
  assign \new_[58008]_  = A201 & ~A200;
  assign \new_[58011]_  = A267 & A202;
  assign \new_[58012]_  = \new_[58011]_  & \new_[58008]_ ;
  assign \new_[58013]_  = \new_[58012]_  & \new_[58005]_ ;
  assign \new_[58017]_  = A298 & ~A269;
  assign \new_[58018]_  = ~A268 & \new_[58017]_ ;
  assign \new_[58021]_  = ~A300 & ~A299;
  assign \new_[58024]_  = ~A302 & ~A301;
  assign \new_[58025]_  = \new_[58024]_  & \new_[58021]_ ;
  assign \new_[58026]_  = \new_[58025]_  & \new_[58018]_ ;
  assign \new_[58030]_  = A199 & ~A166;
  assign \new_[58031]_  = ~A167 & \new_[58030]_ ;
  assign \new_[58034]_  = A201 & ~A200;
  assign \new_[58037]_  = A267 & A202;
  assign \new_[58038]_  = \new_[58037]_  & \new_[58034]_ ;
  assign \new_[58039]_  = \new_[58038]_  & \new_[58031]_ ;
  assign \new_[58043]_  = ~A298 & ~A269;
  assign \new_[58044]_  = ~A268 & \new_[58043]_ ;
  assign \new_[58047]_  = ~A300 & A299;
  assign \new_[58050]_  = ~A302 & ~A301;
  assign \new_[58051]_  = \new_[58050]_  & \new_[58047]_ ;
  assign \new_[58052]_  = \new_[58051]_  & \new_[58044]_ ;
  assign \new_[58056]_  = A199 & ~A166;
  assign \new_[58057]_  = ~A167 & \new_[58056]_ ;
  assign \new_[58060]_  = A201 & ~A200;
  assign \new_[58063]_  = A267 & A203;
  assign \new_[58064]_  = \new_[58063]_  & \new_[58060]_ ;
  assign \new_[58065]_  = \new_[58064]_  & \new_[58057]_ ;
  assign \new_[58069]_  = A298 & ~A269;
  assign \new_[58070]_  = ~A268 & \new_[58069]_ ;
  assign \new_[58073]_  = ~A300 & ~A299;
  assign \new_[58076]_  = ~A302 & ~A301;
  assign \new_[58077]_  = \new_[58076]_  & \new_[58073]_ ;
  assign \new_[58078]_  = \new_[58077]_  & \new_[58070]_ ;
  assign \new_[58082]_  = A199 & ~A166;
  assign \new_[58083]_  = ~A167 & \new_[58082]_ ;
  assign \new_[58086]_  = A201 & ~A200;
  assign \new_[58089]_  = A267 & A203;
  assign \new_[58090]_  = \new_[58089]_  & \new_[58086]_ ;
  assign \new_[58091]_  = \new_[58090]_  & \new_[58083]_ ;
  assign \new_[58095]_  = ~A298 & ~A269;
  assign \new_[58096]_  = ~A268 & \new_[58095]_ ;
  assign \new_[58099]_  = ~A300 & A299;
  assign \new_[58102]_  = ~A302 & ~A301;
  assign \new_[58103]_  = \new_[58102]_  & \new_[58099]_ ;
  assign \new_[58104]_  = \new_[58103]_  & \new_[58096]_ ;
  assign \new_[58108]_  = A199 & ~A166;
  assign \new_[58109]_  = ~A167 & \new_[58108]_ ;
  assign \new_[58112]_  = ~A201 & ~A200;
  assign \new_[58115]_  = ~A203 & ~A202;
  assign \new_[58116]_  = \new_[58115]_  & \new_[58112]_ ;
  assign \new_[58117]_  = \new_[58116]_  & \new_[58109]_ ;
  assign \new_[58121]_  = ~A269 & ~A268;
  assign \new_[58122]_  = A267 & \new_[58121]_ ;
  assign \new_[58125]_  = ~A299 & A298;
  assign \new_[58128]_  = A301 & A300;
  assign \new_[58129]_  = \new_[58128]_  & \new_[58125]_ ;
  assign \new_[58130]_  = \new_[58129]_  & \new_[58122]_ ;
  assign \new_[58134]_  = A199 & ~A166;
  assign \new_[58135]_  = ~A167 & \new_[58134]_ ;
  assign \new_[58138]_  = ~A201 & ~A200;
  assign \new_[58141]_  = ~A203 & ~A202;
  assign \new_[58142]_  = \new_[58141]_  & \new_[58138]_ ;
  assign \new_[58143]_  = \new_[58142]_  & \new_[58135]_ ;
  assign \new_[58147]_  = ~A269 & ~A268;
  assign \new_[58148]_  = A267 & \new_[58147]_ ;
  assign \new_[58151]_  = ~A299 & A298;
  assign \new_[58154]_  = A302 & A300;
  assign \new_[58155]_  = \new_[58154]_  & \new_[58151]_ ;
  assign \new_[58156]_  = \new_[58155]_  & \new_[58148]_ ;
  assign \new_[58160]_  = A199 & ~A166;
  assign \new_[58161]_  = ~A167 & \new_[58160]_ ;
  assign \new_[58164]_  = ~A201 & ~A200;
  assign \new_[58167]_  = ~A203 & ~A202;
  assign \new_[58168]_  = \new_[58167]_  & \new_[58164]_ ;
  assign \new_[58169]_  = \new_[58168]_  & \new_[58161]_ ;
  assign \new_[58173]_  = ~A269 & ~A268;
  assign \new_[58174]_  = A267 & \new_[58173]_ ;
  assign \new_[58177]_  = A299 & ~A298;
  assign \new_[58180]_  = A301 & A300;
  assign \new_[58181]_  = \new_[58180]_  & \new_[58177]_ ;
  assign \new_[58182]_  = \new_[58181]_  & \new_[58174]_ ;
  assign \new_[58186]_  = A199 & ~A166;
  assign \new_[58187]_  = ~A167 & \new_[58186]_ ;
  assign \new_[58190]_  = ~A201 & ~A200;
  assign \new_[58193]_  = ~A203 & ~A202;
  assign \new_[58194]_  = \new_[58193]_  & \new_[58190]_ ;
  assign \new_[58195]_  = \new_[58194]_  & \new_[58187]_ ;
  assign \new_[58199]_  = ~A269 & ~A268;
  assign \new_[58200]_  = A267 & \new_[58199]_ ;
  assign \new_[58203]_  = A299 & ~A298;
  assign \new_[58206]_  = A302 & A300;
  assign \new_[58207]_  = \new_[58206]_  & \new_[58203]_ ;
  assign \new_[58208]_  = \new_[58207]_  & \new_[58200]_ ;
  assign \new_[58212]_  = A199 & ~A166;
  assign \new_[58213]_  = ~A167 & \new_[58212]_ ;
  assign \new_[58216]_  = ~A201 & ~A200;
  assign \new_[58219]_  = ~A203 & ~A202;
  assign \new_[58220]_  = \new_[58219]_  & \new_[58216]_ ;
  assign \new_[58221]_  = \new_[58220]_  & \new_[58213]_ ;
  assign \new_[58225]_  = A298 & A268;
  assign \new_[58226]_  = ~A267 & \new_[58225]_ ;
  assign \new_[58229]_  = ~A300 & ~A299;
  assign \new_[58232]_  = ~A302 & ~A301;
  assign \new_[58233]_  = \new_[58232]_  & \new_[58229]_ ;
  assign \new_[58234]_  = \new_[58233]_  & \new_[58226]_ ;
  assign \new_[58238]_  = A199 & ~A166;
  assign \new_[58239]_  = ~A167 & \new_[58238]_ ;
  assign \new_[58242]_  = ~A201 & ~A200;
  assign \new_[58245]_  = ~A203 & ~A202;
  assign \new_[58246]_  = \new_[58245]_  & \new_[58242]_ ;
  assign \new_[58247]_  = \new_[58246]_  & \new_[58239]_ ;
  assign \new_[58251]_  = ~A298 & A268;
  assign \new_[58252]_  = ~A267 & \new_[58251]_ ;
  assign \new_[58255]_  = ~A300 & A299;
  assign \new_[58258]_  = ~A302 & ~A301;
  assign \new_[58259]_  = \new_[58258]_  & \new_[58255]_ ;
  assign \new_[58260]_  = \new_[58259]_  & \new_[58252]_ ;
  assign \new_[58264]_  = A199 & ~A166;
  assign \new_[58265]_  = ~A167 & \new_[58264]_ ;
  assign \new_[58268]_  = ~A201 & ~A200;
  assign \new_[58271]_  = ~A203 & ~A202;
  assign \new_[58272]_  = \new_[58271]_  & \new_[58268]_ ;
  assign \new_[58273]_  = \new_[58272]_  & \new_[58265]_ ;
  assign \new_[58277]_  = A298 & A269;
  assign \new_[58278]_  = ~A267 & \new_[58277]_ ;
  assign \new_[58281]_  = ~A300 & ~A299;
  assign \new_[58284]_  = ~A302 & ~A301;
  assign \new_[58285]_  = \new_[58284]_  & \new_[58281]_ ;
  assign \new_[58286]_  = \new_[58285]_  & \new_[58278]_ ;
  assign \new_[58290]_  = A199 & ~A166;
  assign \new_[58291]_  = ~A167 & \new_[58290]_ ;
  assign \new_[58294]_  = ~A201 & ~A200;
  assign \new_[58297]_  = ~A203 & ~A202;
  assign \new_[58298]_  = \new_[58297]_  & \new_[58294]_ ;
  assign \new_[58299]_  = \new_[58298]_  & \new_[58291]_ ;
  assign \new_[58303]_  = ~A298 & A269;
  assign \new_[58304]_  = ~A267 & \new_[58303]_ ;
  assign \new_[58307]_  = ~A300 & A299;
  assign \new_[58310]_  = ~A302 & ~A301;
  assign \new_[58311]_  = \new_[58310]_  & \new_[58307]_ ;
  assign \new_[58312]_  = \new_[58311]_  & \new_[58304]_ ;
  assign \new_[58316]_  = A199 & ~A166;
  assign \new_[58317]_  = ~A167 & \new_[58316]_ ;
  assign \new_[58320]_  = ~A201 & ~A200;
  assign \new_[58323]_  = ~A203 & ~A202;
  assign \new_[58324]_  = \new_[58323]_  & \new_[58320]_ ;
  assign \new_[58325]_  = \new_[58324]_  & \new_[58317]_ ;
  assign \new_[58329]_  = A298 & A266;
  assign \new_[58330]_  = A265 & \new_[58329]_ ;
  assign \new_[58333]_  = ~A300 & ~A299;
  assign \new_[58336]_  = ~A302 & ~A301;
  assign \new_[58337]_  = \new_[58336]_  & \new_[58333]_ ;
  assign \new_[58338]_  = \new_[58337]_  & \new_[58330]_ ;
  assign \new_[58342]_  = A199 & ~A166;
  assign \new_[58343]_  = ~A167 & \new_[58342]_ ;
  assign \new_[58346]_  = ~A201 & ~A200;
  assign \new_[58349]_  = ~A203 & ~A202;
  assign \new_[58350]_  = \new_[58349]_  & \new_[58346]_ ;
  assign \new_[58351]_  = \new_[58350]_  & \new_[58343]_ ;
  assign \new_[58355]_  = ~A298 & A266;
  assign \new_[58356]_  = A265 & \new_[58355]_ ;
  assign \new_[58359]_  = ~A300 & A299;
  assign \new_[58362]_  = ~A302 & ~A301;
  assign \new_[58363]_  = \new_[58362]_  & \new_[58359]_ ;
  assign \new_[58364]_  = \new_[58363]_  & \new_[58356]_ ;
  assign \new_[58368]_  = A199 & ~A166;
  assign \new_[58369]_  = ~A167 & \new_[58368]_ ;
  assign \new_[58372]_  = ~A201 & ~A200;
  assign \new_[58375]_  = ~A203 & ~A202;
  assign \new_[58376]_  = \new_[58375]_  & \new_[58372]_ ;
  assign \new_[58377]_  = \new_[58376]_  & \new_[58369]_ ;
  assign \new_[58381]_  = A298 & ~A266;
  assign \new_[58382]_  = ~A265 & \new_[58381]_ ;
  assign \new_[58385]_  = ~A300 & ~A299;
  assign \new_[58388]_  = ~A302 & ~A301;
  assign \new_[58389]_  = \new_[58388]_  & \new_[58385]_ ;
  assign \new_[58390]_  = \new_[58389]_  & \new_[58382]_ ;
  assign \new_[58394]_  = A199 & ~A166;
  assign \new_[58395]_  = ~A167 & \new_[58394]_ ;
  assign \new_[58398]_  = ~A201 & ~A200;
  assign \new_[58401]_  = ~A203 & ~A202;
  assign \new_[58402]_  = \new_[58401]_  & \new_[58398]_ ;
  assign \new_[58403]_  = \new_[58402]_  & \new_[58395]_ ;
  assign \new_[58407]_  = ~A298 & ~A266;
  assign \new_[58408]_  = ~A265 & \new_[58407]_ ;
  assign \new_[58411]_  = ~A300 & A299;
  assign \new_[58414]_  = ~A302 & ~A301;
  assign \new_[58415]_  = \new_[58414]_  & \new_[58411]_ ;
  assign \new_[58416]_  = \new_[58415]_  & \new_[58408]_ ;
  assign \new_[58420]_  = A167 & A168;
  assign \new_[58421]_  = ~A170 & \new_[58420]_ ;
  assign \new_[58424]_  = A201 & ~A166;
  assign \new_[58427]_  = ~A203 & ~A202;
  assign \new_[58428]_  = \new_[58427]_  & \new_[58424]_ ;
  assign \new_[58429]_  = \new_[58428]_  & \new_[58421]_ ;
  assign \new_[58433]_  = ~A269 & ~A268;
  assign \new_[58434]_  = A267 & \new_[58433]_ ;
  assign \new_[58437]_  = ~A299 & A298;
  assign \new_[58440]_  = A301 & A300;
  assign \new_[58441]_  = \new_[58440]_  & \new_[58437]_ ;
  assign \new_[58442]_  = \new_[58441]_  & \new_[58434]_ ;
  assign \new_[58446]_  = A167 & A168;
  assign \new_[58447]_  = ~A170 & \new_[58446]_ ;
  assign \new_[58450]_  = A201 & ~A166;
  assign \new_[58453]_  = ~A203 & ~A202;
  assign \new_[58454]_  = \new_[58453]_  & \new_[58450]_ ;
  assign \new_[58455]_  = \new_[58454]_  & \new_[58447]_ ;
  assign \new_[58459]_  = ~A269 & ~A268;
  assign \new_[58460]_  = A267 & \new_[58459]_ ;
  assign \new_[58463]_  = ~A299 & A298;
  assign \new_[58466]_  = A302 & A300;
  assign \new_[58467]_  = \new_[58466]_  & \new_[58463]_ ;
  assign \new_[58468]_  = \new_[58467]_  & \new_[58460]_ ;
  assign \new_[58472]_  = A167 & A168;
  assign \new_[58473]_  = ~A170 & \new_[58472]_ ;
  assign \new_[58476]_  = A201 & ~A166;
  assign \new_[58479]_  = ~A203 & ~A202;
  assign \new_[58480]_  = \new_[58479]_  & \new_[58476]_ ;
  assign \new_[58481]_  = \new_[58480]_  & \new_[58473]_ ;
  assign \new_[58485]_  = ~A269 & ~A268;
  assign \new_[58486]_  = A267 & \new_[58485]_ ;
  assign \new_[58489]_  = A299 & ~A298;
  assign \new_[58492]_  = A301 & A300;
  assign \new_[58493]_  = \new_[58492]_  & \new_[58489]_ ;
  assign \new_[58494]_  = \new_[58493]_  & \new_[58486]_ ;
  assign \new_[58498]_  = A167 & A168;
  assign \new_[58499]_  = ~A170 & \new_[58498]_ ;
  assign \new_[58502]_  = A201 & ~A166;
  assign \new_[58505]_  = ~A203 & ~A202;
  assign \new_[58506]_  = \new_[58505]_  & \new_[58502]_ ;
  assign \new_[58507]_  = \new_[58506]_  & \new_[58499]_ ;
  assign \new_[58511]_  = ~A269 & ~A268;
  assign \new_[58512]_  = A267 & \new_[58511]_ ;
  assign \new_[58515]_  = A299 & ~A298;
  assign \new_[58518]_  = A302 & A300;
  assign \new_[58519]_  = \new_[58518]_  & \new_[58515]_ ;
  assign \new_[58520]_  = \new_[58519]_  & \new_[58512]_ ;
  assign \new_[58524]_  = A167 & A168;
  assign \new_[58525]_  = ~A170 & \new_[58524]_ ;
  assign \new_[58528]_  = A201 & ~A166;
  assign \new_[58531]_  = ~A203 & ~A202;
  assign \new_[58532]_  = \new_[58531]_  & \new_[58528]_ ;
  assign \new_[58533]_  = \new_[58532]_  & \new_[58525]_ ;
  assign \new_[58537]_  = A298 & A268;
  assign \new_[58538]_  = ~A267 & \new_[58537]_ ;
  assign \new_[58541]_  = ~A300 & ~A299;
  assign \new_[58544]_  = ~A302 & ~A301;
  assign \new_[58545]_  = \new_[58544]_  & \new_[58541]_ ;
  assign \new_[58546]_  = \new_[58545]_  & \new_[58538]_ ;
  assign \new_[58550]_  = A167 & A168;
  assign \new_[58551]_  = ~A170 & \new_[58550]_ ;
  assign \new_[58554]_  = A201 & ~A166;
  assign \new_[58557]_  = ~A203 & ~A202;
  assign \new_[58558]_  = \new_[58557]_  & \new_[58554]_ ;
  assign \new_[58559]_  = \new_[58558]_  & \new_[58551]_ ;
  assign \new_[58563]_  = ~A298 & A268;
  assign \new_[58564]_  = ~A267 & \new_[58563]_ ;
  assign \new_[58567]_  = ~A300 & A299;
  assign \new_[58570]_  = ~A302 & ~A301;
  assign \new_[58571]_  = \new_[58570]_  & \new_[58567]_ ;
  assign \new_[58572]_  = \new_[58571]_  & \new_[58564]_ ;
  assign \new_[58576]_  = A167 & A168;
  assign \new_[58577]_  = ~A170 & \new_[58576]_ ;
  assign \new_[58580]_  = A201 & ~A166;
  assign \new_[58583]_  = ~A203 & ~A202;
  assign \new_[58584]_  = \new_[58583]_  & \new_[58580]_ ;
  assign \new_[58585]_  = \new_[58584]_  & \new_[58577]_ ;
  assign \new_[58589]_  = A298 & A269;
  assign \new_[58590]_  = ~A267 & \new_[58589]_ ;
  assign \new_[58593]_  = ~A300 & ~A299;
  assign \new_[58596]_  = ~A302 & ~A301;
  assign \new_[58597]_  = \new_[58596]_  & \new_[58593]_ ;
  assign \new_[58598]_  = \new_[58597]_  & \new_[58590]_ ;
  assign \new_[58602]_  = A167 & A168;
  assign \new_[58603]_  = ~A170 & \new_[58602]_ ;
  assign \new_[58606]_  = A201 & ~A166;
  assign \new_[58609]_  = ~A203 & ~A202;
  assign \new_[58610]_  = \new_[58609]_  & \new_[58606]_ ;
  assign \new_[58611]_  = \new_[58610]_  & \new_[58603]_ ;
  assign \new_[58615]_  = ~A298 & A269;
  assign \new_[58616]_  = ~A267 & \new_[58615]_ ;
  assign \new_[58619]_  = ~A300 & A299;
  assign \new_[58622]_  = ~A302 & ~A301;
  assign \new_[58623]_  = \new_[58622]_  & \new_[58619]_ ;
  assign \new_[58624]_  = \new_[58623]_  & \new_[58616]_ ;
  assign \new_[58628]_  = A167 & A168;
  assign \new_[58629]_  = ~A170 & \new_[58628]_ ;
  assign \new_[58632]_  = A201 & ~A166;
  assign \new_[58635]_  = ~A203 & ~A202;
  assign \new_[58636]_  = \new_[58635]_  & \new_[58632]_ ;
  assign \new_[58637]_  = \new_[58636]_  & \new_[58629]_ ;
  assign \new_[58641]_  = A298 & A266;
  assign \new_[58642]_  = A265 & \new_[58641]_ ;
  assign \new_[58645]_  = ~A300 & ~A299;
  assign \new_[58648]_  = ~A302 & ~A301;
  assign \new_[58649]_  = \new_[58648]_  & \new_[58645]_ ;
  assign \new_[58650]_  = \new_[58649]_  & \new_[58642]_ ;
  assign \new_[58654]_  = A167 & A168;
  assign \new_[58655]_  = ~A170 & \new_[58654]_ ;
  assign \new_[58658]_  = A201 & ~A166;
  assign \new_[58661]_  = ~A203 & ~A202;
  assign \new_[58662]_  = \new_[58661]_  & \new_[58658]_ ;
  assign \new_[58663]_  = \new_[58662]_  & \new_[58655]_ ;
  assign \new_[58667]_  = ~A298 & A266;
  assign \new_[58668]_  = A265 & \new_[58667]_ ;
  assign \new_[58671]_  = ~A300 & A299;
  assign \new_[58674]_  = ~A302 & ~A301;
  assign \new_[58675]_  = \new_[58674]_  & \new_[58671]_ ;
  assign \new_[58676]_  = \new_[58675]_  & \new_[58668]_ ;
  assign \new_[58680]_  = A167 & A168;
  assign \new_[58681]_  = ~A170 & \new_[58680]_ ;
  assign \new_[58684]_  = A201 & ~A166;
  assign \new_[58687]_  = ~A203 & ~A202;
  assign \new_[58688]_  = \new_[58687]_  & \new_[58684]_ ;
  assign \new_[58689]_  = \new_[58688]_  & \new_[58681]_ ;
  assign \new_[58693]_  = A298 & ~A266;
  assign \new_[58694]_  = ~A265 & \new_[58693]_ ;
  assign \new_[58697]_  = ~A300 & ~A299;
  assign \new_[58700]_  = ~A302 & ~A301;
  assign \new_[58701]_  = \new_[58700]_  & \new_[58697]_ ;
  assign \new_[58702]_  = \new_[58701]_  & \new_[58694]_ ;
  assign \new_[58706]_  = A167 & A168;
  assign \new_[58707]_  = ~A170 & \new_[58706]_ ;
  assign \new_[58710]_  = A201 & ~A166;
  assign \new_[58713]_  = ~A203 & ~A202;
  assign \new_[58714]_  = \new_[58713]_  & \new_[58710]_ ;
  assign \new_[58715]_  = \new_[58714]_  & \new_[58707]_ ;
  assign \new_[58719]_  = ~A298 & ~A266;
  assign \new_[58720]_  = ~A265 & \new_[58719]_ ;
  assign \new_[58723]_  = ~A300 & A299;
  assign \new_[58726]_  = ~A302 & ~A301;
  assign \new_[58727]_  = \new_[58726]_  & \new_[58723]_ ;
  assign \new_[58728]_  = \new_[58727]_  & \new_[58720]_ ;
  assign \new_[58732]_  = A167 & A168;
  assign \new_[58733]_  = ~A170 & \new_[58732]_ ;
  assign \new_[58736]_  = ~A201 & ~A166;
  assign \new_[58739]_  = A267 & A202;
  assign \new_[58740]_  = \new_[58739]_  & \new_[58736]_ ;
  assign \new_[58741]_  = \new_[58740]_  & \new_[58733]_ ;
  assign \new_[58745]_  = A298 & ~A269;
  assign \new_[58746]_  = ~A268 & \new_[58745]_ ;
  assign \new_[58749]_  = ~A300 & ~A299;
  assign \new_[58752]_  = ~A302 & ~A301;
  assign \new_[58753]_  = \new_[58752]_  & \new_[58749]_ ;
  assign \new_[58754]_  = \new_[58753]_  & \new_[58746]_ ;
  assign \new_[58758]_  = A167 & A168;
  assign \new_[58759]_  = ~A170 & \new_[58758]_ ;
  assign \new_[58762]_  = ~A201 & ~A166;
  assign \new_[58765]_  = A267 & A202;
  assign \new_[58766]_  = \new_[58765]_  & \new_[58762]_ ;
  assign \new_[58767]_  = \new_[58766]_  & \new_[58759]_ ;
  assign \new_[58771]_  = ~A298 & ~A269;
  assign \new_[58772]_  = ~A268 & \new_[58771]_ ;
  assign \new_[58775]_  = ~A300 & A299;
  assign \new_[58778]_  = ~A302 & ~A301;
  assign \new_[58779]_  = \new_[58778]_  & \new_[58775]_ ;
  assign \new_[58780]_  = \new_[58779]_  & \new_[58772]_ ;
  assign \new_[58784]_  = A167 & A168;
  assign \new_[58785]_  = ~A170 & \new_[58784]_ ;
  assign \new_[58788]_  = ~A201 & ~A166;
  assign \new_[58791]_  = A267 & A203;
  assign \new_[58792]_  = \new_[58791]_  & \new_[58788]_ ;
  assign \new_[58793]_  = \new_[58792]_  & \new_[58785]_ ;
  assign \new_[58797]_  = A298 & ~A269;
  assign \new_[58798]_  = ~A268 & \new_[58797]_ ;
  assign \new_[58801]_  = ~A300 & ~A299;
  assign \new_[58804]_  = ~A302 & ~A301;
  assign \new_[58805]_  = \new_[58804]_  & \new_[58801]_ ;
  assign \new_[58806]_  = \new_[58805]_  & \new_[58798]_ ;
  assign \new_[58810]_  = A167 & A168;
  assign \new_[58811]_  = ~A170 & \new_[58810]_ ;
  assign \new_[58814]_  = ~A201 & ~A166;
  assign \new_[58817]_  = A267 & A203;
  assign \new_[58818]_  = \new_[58817]_  & \new_[58814]_ ;
  assign \new_[58819]_  = \new_[58818]_  & \new_[58811]_ ;
  assign \new_[58823]_  = ~A298 & ~A269;
  assign \new_[58824]_  = ~A268 & \new_[58823]_ ;
  assign \new_[58827]_  = ~A300 & A299;
  assign \new_[58830]_  = ~A302 & ~A301;
  assign \new_[58831]_  = \new_[58830]_  & \new_[58827]_ ;
  assign \new_[58832]_  = \new_[58831]_  & \new_[58824]_ ;
  assign \new_[58836]_  = A167 & A168;
  assign \new_[58837]_  = ~A170 & \new_[58836]_ ;
  assign \new_[58840]_  = A199 & ~A166;
  assign \new_[58843]_  = A267 & A200;
  assign \new_[58844]_  = \new_[58843]_  & \new_[58840]_ ;
  assign \new_[58845]_  = \new_[58844]_  & \new_[58837]_ ;
  assign \new_[58849]_  = A298 & ~A269;
  assign \new_[58850]_  = ~A268 & \new_[58849]_ ;
  assign \new_[58853]_  = ~A300 & ~A299;
  assign \new_[58856]_  = ~A302 & ~A301;
  assign \new_[58857]_  = \new_[58856]_  & \new_[58853]_ ;
  assign \new_[58858]_  = \new_[58857]_  & \new_[58850]_ ;
  assign \new_[58862]_  = A167 & A168;
  assign \new_[58863]_  = ~A170 & \new_[58862]_ ;
  assign \new_[58866]_  = A199 & ~A166;
  assign \new_[58869]_  = A267 & A200;
  assign \new_[58870]_  = \new_[58869]_  & \new_[58866]_ ;
  assign \new_[58871]_  = \new_[58870]_  & \new_[58863]_ ;
  assign \new_[58875]_  = ~A298 & ~A269;
  assign \new_[58876]_  = ~A268 & \new_[58875]_ ;
  assign \new_[58879]_  = ~A300 & A299;
  assign \new_[58882]_  = ~A302 & ~A301;
  assign \new_[58883]_  = \new_[58882]_  & \new_[58879]_ ;
  assign \new_[58884]_  = \new_[58883]_  & \new_[58876]_ ;
  assign \new_[58888]_  = A167 & A168;
  assign \new_[58889]_  = ~A170 & \new_[58888]_ ;
  assign \new_[58892]_  = ~A199 & ~A166;
  assign \new_[58895]_  = A201 & A200;
  assign \new_[58896]_  = \new_[58895]_  & \new_[58892]_ ;
  assign \new_[58897]_  = \new_[58896]_  & \new_[58889]_ ;
  assign \new_[58901]_  = A266 & ~A265;
  assign \new_[58902]_  = A202 & \new_[58901]_ ;
  assign \new_[58905]_  = A268 & A267;
  assign \new_[58908]_  = A301 & ~A300;
  assign \new_[58909]_  = \new_[58908]_  & \new_[58905]_ ;
  assign \new_[58910]_  = \new_[58909]_  & \new_[58902]_ ;
  assign \new_[58914]_  = A167 & A168;
  assign \new_[58915]_  = ~A170 & \new_[58914]_ ;
  assign \new_[58918]_  = ~A199 & ~A166;
  assign \new_[58921]_  = A201 & A200;
  assign \new_[58922]_  = \new_[58921]_  & \new_[58918]_ ;
  assign \new_[58923]_  = \new_[58922]_  & \new_[58915]_ ;
  assign \new_[58927]_  = A266 & ~A265;
  assign \new_[58928]_  = A202 & \new_[58927]_ ;
  assign \new_[58931]_  = A268 & A267;
  assign \new_[58934]_  = A302 & ~A300;
  assign \new_[58935]_  = \new_[58934]_  & \new_[58931]_ ;
  assign \new_[58936]_  = \new_[58935]_  & \new_[58928]_ ;
  assign \new_[58940]_  = A167 & A168;
  assign \new_[58941]_  = ~A170 & \new_[58940]_ ;
  assign \new_[58944]_  = ~A199 & ~A166;
  assign \new_[58947]_  = A201 & A200;
  assign \new_[58948]_  = \new_[58947]_  & \new_[58944]_ ;
  assign \new_[58949]_  = \new_[58948]_  & \new_[58941]_ ;
  assign \new_[58953]_  = A266 & ~A265;
  assign \new_[58954]_  = A202 & \new_[58953]_ ;
  assign \new_[58957]_  = A268 & A267;
  assign \new_[58960]_  = A299 & A298;
  assign \new_[58961]_  = \new_[58960]_  & \new_[58957]_ ;
  assign \new_[58962]_  = \new_[58961]_  & \new_[58954]_ ;
  assign \new_[58966]_  = A167 & A168;
  assign \new_[58967]_  = ~A170 & \new_[58966]_ ;
  assign \new_[58970]_  = ~A199 & ~A166;
  assign \new_[58973]_  = A201 & A200;
  assign \new_[58974]_  = \new_[58973]_  & \new_[58970]_ ;
  assign \new_[58975]_  = \new_[58974]_  & \new_[58967]_ ;
  assign \new_[58979]_  = A266 & ~A265;
  assign \new_[58980]_  = A202 & \new_[58979]_ ;
  assign \new_[58983]_  = A268 & A267;
  assign \new_[58986]_  = ~A299 & ~A298;
  assign \new_[58987]_  = \new_[58986]_  & \new_[58983]_ ;
  assign \new_[58988]_  = \new_[58987]_  & \new_[58980]_ ;
  assign \new_[58992]_  = A167 & A168;
  assign \new_[58993]_  = ~A170 & \new_[58992]_ ;
  assign \new_[58996]_  = ~A199 & ~A166;
  assign \new_[58999]_  = A201 & A200;
  assign \new_[59000]_  = \new_[58999]_  & \new_[58996]_ ;
  assign \new_[59001]_  = \new_[59000]_  & \new_[58993]_ ;
  assign \new_[59005]_  = A266 & ~A265;
  assign \new_[59006]_  = A202 & \new_[59005]_ ;
  assign \new_[59009]_  = A269 & A267;
  assign \new_[59012]_  = A301 & ~A300;
  assign \new_[59013]_  = \new_[59012]_  & \new_[59009]_ ;
  assign \new_[59014]_  = \new_[59013]_  & \new_[59006]_ ;
  assign \new_[59018]_  = A167 & A168;
  assign \new_[59019]_  = ~A170 & \new_[59018]_ ;
  assign \new_[59022]_  = ~A199 & ~A166;
  assign \new_[59025]_  = A201 & A200;
  assign \new_[59026]_  = \new_[59025]_  & \new_[59022]_ ;
  assign \new_[59027]_  = \new_[59026]_  & \new_[59019]_ ;
  assign \new_[59031]_  = A266 & ~A265;
  assign \new_[59032]_  = A202 & \new_[59031]_ ;
  assign \new_[59035]_  = A269 & A267;
  assign \new_[59038]_  = A302 & ~A300;
  assign \new_[59039]_  = \new_[59038]_  & \new_[59035]_ ;
  assign \new_[59040]_  = \new_[59039]_  & \new_[59032]_ ;
  assign \new_[59044]_  = A167 & A168;
  assign \new_[59045]_  = ~A170 & \new_[59044]_ ;
  assign \new_[59048]_  = ~A199 & ~A166;
  assign \new_[59051]_  = A201 & A200;
  assign \new_[59052]_  = \new_[59051]_  & \new_[59048]_ ;
  assign \new_[59053]_  = \new_[59052]_  & \new_[59045]_ ;
  assign \new_[59057]_  = A266 & ~A265;
  assign \new_[59058]_  = A202 & \new_[59057]_ ;
  assign \new_[59061]_  = A269 & A267;
  assign \new_[59064]_  = A299 & A298;
  assign \new_[59065]_  = \new_[59064]_  & \new_[59061]_ ;
  assign \new_[59066]_  = \new_[59065]_  & \new_[59058]_ ;
  assign \new_[59070]_  = A167 & A168;
  assign \new_[59071]_  = ~A170 & \new_[59070]_ ;
  assign \new_[59074]_  = ~A199 & ~A166;
  assign \new_[59077]_  = A201 & A200;
  assign \new_[59078]_  = \new_[59077]_  & \new_[59074]_ ;
  assign \new_[59079]_  = \new_[59078]_  & \new_[59071]_ ;
  assign \new_[59083]_  = A266 & ~A265;
  assign \new_[59084]_  = A202 & \new_[59083]_ ;
  assign \new_[59087]_  = A269 & A267;
  assign \new_[59090]_  = ~A299 & ~A298;
  assign \new_[59091]_  = \new_[59090]_  & \new_[59087]_ ;
  assign \new_[59092]_  = \new_[59091]_  & \new_[59084]_ ;
  assign \new_[59096]_  = A167 & A168;
  assign \new_[59097]_  = ~A170 & \new_[59096]_ ;
  assign \new_[59100]_  = ~A199 & ~A166;
  assign \new_[59103]_  = A201 & A200;
  assign \new_[59104]_  = \new_[59103]_  & \new_[59100]_ ;
  assign \new_[59105]_  = \new_[59104]_  & \new_[59097]_ ;
  assign \new_[59109]_  = ~A266 & A265;
  assign \new_[59110]_  = A202 & \new_[59109]_ ;
  assign \new_[59113]_  = A268 & A267;
  assign \new_[59116]_  = A301 & ~A300;
  assign \new_[59117]_  = \new_[59116]_  & \new_[59113]_ ;
  assign \new_[59118]_  = \new_[59117]_  & \new_[59110]_ ;
  assign \new_[59122]_  = A167 & A168;
  assign \new_[59123]_  = ~A170 & \new_[59122]_ ;
  assign \new_[59126]_  = ~A199 & ~A166;
  assign \new_[59129]_  = A201 & A200;
  assign \new_[59130]_  = \new_[59129]_  & \new_[59126]_ ;
  assign \new_[59131]_  = \new_[59130]_  & \new_[59123]_ ;
  assign \new_[59135]_  = ~A266 & A265;
  assign \new_[59136]_  = A202 & \new_[59135]_ ;
  assign \new_[59139]_  = A268 & A267;
  assign \new_[59142]_  = A302 & ~A300;
  assign \new_[59143]_  = \new_[59142]_  & \new_[59139]_ ;
  assign \new_[59144]_  = \new_[59143]_  & \new_[59136]_ ;
  assign \new_[59148]_  = A167 & A168;
  assign \new_[59149]_  = ~A170 & \new_[59148]_ ;
  assign \new_[59152]_  = ~A199 & ~A166;
  assign \new_[59155]_  = A201 & A200;
  assign \new_[59156]_  = \new_[59155]_  & \new_[59152]_ ;
  assign \new_[59157]_  = \new_[59156]_  & \new_[59149]_ ;
  assign \new_[59161]_  = ~A266 & A265;
  assign \new_[59162]_  = A202 & \new_[59161]_ ;
  assign \new_[59165]_  = A268 & A267;
  assign \new_[59168]_  = A299 & A298;
  assign \new_[59169]_  = \new_[59168]_  & \new_[59165]_ ;
  assign \new_[59170]_  = \new_[59169]_  & \new_[59162]_ ;
  assign \new_[59174]_  = A167 & A168;
  assign \new_[59175]_  = ~A170 & \new_[59174]_ ;
  assign \new_[59178]_  = ~A199 & ~A166;
  assign \new_[59181]_  = A201 & A200;
  assign \new_[59182]_  = \new_[59181]_  & \new_[59178]_ ;
  assign \new_[59183]_  = \new_[59182]_  & \new_[59175]_ ;
  assign \new_[59187]_  = ~A266 & A265;
  assign \new_[59188]_  = A202 & \new_[59187]_ ;
  assign \new_[59191]_  = A268 & A267;
  assign \new_[59194]_  = ~A299 & ~A298;
  assign \new_[59195]_  = \new_[59194]_  & \new_[59191]_ ;
  assign \new_[59196]_  = \new_[59195]_  & \new_[59188]_ ;
  assign \new_[59200]_  = A167 & A168;
  assign \new_[59201]_  = ~A170 & \new_[59200]_ ;
  assign \new_[59204]_  = ~A199 & ~A166;
  assign \new_[59207]_  = A201 & A200;
  assign \new_[59208]_  = \new_[59207]_  & \new_[59204]_ ;
  assign \new_[59209]_  = \new_[59208]_  & \new_[59201]_ ;
  assign \new_[59213]_  = ~A266 & A265;
  assign \new_[59214]_  = A202 & \new_[59213]_ ;
  assign \new_[59217]_  = A269 & A267;
  assign \new_[59220]_  = A301 & ~A300;
  assign \new_[59221]_  = \new_[59220]_  & \new_[59217]_ ;
  assign \new_[59222]_  = \new_[59221]_  & \new_[59214]_ ;
  assign \new_[59226]_  = A167 & A168;
  assign \new_[59227]_  = ~A170 & \new_[59226]_ ;
  assign \new_[59230]_  = ~A199 & ~A166;
  assign \new_[59233]_  = A201 & A200;
  assign \new_[59234]_  = \new_[59233]_  & \new_[59230]_ ;
  assign \new_[59235]_  = \new_[59234]_  & \new_[59227]_ ;
  assign \new_[59239]_  = ~A266 & A265;
  assign \new_[59240]_  = A202 & \new_[59239]_ ;
  assign \new_[59243]_  = A269 & A267;
  assign \new_[59246]_  = A302 & ~A300;
  assign \new_[59247]_  = \new_[59246]_  & \new_[59243]_ ;
  assign \new_[59248]_  = \new_[59247]_  & \new_[59240]_ ;
  assign \new_[59252]_  = A167 & A168;
  assign \new_[59253]_  = ~A170 & \new_[59252]_ ;
  assign \new_[59256]_  = ~A199 & ~A166;
  assign \new_[59259]_  = A201 & A200;
  assign \new_[59260]_  = \new_[59259]_  & \new_[59256]_ ;
  assign \new_[59261]_  = \new_[59260]_  & \new_[59253]_ ;
  assign \new_[59265]_  = ~A266 & A265;
  assign \new_[59266]_  = A202 & \new_[59265]_ ;
  assign \new_[59269]_  = A269 & A267;
  assign \new_[59272]_  = A299 & A298;
  assign \new_[59273]_  = \new_[59272]_  & \new_[59269]_ ;
  assign \new_[59274]_  = \new_[59273]_  & \new_[59266]_ ;
  assign \new_[59278]_  = A167 & A168;
  assign \new_[59279]_  = ~A170 & \new_[59278]_ ;
  assign \new_[59282]_  = ~A199 & ~A166;
  assign \new_[59285]_  = A201 & A200;
  assign \new_[59286]_  = \new_[59285]_  & \new_[59282]_ ;
  assign \new_[59287]_  = \new_[59286]_  & \new_[59279]_ ;
  assign \new_[59291]_  = ~A266 & A265;
  assign \new_[59292]_  = A202 & \new_[59291]_ ;
  assign \new_[59295]_  = A269 & A267;
  assign \new_[59298]_  = ~A299 & ~A298;
  assign \new_[59299]_  = \new_[59298]_  & \new_[59295]_ ;
  assign \new_[59300]_  = \new_[59299]_  & \new_[59292]_ ;
  assign \new_[59304]_  = A167 & A168;
  assign \new_[59305]_  = ~A170 & \new_[59304]_ ;
  assign \new_[59308]_  = ~A199 & ~A166;
  assign \new_[59311]_  = A201 & A200;
  assign \new_[59312]_  = \new_[59311]_  & \new_[59308]_ ;
  assign \new_[59313]_  = \new_[59312]_  & \new_[59305]_ ;
  assign \new_[59317]_  = A266 & ~A265;
  assign \new_[59318]_  = A203 & \new_[59317]_ ;
  assign \new_[59321]_  = A268 & A267;
  assign \new_[59324]_  = A301 & ~A300;
  assign \new_[59325]_  = \new_[59324]_  & \new_[59321]_ ;
  assign \new_[59326]_  = \new_[59325]_  & \new_[59318]_ ;
  assign \new_[59330]_  = A167 & A168;
  assign \new_[59331]_  = ~A170 & \new_[59330]_ ;
  assign \new_[59334]_  = ~A199 & ~A166;
  assign \new_[59337]_  = A201 & A200;
  assign \new_[59338]_  = \new_[59337]_  & \new_[59334]_ ;
  assign \new_[59339]_  = \new_[59338]_  & \new_[59331]_ ;
  assign \new_[59343]_  = A266 & ~A265;
  assign \new_[59344]_  = A203 & \new_[59343]_ ;
  assign \new_[59347]_  = A268 & A267;
  assign \new_[59350]_  = A302 & ~A300;
  assign \new_[59351]_  = \new_[59350]_  & \new_[59347]_ ;
  assign \new_[59352]_  = \new_[59351]_  & \new_[59344]_ ;
  assign \new_[59356]_  = A167 & A168;
  assign \new_[59357]_  = ~A170 & \new_[59356]_ ;
  assign \new_[59360]_  = ~A199 & ~A166;
  assign \new_[59363]_  = A201 & A200;
  assign \new_[59364]_  = \new_[59363]_  & \new_[59360]_ ;
  assign \new_[59365]_  = \new_[59364]_  & \new_[59357]_ ;
  assign \new_[59369]_  = A266 & ~A265;
  assign \new_[59370]_  = A203 & \new_[59369]_ ;
  assign \new_[59373]_  = A268 & A267;
  assign \new_[59376]_  = A299 & A298;
  assign \new_[59377]_  = \new_[59376]_  & \new_[59373]_ ;
  assign \new_[59378]_  = \new_[59377]_  & \new_[59370]_ ;
  assign \new_[59382]_  = A167 & A168;
  assign \new_[59383]_  = ~A170 & \new_[59382]_ ;
  assign \new_[59386]_  = ~A199 & ~A166;
  assign \new_[59389]_  = A201 & A200;
  assign \new_[59390]_  = \new_[59389]_  & \new_[59386]_ ;
  assign \new_[59391]_  = \new_[59390]_  & \new_[59383]_ ;
  assign \new_[59395]_  = A266 & ~A265;
  assign \new_[59396]_  = A203 & \new_[59395]_ ;
  assign \new_[59399]_  = A268 & A267;
  assign \new_[59402]_  = ~A299 & ~A298;
  assign \new_[59403]_  = \new_[59402]_  & \new_[59399]_ ;
  assign \new_[59404]_  = \new_[59403]_  & \new_[59396]_ ;
  assign \new_[59408]_  = A167 & A168;
  assign \new_[59409]_  = ~A170 & \new_[59408]_ ;
  assign \new_[59412]_  = ~A199 & ~A166;
  assign \new_[59415]_  = A201 & A200;
  assign \new_[59416]_  = \new_[59415]_  & \new_[59412]_ ;
  assign \new_[59417]_  = \new_[59416]_  & \new_[59409]_ ;
  assign \new_[59421]_  = A266 & ~A265;
  assign \new_[59422]_  = A203 & \new_[59421]_ ;
  assign \new_[59425]_  = A269 & A267;
  assign \new_[59428]_  = A301 & ~A300;
  assign \new_[59429]_  = \new_[59428]_  & \new_[59425]_ ;
  assign \new_[59430]_  = \new_[59429]_  & \new_[59422]_ ;
  assign \new_[59434]_  = A167 & A168;
  assign \new_[59435]_  = ~A170 & \new_[59434]_ ;
  assign \new_[59438]_  = ~A199 & ~A166;
  assign \new_[59441]_  = A201 & A200;
  assign \new_[59442]_  = \new_[59441]_  & \new_[59438]_ ;
  assign \new_[59443]_  = \new_[59442]_  & \new_[59435]_ ;
  assign \new_[59447]_  = A266 & ~A265;
  assign \new_[59448]_  = A203 & \new_[59447]_ ;
  assign \new_[59451]_  = A269 & A267;
  assign \new_[59454]_  = A302 & ~A300;
  assign \new_[59455]_  = \new_[59454]_  & \new_[59451]_ ;
  assign \new_[59456]_  = \new_[59455]_  & \new_[59448]_ ;
  assign \new_[59460]_  = A167 & A168;
  assign \new_[59461]_  = ~A170 & \new_[59460]_ ;
  assign \new_[59464]_  = ~A199 & ~A166;
  assign \new_[59467]_  = A201 & A200;
  assign \new_[59468]_  = \new_[59467]_  & \new_[59464]_ ;
  assign \new_[59469]_  = \new_[59468]_  & \new_[59461]_ ;
  assign \new_[59473]_  = A266 & ~A265;
  assign \new_[59474]_  = A203 & \new_[59473]_ ;
  assign \new_[59477]_  = A269 & A267;
  assign \new_[59480]_  = A299 & A298;
  assign \new_[59481]_  = \new_[59480]_  & \new_[59477]_ ;
  assign \new_[59482]_  = \new_[59481]_  & \new_[59474]_ ;
  assign \new_[59486]_  = A167 & A168;
  assign \new_[59487]_  = ~A170 & \new_[59486]_ ;
  assign \new_[59490]_  = ~A199 & ~A166;
  assign \new_[59493]_  = A201 & A200;
  assign \new_[59494]_  = \new_[59493]_  & \new_[59490]_ ;
  assign \new_[59495]_  = \new_[59494]_  & \new_[59487]_ ;
  assign \new_[59499]_  = A266 & ~A265;
  assign \new_[59500]_  = A203 & \new_[59499]_ ;
  assign \new_[59503]_  = A269 & A267;
  assign \new_[59506]_  = ~A299 & ~A298;
  assign \new_[59507]_  = \new_[59506]_  & \new_[59503]_ ;
  assign \new_[59508]_  = \new_[59507]_  & \new_[59500]_ ;
  assign \new_[59512]_  = A167 & A168;
  assign \new_[59513]_  = ~A170 & \new_[59512]_ ;
  assign \new_[59516]_  = ~A199 & ~A166;
  assign \new_[59519]_  = A201 & A200;
  assign \new_[59520]_  = \new_[59519]_  & \new_[59516]_ ;
  assign \new_[59521]_  = \new_[59520]_  & \new_[59513]_ ;
  assign \new_[59525]_  = ~A266 & A265;
  assign \new_[59526]_  = A203 & \new_[59525]_ ;
  assign \new_[59529]_  = A268 & A267;
  assign \new_[59532]_  = A301 & ~A300;
  assign \new_[59533]_  = \new_[59532]_  & \new_[59529]_ ;
  assign \new_[59534]_  = \new_[59533]_  & \new_[59526]_ ;
  assign \new_[59538]_  = A167 & A168;
  assign \new_[59539]_  = ~A170 & \new_[59538]_ ;
  assign \new_[59542]_  = ~A199 & ~A166;
  assign \new_[59545]_  = A201 & A200;
  assign \new_[59546]_  = \new_[59545]_  & \new_[59542]_ ;
  assign \new_[59547]_  = \new_[59546]_  & \new_[59539]_ ;
  assign \new_[59551]_  = ~A266 & A265;
  assign \new_[59552]_  = A203 & \new_[59551]_ ;
  assign \new_[59555]_  = A268 & A267;
  assign \new_[59558]_  = A302 & ~A300;
  assign \new_[59559]_  = \new_[59558]_  & \new_[59555]_ ;
  assign \new_[59560]_  = \new_[59559]_  & \new_[59552]_ ;
  assign \new_[59564]_  = A167 & A168;
  assign \new_[59565]_  = ~A170 & \new_[59564]_ ;
  assign \new_[59568]_  = ~A199 & ~A166;
  assign \new_[59571]_  = A201 & A200;
  assign \new_[59572]_  = \new_[59571]_  & \new_[59568]_ ;
  assign \new_[59573]_  = \new_[59572]_  & \new_[59565]_ ;
  assign \new_[59577]_  = ~A266 & A265;
  assign \new_[59578]_  = A203 & \new_[59577]_ ;
  assign \new_[59581]_  = A268 & A267;
  assign \new_[59584]_  = A299 & A298;
  assign \new_[59585]_  = \new_[59584]_  & \new_[59581]_ ;
  assign \new_[59586]_  = \new_[59585]_  & \new_[59578]_ ;
  assign \new_[59590]_  = A167 & A168;
  assign \new_[59591]_  = ~A170 & \new_[59590]_ ;
  assign \new_[59594]_  = ~A199 & ~A166;
  assign \new_[59597]_  = A201 & A200;
  assign \new_[59598]_  = \new_[59597]_  & \new_[59594]_ ;
  assign \new_[59599]_  = \new_[59598]_  & \new_[59591]_ ;
  assign \new_[59603]_  = ~A266 & A265;
  assign \new_[59604]_  = A203 & \new_[59603]_ ;
  assign \new_[59607]_  = A268 & A267;
  assign \new_[59610]_  = ~A299 & ~A298;
  assign \new_[59611]_  = \new_[59610]_  & \new_[59607]_ ;
  assign \new_[59612]_  = \new_[59611]_  & \new_[59604]_ ;
  assign \new_[59616]_  = A167 & A168;
  assign \new_[59617]_  = ~A170 & \new_[59616]_ ;
  assign \new_[59620]_  = ~A199 & ~A166;
  assign \new_[59623]_  = A201 & A200;
  assign \new_[59624]_  = \new_[59623]_  & \new_[59620]_ ;
  assign \new_[59625]_  = \new_[59624]_  & \new_[59617]_ ;
  assign \new_[59629]_  = ~A266 & A265;
  assign \new_[59630]_  = A203 & \new_[59629]_ ;
  assign \new_[59633]_  = A269 & A267;
  assign \new_[59636]_  = A301 & ~A300;
  assign \new_[59637]_  = \new_[59636]_  & \new_[59633]_ ;
  assign \new_[59638]_  = \new_[59637]_  & \new_[59630]_ ;
  assign \new_[59642]_  = A167 & A168;
  assign \new_[59643]_  = ~A170 & \new_[59642]_ ;
  assign \new_[59646]_  = ~A199 & ~A166;
  assign \new_[59649]_  = A201 & A200;
  assign \new_[59650]_  = \new_[59649]_  & \new_[59646]_ ;
  assign \new_[59651]_  = \new_[59650]_  & \new_[59643]_ ;
  assign \new_[59655]_  = ~A266 & A265;
  assign \new_[59656]_  = A203 & \new_[59655]_ ;
  assign \new_[59659]_  = A269 & A267;
  assign \new_[59662]_  = A302 & ~A300;
  assign \new_[59663]_  = \new_[59662]_  & \new_[59659]_ ;
  assign \new_[59664]_  = \new_[59663]_  & \new_[59656]_ ;
  assign \new_[59668]_  = A167 & A168;
  assign \new_[59669]_  = ~A170 & \new_[59668]_ ;
  assign \new_[59672]_  = ~A199 & ~A166;
  assign \new_[59675]_  = A201 & A200;
  assign \new_[59676]_  = \new_[59675]_  & \new_[59672]_ ;
  assign \new_[59677]_  = \new_[59676]_  & \new_[59669]_ ;
  assign \new_[59681]_  = ~A266 & A265;
  assign \new_[59682]_  = A203 & \new_[59681]_ ;
  assign \new_[59685]_  = A269 & A267;
  assign \new_[59688]_  = A299 & A298;
  assign \new_[59689]_  = \new_[59688]_  & \new_[59685]_ ;
  assign \new_[59690]_  = \new_[59689]_  & \new_[59682]_ ;
  assign \new_[59694]_  = A167 & A168;
  assign \new_[59695]_  = ~A170 & \new_[59694]_ ;
  assign \new_[59698]_  = ~A199 & ~A166;
  assign \new_[59701]_  = A201 & A200;
  assign \new_[59702]_  = \new_[59701]_  & \new_[59698]_ ;
  assign \new_[59703]_  = \new_[59702]_  & \new_[59695]_ ;
  assign \new_[59707]_  = ~A266 & A265;
  assign \new_[59708]_  = A203 & \new_[59707]_ ;
  assign \new_[59711]_  = A269 & A267;
  assign \new_[59714]_  = ~A299 & ~A298;
  assign \new_[59715]_  = \new_[59714]_  & \new_[59711]_ ;
  assign \new_[59716]_  = \new_[59715]_  & \new_[59708]_ ;
  assign \new_[59720]_  = A167 & A168;
  assign \new_[59721]_  = ~A170 & \new_[59720]_ ;
  assign \new_[59724]_  = A199 & ~A166;
  assign \new_[59727]_  = A201 & ~A200;
  assign \new_[59728]_  = \new_[59727]_  & \new_[59724]_ ;
  assign \new_[59729]_  = \new_[59728]_  & \new_[59721]_ ;
  assign \new_[59733]_  = A266 & ~A265;
  assign \new_[59734]_  = A202 & \new_[59733]_ ;
  assign \new_[59737]_  = A268 & A267;
  assign \new_[59740]_  = A301 & ~A300;
  assign \new_[59741]_  = \new_[59740]_  & \new_[59737]_ ;
  assign \new_[59742]_  = \new_[59741]_  & \new_[59734]_ ;
  assign \new_[59746]_  = A167 & A168;
  assign \new_[59747]_  = ~A170 & \new_[59746]_ ;
  assign \new_[59750]_  = A199 & ~A166;
  assign \new_[59753]_  = A201 & ~A200;
  assign \new_[59754]_  = \new_[59753]_  & \new_[59750]_ ;
  assign \new_[59755]_  = \new_[59754]_  & \new_[59747]_ ;
  assign \new_[59759]_  = A266 & ~A265;
  assign \new_[59760]_  = A202 & \new_[59759]_ ;
  assign \new_[59763]_  = A268 & A267;
  assign \new_[59766]_  = A302 & ~A300;
  assign \new_[59767]_  = \new_[59766]_  & \new_[59763]_ ;
  assign \new_[59768]_  = \new_[59767]_  & \new_[59760]_ ;
  assign \new_[59772]_  = A167 & A168;
  assign \new_[59773]_  = ~A170 & \new_[59772]_ ;
  assign \new_[59776]_  = A199 & ~A166;
  assign \new_[59779]_  = A201 & ~A200;
  assign \new_[59780]_  = \new_[59779]_  & \new_[59776]_ ;
  assign \new_[59781]_  = \new_[59780]_  & \new_[59773]_ ;
  assign \new_[59785]_  = A266 & ~A265;
  assign \new_[59786]_  = A202 & \new_[59785]_ ;
  assign \new_[59789]_  = A268 & A267;
  assign \new_[59792]_  = A299 & A298;
  assign \new_[59793]_  = \new_[59792]_  & \new_[59789]_ ;
  assign \new_[59794]_  = \new_[59793]_  & \new_[59786]_ ;
  assign \new_[59798]_  = A167 & A168;
  assign \new_[59799]_  = ~A170 & \new_[59798]_ ;
  assign \new_[59802]_  = A199 & ~A166;
  assign \new_[59805]_  = A201 & ~A200;
  assign \new_[59806]_  = \new_[59805]_  & \new_[59802]_ ;
  assign \new_[59807]_  = \new_[59806]_  & \new_[59799]_ ;
  assign \new_[59811]_  = A266 & ~A265;
  assign \new_[59812]_  = A202 & \new_[59811]_ ;
  assign \new_[59815]_  = A268 & A267;
  assign \new_[59818]_  = ~A299 & ~A298;
  assign \new_[59819]_  = \new_[59818]_  & \new_[59815]_ ;
  assign \new_[59820]_  = \new_[59819]_  & \new_[59812]_ ;
  assign \new_[59824]_  = A167 & A168;
  assign \new_[59825]_  = ~A170 & \new_[59824]_ ;
  assign \new_[59828]_  = A199 & ~A166;
  assign \new_[59831]_  = A201 & ~A200;
  assign \new_[59832]_  = \new_[59831]_  & \new_[59828]_ ;
  assign \new_[59833]_  = \new_[59832]_  & \new_[59825]_ ;
  assign \new_[59837]_  = A266 & ~A265;
  assign \new_[59838]_  = A202 & \new_[59837]_ ;
  assign \new_[59841]_  = A269 & A267;
  assign \new_[59844]_  = A301 & ~A300;
  assign \new_[59845]_  = \new_[59844]_  & \new_[59841]_ ;
  assign \new_[59846]_  = \new_[59845]_  & \new_[59838]_ ;
  assign \new_[59850]_  = A167 & A168;
  assign \new_[59851]_  = ~A170 & \new_[59850]_ ;
  assign \new_[59854]_  = A199 & ~A166;
  assign \new_[59857]_  = A201 & ~A200;
  assign \new_[59858]_  = \new_[59857]_  & \new_[59854]_ ;
  assign \new_[59859]_  = \new_[59858]_  & \new_[59851]_ ;
  assign \new_[59863]_  = A266 & ~A265;
  assign \new_[59864]_  = A202 & \new_[59863]_ ;
  assign \new_[59867]_  = A269 & A267;
  assign \new_[59870]_  = A302 & ~A300;
  assign \new_[59871]_  = \new_[59870]_  & \new_[59867]_ ;
  assign \new_[59872]_  = \new_[59871]_  & \new_[59864]_ ;
  assign \new_[59876]_  = A167 & A168;
  assign \new_[59877]_  = ~A170 & \new_[59876]_ ;
  assign \new_[59880]_  = A199 & ~A166;
  assign \new_[59883]_  = A201 & ~A200;
  assign \new_[59884]_  = \new_[59883]_  & \new_[59880]_ ;
  assign \new_[59885]_  = \new_[59884]_  & \new_[59877]_ ;
  assign \new_[59889]_  = A266 & ~A265;
  assign \new_[59890]_  = A202 & \new_[59889]_ ;
  assign \new_[59893]_  = A269 & A267;
  assign \new_[59896]_  = A299 & A298;
  assign \new_[59897]_  = \new_[59896]_  & \new_[59893]_ ;
  assign \new_[59898]_  = \new_[59897]_  & \new_[59890]_ ;
  assign \new_[59902]_  = A167 & A168;
  assign \new_[59903]_  = ~A170 & \new_[59902]_ ;
  assign \new_[59906]_  = A199 & ~A166;
  assign \new_[59909]_  = A201 & ~A200;
  assign \new_[59910]_  = \new_[59909]_  & \new_[59906]_ ;
  assign \new_[59911]_  = \new_[59910]_  & \new_[59903]_ ;
  assign \new_[59915]_  = A266 & ~A265;
  assign \new_[59916]_  = A202 & \new_[59915]_ ;
  assign \new_[59919]_  = A269 & A267;
  assign \new_[59922]_  = ~A299 & ~A298;
  assign \new_[59923]_  = \new_[59922]_  & \new_[59919]_ ;
  assign \new_[59924]_  = \new_[59923]_  & \new_[59916]_ ;
  assign \new_[59928]_  = A167 & A168;
  assign \new_[59929]_  = ~A170 & \new_[59928]_ ;
  assign \new_[59932]_  = A199 & ~A166;
  assign \new_[59935]_  = A201 & ~A200;
  assign \new_[59936]_  = \new_[59935]_  & \new_[59932]_ ;
  assign \new_[59937]_  = \new_[59936]_  & \new_[59929]_ ;
  assign \new_[59941]_  = ~A266 & A265;
  assign \new_[59942]_  = A202 & \new_[59941]_ ;
  assign \new_[59945]_  = A268 & A267;
  assign \new_[59948]_  = A301 & ~A300;
  assign \new_[59949]_  = \new_[59948]_  & \new_[59945]_ ;
  assign \new_[59950]_  = \new_[59949]_  & \new_[59942]_ ;
  assign \new_[59954]_  = A167 & A168;
  assign \new_[59955]_  = ~A170 & \new_[59954]_ ;
  assign \new_[59958]_  = A199 & ~A166;
  assign \new_[59961]_  = A201 & ~A200;
  assign \new_[59962]_  = \new_[59961]_  & \new_[59958]_ ;
  assign \new_[59963]_  = \new_[59962]_  & \new_[59955]_ ;
  assign \new_[59967]_  = ~A266 & A265;
  assign \new_[59968]_  = A202 & \new_[59967]_ ;
  assign \new_[59971]_  = A268 & A267;
  assign \new_[59974]_  = A302 & ~A300;
  assign \new_[59975]_  = \new_[59974]_  & \new_[59971]_ ;
  assign \new_[59976]_  = \new_[59975]_  & \new_[59968]_ ;
  assign \new_[59980]_  = A167 & A168;
  assign \new_[59981]_  = ~A170 & \new_[59980]_ ;
  assign \new_[59984]_  = A199 & ~A166;
  assign \new_[59987]_  = A201 & ~A200;
  assign \new_[59988]_  = \new_[59987]_  & \new_[59984]_ ;
  assign \new_[59989]_  = \new_[59988]_  & \new_[59981]_ ;
  assign \new_[59993]_  = ~A266 & A265;
  assign \new_[59994]_  = A202 & \new_[59993]_ ;
  assign \new_[59997]_  = A268 & A267;
  assign \new_[60000]_  = A299 & A298;
  assign \new_[60001]_  = \new_[60000]_  & \new_[59997]_ ;
  assign \new_[60002]_  = \new_[60001]_  & \new_[59994]_ ;
  assign \new_[60006]_  = A167 & A168;
  assign \new_[60007]_  = ~A170 & \new_[60006]_ ;
  assign \new_[60010]_  = A199 & ~A166;
  assign \new_[60013]_  = A201 & ~A200;
  assign \new_[60014]_  = \new_[60013]_  & \new_[60010]_ ;
  assign \new_[60015]_  = \new_[60014]_  & \new_[60007]_ ;
  assign \new_[60019]_  = ~A266 & A265;
  assign \new_[60020]_  = A202 & \new_[60019]_ ;
  assign \new_[60023]_  = A268 & A267;
  assign \new_[60026]_  = ~A299 & ~A298;
  assign \new_[60027]_  = \new_[60026]_  & \new_[60023]_ ;
  assign \new_[60028]_  = \new_[60027]_  & \new_[60020]_ ;
  assign \new_[60032]_  = A167 & A168;
  assign \new_[60033]_  = ~A170 & \new_[60032]_ ;
  assign \new_[60036]_  = A199 & ~A166;
  assign \new_[60039]_  = A201 & ~A200;
  assign \new_[60040]_  = \new_[60039]_  & \new_[60036]_ ;
  assign \new_[60041]_  = \new_[60040]_  & \new_[60033]_ ;
  assign \new_[60045]_  = ~A266 & A265;
  assign \new_[60046]_  = A202 & \new_[60045]_ ;
  assign \new_[60049]_  = A269 & A267;
  assign \new_[60052]_  = A301 & ~A300;
  assign \new_[60053]_  = \new_[60052]_  & \new_[60049]_ ;
  assign \new_[60054]_  = \new_[60053]_  & \new_[60046]_ ;
  assign \new_[60058]_  = A167 & A168;
  assign \new_[60059]_  = ~A170 & \new_[60058]_ ;
  assign \new_[60062]_  = A199 & ~A166;
  assign \new_[60065]_  = A201 & ~A200;
  assign \new_[60066]_  = \new_[60065]_  & \new_[60062]_ ;
  assign \new_[60067]_  = \new_[60066]_  & \new_[60059]_ ;
  assign \new_[60071]_  = ~A266 & A265;
  assign \new_[60072]_  = A202 & \new_[60071]_ ;
  assign \new_[60075]_  = A269 & A267;
  assign \new_[60078]_  = A302 & ~A300;
  assign \new_[60079]_  = \new_[60078]_  & \new_[60075]_ ;
  assign \new_[60080]_  = \new_[60079]_  & \new_[60072]_ ;
  assign \new_[60084]_  = A167 & A168;
  assign \new_[60085]_  = ~A170 & \new_[60084]_ ;
  assign \new_[60088]_  = A199 & ~A166;
  assign \new_[60091]_  = A201 & ~A200;
  assign \new_[60092]_  = \new_[60091]_  & \new_[60088]_ ;
  assign \new_[60093]_  = \new_[60092]_  & \new_[60085]_ ;
  assign \new_[60097]_  = ~A266 & A265;
  assign \new_[60098]_  = A202 & \new_[60097]_ ;
  assign \new_[60101]_  = A269 & A267;
  assign \new_[60104]_  = A299 & A298;
  assign \new_[60105]_  = \new_[60104]_  & \new_[60101]_ ;
  assign \new_[60106]_  = \new_[60105]_  & \new_[60098]_ ;
  assign \new_[60110]_  = A167 & A168;
  assign \new_[60111]_  = ~A170 & \new_[60110]_ ;
  assign \new_[60114]_  = A199 & ~A166;
  assign \new_[60117]_  = A201 & ~A200;
  assign \new_[60118]_  = \new_[60117]_  & \new_[60114]_ ;
  assign \new_[60119]_  = \new_[60118]_  & \new_[60111]_ ;
  assign \new_[60123]_  = ~A266 & A265;
  assign \new_[60124]_  = A202 & \new_[60123]_ ;
  assign \new_[60127]_  = A269 & A267;
  assign \new_[60130]_  = ~A299 & ~A298;
  assign \new_[60131]_  = \new_[60130]_  & \new_[60127]_ ;
  assign \new_[60132]_  = \new_[60131]_  & \new_[60124]_ ;
  assign \new_[60136]_  = A167 & A168;
  assign \new_[60137]_  = ~A170 & \new_[60136]_ ;
  assign \new_[60140]_  = A199 & ~A166;
  assign \new_[60143]_  = A201 & ~A200;
  assign \new_[60144]_  = \new_[60143]_  & \new_[60140]_ ;
  assign \new_[60145]_  = \new_[60144]_  & \new_[60137]_ ;
  assign \new_[60149]_  = A266 & ~A265;
  assign \new_[60150]_  = A203 & \new_[60149]_ ;
  assign \new_[60153]_  = A268 & A267;
  assign \new_[60156]_  = A301 & ~A300;
  assign \new_[60157]_  = \new_[60156]_  & \new_[60153]_ ;
  assign \new_[60158]_  = \new_[60157]_  & \new_[60150]_ ;
  assign \new_[60162]_  = A167 & A168;
  assign \new_[60163]_  = ~A170 & \new_[60162]_ ;
  assign \new_[60166]_  = A199 & ~A166;
  assign \new_[60169]_  = A201 & ~A200;
  assign \new_[60170]_  = \new_[60169]_  & \new_[60166]_ ;
  assign \new_[60171]_  = \new_[60170]_  & \new_[60163]_ ;
  assign \new_[60175]_  = A266 & ~A265;
  assign \new_[60176]_  = A203 & \new_[60175]_ ;
  assign \new_[60179]_  = A268 & A267;
  assign \new_[60182]_  = A302 & ~A300;
  assign \new_[60183]_  = \new_[60182]_  & \new_[60179]_ ;
  assign \new_[60184]_  = \new_[60183]_  & \new_[60176]_ ;
  assign \new_[60188]_  = A167 & A168;
  assign \new_[60189]_  = ~A170 & \new_[60188]_ ;
  assign \new_[60192]_  = A199 & ~A166;
  assign \new_[60195]_  = A201 & ~A200;
  assign \new_[60196]_  = \new_[60195]_  & \new_[60192]_ ;
  assign \new_[60197]_  = \new_[60196]_  & \new_[60189]_ ;
  assign \new_[60201]_  = A266 & ~A265;
  assign \new_[60202]_  = A203 & \new_[60201]_ ;
  assign \new_[60205]_  = A268 & A267;
  assign \new_[60208]_  = A299 & A298;
  assign \new_[60209]_  = \new_[60208]_  & \new_[60205]_ ;
  assign \new_[60210]_  = \new_[60209]_  & \new_[60202]_ ;
  assign \new_[60214]_  = A167 & A168;
  assign \new_[60215]_  = ~A170 & \new_[60214]_ ;
  assign \new_[60218]_  = A199 & ~A166;
  assign \new_[60221]_  = A201 & ~A200;
  assign \new_[60222]_  = \new_[60221]_  & \new_[60218]_ ;
  assign \new_[60223]_  = \new_[60222]_  & \new_[60215]_ ;
  assign \new_[60227]_  = A266 & ~A265;
  assign \new_[60228]_  = A203 & \new_[60227]_ ;
  assign \new_[60231]_  = A268 & A267;
  assign \new_[60234]_  = ~A299 & ~A298;
  assign \new_[60235]_  = \new_[60234]_  & \new_[60231]_ ;
  assign \new_[60236]_  = \new_[60235]_  & \new_[60228]_ ;
  assign \new_[60240]_  = A167 & A168;
  assign \new_[60241]_  = ~A170 & \new_[60240]_ ;
  assign \new_[60244]_  = A199 & ~A166;
  assign \new_[60247]_  = A201 & ~A200;
  assign \new_[60248]_  = \new_[60247]_  & \new_[60244]_ ;
  assign \new_[60249]_  = \new_[60248]_  & \new_[60241]_ ;
  assign \new_[60253]_  = A266 & ~A265;
  assign \new_[60254]_  = A203 & \new_[60253]_ ;
  assign \new_[60257]_  = A269 & A267;
  assign \new_[60260]_  = A301 & ~A300;
  assign \new_[60261]_  = \new_[60260]_  & \new_[60257]_ ;
  assign \new_[60262]_  = \new_[60261]_  & \new_[60254]_ ;
  assign \new_[60266]_  = A167 & A168;
  assign \new_[60267]_  = ~A170 & \new_[60266]_ ;
  assign \new_[60270]_  = A199 & ~A166;
  assign \new_[60273]_  = A201 & ~A200;
  assign \new_[60274]_  = \new_[60273]_  & \new_[60270]_ ;
  assign \new_[60275]_  = \new_[60274]_  & \new_[60267]_ ;
  assign \new_[60279]_  = A266 & ~A265;
  assign \new_[60280]_  = A203 & \new_[60279]_ ;
  assign \new_[60283]_  = A269 & A267;
  assign \new_[60286]_  = A302 & ~A300;
  assign \new_[60287]_  = \new_[60286]_  & \new_[60283]_ ;
  assign \new_[60288]_  = \new_[60287]_  & \new_[60280]_ ;
  assign \new_[60292]_  = A167 & A168;
  assign \new_[60293]_  = ~A170 & \new_[60292]_ ;
  assign \new_[60296]_  = A199 & ~A166;
  assign \new_[60299]_  = A201 & ~A200;
  assign \new_[60300]_  = \new_[60299]_  & \new_[60296]_ ;
  assign \new_[60301]_  = \new_[60300]_  & \new_[60293]_ ;
  assign \new_[60305]_  = A266 & ~A265;
  assign \new_[60306]_  = A203 & \new_[60305]_ ;
  assign \new_[60309]_  = A269 & A267;
  assign \new_[60312]_  = A299 & A298;
  assign \new_[60313]_  = \new_[60312]_  & \new_[60309]_ ;
  assign \new_[60314]_  = \new_[60313]_  & \new_[60306]_ ;
  assign \new_[60318]_  = A167 & A168;
  assign \new_[60319]_  = ~A170 & \new_[60318]_ ;
  assign \new_[60322]_  = A199 & ~A166;
  assign \new_[60325]_  = A201 & ~A200;
  assign \new_[60326]_  = \new_[60325]_  & \new_[60322]_ ;
  assign \new_[60327]_  = \new_[60326]_  & \new_[60319]_ ;
  assign \new_[60331]_  = A266 & ~A265;
  assign \new_[60332]_  = A203 & \new_[60331]_ ;
  assign \new_[60335]_  = A269 & A267;
  assign \new_[60338]_  = ~A299 & ~A298;
  assign \new_[60339]_  = \new_[60338]_  & \new_[60335]_ ;
  assign \new_[60340]_  = \new_[60339]_  & \new_[60332]_ ;
  assign \new_[60344]_  = A167 & A168;
  assign \new_[60345]_  = ~A170 & \new_[60344]_ ;
  assign \new_[60348]_  = A199 & ~A166;
  assign \new_[60351]_  = A201 & ~A200;
  assign \new_[60352]_  = \new_[60351]_  & \new_[60348]_ ;
  assign \new_[60353]_  = \new_[60352]_  & \new_[60345]_ ;
  assign \new_[60357]_  = ~A266 & A265;
  assign \new_[60358]_  = A203 & \new_[60357]_ ;
  assign \new_[60361]_  = A268 & A267;
  assign \new_[60364]_  = A301 & ~A300;
  assign \new_[60365]_  = \new_[60364]_  & \new_[60361]_ ;
  assign \new_[60366]_  = \new_[60365]_  & \new_[60358]_ ;
  assign \new_[60370]_  = A167 & A168;
  assign \new_[60371]_  = ~A170 & \new_[60370]_ ;
  assign \new_[60374]_  = A199 & ~A166;
  assign \new_[60377]_  = A201 & ~A200;
  assign \new_[60378]_  = \new_[60377]_  & \new_[60374]_ ;
  assign \new_[60379]_  = \new_[60378]_  & \new_[60371]_ ;
  assign \new_[60383]_  = ~A266 & A265;
  assign \new_[60384]_  = A203 & \new_[60383]_ ;
  assign \new_[60387]_  = A268 & A267;
  assign \new_[60390]_  = A302 & ~A300;
  assign \new_[60391]_  = \new_[60390]_  & \new_[60387]_ ;
  assign \new_[60392]_  = \new_[60391]_  & \new_[60384]_ ;
  assign \new_[60396]_  = A167 & A168;
  assign \new_[60397]_  = ~A170 & \new_[60396]_ ;
  assign \new_[60400]_  = A199 & ~A166;
  assign \new_[60403]_  = A201 & ~A200;
  assign \new_[60404]_  = \new_[60403]_  & \new_[60400]_ ;
  assign \new_[60405]_  = \new_[60404]_  & \new_[60397]_ ;
  assign \new_[60409]_  = ~A266 & A265;
  assign \new_[60410]_  = A203 & \new_[60409]_ ;
  assign \new_[60413]_  = A268 & A267;
  assign \new_[60416]_  = A299 & A298;
  assign \new_[60417]_  = \new_[60416]_  & \new_[60413]_ ;
  assign \new_[60418]_  = \new_[60417]_  & \new_[60410]_ ;
  assign \new_[60422]_  = A167 & A168;
  assign \new_[60423]_  = ~A170 & \new_[60422]_ ;
  assign \new_[60426]_  = A199 & ~A166;
  assign \new_[60429]_  = A201 & ~A200;
  assign \new_[60430]_  = \new_[60429]_  & \new_[60426]_ ;
  assign \new_[60431]_  = \new_[60430]_  & \new_[60423]_ ;
  assign \new_[60435]_  = ~A266 & A265;
  assign \new_[60436]_  = A203 & \new_[60435]_ ;
  assign \new_[60439]_  = A268 & A267;
  assign \new_[60442]_  = ~A299 & ~A298;
  assign \new_[60443]_  = \new_[60442]_  & \new_[60439]_ ;
  assign \new_[60444]_  = \new_[60443]_  & \new_[60436]_ ;
  assign \new_[60448]_  = A167 & A168;
  assign \new_[60449]_  = ~A170 & \new_[60448]_ ;
  assign \new_[60452]_  = A199 & ~A166;
  assign \new_[60455]_  = A201 & ~A200;
  assign \new_[60456]_  = \new_[60455]_  & \new_[60452]_ ;
  assign \new_[60457]_  = \new_[60456]_  & \new_[60449]_ ;
  assign \new_[60461]_  = ~A266 & A265;
  assign \new_[60462]_  = A203 & \new_[60461]_ ;
  assign \new_[60465]_  = A269 & A267;
  assign \new_[60468]_  = A301 & ~A300;
  assign \new_[60469]_  = \new_[60468]_  & \new_[60465]_ ;
  assign \new_[60470]_  = \new_[60469]_  & \new_[60462]_ ;
  assign \new_[60474]_  = A167 & A168;
  assign \new_[60475]_  = ~A170 & \new_[60474]_ ;
  assign \new_[60478]_  = A199 & ~A166;
  assign \new_[60481]_  = A201 & ~A200;
  assign \new_[60482]_  = \new_[60481]_  & \new_[60478]_ ;
  assign \new_[60483]_  = \new_[60482]_  & \new_[60475]_ ;
  assign \new_[60487]_  = ~A266 & A265;
  assign \new_[60488]_  = A203 & \new_[60487]_ ;
  assign \new_[60491]_  = A269 & A267;
  assign \new_[60494]_  = A302 & ~A300;
  assign \new_[60495]_  = \new_[60494]_  & \new_[60491]_ ;
  assign \new_[60496]_  = \new_[60495]_  & \new_[60488]_ ;
  assign \new_[60500]_  = A167 & A168;
  assign \new_[60501]_  = ~A170 & \new_[60500]_ ;
  assign \new_[60504]_  = A199 & ~A166;
  assign \new_[60507]_  = A201 & ~A200;
  assign \new_[60508]_  = \new_[60507]_  & \new_[60504]_ ;
  assign \new_[60509]_  = \new_[60508]_  & \new_[60501]_ ;
  assign \new_[60513]_  = ~A266 & A265;
  assign \new_[60514]_  = A203 & \new_[60513]_ ;
  assign \new_[60517]_  = A269 & A267;
  assign \new_[60520]_  = A299 & A298;
  assign \new_[60521]_  = \new_[60520]_  & \new_[60517]_ ;
  assign \new_[60522]_  = \new_[60521]_  & \new_[60514]_ ;
  assign \new_[60526]_  = A167 & A168;
  assign \new_[60527]_  = ~A170 & \new_[60526]_ ;
  assign \new_[60530]_  = A199 & ~A166;
  assign \new_[60533]_  = A201 & ~A200;
  assign \new_[60534]_  = \new_[60533]_  & \new_[60530]_ ;
  assign \new_[60535]_  = \new_[60534]_  & \new_[60527]_ ;
  assign \new_[60539]_  = ~A266 & A265;
  assign \new_[60540]_  = A203 & \new_[60539]_ ;
  assign \new_[60543]_  = A269 & A267;
  assign \new_[60546]_  = ~A299 & ~A298;
  assign \new_[60547]_  = \new_[60546]_  & \new_[60543]_ ;
  assign \new_[60548]_  = \new_[60547]_  & \new_[60540]_ ;
  assign \new_[60552]_  = A167 & A168;
  assign \new_[60553]_  = ~A170 & \new_[60552]_ ;
  assign \new_[60556]_  = ~A199 & ~A166;
  assign \new_[60559]_  = A267 & ~A200;
  assign \new_[60560]_  = \new_[60559]_  & \new_[60556]_ ;
  assign \new_[60561]_  = \new_[60560]_  & \new_[60553]_ ;
  assign \new_[60565]_  = A298 & ~A269;
  assign \new_[60566]_  = ~A268 & \new_[60565]_ ;
  assign \new_[60569]_  = ~A300 & ~A299;
  assign \new_[60572]_  = ~A302 & ~A301;
  assign \new_[60573]_  = \new_[60572]_  & \new_[60569]_ ;
  assign \new_[60574]_  = \new_[60573]_  & \new_[60566]_ ;
  assign \new_[60578]_  = A167 & A168;
  assign \new_[60579]_  = ~A170 & \new_[60578]_ ;
  assign \new_[60582]_  = ~A199 & ~A166;
  assign \new_[60585]_  = A267 & ~A200;
  assign \new_[60586]_  = \new_[60585]_  & \new_[60582]_ ;
  assign \new_[60587]_  = \new_[60586]_  & \new_[60579]_ ;
  assign \new_[60591]_  = ~A298 & ~A269;
  assign \new_[60592]_  = ~A268 & \new_[60591]_ ;
  assign \new_[60595]_  = ~A300 & A299;
  assign \new_[60598]_  = ~A302 & ~A301;
  assign \new_[60599]_  = \new_[60598]_  & \new_[60595]_ ;
  assign \new_[60600]_  = \new_[60599]_  & \new_[60592]_ ;
  assign \new_[60604]_  = ~A167 & A168;
  assign \new_[60605]_  = ~A170 & \new_[60604]_ ;
  assign \new_[60608]_  = A201 & A166;
  assign \new_[60611]_  = ~A203 & ~A202;
  assign \new_[60612]_  = \new_[60611]_  & \new_[60608]_ ;
  assign \new_[60613]_  = \new_[60612]_  & \new_[60605]_ ;
  assign \new_[60617]_  = ~A269 & ~A268;
  assign \new_[60618]_  = A267 & \new_[60617]_ ;
  assign \new_[60621]_  = ~A299 & A298;
  assign \new_[60624]_  = A301 & A300;
  assign \new_[60625]_  = \new_[60624]_  & \new_[60621]_ ;
  assign \new_[60626]_  = \new_[60625]_  & \new_[60618]_ ;
  assign \new_[60630]_  = ~A167 & A168;
  assign \new_[60631]_  = ~A170 & \new_[60630]_ ;
  assign \new_[60634]_  = A201 & A166;
  assign \new_[60637]_  = ~A203 & ~A202;
  assign \new_[60638]_  = \new_[60637]_  & \new_[60634]_ ;
  assign \new_[60639]_  = \new_[60638]_  & \new_[60631]_ ;
  assign \new_[60643]_  = ~A269 & ~A268;
  assign \new_[60644]_  = A267 & \new_[60643]_ ;
  assign \new_[60647]_  = ~A299 & A298;
  assign \new_[60650]_  = A302 & A300;
  assign \new_[60651]_  = \new_[60650]_  & \new_[60647]_ ;
  assign \new_[60652]_  = \new_[60651]_  & \new_[60644]_ ;
  assign \new_[60656]_  = ~A167 & A168;
  assign \new_[60657]_  = ~A170 & \new_[60656]_ ;
  assign \new_[60660]_  = A201 & A166;
  assign \new_[60663]_  = ~A203 & ~A202;
  assign \new_[60664]_  = \new_[60663]_  & \new_[60660]_ ;
  assign \new_[60665]_  = \new_[60664]_  & \new_[60657]_ ;
  assign \new_[60669]_  = ~A269 & ~A268;
  assign \new_[60670]_  = A267 & \new_[60669]_ ;
  assign \new_[60673]_  = A299 & ~A298;
  assign \new_[60676]_  = A301 & A300;
  assign \new_[60677]_  = \new_[60676]_  & \new_[60673]_ ;
  assign \new_[60678]_  = \new_[60677]_  & \new_[60670]_ ;
  assign \new_[60682]_  = ~A167 & A168;
  assign \new_[60683]_  = ~A170 & \new_[60682]_ ;
  assign \new_[60686]_  = A201 & A166;
  assign \new_[60689]_  = ~A203 & ~A202;
  assign \new_[60690]_  = \new_[60689]_  & \new_[60686]_ ;
  assign \new_[60691]_  = \new_[60690]_  & \new_[60683]_ ;
  assign \new_[60695]_  = ~A269 & ~A268;
  assign \new_[60696]_  = A267 & \new_[60695]_ ;
  assign \new_[60699]_  = A299 & ~A298;
  assign \new_[60702]_  = A302 & A300;
  assign \new_[60703]_  = \new_[60702]_  & \new_[60699]_ ;
  assign \new_[60704]_  = \new_[60703]_  & \new_[60696]_ ;
  assign \new_[60708]_  = ~A167 & A168;
  assign \new_[60709]_  = ~A170 & \new_[60708]_ ;
  assign \new_[60712]_  = A201 & A166;
  assign \new_[60715]_  = ~A203 & ~A202;
  assign \new_[60716]_  = \new_[60715]_  & \new_[60712]_ ;
  assign \new_[60717]_  = \new_[60716]_  & \new_[60709]_ ;
  assign \new_[60721]_  = A298 & A268;
  assign \new_[60722]_  = ~A267 & \new_[60721]_ ;
  assign \new_[60725]_  = ~A300 & ~A299;
  assign \new_[60728]_  = ~A302 & ~A301;
  assign \new_[60729]_  = \new_[60728]_  & \new_[60725]_ ;
  assign \new_[60730]_  = \new_[60729]_  & \new_[60722]_ ;
  assign \new_[60734]_  = ~A167 & A168;
  assign \new_[60735]_  = ~A170 & \new_[60734]_ ;
  assign \new_[60738]_  = A201 & A166;
  assign \new_[60741]_  = ~A203 & ~A202;
  assign \new_[60742]_  = \new_[60741]_  & \new_[60738]_ ;
  assign \new_[60743]_  = \new_[60742]_  & \new_[60735]_ ;
  assign \new_[60747]_  = ~A298 & A268;
  assign \new_[60748]_  = ~A267 & \new_[60747]_ ;
  assign \new_[60751]_  = ~A300 & A299;
  assign \new_[60754]_  = ~A302 & ~A301;
  assign \new_[60755]_  = \new_[60754]_  & \new_[60751]_ ;
  assign \new_[60756]_  = \new_[60755]_  & \new_[60748]_ ;
  assign \new_[60760]_  = ~A167 & A168;
  assign \new_[60761]_  = ~A170 & \new_[60760]_ ;
  assign \new_[60764]_  = A201 & A166;
  assign \new_[60767]_  = ~A203 & ~A202;
  assign \new_[60768]_  = \new_[60767]_  & \new_[60764]_ ;
  assign \new_[60769]_  = \new_[60768]_  & \new_[60761]_ ;
  assign \new_[60773]_  = A298 & A269;
  assign \new_[60774]_  = ~A267 & \new_[60773]_ ;
  assign \new_[60777]_  = ~A300 & ~A299;
  assign \new_[60780]_  = ~A302 & ~A301;
  assign \new_[60781]_  = \new_[60780]_  & \new_[60777]_ ;
  assign \new_[60782]_  = \new_[60781]_  & \new_[60774]_ ;
  assign \new_[60786]_  = ~A167 & A168;
  assign \new_[60787]_  = ~A170 & \new_[60786]_ ;
  assign \new_[60790]_  = A201 & A166;
  assign \new_[60793]_  = ~A203 & ~A202;
  assign \new_[60794]_  = \new_[60793]_  & \new_[60790]_ ;
  assign \new_[60795]_  = \new_[60794]_  & \new_[60787]_ ;
  assign \new_[60799]_  = ~A298 & A269;
  assign \new_[60800]_  = ~A267 & \new_[60799]_ ;
  assign \new_[60803]_  = ~A300 & A299;
  assign \new_[60806]_  = ~A302 & ~A301;
  assign \new_[60807]_  = \new_[60806]_  & \new_[60803]_ ;
  assign \new_[60808]_  = \new_[60807]_  & \new_[60800]_ ;
  assign \new_[60812]_  = ~A167 & A168;
  assign \new_[60813]_  = ~A170 & \new_[60812]_ ;
  assign \new_[60816]_  = A201 & A166;
  assign \new_[60819]_  = ~A203 & ~A202;
  assign \new_[60820]_  = \new_[60819]_  & \new_[60816]_ ;
  assign \new_[60821]_  = \new_[60820]_  & \new_[60813]_ ;
  assign \new_[60825]_  = A298 & A266;
  assign \new_[60826]_  = A265 & \new_[60825]_ ;
  assign \new_[60829]_  = ~A300 & ~A299;
  assign \new_[60832]_  = ~A302 & ~A301;
  assign \new_[60833]_  = \new_[60832]_  & \new_[60829]_ ;
  assign \new_[60834]_  = \new_[60833]_  & \new_[60826]_ ;
  assign \new_[60838]_  = ~A167 & A168;
  assign \new_[60839]_  = ~A170 & \new_[60838]_ ;
  assign \new_[60842]_  = A201 & A166;
  assign \new_[60845]_  = ~A203 & ~A202;
  assign \new_[60846]_  = \new_[60845]_  & \new_[60842]_ ;
  assign \new_[60847]_  = \new_[60846]_  & \new_[60839]_ ;
  assign \new_[60851]_  = ~A298 & A266;
  assign \new_[60852]_  = A265 & \new_[60851]_ ;
  assign \new_[60855]_  = ~A300 & A299;
  assign \new_[60858]_  = ~A302 & ~A301;
  assign \new_[60859]_  = \new_[60858]_  & \new_[60855]_ ;
  assign \new_[60860]_  = \new_[60859]_  & \new_[60852]_ ;
  assign \new_[60864]_  = ~A167 & A168;
  assign \new_[60865]_  = ~A170 & \new_[60864]_ ;
  assign \new_[60868]_  = A201 & A166;
  assign \new_[60871]_  = ~A203 & ~A202;
  assign \new_[60872]_  = \new_[60871]_  & \new_[60868]_ ;
  assign \new_[60873]_  = \new_[60872]_  & \new_[60865]_ ;
  assign \new_[60877]_  = A298 & ~A266;
  assign \new_[60878]_  = ~A265 & \new_[60877]_ ;
  assign \new_[60881]_  = ~A300 & ~A299;
  assign \new_[60884]_  = ~A302 & ~A301;
  assign \new_[60885]_  = \new_[60884]_  & \new_[60881]_ ;
  assign \new_[60886]_  = \new_[60885]_  & \new_[60878]_ ;
  assign \new_[60890]_  = ~A167 & A168;
  assign \new_[60891]_  = ~A170 & \new_[60890]_ ;
  assign \new_[60894]_  = A201 & A166;
  assign \new_[60897]_  = ~A203 & ~A202;
  assign \new_[60898]_  = \new_[60897]_  & \new_[60894]_ ;
  assign \new_[60899]_  = \new_[60898]_  & \new_[60891]_ ;
  assign \new_[60903]_  = ~A298 & ~A266;
  assign \new_[60904]_  = ~A265 & \new_[60903]_ ;
  assign \new_[60907]_  = ~A300 & A299;
  assign \new_[60910]_  = ~A302 & ~A301;
  assign \new_[60911]_  = \new_[60910]_  & \new_[60907]_ ;
  assign \new_[60912]_  = \new_[60911]_  & \new_[60904]_ ;
  assign \new_[60916]_  = ~A167 & A168;
  assign \new_[60917]_  = ~A170 & \new_[60916]_ ;
  assign \new_[60920]_  = ~A201 & A166;
  assign \new_[60923]_  = A267 & A202;
  assign \new_[60924]_  = \new_[60923]_  & \new_[60920]_ ;
  assign \new_[60925]_  = \new_[60924]_  & \new_[60917]_ ;
  assign \new_[60929]_  = A298 & ~A269;
  assign \new_[60930]_  = ~A268 & \new_[60929]_ ;
  assign \new_[60933]_  = ~A300 & ~A299;
  assign \new_[60936]_  = ~A302 & ~A301;
  assign \new_[60937]_  = \new_[60936]_  & \new_[60933]_ ;
  assign \new_[60938]_  = \new_[60937]_  & \new_[60930]_ ;
  assign \new_[60942]_  = ~A167 & A168;
  assign \new_[60943]_  = ~A170 & \new_[60942]_ ;
  assign \new_[60946]_  = ~A201 & A166;
  assign \new_[60949]_  = A267 & A202;
  assign \new_[60950]_  = \new_[60949]_  & \new_[60946]_ ;
  assign \new_[60951]_  = \new_[60950]_  & \new_[60943]_ ;
  assign \new_[60955]_  = ~A298 & ~A269;
  assign \new_[60956]_  = ~A268 & \new_[60955]_ ;
  assign \new_[60959]_  = ~A300 & A299;
  assign \new_[60962]_  = ~A302 & ~A301;
  assign \new_[60963]_  = \new_[60962]_  & \new_[60959]_ ;
  assign \new_[60964]_  = \new_[60963]_  & \new_[60956]_ ;
  assign \new_[60968]_  = ~A167 & A168;
  assign \new_[60969]_  = ~A170 & \new_[60968]_ ;
  assign \new_[60972]_  = ~A201 & A166;
  assign \new_[60975]_  = A267 & A203;
  assign \new_[60976]_  = \new_[60975]_  & \new_[60972]_ ;
  assign \new_[60977]_  = \new_[60976]_  & \new_[60969]_ ;
  assign \new_[60981]_  = A298 & ~A269;
  assign \new_[60982]_  = ~A268 & \new_[60981]_ ;
  assign \new_[60985]_  = ~A300 & ~A299;
  assign \new_[60988]_  = ~A302 & ~A301;
  assign \new_[60989]_  = \new_[60988]_  & \new_[60985]_ ;
  assign \new_[60990]_  = \new_[60989]_  & \new_[60982]_ ;
  assign \new_[60994]_  = ~A167 & A168;
  assign \new_[60995]_  = ~A170 & \new_[60994]_ ;
  assign \new_[60998]_  = ~A201 & A166;
  assign \new_[61001]_  = A267 & A203;
  assign \new_[61002]_  = \new_[61001]_  & \new_[60998]_ ;
  assign \new_[61003]_  = \new_[61002]_  & \new_[60995]_ ;
  assign \new_[61007]_  = ~A298 & ~A269;
  assign \new_[61008]_  = ~A268 & \new_[61007]_ ;
  assign \new_[61011]_  = ~A300 & A299;
  assign \new_[61014]_  = ~A302 & ~A301;
  assign \new_[61015]_  = \new_[61014]_  & \new_[61011]_ ;
  assign \new_[61016]_  = \new_[61015]_  & \new_[61008]_ ;
  assign \new_[61020]_  = ~A167 & A168;
  assign \new_[61021]_  = ~A170 & \new_[61020]_ ;
  assign \new_[61024]_  = A199 & A166;
  assign \new_[61027]_  = A267 & A200;
  assign \new_[61028]_  = \new_[61027]_  & \new_[61024]_ ;
  assign \new_[61029]_  = \new_[61028]_  & \new_[61021]_ ;
  assign \new_[61033]_  = A298 & ~A269;
  assign \new_[61034]_  = ~A268 & \new_[61033]_ ;
  assign \new_[61037]_  = ~A300 & ~A299;
  assign \new_[61040]_  = ~A302 & ~A301;
  assign \new_[61041]_  = \new_[61040]_  & \new_[61037]_ ;
  assign \new_[61042]_  = \new_[61041]_  & \new_[61034]_ ;
  assign \new_[61046]_  = ~A167 & A168;
  assign \new_[61047]_  = ~A170 & \new_[61046]_ ;
  assign \new_[61050]_  = A199 & A166;
  assign \new_[61053]_  = A267 & A200;
  assign \new_[61054]_  = \new_[61053]_  & \new_[61050]_ ;
  assign \new_[61055]_  = \new_[61054]_  & \new_[61047]_ ;
  assign \new_[61059]_  = ~A298 & ~A269;
  assign \new_[61060]_  = ~A268 & \new_[61059]_ ;
  assign \new_[61063]_  = ~A300 & A299;
  assign \new_[61066]_  = ~A302 & ~A301;
  assign \new_[61067]_  = \new_[61066]_  & \new_[61063]_ ;
  assign \new_[61068]_  = \new_[61067]_  & \new_[61060]_ ;
  assign \new_[61072]_  = ~A167 & A168;
  assign \new_[61073]_  = ~A170 & \new_[61072]_ ;
  assign \new_[61076]_  = ~A199 & A166;
  assign \new_[61079]_  = A201 & A200;
  assign \new_[61080]_  = \new_[61079]_  & \new_[61076]_ ;
  assign \new_[61081]_  = \new_[61080]_  & \new_[61073]_ ;
  assign \new_[61085]_  = A266 & ~A265;
  assign \new_[61086]_  = A202 & \new_[61085]_ ;
  assign \new_[61089]_  = A268 & A267;
  assign \new_[61092]_  = A301 & ~A300;
  assign \new_[61093]_  = \new_[61092]_  & \new_[61089]_ ;
  assign \new_[61094]_  = \new_[61093]_  & \new_[61086]_ ;
  assign \new_[61098]_  = ~A167 & A168;
  assign \new_[61099]_  = ~A170 & \new_[61098]_ ;
  assign \new_[61102]_  = ~A199 & A166;
  assign \new_[61105]_  = A201 & A200;
  assign \new_[61106]_  = \new_[61105]_  & \new_[61102]_ ;
  assign \new_[61107]_  = \new_[61106]_  & \new_[61099]_ ;
  assign \new_[61111]_  = A266 & ~A265;
  assign \new_[61112]_  = A202 & \new_[61111]_ ;
  assign \new_[61115]_  = A268 & A267;
  assign \new_[61118]_  = A302 & ~A300;
  assign \new_[61119]_  = \new_[61118]_  & \new_[61115]_ ;
  assign \new_[61120]_  = \new_[61119]_  & \new_[61112]_ ;
  assign \new_[61124]_  = ~A167 & A168;
  assign \new_[61125]_  = ~A170 & \new_[61124]_ ;
  assign \new_[61128]_  = ~A199 & A166;
  assign \new_[61131]_  = A201 & A200;
  assign \new_[61132]_  = \new_[61131]_  & \new_[61128]_ ;
  assign \new_[61133]_  = \new_[61132]_  & \new_[61125]_ ;
  assign \new_[61137]_  = A266 & ~A265;
  assign \new_[61138]_  = A202 & \new_[61137]_ ;
  assign \new_[61141]_  = A268 & A267;
  assign \new_[61144]_  = A299 & A298;
  assign \new_[61145]_  = \new_[61144]_  & \new_[61141]_ ;
  assign \new_[61146]_  = \new_[61145]_  & \new_[61138]_ ;
  assign \new_[61150]_  = ~A167 & A168;
  assign \new_[61151]_  = ~A170 & \new_[61150]_ ;
  assign \new_[61154]_  = ~A199 & A166;
  assign \new_[61157]_  = A201 & A200;
  assign \new_[61158]_  = \new_[61157]_  & \new_[61154]_ ;
  assign \new_[61159]_  = \new_[61158]_  & \new_[61151]_ ;
  assign \new_[61163]_  = A266 & ~A265;
  assign \new_[61164]_  = A202 & \new_[61163]_ ;
  assign \new_[61167]_  = A268 & A267;
  assign \new_[61170]_  = ~A299 & ~A298;
  assign \new_[61171]_  = \new_[61170]_  & \new_[61167]_ ;
  assign \new_[61172]_  = \new_[61171]_  & \new_[61164]_ ;
  assign \new_[61176]_  = ~A167 & A168;
  assign \new_[61177]_  = ~A170 & \new_[61176]_ ;
  assign \new_[61180]_  = ~A199 & A166;
  assign \new_[61183]_  = A201 & A200;
  assign \new_[61184]_  = \new_[61183]_  & \new_[61180]_ ;
  assign \new_[61185]_  = \new_[61184]_  & \new_[61177]_ ;
  assign \new_[61189]_  = A266 & ~A265;
  assign \new_[61190]_  = A202 & \new_[61189]_ ;
  assign \new_[61193]_  = A269 & A267;
  assign \new_[61196]_  = A301 & ~A300;
  assign \new_[61197]_  = \new_[61196]_  & \new_[61193]_ ;
  assign \new_[61198]_  = \new_[61197]_  & \new_[61190]_ ;
  assign \new_[61202]_  = ~A167 & A168;
  assign \new_[61203]_  = ~A170 & \new_[61202]_ ;
  assign \new_[61206]_  = ~A199 & A166;
  assign \new_[61209]_  = A201 & A200;
  assign \new_[61210]_  = \new_[61209]_  & \new_[61206]_ ;
  assign \new_[61211]_  = \new_[61210]_  & \new_[61203]_ ;
  assign \new_[61215]_  = A266 & ~A265;
  assign \new_[61216]_  = A202 & \new_[61215]_ ;
  assign \new_[61219]_  = A269 & A267;
  assign \new_[61222]_  = A302 & ~A300;
  assign \new_[61223]_  = \new_[61222]_  & \new_[61219]_ ;
  assign \new_[61224]_  = \new_[61223]_  & \new_[61216]_ ;
  assign \new_[61228]_  = ~A167 & A168;
  assign \new_[61229]_  = ~A170 & \new_[61228]_ ;
  assign \new_[61232]_  = ~A199 & A166;
  assign \new_[61235]_  = A201 & A200;
  assign \new_[61236]_  = \new_[61235]_  & \new_[61232]_ ;
  assign \new_[61237]_  = \new_[61236]_  & \new_[61229]_ ;
  assign \new_[61241]_  = A266 & ~A265;
  assign \new_[61242]_  = A202 & \new_[61241]_ ;
  assign \new_[61245]_  = A269 & A267;
  assign \new_[61248]_  = A299 & A298;
  assign \new_[61249]_  = \new_[61248]_  & \new_[61245]_ ;
  assign \new_[61250]_  = \new_[61249]_  & \new_[61242]_ ;
  assign \new_[61254]_  = ~A167 & A168;
  assign \new_[61255]_  = ~A170 & \new_[61254]_ ;
  assign \new_[61258]_  = ~A199 & A166;
  assign \new_[61261]_  = A201 & A200;
  assign \new_[61262]_  = \new_[61261]_  & \new_[61258]_ ;
  assign \new_[61263]_  = \new_[61262]_  & \new_[61255]_ ;
  assign \new_[61267]_  = A266 & ~A265;
  assign \new_[61268]_  = A202 & \new_[61267]_ ;
  assign \new_[61271]_  = A269 & A267;
  assign \new_[61274]_  = ~A299 & ~A298;
  assign \new_[61275]_  = \new_[61274]_  & \new_[61271]_ ;
  assign \new_[61276]_  = \new_[61275]_  & \new_[61268]_ ;
  assign \new_[61280]_  = ~A167 & A168;
  assign \new_[61281]_  = ~A170 & \new_[61280]_ ;
  assign \new_[61284]_  = ~A199 & A166;
  assign \new_[61287]_  = A201 & A200;
  assign \new_[61288]_  = \new_[61287]_  & \new_[61284]_ ;
  assign \new_[61289]_  = \new_[61288]_  & \new_[61281]_ ;
  assign \new_[61293]_  = ~A266 & A265;
  assign \new_[61294]_  = A202 & \new_[61293]_ ;
  assign \new_[61297]_  = A268 & A267;
  assign \new_[61300]_  = A301 & ~A300;
  assign \new_[61301]_  = \new_[61300]_  & \new_[61297]_ ;
  assign \new_[61302]_  = \new_[61301]_  & \new_[61294]_ ;
  assign \new_[61306]_  = ~A167 & A168;
  assign \new_[61307]_  = ~A170 & \new_[61306]_ ;
  assign \new_[61310]_  = ~A199 & A166;
  assign \new_[61313]_  = A201 & A200;
  assign \new_[61314]_  = \new_[61313]_  & \new_[61310]_ ;
  assign \new_[61315]_  = \new_[61314]_  & \new_[61307]_ ;
  assign \new_[61319]_  = ~A266 & A265;
  assign \new_[61320]_  = A202 & \new_[61319]_ ;
  assign \new_[61323]_  = A268 & A267;
  assign \new_[61326]_  = A302 & ~A300;
  assign \new_[61327]_  = \new_[61326]_  & \new_[61323]_ ;
  assign \new_[61328]_  = \new_[61327]_  & \new_[61320]_ ;
  assign \new_[61332]_  = ~A167 & A168;
  assign \new_[61333]_  = ~A170 & \new_[61332]_ ;
  assign \new_[61336]_  = ~A199 & A166;
  assign \new_[61339]_  = A201 & A200;
  assign \new_[61340]_  = \new_[61339]_  & \new_[61336]_ ;
  assign \new_[61341]_  = \new_[61340]_  & \new_[61333]_ ;
  assign \new_[61345]_  = ~A266 & A265;
  assign \new_[61346]_  = A202 & \new_[61345]_ ;
  assign \new_[61349]_  = A268 & A267;
  assign \new_[61352]_  = A299 & A298;
  assign \new_[61353]_  = \new_[61352]_  & \new_[61349]_ ;
  assign \new_[61354]_  = \new_[61353]_  & \new_[61346]_ ;
  assign \new_[61358]_  = ~A167 & A168;
  assign \new_[61359]_  = ~A170 & \new_[61358]_ ;
  assign \new_[61362]_  = ~A199 & A166;
  assign \new_[61365]_  = A201 & A200;
  assign \new_[61366]_  = \new_[61365]_  & \new_[61362]_ ;
  assign \new_[61367]_  = \new_[61366]_  & \new_[61359]_ ;
  assign \new_[61371]_  = ~A266 & A265;
  assign \new_[61372]_  = A202 & \new_[61371]_ ;
  assign \new_[61375]_  = A268 & A267;
  assign \new_[61378]_  = ~A299 & ~A298;
  assign \new_[61379]_  = \new_[61378]_  & \new_[61375]_ ;
  assign \new_[61380]_  = \new_[61379]_  & \new_[61372]_ ;
  assign \new_[61384]_  = ~A167 & A168;
  assign \new_[61385]_  = ~A170 & \new_[61384]_ ;
  assign \new_[61388]_  = ~A199 & A166;
  assign \new_[61391]_  = A201 & A200;
  assign \new_[61392]_  = \new_[61391]_  & \new_[61388]_ ;
  assign \new_[61393]_  = \new_[61392]_  & \new_[61385]_ ;
  assign \new_[61397]_  = ~A266 & A265;
  assign \new_[61398]_  = A202 & \new_[61397]_ ;
  assign \new_[61401]_  = A269 & A267;
  assign \new_[61404]_  = A301 & ~A300;
  assign \new_[61405]_  = \new_[61404]_  & \new_[61401]_ ;
  assign \new_[61406]_  = \new_[61405]_  & \new_[61398]_ ;
  assign \new_[61410]_  = ~A167 & A168;
  assign \new_[61411]_  = ~A170 & \new_[61410]_ ;
  assign \new_[61414]_  = ~A199 & A166;
  assign \new_[61417]_  = A201 & A200;
  assign \new_[61418]_  = \new_[61417]_  & \new_[61414]_ ;
  assign \new_[61419]_  = \new_[61418]_  & \new_[61411]_ ;
  assign \new_[61423]_  = ~A266 & A265;
  assign \new_[61424]_  = A202 & \new_[61423]_ ;
  assign \new_[61427]_  = A269 & A267;
  assign \new_[61430]_  = A302 & ~A300;
  assign \new_[61431]_  = \new_[61430]_  & \new_[61427]_ ;
  assign \new_[61432]_  = \new_[61431]_  & \new_[61424]_ ;
  assign \new_[61436]_  = ~A167 & A168;
  assign \new_[61437]_  = ~A170 & \new_[61436]_ ;
  assign \new_[61440]_  = ~A199 & A166;
  assign \new_[61443]_  = A201 & A200;
  assign \new_[61444]_  = \new_[61443]_  & \new_[61440]_ ;
  assign \new_[61445]_  = \new_[61444]_  & \new_[61437]_ ;
  assign \new_[61449]_  = ~A266 & A265;
  assign \new_[61450]_  = A202 & \new_[61449]_ ;
  assign \new_[61453]_  = A269 & A267;
  assign \new_[61456]_  = A299 & A298;
  assign \new_[61457]_  = \new_[61456]_  & \new_[61453]_ ;
  assign \new_[61458]_  = \new_[61457]_  & \new_[61450]_ ;
  assign \new_[61462]_  = ~A167 & A168;
  assign \new_[61463]_  = ~A170 & \new_[61462]_ ;
  assign \new_[61466]_  = ~A199 & A166;
  assign \new_[61469]_  = A201 & A200;
  assign \new_[61470]_  = \new_[61469]_  & \new_[61466]_ ;
  assign \new_[61471]_  = \new_[61470]_  & \new_[61463]_ ;
  assign \new_[61475]_  = ~A266 & A265;
  assign \new_[61476]_  = A202 & \new_[61475]_ ;
  assign \new_[61479]_  = A269 & A267;
  assign \new_[61482]_  = ~A299 & ~A298;
  assign \new_[61483]_  = \new_[61482]_  & \new_[61479]_ ;
  assign \new_[61484]_  = \new_[61483]_  & \new_[61476]_ ;
  assign \new_[61488]_  = ~A167 & A168;
  assign \new_[61489]_  = ~A170 & \new_[61488]_ ;
  assign \new_[61492]_  = ~A199 & A166;
  assign \new_[61495]_  = A201 & A200;
  assign \new_[61496]_  = \new_[61495]_  & \new_[61492]_ ;
  assign \new_[61497]_  = \new_[61496]_  & \new_[61489]_ ;
  assign \new_[61501]_  = A266 & ~A265;
  assign \new_[61502]_  = A203 & \new_[61501]_ ;
  assign \new_[61505]_  = A268 & A267;
  assign \new_[61508]_  = A301 & ~A300;
  assign \new_[61509]_  = \new_[61508]_  & \new_[61505]_ ;
  assign \new_[61510]_  = \new_[61509]_  & \new_[61502]_ ;
  assign \new_[61514]_  = ~A167 & A168;
  assign \new_[61515]_  = ~A170 & \new_[61514]_ ;
  assign \new_[61518]_  = ~A199 & A166;
  assign \new_[61521]_  = A201 & A200;
  assign \new_[61522]_  = \new_[61521]_  & \new_[61518]_ ;
  assign \new_[61523]_  = \new_[61522]_  & \new_[61515]_ ;
  assign \new_[61527]_  = A266 & ~A265;
  assign \new_[61528]_  = A203 & \new_[61527]_ ;
  assign \new_[61531]_  = A268 & A267;
  assign \new_[61534]_  = A302 & ~A300;
  assign \new_[61535]_  = \new_[61534]_  & \new_[61531]_ ;
  assign \new_[61536]_  = \new_[61535]_  & \new_[61528]_ ;
  assign \new_[61540]_  = ~A167 & A168;
  assign \new_[61541]_  = ~A170 & \new_[61540]_ ;
  assign \new_[61544]_  = ~A199 & A166;
  assign \new_[61547]_  = A201 & A200;
  assign \new_[61548]_  = \new_[61547]_  & \new_[61544]_ ;
  assign \new_[61549]_  = \new_[61548]_  & \new_[61541]_ ;
  assign \new_[61553]_  = A266 & ~A265;
  assign \new_[61554]_  = A203 & \new_[61553]_ ;
  assign \new_[61557]_  = A268 & A267;
  assign \new_[61560]_  = A299 & A298;
  assign \new_[61561]_  = \new_[61560]_  & \new_[61557]_ ;
  assign \new_[61562]_  = \new_[61561]_  & \new_[61554]_ ;
  assign \new_[61566]_  = ~A167 & A168;
  assign \new_[61567]_  = ~A170 & \new_[61566]_ ;
  assign \new_[61570]_  = ~A199 & A166;
  assign \new_[61573]_  = A201 & A200;
  assign \new_[61574]_  = \new_[61573]_  & \new_[61570]_ ;
  assign \new_[61575]_  = \new_[61574]_  & \new_[61567]_ ;
  assign \new_[61579]_  = A266 & ~A265;
  assign \new_[61580]_  = A203 & \new_[61579]_ ;
  assign \new_[61583]_  = A268 & A267;
  assign \new_[61586]_  = ~A299 & ~A298;
  assign \new_[61587]_  = \new_[61586]_  & \new_[61583]_ ;
  assign \new_[61588]_  = \new_[61587]_  & \new_[61580]_ ;
  assign \new_[61592]_  = ~A167 & A168;
  assign \new_[61593]_  = ~A170 & \new_[61592]_ ;
  assign \new_[61596]_  = ~A199 & A166;
  assign \new_[61599]_  = A201 & A200;
  assign \new_[61600]_  = \new_[61599]_  & \new_[61596]_ ;
  assign \new_[61601]_  = \new_[61600]_  & \new_[61593]_ ;
  assign \new_[61605]_  = A266 & ~A265;
  assign \new_[61606]_  = A203 & \new_[61605]_ ;
  assign \new_[61609]_  = A269 & A267;
  assign \new_[61612]_  = A301 & ~A300;
  assign \new_[61613]_  = \new_[61612]_  & \new_[61609]_ ;
  assign \new_[61614]_  = \new_[61613]_  & \new_[61606]_ ;
  assign \new_[61618]_  = ~A167 & A168;
  assign \new_[61619]_  = ~A170 & \new_[61618]_ ;
  assign \new_[61622]_  = ~A199 & A166;
  assign \new_[61625]_  = A201 & A200;
  assign \new_[61626]_  = \new_[61625]_  & \new_[61622]_ ;
  assign \new_[61627]_  = \new_[61626]_  & \new_[61619]_ ;
  assign \new_[61631]_  = A266 & ~A265;
  assign \new_[61632]_  = A203 & \new_[61631]_ ;
  assign \new_[61635]_  = A269 & A267;
  assign \new_[61638]_  = A302 & ~A300;
  assign \new_[61639]_  = \new_[61638]_  & \new_[61635]_ ;
  assign \new_[61640]_  = \new_[61639]_  & \new_[61632]_ ;
  assign \new_[61644]_  = ~A167 & A168;
  assign \new_[61645]_  = ~A170 & \new_[61644]_ ;
  assign \new_[61648]_  = ~A199 & A166;
  assign \new_[61651]_  = A201 & A200;
  assign \new_[61652]_  = \new_[61651]_  & \new_[61648]_ ;
  assign \new_[61653]_  = \new_[61652]_  & \new_[61645]_ ;
  assign \new_[61657]_  = A266 & ~A265;
  assign \new_[61658]_  = A203 & \new_[61657]_ ;
  assign \new_[61661]_  = A269 & A267;
  assign \new_[61664]_  = A299 & A298;
  assign \new_[61665]_  = \new_[61664]_  & \new_[61661]_ ;
  assign \new_[61666]_  = \new_[61665]_  & \new_[61658]_ ;
  assign \new_[61670]_  = ~A167 & A168;
  assign \new_[61671]_  = ~A170 & \new_[61670]_ ;
  assign \new_[61674]_  = ~A199 & A166;
  assign \new_[61677]_  = A201 & A200;
  assign \new_[61678]_  = \new_[61677]_  & \new_[61674]_ ;
  assign \new_[61679]_  = \new_[61678]_  & \new_[61671]_ ;
  assign \new_[61683]_  = A266 & ~A265;
  assign \new_[61684]_  = A203 & \new_[61683]_ ;
  assign \new_[61687]_  = A269 & A267;
  assign \new_[61690]_  = ~A299 & ~A298;
  assign \new_[61691]_  = \new_[61690]_  & \new_[61687]_ ;
  assign \new_[61692]_  = \new_[61691]_  & \new_[61684]_ ;
  assign \new_[61696]_  = ~A167 & A168;
  assign \new_[61697]_  = ~A170 & \new_[61696]_ ;
  assign \new_[61700]_  = ~A199 & A166;
  assign \new_[61703]_  = A201 & A200;
  assign \new_[61704]_  = \new_[61703]_  & \new_[61700]_ ;
  assign \new_[61705]_  = \new_[61704]_  & \new_[61697]_ ;
  assign \new_[61709]_  = ~A266 & A265;
  assign \new_[61710]_  = A203 & \new_[61709]_ ;
  assign \new_[61713]_  = A268 & A267;
  assign \new_[61716]_  = A301 & ~A300;
  assign \new_[61717]_  = \new_[61716]_  & \new_[61713]_ ;
  assign \new_[61718]_  = \new_[61717]_  & \new_[61710]_ ;
  assign \new_[61722]_  = ~A167 & A168;
  assign \new_[61723]_  = ~A170 & \new_[61722]_ ;
  assign \new_[61726]_  = ~A199 & A166;
  assign \new_[61729]_  = A201 & A200;
  assign \new_[61730]_  = \new_[61729]_  & \new_[61726]_ ;
  assign \new_[61731]_  = \new_[61730]_  & \new_[61723]_ ;
  assign \new_[61735]_  = ~A266 & A265;
  assign \new_[61736]_  = A203 & \new_[61735]_ ;
  assign \new_[61739]_  = A268 & A267;
  assign \new_[61742]_  = A302 & ~A300;
  assign \new_[61743]_  = \new_[61742]_  & \new_[61739]_ ;
  assign \new_[61744]_  = \new_[61743]_  & \new_[61736]_ ;
  assign \new_[61748]_  = ~A167 & A168;
  assign \new_[61749]_  = ~A170 & \new_[61748]_ ;
  assign \new_[61752]_  = ~A199 & A166;
  assign \new_[61755]_  = A201 & A200;
  assign \new_[61756]_  = \new_[61755]_  & \new_[61752]_ ;
  assign \new_[61757]_  = \new_[61756]_  & \new_[61749]_ ;
  assign \new_[61761]_  = ~A266 & A265;
  assign \new_[61762]_  = A203 & \new_[61761]_ ;
  assign \new_[61765]_  = A268 & A267;
  assign \new_[61768]_  = A299 & A298;
  assign \new_[61769]_  = \new_[61768]_  & \new_[61765]_ ;
  assign \new_[61770]_  = \new_[61769]_  & \new_[61762]_ ;
  assign \new_[61774]_  = ~A167 & A168;
  assign \new_[61775]_  = ~A170 & \new_[61774]_ ;
  assign \new_[61778]_  = ~A199 & A166;
  assign \new_[61781]_  = A201 & A200;
  assign \new_[61782]_  = \new_[61781]_  & \new_[61778]_ ;
  assign \new_[61783]_  = \new_[61782]_  & \new_[61775]_ ;
  assign \new_[61787]_  = ~A266 & A265;
  assign \new_[61788]_  = A203 & \new_[61787]_ ;
  assign \new_[61791]_  = A268 & A267;
  assign \new_[61794]_  = ~A299 & ~A298;
  assign \new_[61795]_  = \new_[61794]_  & \new_[61791]_ ;
  assign \new_[61796]_  = \new_[61795]_  & \new_[61788]_ ;
  assign \new_[61800]_  = ~A167 & A168;
  assign \new_[61801]_  = ~A170 & \new_[61800]_ ;
  assign \new_[61804]_  = ~A199 & A166;
  assign \new_[61807]_  = A201 & A200;
  assign \new_[61808]_  = \new_[61807]_  & \new_[61804]_ ;
  assign \new_[61809]_  = \new_[61808]_  & \new_[61801]_ ;
  assign \new_[61813]_  = ~A266 & A265;
  assign \new_[61814]_  = A203 & \new_[61813]_ ;
  assign \new_[61817]_  = A269 & A267;
  assign \new_[61820]_  = A301 & ~A300;
  assign \new_[61821]_  = \new_[61820]_  & \new_[61817]_ ;
  assign \new_[61822]_  = \new_[61821]_  & \new_[61814]_ ;
  assign \new_[61826]_  = ~A167 & A168;
  assign \new_[61827]_  = ~A170 & \new_[61826]_ ;
  assign \new_[61830]_  = ~A199 & A166;
  assign \new_[61833]_  = A201 & A200;
  assign \new_[61834]_  = \new_[61833]_  & \new_[61830]_ ;
  assign \new_[61835]_  = \new_[61834]_  & \new_[61827]_ ;
  assign \new_[61839]_  = ~A266 & A265;
  assign \new_[61840]_  = A203 & \new_[61839]_ ;
  assign \new_[61843]_  = A269 & A267;
  assign \new_[61846]_  = A302 & ~A300;
  assign \new_[61847]_  = \new_[61846]_  & \new_[61843]_ ;
  assign \new_[61848]_  = \new_[61847]_  & \new_[61840]_ ;
  assign \new_[61852]_  = ~A167 & A168;
  assign \new_[61853]_  = ~A170 & \new_[61852]_ ;
  assign \new_[61856]_  = ~A199 & A166;
  assign \new_[61859]_  = A201 & A200;
  assign \new_[61860]_  = \new_[61859]_  & \new_[61856]_ ;
  assign \new_[61861]_  = \new_[61860]_  & \new_[61853]_ ;
  assign \new_[61865]_  = ~A266 & A265;
  assign \new_[61866]_  = A203 & \new_[61865]_ ;
  assign \new_[61869]_  = A269 & A267;
  assign \new_[61872]_  = A299 & A298;
  assign \new_[61873]_  = \new_[61872]_  & \new_[61869]_ ;
  assign \new_[61874]_  = \new_[61873]_  & \new_[61866]_ ;
  assign \new_[61878]_  = ~A167 & A168;
  assign \new_[61879]_  = ~A170 & \new_[61878]_ ;
  assign \new_[61882]_  = ~A199 & A166;
  assign \new_[61885]_  = A201 & A200;
  assign \new_[61886]_  = \new_[61885]_  & \new_[61882]_ ;
  assign \new_[61887]_  = \new_[61886]_  & \new_[61879]_ ;
  assign \new_[61891]_  = ~A266 & A265;
  assign \new_[61892]_  = A203 & \new_[61891]_ ;
  assign \new_[61895]_  = A269 & A267;
  assign \new_[61898]_  = ~A299 & ~A298;
  assign \new_[61899]_  = \new_[61898]_  & \new_[61895]_ ;
  assign \new_[61900]_  = \new_[61899]_  & \new_[61892]_ ;
  assign \new_[61904]_  = ~A167 & A168;
  assign \new_[61905]_  = ~A170 & \new_[61904]_ ;
  assign \new_[61908]_  = A199 & A166;
  assign \new_[61911]_  = A201 & ~A200;
  assign \new_[61912]_  = \new_[61911]_  & \new_[61908]_ ;
  assign \new_[61913]_  = \new_[61912]_  & \new_[61905]_ ;
  assign \new_[61917]_  = A266 & ~A265;
  assign \new_[61918]_  = A202 & \new_[61917]_ ;
  assign \new_[61921]_  = A268 & A267;
  assign \new_[61924]_  = A301 & ~A300;
  assign \new_[61925]_  = \new_[61924]_  & \new_[61921]_ ;
  assign \new_[61926]_  = \new_[61925]_  & \new_[61918]_ ;
  assign \new_[61930]_  = ~A167 & A168;
  assign \new_[61931]_  = ~A170 & \new_[61930]_ ;
  assign \new_[61934]_  = A199 & A166;
  assign \new_[61937]_  = A201 & ~A200;
  assign \new_[61938]_  = \new_[61937]_  & \new_[61934]_ ;
  assign \new_[61939]_  = \new_[61938]_  & \new_[61931]_ ;
  assign \new_[61943]_  = A266 & ~A265;
  assign \new_[61944]_  = A202 & \new_[61943]_ ;
  assign \new_[61947]_  = A268 & A267;
  assign \new_[61950]_  = A302 & ~A300;
  assign \new_[61951]_  = \new_[61950]_  & \new_[61947]_ ;
  assign \new_[61952]_  = \new_[61951]_  & \new_[61944]_ ;
  assign \new_[61956]_  = ~A167 & A168;
  assign \new_[61957]_  = ~A170 & \new_[61956]_ ;
  assign \new_[61960]_  = A199 & A166;
  assign \new_[61963]_  = A201 & ~A200;
  assign \new_[61964]_  = \new_[61963]_  & \new_[61960]_ ;
  assign \new_[61965]_  = \new_[61964]_  & \new_[61957]_ ;
  assign \new_[61969]_  = A266 & ~A265;
  assign \new_[61970]_  = A202 & \new_[61969]_ ;
  assign \new_[61973]_  = A268 & A267;
  assign \new_[61976]_  = A299 & A298;
  assign \new_[61977]_  = \new_[61976]_  & \new_[61973]_ ;
  assign \new_[61978]_  = \new_[61977]_  & \new_[61970]_ ;
  assign \new_[61982]_  = ~A167 & A168;
  assign \new_[61983]_  = ~A170 & \new_[61982]_ ;
  assign \new_[61986]_  = A199 & A166;
  assign \new_[61989]_  = A201 & ~A200;
  assign \new_[61990]_  = \new_[61989]_  & \new_[61986]_ ;
  assign \new_[61991]_  = \new_[61990]_  & \new_[61983]_ ;
  assign \new_[61995]_  = A266 & ~A265;
  assign \new_[61996]_  = A202 & \new_[61995]_ ;
  assign \new_[61999]_  = A268 & A267;
  assign \new_[62002]_  = ~A299 & ~A298;
  assign \new_[62003]_  = \new_[62002]_  & \new_[61999]_ ;
  assign \new_[62004]_  = \new_[62003]_  & \new_[61996]_ ;
  assign \new_[62008]_  = ~A167 & A168;
  assign \new_[62009]_  = ~A170 & \new_[62008]_ ;
  assign \new_[62012]_  = A199 & A166;
  assign \new_[62015]_  = A201 & ~A200;
  assign \new_[62016]_  = \new_[62015]_  & \new_[62012]_ ;
  assign \new_[62017]_  = \new_[62016]_  & \new_[62009]_ ;
  assign \new_[62021]_  = A266 & ~A265;
  assign \new_[62022]_  = A202 & \new_[62021]_ ;
  assign \new_[62025]_  = A269 & A267;
  assign \new_[62028]_  = A301 & ~A300;
  assign \new_[62029]_  = \new_[62028]_  & \new_[62025]_ ;
  assign \new_[62030]_  = \new_[62029]_  & \new_[62022]_ ;
  assign \new_[62034]_  = ~A167 & A168;
  assign \new_[62035]_  = ~A170 & \new_[62034]_ ;
  assign \new_[62038]_  = A199 & A166;
  assign \new_[62041]_  = A201 & ~A200;
  assign \new_[62042]_  = \new_[62041]_  & \new_[62038]_ ;
  assign \new_[62043]_  = \new_[62042]_  & \new_[62035]_ ;
  assign \new_[62047]_  = A266 & ~A265;
  assign \new_[62048]_  = A202 & \new_[62047]_ ;
  assign \new_[62051]_  = A269 & A267;
  assign \new_[62054]_  = A302 & ~A300;
  assign \new_[62055]_  = \new_[62054]_  & \new_[62051]_ ;
  assign \new_[62056]_  = \new_[62055]_  & \new_[62048]_ ;
  assign \new_[62060]_  = ~A167 & A168;
  assign \new_[62061]_  = ~A170 & \new_[62060]_ ;
  assign \new_[62064]_  = A199 & A166;
  assign \new_[62067]_  = A201 & ~A200;
  assign \new_[62068]_  = \new_[62067]_  & \new_[62064]_ ;
  assign \new_[62069]_  = \new_[62068]_  & \new_[62061]_ ;
  assign \new_[62073]_  = A266 & ~A265;
  assign \new_[62074]_  = A202 & \new_[62073]_ ;
  assign \new_[62077]_  = A269 & A267;
  assign \new_[62080]_  = A299 & A298;
  assign \new_[62081]_  = \new_[62080]_  & \new_[62077]_ ;
  assign \new_[62082]_  = \new_[62081]_  & \new_[62074]_ ;
  assign \new_[62086]_  = ~A167 & A168;
  assign \new_[62087]_  = ~A170 & \new_[62086]_ ;
  assign \new_[62090]_  = A199 & A166;
  assign \new_[62093]_  = A201 & ~A200;
  assign \new_[62094]_  = \new_[62093]_  & \new_[62090]_ ;
  assign \new_[62095]_  = \new_[62094]_  & \new_[62087]_ ;
  assign \new_[62099]_  = A266 & ~A265;
  assign \new_[62100]_  = A202 & \new_[62099]_ ;
  assign \new_[62103]_  = A269 & A267;
  assign \new_[62106]_  = ~A299 & ~A298;
  assign \new_[62107]_  = \new_[62106]_  & \new_[62103]_ ;
  assign \new_[62108]_  = \new_[62107]_  & \new_[62100]_ ;
  assign \new_[62112]_  = ~A167 & A168;
  assign \new_[62113]_  = ~A170 & \new_[62112]_ ;
  assign \new_[62116]_  = A199 & A166;
  assign \new_[62119]_  = A201 & ~A200;
  assign \new_[62120]_  = \new_[62119]_  & \new_[62116]_ ;
  assign \new_[62121]_  = \new_[62120]_  & \new_[62113]_ ;
  assign \new_[62125]_  = ~A266 & A265;
  assign \new_[62126]_  = A202 & \new_[62125]_ ;
  assign \new_[62129]_  = A268 & A267;
  assign \new_[62132]_  = A301 & ~A300;
  assign \new_[62133]_  = \new_[62132]_  & \new_[62129]_ ;
  assign \new_[62134]_  = \new_[62133]_  & \new_[62126]_ ;
  assign \new_[62138]_  = ~A167 & A168;
  assign \new_[62139]_  = ~A170 & \new_[62138]_ ;
  assign \new_[62142]_  = A199 & A166;
  assign \new_[62145]_  = A201 & ~A200;
  assign \new_[62146]_  = \new_[62145]_  & \new_[62142]_ ;
  assign \new_[62147]_  = \new_[62146]_  & \new_[62139]_ ;
  assign \new_[62151]_  = ~A266 & A265;
  assign \new_[62152]_  = A202 & \new_[62151]_ ;
  assign \new_[62155]_  = A268 & A267;
  assign \new_[62158]_  = A302 & ~A300;
  assign \new_[62159]_  = \new_[62158]_  & \new_[62155]_ ;
  assign \new_[62160]_  = \new_[62159]_  & \new_[62152]_ ;
  assign \new_[62164]_  = ~A167 & A168;
  assign \new_[62165]_  = ~A170 & \new_[62164]_ ;
  assign \new_[62168]_  = A199 & A166;
  assign \new_[62171]_  = A201 & ~A200;
  assign \new_[62172]_  = \new_[62171]_  & \new_[62168]_ ;
  assign \new_[62173]_  = \new_[62172]_  & \new_[62165]_ ;
  assign \new_[62177]_  = ~A266 & A265;
  assign \new_[62178]_  = A202 & \new_[62177]_ ;
  assign \new_[62181]_  = A268 & A267;
  assign \new_[62184]_  = A299 & A298;
  assign \new_[62185]_  = \new_[62184]_  & \new_[62181]_ ;
  assign \new_[62186]_  = \new_[62185]_  & \new_[62178]_ ;
  assign \new_[62190]_  = ~A167 & A168;
  assign \new_[62191]_  = ~A170 & \new_[62190]_ ;
  assign \new_[62194]_  = A199 & A166;
  assign \new_[62197]_  = A201 & ~A200;
  assign \new_[62198]_  = \new_[62197]_  & \new_[62194]_ ;
  assign \new_[62199]_  = \new_[62198]_  & \new_[62191]_ ;
  assign \new_[62203]_  = ~A266 & A265;
  assign \new_[62204]_  = A202 & \new_[62203]_ ;
  assign \new_[62207]_  = A268 & A267;
  assign \new_[62210]_  = ~A299 & ~A298;
  assign \new_[62211]_  = \new_[62210]_  & \new_[62207]_ ;
  assign \new_[62212]_  = \new_[62211]_  & \new_[62204]_ ;
  assign \new_[62216]_  = ~A167 & A168;
  assign \new_[62217]_  = ~A170 & \new_[62216]_ ;
  assign \new_[62220]_  = A199 & A166;
  assign \new_[62223]_  = A201 & ~A200;
  assign \new_[62224]_  = \new_[62223]_  & \new_[62220]_ ;
  assign \new_[62225]_  = \new_[62224]_  & \new_[62217]_ ;
  assign \new_[62229]_  = ~A266 & A265;
  assign \new_[62230]_  = A202 & \new_[62229]_ ;
  assign \new_[62233]_  = A269 & A267;
  assign \new_[62236]_  = A301 & ~A300;
  assign \new_[62237]_  = \new_[62236]_  & \new_[62233]_ ;
  assign \new_[62238]_  = \new_[62237]_  & \new_[62230]_ ;
  assign \new_[62242]_  = ~A167 & A168;
  assign \new_[62243]_  = ~A170 & \new_[62242]_ ;
  assign \new_[62246]_  = A199 & A166;
  assign \new_[62249]_  = A201 & ~A200;
  assign \new_[62250]_  = \new_[62249]_  & \new_[62246]_ ;
  assign \new_[62251]_  = \new_[62250]_  & \new_[62243]_ ;
  assign \new_[62255]_  = ~A266 & A265;
  assign \new_[62256]_  = A202 & \new_[62255]_ ;
  assign \new_[62259]_  = A269 & A267;
  assign \new_[62262]_  = A302 & ~A300;
  assign \new_[62263]_  = \new_[62262]_  & \new_[62259]_ ;
  assign \new_[62264]_  = \new_[62263]_  & \new_[62256]_ ;
  assign \new_[62268]_  = ~A167 & A168;
  assign \new_[62269]_  = ~A170 & \new_[62268]_ ;
  assign \new_[62272]_  = A199 & A166;
  assign \new_[62275]_  = A201 & ~A200;
  assign \new_[62276]_  = \new_[62275]_  & \new_[62272]_ ;
  assign \new_[62277]_  = \new_[62276]_  & \new_[62269]_ ;
  assign \new_[62281]_  = ~A266 & A265;
  assign \new_[62282]_  = A202 & \new_[62281]_ ;
  assign \new_[62285]_  = A269 & A267;
  assign \new_[62288]_  = A299 & A298;
  assign \new_[62289]_  = \new_[62288]_  & \new_[62285]_ ;
  assign \new_[62290]_  = \new_[62289]_  & \new_[62282]_ ;
  assign \new_[62294]_  = ~A167 & A168;
  assign \new_[62295]_  = ~A170 & \new_[62294]_ ;
  assign \new_[62298]_  = A199 & A166;
  assign \new_[62301]_  = A201 & ~A200;
  assign \new_[62302]_  = \new_[62301]_  & \new_[62298]_ ;
  assign \new_[62303]_  = \new_[62302]_  & \new_[62295]_ ;
  assign \new_[62307]_  = ~A266 & A265;
  assign \new_[62308]_  = A202 & \new_[62307]_ ;
  assign \new_[62311]_  = A269 & A267;
  assign \new_[62314]_  = ~A299 & ~A298;
  assign \new_[62315]_  = \new_[62314]_  & \new_[62311]_ ;
  assign \new_[62316]_  = \new_[62315]_  & \new_[62308]_ ;
  assign \new_[62320]_  = ~A167 & A168;
  assign \new_[62321]_  = ~A170 & \new_[62320]_ ;
  assign \new_[62324]_  = A199 & A166;
  assign \new_[62327]_  = A201 & ~A200;
  assign \new_[62328]_  = \new_[62327]_  & \new_[62324]_ ;
  assign \new_[62329]_  = \new_[62328]_  & \new_[62321]_ ;
  assign \new_[62333]_  = A266 & ~A265;
  assign \new_[62334]_  = A203 & \new_[62333]_ ;
  assign \new_[62337]_  = A268 & A267;
  assign \new_[62340]_  = A301 & ~A300;
  assign \new_[62341]_  = \new_[62340]_  & \new_[62337]_ ;
  assign \new_[62342]_  = \new_[62341]_  & \new_[62334]_ ;
  assign \new_[62346]_  = ~A167 & A168;
  assign \new_[62347]_  = ~A170 & \new_[62346]_ ;
  assign \new_[62350]_  = A199 & A166;
  assign \new_[62353]_  = A201 & ~A200;
  assign \new_[62354]_  = \new_[62353]_  & \new_[62350]_ ;
  assign \new_[62355]_  = \new_[62354]_  & \new_[62347]_ ;
  assign \new_[62359]_  = A266 & ~A265;
  assign \new_[62360]_  = A203 & \new_[62359]_ ;
  assign \new_[62363]_  = A268 & A267;
  assign \new_[62366]_  = A302 & ~A300;
  assign \new_[62367]_  = \new_[62366]_  & \new_[62363]_ ;
  assign \new_[62368]_  = \new_[62367]_  & \new_[62360]_ ;
  assign \new_[62372]_  = ~A167 & A168;
  assign \new_[62373]_  = ~A170 & \new_[62372]_ ;
  assign \new_[62376]_  = A199 & A166;
  assign \new_[62379]_  = A201 & ~A200;
  assign \new_[62380]_  = \new_[62379]_  & \new_[62376]_ ;
  assign \new_[62381]_  = \new_[62380]_  & \new_[62373]_ ;
  assign \new_[62385]_  = A266 & ~A265;
  assign \new_[62386]_  = A203 & \new_[62385]_ ;
  assign \new_[62389]_  = A268 & A267;
  assign \new_[62392]_  = A299 & A298;
  assign \new_[62393]_  = \new_[62392]_  & \new_[62389]_ ;
  assign \new_[62394]_  = \new_[62393]_  & \new_[62386]_ ;
  assign \new_[62398]_  = ~A167 & A168;
  assign \new_[62399]_  = ~A170 & \new_[62398]_ ;
  assign \new_[62402]_  = A199 & A166;
  assign \new_[62405]_  = A201 & ~A200;
  assign \new_[62406]_  = \new_[62405]_  & \new_[62402]_ ;
  assign \new_[62407]_  = \new_[62406]_  & \new_[62399]_ ;
  assign \new_[62411]_  = A266 & ~A265;
  assign \new_[62412]_  = A203 & \new_[62411]_ ;
  assign \new_[62415]_  = A268 & A267;
  assign \new_[62418]_  = ~A299 & ~A298;
  assign \new_[62419]_  = \new_[62418]_  & \new_[62415]_ ;
  assign \new_[62420]_  = \new_[62419]_  & \new_[62412]_ ;
  assign \new_[62424]_  = ~A167 & A168;
  assign \new_[62425]_  = ~A170 & \new_[62424]_ ;
  assign \new_[62428]_  = A199 & A166;
  assign \new_[62431]_  = A201 & ~A200;
  assign \new_[62432]_  = \new_[62431]_  & \new_[62428]_ ;
  assign \new_[62433]_  = \new_[62432]_  & \new_[62425]_ ;
  assign \new_[62437]_  = A266 & ~A265;
  assign \new_[62438]_  = A203 & \new_[62437]_ ;
  assign \new_[62441]_  = A269 & A267;
  assign \new_[62444]_  = A301 & ~A300;
  assign \new_[62445]_  = \new_[62444]_  & \new_[62441]_ ;
  assign \new_[62446]_  = \new_[62445]_  & \new_[62438]_ ;
  assign \new_[62450]_  = ~A167 & A168;
  assign \new_[62451]_  = ~A170 & \new_[62450]_ ;
  assign \new_[62454]_  = A199 & A166;
  assign \new_[62457]_  = A201 & ~A200;
  assign \new_[62458]_  = \new_[62457]_  & \new_[62454]_ ;
  assign \new_[62459]_  = \new_[62458]_  & \new_[62451]_ ;
  assign \new_[62463]_  = A266 & ~A265;
  assign \new_[62464]_  = A203 & \new_[62463]_ ;
  assign \new_[62467]_  = A269 & A267;
  assign \new_[62470]_  = A302 & ~A300;
  assign \new_[62471]_  = \new_[62470]_  & \new_[62467]_ ;
  assign \new_[62472]_  = \new_[62471]_  & \new_[62464]_ ;
  assign \new_[62476]_  = ~A167 & A168;
  assign \new_[62477]_  = ~A170 & \new_[62476]_ ;
  assign \new_[62480]_  = A199 & A166;
  assign \new_[62483]_  = A201 & ~A200;
  assign \new_[62484]_  = \new_[62483]_  & \new_[62480]_ ;
  assign \new_[62485]_  = \new_[62484]_  & \new_[62477]_ ;
  assign \new_[62489]_  = A266 & ~A265;
  assign \new_[62490]_  = A203 & \new_[62489]_ ;
  assign \new_[62493]_  = A269 & A267;
  assign \new_[62496]_  = A299 & A298;
  assign \new_[62497]_  = \new_[62496]_  & \new_[62493]_ ;
  assign \new_[62498]_  = \new_[62497]_  & \new_[62490]_ ;
  assign \new_[62502]_  = ~A167 & A168;
  assign \new_[62503]_  = ~A170 & \new_[62502]_ ;
  assign \new_[62506]_  = A199 & A166;
  assign \new_[62509]_  = A201 & ~A200;
  assign \new_[62510]_  = \new_[62509]_  & \new_[62506]_ ;
  assign \new_[62511]_  = \new_[62510]_  & \new_[62503]_ ;
  assign \new_[62515]_  = A266 & ~A265;
  assign \new_[62516]_  = A203 & \new_[62515]_ ;
  assign \new_[62519]_  = A269 & A267;
  assign \new_[62522]_  = ~A299 & ~A298;
  assign \new_[62523]_  = \new_[62522]_  & \new_[62519]_ ;
  assign \new_[62524]_  = \new_[62523]_  & \new_[62516]_ ;
  assign \new_[62528]_  = ~A167 & A168;
  assign \new_[62529]_  = ~A170 & \new_[62528]_ ;
  assign \new_[62532]_  = A199 & A166;
  assign \new_[62535]_  = A201 & ~A200;
  assign \new_[62536]_  = \new_[62535]_  & \new_[62532]_ ;
  assign \new_[62537]_  = \new_[62536]_  & \new_[62529]_ ;
  assign \new_[62541]_  = ~A266 & A265;
  assign \new_[62542]_  = A203 & \new_[62541]_ ;
  assign \new_[62545]_  = A268 & A267;
  assign \new_[62548]_  = A301 & ~A300;
  assign \new_[62549]_  = \new_[62548]_  & \new_[62545]_ ;
  assign \new_[62550]_  = \new_[62549]_  & \new_[62542]_ ;
  assign \new_[62554]_  = ~A167 & A168;
  assign \new_[62555]_  = ~A170 & \new_[62554]_ ;
  assign \new_[62558]_  = A199 & A166;
  assign \new_[62561]_  = A201 & ~A200;
  assign \new_[62562]_  = \new_[62561]_  & \new_[62558]_ ;
  assign \new_[62563]_  = \new_[62562]_  & \new_[62555]_ ;
  assign \new_[62567]_  = ~A266 & A265;
  assign \new_[62568]_  = A203 & \new_[62567]_ ;
  assign \new_[62571]_  = A268 & A267;
  assign \new_[62574]_  = A302 & ~A300;
  assign \new_[62575]_  = \new_[62574]_  & \new_[62571]_ ;
  assign \new_[62576]_  = \new_[62575]_  & \new_[62568]_ ;
  assign \new_[62580]_  = ~A167 & A168;
  assign \new_[62581]_  = ~A170 & \new_[62580]_ ;
  assign \new_[62584]_  = A199 & A166;
  assign \new_[62587]_  = A201 & ~A200;
  assign \new_[62588]_  = \new_[62587]_  & \new_[62584]_ ;
  assign \new_[62589]_  = \new_[62588]_  & \new_[62581]_ ;
  assign \new_[62593]_  = ~A266 & A265;
  assign \new_[62594]_  = A203 & \new_[62593]_ ;
  assign \new_[62597]_  = A268 & A267;
  assign \new_[62600]_  = A299 & A298;
  assign \new_[62601]_  = \new_[62600]_  & \new_[62597]_ ;
  assign \new_[62602]_  = \new_[62601]_  & \new_[62594]_ ;
  assign \new_[62606]_  = ~A167 & A168;
  assign \new_[62607]_  = ~A170 & \new_[62606]_ ;
  assign \new_[62610]_  = A199 & A166;
  assign \new_[62613]_  = A201 & ~A200;
  assign \new_[62614]_  = \new_[62613]_  & \new_[62610]_ ;
  assign \new_[62615]_  = \new_[62614]_  & \new_[62607]_ ;
  assign \new_[62619]_  = ~A266 & A265;
  assign \new_[62620]_  = A203 & \new_[62619]_ ;
  assign \new_[62623]_  = A268 & A267;
  assign \new_[62626]_  = ~A299 & ~A298;
  assign \new_[62627]_  = \new_[62626]_  & \new_[62623]_ ;
  assign \new_[62628]_  = \new_[62627]_  & \new_[62620]_ ;
  assign \new_[62632]_  = ~A167 & A168;
  assign \new_[62633]_  = ~A170 & \new_[62632]_ ;
  assign \new_[62636]_  = A199 & A166;
  assign \new_[62639]_  = A201 & ~A200;
  assign \new_[62640]_  = \new_[62639]_  & \new_[62636]_ ;
  assign \new_[62641]_  = \new_[62640]_  & \new_[62633]_ ;
  assign \new_[62645]_  = ~A266 & A265;
  assign \new_[62646]_  = A203 & \new_[62645]_ ;
  assign \new_[62649]_  = A269 & A267;
  assign \new_[62652]_  = A301 & ~A300;
  assign \new_[62653]_  = \new_[62652]_  & \new_[62649]_ ;
  assign \new_[62654]_  = \new_[62653]_  & \new_[62646]_ ;
  assign \new_[62658]_  = ~A167 & A168;
  assign \new_[62659]_  = ~A170 & \new_[62658]_ ;
  assign \new_[62662]_  = A199 & A166;
  assign \new_[62665]_  = A201 & ~A200;
  assign \new_[62666]_  = \new_[62665]_  & \new_[62662]_ ;
  assign \new_[62667]_  = \new_[62666]_  & \new_[62659]_ ;
  assign \new_[62671]_  = ~A266 & A265;
  assign \new_[62672]_  = A203 & \new_[62671]_ ;
  assign \new_[62675]_  = A269 & A267;
  assign \new_[62678]_  = A302 & ~A300;
  assign \new_[62679]_  = \new_[62678]_  & \new_[62675]_ ;
  assign \new_[62680]_  = \new_[62679]_  & \new_[62672]_ ;
  assign \new_[62684]_  = ~A167 & A168;
  assign \new_[62685]_  = ~A170 & \new_[62684]_ ;
  assign \new_[62688]_  = A199 & A166;
  assign \new_[62691]_  = A201 & ~A200;
  assign \new_[62692]_  = \new_[62691]_  & \new_[62688]_ ;
  assign \new_[62693]_  = \new_[62692]_  & \new_[62685]_ ;
  assign \new_[62697]_  = ~A266 & A265;
  assign \new_[62698]_  = A203 & \new_[62697]_ ;
  assign \new_[62701]_  = A269 & A267;
  assign \new_[62704]_  = A299 & A298;
  assign \new_[62705]_  = \new_[62704]_  & \new_[62701]_ ;
  assign \new_[62706]_  = \new_[62705]_  & \new_[62698]_ ;
  assign \new_[62710]_  = ~A167 & A168;
  assign \new_[62711]_  = ~A170 & \new_[62710]_ ;
  assign \new_[62714]_  = A199 & A166;
  assign \new_[62717]_  = A201 & ~A200;
  assign \new_[62718]_  = \new_[62717]_  & \new_[62714]_ ;
  assign \new_[62719]_  = \new_[62718]_  & \new_[62711]_ ;
  assign \new_[62723]_  = ~A266 & A265;
  assign \new_[62724]_  = A203 & \new_[62723]_ ;
  assign \new_[62727]_  = A269 & A267;
  assign \new_[62730]_  = ~A299 & ~A298;
  assign \new_[62731]_  = \new_[62730]_  & \new_[62727]_ ;
  assign \new_[62732]_  = \new_[62731]_  & \new_[62724]_ ;
  assign \new_[62736]_  = ~A167 & A168;
  assign \new_[62737]_  = ~A170 & \new_[62736]_ ;
  assign \new_[62740]_  = ~A199 & A166;
  assign \new_[62743]_  = A267 & ~A200;
  assign \new_[62744]_  = \new_[62743]_  & \new_[62740]_ ;
  assign \new_[62745]_  = \new_[62744]_  & \new_[62737]_ ;
  assign \new_[62749]_  = A298 & ~A269;
  assign \new_[62750]_  = ~A268 & \new_[62749]_ ;
  assign \new_[62753]_  = ~A300 & ~A299;
  assign \new_[62756]_  = ~A302 & ~A301;
  assign \new_[62757]_  = \new_[62756]_  & \new_[62753]_ ;
  assign \new_[62758]_  = \new_[62757]_  & \new_[62750]_ ;
  assign \new_[62762]_  = ~A167 & A168;
  assign \new_[62763]_  = ~A170 & \new_[62762]_ ;
  assign \new_[62766]_  = ~A199 & A166;
  assign \new_[62769]_  = A267 & ~A200;
  assign \new_[62770]_  = \new_[62769]_  & \new_[62766]_ ;
  assign \new_[62771]_  = \new_[62770]_  & \new_[62763]_ ;
  assign \new_[62775]_  = ~A298 & ~A269;
  assign \new_[62776]_  = ~A268 & \new_[62775]_ ;
  assign \new_[62779]_  = ~A300 & A299;
  assign \new_[62782]_  = ~A302 & ~A301;
  assign \new_[62783]_  = \new_[62782]_  & \new_[62779]_ ;
  assign \new_[62784]_  = \new_[62783]_  & \new_[62776]_ ;
  assign \new_[62788]_  = ~A199 & ~A168;
  assign \new_[62789]_  = ~A170 & \new_[62788]_ ;
  assign \new_[62792]_  = A201 & A200;
  assign \new_[62795]_  = A267 & A202;
  assign \new_[62796]_  = \new_[62795]_  & \new_[62792]_ ;
  assign \new_[62797]_  = \new_[62796]_  & \new_[62789]_ ;
  assign \new_[62801]_  = A298 & ~A269;
  assign \new_[62802]_  = ~A268 & \new_[62801]_ ;
  assign \new_[62805]_  = ~A300 & ~A299;
  assign \new_[62808]_  = ~A302 & ~A301;
  assign \new_[62809]_  = \new_[62808]_  & \new_[62805]_ ;
  assign \new_[62810]_  = \new_[62809]_  & \new_[62802]_ ;
  assign \new_[62814]_  = ~A199 & ~A168;
  assign \new_[62815]_  = ~A170 & \new_[62814]_ ;
  assign \new_[62818]_  = A201 & A200;
  assign \new_[62821]_  = A267 & A202;
  assign \new_[62822]_  = \new_[62821]_  & \new_[62818]_ ;
  assign \new_[62823]_  = \new_[62822]_  & \new_[62815]_ ;
  assign \new_[62827]_  = ~A298 & ~A269;
  assign \new_[62828]_  = ~A268 & \new_[62827]_ ;
  assign \new_[62831]_  = ~A300 & A299;
  assign \new_[62834]_  = ~A302 & ~A301;
  assign \new_[62835]_  = \new_[62834]_  & \new_[62831]_ ;
  assign \new_[62836]_  = \new_[62835]_  & \new_[62828]_ ;
  assign \new_[62840]_  = ~A199 & ~A168;
  assign \new_[62841]_  = ~A170 & \new_[62840]_ ;
  assign \new_[62844]_  = A201 & A200;
  assign \new_[62847]_  = A267 & A203;
  assign \new_[62848]_  = \new_[62847]_  & \new_[62844]_ ;
  assign \new_[62849]_  = \new_[62848]_  & \new_[62841]_ ;
  assign \new_[62853]_  = A298 & ~A269;
  assign \new_[62854]_  = ~A268 & \new_[62853]_ ;
  assign \new_[62857]_  = ~A300 & ~A299;
  assign \new_[62860]_  = ~A302 & ~A301;
  assign \new_[62861]_  = \new_[62860]_  & \new_[62857]_ ;
  assign \new_[62862]_  = \new_[62861]_  & \new_[62854]_ ;
  assign \new_[62866]_  = ~A199 & ~A168;
  assign \new_[62867]_  = ~A170 & \new_[62866]_ ;
  assign \new_[62870]_  = A201 & A200;
  assign \new_[62873]_  = A267 & A203;
  assign \new_[62874]_  = \new_[62873]_  & \new_[62870]_ ;
  assign \new_[62875]_  = \new_[62874]_  & \new_[62867]_ ;
  assign \new_[62879]_  = ~A298 & ~A269;
  assign \new_[62880]_  = ~A268 & \new_[62879]_ ;
  assign \new_[62883]_  = ~A300 & A299;
  assign \new_[62886]_  = ~A302 & ~A301;
  assign \new_[62887]_  = \new_[62886]_  & \new_[62883]_ ;
  assign \new_[62888]_  = \new_[62887]_  & \new_[62880]_ ;
  assign \new_[62892]_  = ~A199 & ~A168;
  assign \new_[62893]_  = ~A170 & \new_[62892]_ ;
  assign \new_[62896]_  = ~A201 & A200;
  assign \new_[62899]_  = ~A203 & ~A202;
  assign \new_[62900]_  = \new_[62899]_  & \new_[62896]_ ;
  assign \new_[62901]_  = \new_[62900]_  & \new_[62893]_ ;
  assign \new_[62905]_  = ~A269 & ~A268;
  assign \new_[62906]_  = A267 & \new_[62905]_ ;
  assign \new_[62909]_  = ~A299 & A298;
  assign \new_[62912]_  = A301 & A300;
  assign \new_[62913]_  = \new_[62912]_  & \new_[62909]_ ;
  assign \new_[62914]_  = \new_[62913]_  & \new_[62906]_ ;
  assign \new_[62918]_  = ~A199 & ~A168;
  assign \new_[62919]_  = ~A170 & \new_[62918]_ ;
  assign \new_[62922]_  = ~A201 & A200;
  assign \new_[62925]_  = ~A203 & ~A202;
  assign \new_[62926]_  = \new_[62925]_  & \new_[62922]_ ;
  assign \new_[62927]_  = \new_[62926]_  & \new_[62919]_ ;
  assign \new_[62931]_  = ~A269 & ~A268;
  assign \new_[62932]_  = A267 & \new_[62931]_ ;
  assign \new_[62935]_  = ~A299 & A298;
  assign \new_[62938]_  = A302 & A300;
  assign \new_[62939]_  = \new_[62938]_  & \new_[62935]_ ;
  assign \new_[62940]_  = \new_[62939]_  & \new_[62932]_ ;
  assign \new_[62944]_  = ~A199 & ~A168;
  assign \new_[62945]_  = ~A170 & \new_[62944]_ ;
  assign \new_[62948]_  = ~A201 & A200;
  assign \new_[62951]_  = ~A203 & ~A202;
  assign \new_[62952]_  = \new_[62951]_  & \new_[62948]_ ;
  assign \new_[62953]_  = \new_[62952]_  & \new_[62945]_ ;
  assign \new_[62957]_  = ~A269 & ~A268;
  assign \new_[62958]_  = A267 & \new_[62957]_ ;
  assign \new_[62961]_  = A299 & ~A298;
  assign \new_[62964]_  = A301 & A300;
  assign \new_[62965]_  = \new_[62964]_  & \new_[62961]_ ;
  assign \new_[62966]_  = \new_[62965]_  & \new_[62958]_ ;
  assign \new_[62970]_  = ~A199 & ~A168;
  assign \new_[62971]_  = ~A170 & \new_[62970]_ ;
  assign \new_[62974]_  = ~A201 & A200;
  assign \new_[62977]_  = ~A203 & ~A202;
  assign \new_[62978]_  = \new_[62977]_  & \new_[62974]_ ;
  assign \new_[62979]_  = \new_[62978]_  & \new_[62971]_ ;
  assign \new_[62983]_  = ~A269 & ~A268;
  assign \new_[62984]_  = A267 & \new_[62983]_ ;
  assign \new_[62987]_  = A299 & ~A298;
  assign \new_[62990]_  = A302 & A300;
  assign \new_[62991]_  = \new_[62990]_  & \new_[62987]_ ;
  assign \new_[62992]_  = \new_[62991]_  & \new_[62984]_ ;
  assign \new_[62996]_  = ~A199 & ~A168;
  assign \new_[62997]_  = ~A170 & \new_[62996]_ ;
  assign \new_[63000]_  = ~A201 & A200;
  assign \new_[63003]_  = ~A203 & ~A202;
  assign \new_[63004]_  = \new_[63003]_  & \new_[63000]_ ;
  assign \new_[63005]_  = \new_[63004]_  & \new_[62997]_ ;
  assign \new_[63009]_  = A298 & A268;
  assign \new_[63010]_  = ~A267 & \new_[63009]_ ;
  assign \new_[63013]_  = ~A300 & ~A299;
  assign \new_[63016]_  = ~A302 & ~A301;
  assign \new_[63017]_  = \new_[63016]_  & \new_[63013]_ ;
  assign \new_[63018]_  = \new_[63017]_  & \new_[63010]_ ;
  assign \new_[63022]_  = ~A199 & ~A168;
  assign \new_[63023]_  = ~A170 & \new_[63022]_ ;
  assign \new_[63026]_  = ~A201 & A200;
  assign \new_[63029]_  = ~A203 & ~A202;
  assign \new_[63030]_  = \new_[63029]_  & \new_[63026]_ ;
  assign \new_[63031]_  = \new_[63030]_  & \new_[63023]_ ;
  assign \new_[63035]_  = ~A298 & A268;
  assign \new_[63036]_  = ~A267 & \new_[63035]_ ;
  assign \new_[63039]_  = ~A300 & A299;
  assign \new_[63042]_  = ~A302 & ~A301;
  assign \new_[63043]_  = \new_[63042]_  & \new_[63039]_ ;
  assign \new_[63044]_  = \new_[63043]_  & \new_[63036]_ ;
  assign \new_[63048]_  = ~A199 & ~A168;
  assign \new_[63049]_  = ~A170 & \new_[63048]_ ;
  assign \new_[63052]_  = ~A201 & A200;
  assign \new_[63055]_  = ~A203 & ~A202;
  assign \new_[63056]_  = \new_[63055]_  & \new_[63052]_ ;
  assign \new_[63057]_  = \new_[63056]_  & \new_[63049]_ ;
  assign \new_[63061]_  = A298 & A269;
  assign \new_[63062]_  = ~A267 & \new_[63061]_ ;
  assign \new_[63065]_  = ~A300 & ~A299;
  assign \new_[63068]_  = ~A302 & ~A301;
  assign \new_[63069]_  = \new_[63068]_  & \new_[63065]_ ;
  assign \new_[63070]_  = \new_[63069]_  & \new_[63062]_ ;
  assign \new_[63074]_  = ~A199 & ~A168;
  assign \new_[63075]_  = ~A170 & \new_[63074]_ ;
  assign \new_[63078]_  = ~A201 & A200;
  assign \new_[63081]_  = ~A203 & ~A202;
  assign \new_[63082]_  = \new_[63081]_  & \new_[63078]_ ;
  assign \new_[63083]_  = \new_[63082]_  & \new_[63075]_ ;
  assign \new_[63087]_  = ~A298 & A269;
  assign \new_[63088]_  = ~A267 & \new_[63087]_ ;
  assign \new_[63091]_  = ~A300 & A299;
  assign \new_[63094]_  = ~A302 & ~A301;
  assign \new_[63095]_  = \new_[63094]_  & \new_[63091]_ ;
  assign \new_[63096]_  = \new_[63095]_  & \new_[63088]_ ;
  assign \new_[63100]_  = ~A199 & ~A168;
  assign \new_[63101]_  = ~A170 & \new_[63100]_ ;
  assign \new_[63104]_  = ~A201 & A200;
  assign \new_[63107]_  = ~A203 & ~A202;
  assign \new_[63108]_  = \new_[63107]_  & \new_[63104]_ ;
  assign \new_[63109]_  = \new_[63108]_  & \new_[63101]_ ;
  assign \new_[63113]_  = A298 & A266;
  assign \new_[63114]_  = A265 & \new_[63113]_ ;
  assign \new_[63117]_  = ~A300 & ~A299;
  assign \new_[63120]_  = ~A302 & ~A301;
  assign \new_[63121]_  = \new_[63120]_  & \new_[63117]_ ;
  assign \new_[63122]_  = \new_[63121]_  & \new_[63114]_ ;
  assign \new_[63126]_  = ~A199 & ~A168;
  assign \new_[63127]_  = ~A170 & \new_[63126]_ ;
  assign \new_[63130]_  = ~A201 & A200;
  assign \new_[63133]_  = ~A203 & ~A202;
  assign \new_[63134]_  = \new_[63133]_  & \new_[63130]_ ;
  assign \new_[63135]_  = \new_[63134]_  & \new_[63127]_ ;
  assign \new_[63139]_  = ~A298 & A266;
  assign \new_[63140]_  = A265 & \new_[63139]_ ;
  assign \new_[63143]_  = ~A300 & A299;
  assign \new_[63146]_  = ~A302 & ~A301;
  assign \new_[63147]_  = \new_[63146]_  & \new_[63143]_ ;
  assign \new_[63148]_  = \new_[63147]_  & \new_[63140]_ ;
  assign \new_[63152]_  = ~A199 & ~A168;
  assign \new_[63153]_  = ~A170 & \new_[63152]_ ;
  assign \new_[63156]_  = ~A201 & A200;
  assign \new_[63159]_  = ~A203 & ~A202;
  assign \new_[63160]_  = \new_[63159]_  & \new_[63156]_ ;
  assign \new_[63161]_  = \new_[63160]_  & \new_[63153]_ ;
  assign \new_[63165]_  = A298 & ~A266;
  assign \new_[63166]_  = ~A265 & \new_[63165]_ ;
  assign \new_[63169]_  = ~A300 & ~A299;
  assign \new_[63172]_  = ~A302 & ~A301;
  assign \new_[63173]_  = \new_[63172]_  & \new_[63169]_ ;
  assign \new_[63174]_  = \new_[63173]_  & \new_[63166]_ ;
  assign \new_[63178]_  = ~A199 & ~A168;
  assign \new_[63179]_  = ~A170 & \new_[63178]_ ;
  assign \new_[63182]_  = ~A201 & A200;
  assign \new_[63185]_  = ~A203 & ~A202;
  assign \new_[63186]_  = \new_[63185]_  & \new_[63182]_ ;
  assign \new_[63187]_  = \new_[63186]_  & \new_[63179]_ ;
  assign \new_[63191]_  = ~A298 & ~A266;
  assign \new_[63192]_  = ~A265 & \new_[63191]_ ;
  assign \new_[63195]_  = ~A300 & A299;
  assign \new_[63198]_  = ~A302 & ~A301;
  assign \new_[63199]_  = \new_[63198]_  & \new_[63195]_ ;
  assign \new_[63200]_  = \new_[63199]_  & \new_[63192]_ ;
  assign \new_[63204]_  = A199 & ~A168;
  assign \new_[63205]_  = ~A170 & \new_[63204]_ ;
  assign \new_[63208]_  = A201 & ~A200;
  assign \new_[63211]_  = A267 & A202;
  assign \new_[63212]_  = \new_[63211]_  & \new_[63208]_ ;
  assign \new_[63213]_  = \new_[63212]_  & \new_[63205]_ ;
  assign \new_[63217]_  = A298 & ~A269;
  assign \new_[63218]_  = ~A268 & \new_[63217]_ ;
  assign \new_[63221]_  = ~A300 & ~A299;
  assign \new_[63224]_  = ~A302 & ~A301;
  assign \new_[63225]_  = \new_[63224]_  & \new_[63221]_ ;
  assign \new_[63226]_  = \new_[63225]_  & \new_[63218]_ ;
  assign \new_[63230]_  = A199 & ~A168;
  assign \new_[63231]_  = ~A170 & \new_[63230]_ ;
  assign \new_[63234]_  = A201 & ~A200;
  assign \new_[63237]_  = A267 & A202;
  assign \new_[63238]_  = \new_[63237]_  & \new_[63234]_ ;
  assign \new_[63239]_  = \new_[63238]_  & \new_[63231]_ ;
  assign \new_[63243]_  = ~A298 & ~A269;
  assign \new_[63244]_  = ~A268 & \new_[63243]_ ;
  assign \new_[63247]_  = ~A300 & A299;
  assign \new_[63250]_  = ~A302 & ~A301;
  assign \new_[63251]_  = \new_[63250]_  & \new_[63247]_ ;
  assign \new_[63252]_  = \new_[63251]_  & \new_[63244]_ ;
  assign \new_[63256]_  = A199 & ~A168;
  assign \new_[63257]_  = ~A170 & \new_[63256]_ ;
  assign \new_[63260]_  = A201 & ~A200;
  assign \new_[63263]_  = A267 & A203;
  assign \new_[63264]_  = \new_[63263]_  & \new_[63260]_ ;
  assign \new_[63265]_  = \new_[63264]_  & \new_[63257]_ ;
  assign \new_[63269]_  = A298 & ~A269;
  assign \new_[63270]_  = ~A268 & \new_[63269]_ ;
  assign \new_[63273]_  = ~A300 & ~A299;
  assign \new_[63276]_  = ~A302 & ~A301;
  assign \new_[63277]_  = \new_[63276]_  & \new_[63273]_ ;
  assign \new_[63278]_  = \new_[63277]_  & \new_[63270]_ ;
  assign \new_[63282]_  = A199 & ~A168;
  assign \new_[63283]_  = ~A170 & \new_[63282]_ ;
  assign \new_[63286]_  = A201 & ~A200;
  assign \new_[63289]_  = A267 & A203;
  assign \new_[63290]_  = \new_[63289]_  & \new_[63286]_ ;
  assign \new_[63291]_  = \new_[63290]_  & \new_[63283]_ ;
  assign \new_[63295]_  = ~A298 & ~A269;
  assign \new_[63296]_  = ~A268 & \new_[63295]_ ;
  assign \new_[63299]_  = ~A300 & A299;
  assign \new_[63302]_  = ~A302 & ~A301;
  assign \new_[63303]_  = \new_[63302]_  & \new_[63299]_ ;
  assign \new_[63304]_  = \new_[63303]_  & \new_[63296]_ ;
  assign \new_[63308]_  = A199 & ~A168;
  assign \new_[63309]_  = ~A170 & \new_[63308]_ ;
  assign \new_[63312]_  = ~A201 & ~A200;
  assign \new_[63315]_  = ~A203 & ~A202;
  assign \new_[63316]_  = \new_[63315]_  & \new_[63312]_ ;
  assign \new_[63317]_  = \new_[63316]_  & \new_[63309]_ ;
  assign \new_[63321]_  = ~A269 & ~A268;
  assign \new_[63322]_  = A267 & \new_[63321]_ ;
  assign \new_[63325]_  = ~A299 & A298;
  assign \new_[63328]_  = A301 & A300;
  assign \new_[63329]_  = \new_[63328]_  & \new_[63325]_ ;
  assign \new_[63330]_  = \new_[63329]_  & \new_[63322]_ ;
  assign \new_[63334]_  = A199 & ~A168;
  assign \new_[63335]_  = ~A170 & \new_[63334]_ ;
  assign \new_[63338]_  = ~A201 & ~A200;
  assign \new_[63341]_  = ~A203 & ~A202;
  assign \new_[63342]_  = \new_[63341]_  & \new_[63338]_ ;
  assign \new_[63343]_  = \new_[63342]_  & \new_[63335]_ ;
  assign \new_[63347]_  = ~A269 & ~A268;
  assign \new_[63348]_  = A267 & \new_[63347]_ ;
  assign \new_[63351]_  = ~A299 & A298;
  assign \new_[63354]_  = A302 & A300;
  assign \new_[63355]_  = \new_[63354]_  & \new_[63351]_ ;
  assign \new_[63356]_  = \new_[63355]_  & \new_[63348]_ ;
  assign \new_[63360]_  = A199 & ~A168;
  assign \new_[63361]_  = ~A170 & \new_[63360]_ ;
  assign \new_[63364]_  = ~A201 & ~A200;
  assign \new_[63367]_  = ~A203 & ~A202;
  assign \new_[63368]_  = \new_[63367]_  & \new_[63364]_ ;
  assign \new_[63369]_  = \new_[63368]_  & \new_[63361]_ ;
  assign \new_[63373]_  = ~A269 & ~A268;
  assign \new_[63374]_  = A267 & \new_[63373]_ ;
  assign \new_[63377]_  = A299 & ~A298;
  assign \new_[63380]_  = A301 & A300;
  assign \new_[63381]_  = \new_[63380]_  & \new_[63377]_ ;
  assign \new_[63382]_  = \new_[63381]_  & \new_[63374]_ ;
  assign \new_[63386]_  = A199 & ~A168;
  assign \new_[63387]_  = ~A170 & \new_[63386]_ ;
  assign \new_[63390]_  = ~A201 & ~A200;
  assign \new_[63393]_  = ~A203 & ~A202;
  assign \new_[63394]_  = \new_[63393]_  & \new_[63390]_ ;
  assign \new_[63395]_  = \new_[63394]_  & \new_[63387]_ ;
  assign \new_[63399]_  = ~A269 & ~A268;
  assign \new_[63400]_  = A267 & \new_[63399]_ ;
  assign \new_[63403]_  = A299 & ~A298;
  assign \new_[63406]_  = A302 & A300;
  assign \new_[63407]_  = \new_[63406]_  & \new_[63403]_ ;
  assign \new_[63408]_  = \new_[63407]_  & \new_[63400]_ ;
  assign \new_[63412]_  = A199 & ~A168;
  assign \new_[63413]_  = ~A170 & \new_[63412]_ ;
  assign \new_[63416]_  = ~A201 & ~A200;
  assign \new_[63419]_  = ~A203 & ~A202;
  assign \new_[63420]_  = \new_[63419]_  & \new_[63416]_ ;
  assign \new_[63421]_  = \new_[63420]_  & \new_[63413]_ ;
  assign \new_[63425]_  = A298 & A268;
  assign \new_[63426]_  = ~A267 & \new_[63425]_ ;
  assign \new_[63429]_  = ~A300 & ~A299;
  assign \new_[63432]_  = ~A302 & ~A301;
  assign \new_[63433]_  = \new_[63432]_  & \new_[63429]_ ;
  assign \new_[63434]_  = \new_[63433]_  & \new_[63426]_ ;
  assign \new_[63438]_  = A199 & ~A168;
  assign \new_[63439]_  = ~A170 & \new_[63438]_ ;
  assign \new_[63442]_  = ~A201 & ~A200;
  assign \new_[63445]_  = ~A203 & ~A202;
  assign \new_[63446]_  = \new_[63445]_  & \new_[63442]_ ;
  assign \new_[63447]_  = \new_[63446]_  & \new_[63439]_ ;
  assign \new_[63451]_  = ~A298 & A268;
  assign \new_[63452]_  = ~A267 & \new_[63451]_ ;
  assign \new_[63455]_  = ~A300 & A299;
  assign \new_[63458]_  = ~A302 & ~A301;
  assign \new_[63459]_  = \new_[63458]_  & \new_[63455]_ ;
  assign \new_[63460]_  = \new_[63459]_  & \new_[63452]_ ;
  assign \new_[63464]_  = A199 & ~A168;
  assign \new_[63465]_  = ~A170 & \new_[63464]_ ;
  assign \new_[63468]_  = ~A201 & ~A200;
  assign \new_[63471]_  = ~A203 & ~A202;
  assign \new_[63472]_  = \new_[63471]_  & \new_[63468]_ ;
  assign \new_[63473]_  = \new_[63472]_  & \new_[63465]_ ;
  assign \new_[63477]_  = A298 & A269;
  assign \new_[63478]_  = ~A267 & \new_[63477]_ ;
  assign \new_[63481]_  = ~A300 & ~A299;
  assign \new_[63484]_  = ~A302 & ~A301;
  assign \new_[63485]_  = \new_[63484]_  & \new_[63481]_ ;
  assign \new_[63486]_  = \new_[63485]_  & \new_[63478]_ ;
  assign \new_[63490]_  = A199 & ~A168;
  assign \new_[63491]_  = ~A170 & \new_[63490]_ ;
  assign \new_[63494]_  = ~A201 & ~A200;
  assign \new_[63497]_  = ~A203 & ~A202;
  assign \new_[63498]_  = \new_[63497]_  & \new_[63494]_ ;
  assign \new_[63499]_  = \new_[63498]_  & \new_[63491]_ ;
  assign \new_[63503]_  = ~A298 & A269;
  assign \new_[63504]_  = ~A267 & \new_[63503]_ ;
  assign \new_[63507]_  = ~A300 & A299;
  assign \new_[63510]_  = ~A302 & ~A301;
  assign \new_[63511]_  = \new_[63510]_  & \new_[63507]_ ;
  assign \new_[63512]_  = \new_[63511]_  & \new_[63504]_ ;
  assign \new_[63516]_  = A199 & ~A168;
  assign \new_[63517]_  = ~A170 & \new_[63516]_ ;
  assign \new_[63520]_  = ~A201 & ~A200;
  assign \new_[63523]_  = ~A203 & ~A202;
  assign \new_[63524]_  = \new_[63523]_  & \new_[63520]_ ;
  assign \new_[63525]_  = \new_[63524]_  & \new_[63517]_ ;
  assign \new_[63529]_  = A298 & A266;
  assign \new_[63530]_  = A265 & \new_[63529]_ ;
  assign \new_[63533]_  = ~A300 & ~A299;
  assign \new_[63536]_  = ~A302 & ~A301;
  assign \new_[63537]_  = \new_[63536]_  & \new_[63533]_ ;
  assign \new_[63538]_  = \new_[63537]_  & \new_[63530]_ ;
  assign \new_[63542]_  = A199 & ~A168;
  assign \new_[63543]_  = ~A170 & \new_[63542]_ ;
  assign \new_[63546]_  = ~A201 & ~A200;
  assign \new_[63549]_  = ~A203 & ~A202;
  assign \new_[63550]_  = \new_[63549]_  & \new_[63546]_ ;
  assign \new_[63551]_  = \new_[63550]_  & \new_[63543]_ ;
  assign \new_[63555]_  = ~A298 & A266;
  assign \new_[63556]_  = A265 & \new_[63555]_ ;
  assign \new_[63559]_  = ~A300 & A299;
  assign \new_[63562]_  = ~A302 & ~A301;
  assign \new_[63563]_  = \new_[63562]_  & \new_[63559]_ ;
  assign \new_[63564]_  = \new_[63563]_  & \new_[63556]_ ;
  assign \new_[63568]_  = A199 & ~A168;
  assign \new_[63569]_  = ~A170 & \new_[63568]_ ;
  assign \new_[63572]_  = ~A201 & ~A200;
  assign \new_[63575]_  = ~A203 & ~A202;
  assign \new_[63576]_  = \new_[63575]_  & \new_[63572]_ ;
  assign \new_[63577]_  = \new_[63576]_  & \new_[63569]_ ;
  assign \new_[63581]_  = A298 & ~A266;
  assign \new_[63582]_  = ~A265 & \new_[63581]_ ;
  assign \new_[63585]_  = ~A300 & ~A299;
  assign \new_[63588]_  = ~A302 & ~A301;
  assign \new_[63589]_  = \new_[63588]_  & \new_[63585]_ ;
  assign \new_[63590]_  = \new_[63589]_  & \new_[63582]_ ;
  assign \new_[63594]_  = A199 & ~A168;
  assign \new_[63595]_  = ~A170 & \new_[63594]_ ;
  assign \new_[63598]_  = ~A201 & ~A200;
  assign \new_[63601]_  = ~A203 & ~A202;
  assign \new_[63602]_  = \new_[63601]_  & \new_[63598]_ ;
  assign \new_[63603]_  = \new_[63602]_  & \new_[63595]_ ;
  assign \new_[63607]_  = ~A298 & ~A266;
  assign \new_[63608]_  = ~A265 & \new_[63607]_ ;
  assign \new_[63611]_  = ~A300 & A299;
  assign \new_[63614]_  = ~A302 & ~A301;
  assign \new_[63615]_  = \new_[63614]_  & \new_[63611]_ ;
  assign \new_[63616]_  = \new_[63615]_  & \new_[63608]_ ;
  assign \new_[63620]_  = A167 & A168;
  assign \new_[63621]_  = A169 & \new_[63620]_ ;
  assign \new_[63624]_  = A201 & ~A166;
  assign \new_[63627]_  = ~A203 & ~A202;
  assign \new_[63628]_  = \new_[63627]_  & \new_[63624]_ ;
  assign \new_[63629]_  = \new_[63628]_  & \new_[63621]_ ;
  assign \new_[63633]_  = ~A269 & ~A268;
  assign \new_[63634]_  = A267 & \new_[63633]_ ;
  assign \new_[63637]_  = ~A299 & A298;
  assign \new_[63640]_  = A301 & A300;
  assign \new_[63641]_  = \new_[63640]_  & \new_[63637]_ ;
  assign \new_[63642]_  = \new_[63641]_  & \new_[63634]_ ;
  assign \new_[63646]_  = A167 & A168;
  assign \new_[63647]_  = A169 & \new_[63646]_ ;
  assign \new_[63650]_  = A201 & ~A166;
  assign \new_[63653]_  = ~A203 & ~A202;
  assign \new_[63654]_  = \new_[63653]_  & \new_[63650]_ ;
  assign \new_[63655]_  = \new_[63654]_  & \new_[63647]_ ;
  assign \new_[63659]_  = ~A269 & ~A268;
  assign \new_[63660]_  = A267 & \new_[63659]_ ;
  assign \new_[63663]_  = ~A299 & A298;
  assign \new_[63666]_  = A302 & A300;
  assign \new_[63667]_  = \new_[63666]_  & \new_[63663]_ ;
  assign \new_[63668]_  = \new_[63667]_  & \new_[63660]_ ;
  assign \new_[63672]_  = A167 & A168;
  assign \new_[63673]_  = A169 & \new_[63672]_ ;
  assign \new_[63676]_  = A201 & ~A166;
  assign \new_[63679]_  = ~A203 & ~A202;
  assign \new_[63680]_  = \new_[63679]_  & \new_[63676]_ ;
  assign \new_[63681]_  = \new_[63680]_  & \new_[63673]_ ;
  assign \new_[63685]_  = ~A269 & ~A268;
  assign \new_[63686]_  = A267 & \new_[63685]_ ;
  assign \new_[63689]_  = A299 & ~A298;
  assign \new_[63692]_  = A301 & A300;
  assign \new_[63693]_  = \new_[63692]_  & \new_[63689]_ ;
  assign \new_[63694]_  = \new_[63693]_  & \new_[63686]_ ;
  assign \new_[63698]_  = A167 & A168;
  assign \new_[63699]_  = A169 & \new_[63698]_ ;
  assign \new_[63702]_  = A201 & ~A166;
  assign \new_[63705]_  = ~A203 & ~A202;
  assign \new_[63706]_  = \new_[63705]_  & \new_[63702]_ ;
  assign \new_[63707]_  = \new_[63706]_  & \new_[63699]_ ;
  assign \new_[63711]_  = ~A269 & ~A268;
  assign \new_[63712]_  = A267 & \new_[63711]_ ;
  assign \new_[63715]_  = A299 & ~A298;
  assign \new_[63718]_  = A302 & A300;
  assign \new_[63719]_  = \new_[63718]_  & \new_[63715]_ ;
  assign \new_[63720]_  = \new_[63719]_  & \new_[63712]_ ;
  assign \new_[63724]_  = A167 & A168;
  assign \new_[63725]_  = A169 & \new_[63724]_ ;
  assign \new_[63728]_  = A201 & ~A166;
  assign \new_[63731]_  = ~A203 & ~A202;
  assign \new_[63732]_  = \new_[63731]_  & \new_[63728]_ ;
  assign \new_[63733]_  = \new_[63732]_  & \new_[63725]_ ;
  assign \new_[63737]_  = A298 & A268;
  assign \new_[63738]_  = ~A267 & \new_[63737]_ ;
  assign \new_[63741]_  = ~A300 & ~A299;
  assign \new_[63744]_  = ~A302 & ~A301;
  assign \new_[63745]_  = \new_[63744]_  & \new_[63741]_ ;
  assign \new_[63746]_  = \new_[63745]_  & \new_[63738]_ ;
  assign \new_[63750]_  = A167 & A168;
  assign \new_[63751]_  = A169 & \new_[63750]_ ;
  assign \new_[63754]_  = A201 & ~A166;
  assign \new_[63757]_  = ~A203 & ~A202;
  assign \new_[63758]_  = \new_[63757]_  & \new_[63754]_ ;
  assign \new_[63759]_  = \new_[63758]_  & \new_[63751]_ ;
  assign \new_[63763]_  = ~A298 & A268;
  assign \new_[63764]_  = ~A267 & \new_[63763]_ ;
  assign \new_[63767]_  = ~A300 & A299;
  assign \new_[63770]_  = ~A302 & ~A301;
  assign \new_[63771]_  = \new_[63770]_  & \new_[63767]_ ;
  assign \new_[63772]_  = \new_[63771]_  & \new_[63764]_ ;
  assign \new_[63776]_  = A167 & A168;
  assign \new_[63777]_  = A169 & \new_[63776]_ ;
  assign \new_[63780]_  = A201 & ~A166;
  assign \new_[63783]_  = ~A203 & ~A202;
  assign \new_[63784]_  = \new_[63783]_  & \new_[63780]_ ;
  assign \new_[63785]_  = \new_[63784]_  & \new_[63777]_ ;
  assign \new_[63789]_  = A298 & A269;
  assign \new_[63790]_  = ~A267 & \new_[63789]_ ;
  assign \new_[63793]_  = ~A300 & ~A299;
  assign \new_[63796]_  = ~A302 & ~A301;
  assign \new_[63797]_  = \new_[63796]_  & \new_[63793]_ ;
  assign \new_[63798]_  = \new_[63797]_  & \new_[63790]_ ;
  assign \new_[63802]_  = A167 & A168;
  assign \new_[63803]_  = A169 & \new_[63802]_ ;
  assign \new_[63806]_  = A201 & ~A166;
  assign \new_[63809]_  = ~A203 & ~A202;
  assign \new_[63810]_  = \new_[63809]_  & \new_[63806]_ ;
  assign \new_[63811]_  = \new_[63810]_  & \new_[63803]_ ;
  assign \new_[63815]_  = ~A298 & A269;
  assign \new_[63816]_  = ~A267 & \new_[63815]_ ;
  assign \new_[63819]_  = ~A300 & A299;
  assign \new_[63822]_  = ~A302 & ~A301;
  assign \new_[63823]_  = \new_[63822]_  & \new_[63819]_ ;
  assign \new_[63824]_  = \new_[63823]_  & \new_[63816]_ ;
  assign \new_[63828]_  = A167 & A168;
  assign \new_[63829]_  = A169 & \new_[63828]_ ;
  assign \new_[63832]_  = A201 & ~A166;
  assign \new_[63835]_  = ~A203 & ~A202;
  assign \new_[63836]_  = \new_[63835]_  & \new_[63832]_ ;
  assign \new_[63837]_  = \new_[63836]_  & \new_[63829]_ ;
  assign \new_[63841]_  = A298 & A266;
  assign \new_[63842]_  = A265 & \new_[63841]_ ;
  assign \new_[63845]_  = ~A300 & ~A299;
  assign \new_[63848]_  = ~A302 & ~A301;
  assign \new_[63849]_  = \new_[63848]_  & \new_[63845]_ ;
  assign \new_[63850]_  = \new_[63849]_  & \new_[63842]_ ;
  assign \new_[63854]_  = A167 & A168;
  assign \new_[63855]_  = A169 & \new_[63854]_ ;
  assign \new_[63858]_  = A201 & ~A166;
  assign \new_[63861]_  = ~A203 & ~A202;
  assign \new_[63862]_  = \new_[63861]_  & \new_[63858]_ ;
  assign \new_[63863]_  = \new_[63862]_  & \new_[63855]_ ;
  assign \new_[63867]_  = ~A298 & A266;
  assign \new_[63868]_  = A265 & \new_[63867]_ ;
  assign \new_[63871]_  = ~A300 & A299;
  assign \new_[63874]_  = ~A302 & ~A301;
  assign \new_[63875]_  = \new_[63874]_  & \new_[63871]_ ;
  assign \new_[63876]_  = \new_[63875]_  & \new_[63868]_ ;
  assign \new_[63880]_  = A167 & A168;
  assign \new_[63881]_  = A169 & \new_[63880]_ ;
  assign \new_[63884]_  = A201 & ~A166;
  assign \new_[63887]_  = ~A203 & ~A202;
  assign \new_[63888]_  = \new_[63887]_  & \new_[63884]_ ;
  assign \new_[63889]_  = \new_[63888]_  & \new_[63881]_ ;
  assign \new_[63893]_  = A298 & ~A266;
  assign \new_[63894]_  = ~A265 & \new_[63893]_ ;
  assign \new_[63897]_  = ~A300 & ~A299;
  assign \new_[63900]_  = ~A302 & ~A301;
  assign \new_[63901]_  = \new_[63900]_  & \new_[63897]_ ;
  assign \new_[63902]_  = \new_[63901]_  & \new_[63894]_ ;
  assign \new_[63906]_  = A167 & A168;
  assign \new_[63907]_  = A169 & \new_[63906]_ ;
  assign \new_[63910]_  = A201 & ~A166;
  assign \new_[63913]_  = ~A203 & ~A202;
  assign \new_[63914]_  = \new_[63913]_  & \new_[63910]_ ;
  assign \new_[63915]_  = \new_[63914]_  & \new_[63907]_ ;
  assign \new_[63919]_  = ~A298 & ~A266;
  assign \new_[63920]_  = ~A265 & \new_[63919]_ ;
  assign \new_[63923]_  = ~A300 & A299;
  assign \new_[63926]_  = ~A302 & ~A301;
  assign \new_[63927]_  = \new_[63926]_  & \new_[63923]_ ;
  assign \new_[63928]_  = \new_[63927]_  & \new_[63920]_ ;
  assign \new_[63932]_  = A167 & A168;
  assign \new_[63933]_  = A169 & \new_[63932]_ ;
  assign \new_[63936]_  = ~A201 & ~A166;
  assign \new_[63939]_  = A267 & A202;
  assign \new_[63940]_  = \new_[63939]_  & \new_[63936]_ ;
  assign \new_[63941]_  = \new_[63940]_  & \new_[63933]_ ;
  assign \new_[63945]_  = A298 & ~A269;
  assign \new_[63946]_  = ~A268 & \new_[63945]_ ;
  assign \new_[63949]_  = ~A300 & ~A299;
  assign \new_[63952]_  = ~A302 & ~A301;
  assign \new_[63953]_  = \new_[63952]_  & \new_[63949]_ ;
  assign \new_[63954]_  = \new_[63953]_  & \new_[63946]_ ;
  assign \new_[63958]_  = A167 & A168;
  assign \new_[63959]_  = A169 & \new_[63958]_ ;
  assign \new_[63962]_  = ~A201 & ~A166;
  assign \new_[63965]_  = A267 & A202;
  assign \new_[63966]_  = \new_[63965]_  & \new_[63962]_ ;
  assign \new_[63967]_  = \new_[63966]_  & \new_[63959]_ ;
  assign \new_[63971]_  = ~A298 & ~A269;
  assign \new_[63972]_  = ~A268 & \new_[63971]_ ;
  assign \new_[63975]_  = ~A300 & A299;
  assign \new_[63978]_  = ~A302 & ~A301;
  assign \new_[63979]_  = \new_[63978]_  & \new_[63975]_ ;
  assign \new_[63980]_  = \new_[63979]_  & \new_[63972]_ ;
  assign \new_[63984]_  = A167 & A168;
  assign \new_[63985]_  = A169 & \new_[63984]_ ;
  assign \new_[63988]_  = ~A201 & ~A166;
  assign \new_[63991]_  = A267 & A203;
  assign \new_[63992]_  = \new_[63991]_  & \new_[63988]_ ;
  assign \new_[63993]_  = \new_[63992]_  & \new_[63985]_ ;
  assign \new_[63997]_  = A298 & ~A269;
  assign \new_[63998]_  = ~A268 & \new_[63997]_ ;
  assign \new_[64001]_  = ~A300 & ~A299;
  assign \new_[64004]_  = ~A302 & ~A301;
  assign \new_[64005]_  = \new_[64004]_  & \new_[64001]_ ;
  assign \new_[64006]_  = \new_[64005]_  & \new_[63998]_ ;
  assign \new_[64010]_  = A167 & A168;
  assign \new_[64011]_  = A169 & \new_[64010]_ ;
  assign \new_[64014]_  = ~A201 & ~A166;
  assign \new_[64017]_  = A267 & A203;
  assign \new_[64018]_  = \new_[64017]_  & \new_[64014]_ ;
  assign \new_[64019]_  = \new_[64018]_  & \new_[64011]_ ;
  assign \new_[64023]_  = ~A298 & ~A269;
  assign \new_[64024]_  = ~A268 & \new_[64023]_ ;
  assign \new_[64027]_  = ~A300 & A299;
  assign \new_[64030]_  = ~A302 & ~A301;
  assign \new_[64031]_  = \new_[64030]_  & \new_[64027]_ ;
  assign \new_[64032]_  = \new_[64031]_  & \new_[64024]_ ;
  assign \new_[64036]_  = A167 & A168;
  assign \new_[64037]_  = A169 & \new_[64036]_ ;
  assign \new_[64040]_  = A199 & ~A166;
  assign \new_[64043]_  = A267 & A200;
  assign \new_[64044]_  = \new_[64043]_  & \new_[64040]_ ;
  assign \new_[64045]_  = \new_[64044]_  & \new_[64037]_ ;
  assign \new_[64049]_  = A298 & ~A269;
  assign \new_[64050]_  = ~A268 & \new_[64049]_ ;
  assign \new_[64053]_  = ~A300 & ~A299;
  assign \new_[64056]_  = ~A302 & ~A301;
  assign \new_[64057]_  = \new_[64056]_  & \new_[64053]_ ;
  assign \new_[64058]_  = \new_[64057]_  & \new_[64050]_ ;
  assign \new_[64062]_  = A167 & A168;
  assign \new_[64063]_  = A169 & \new_[64062]_ ;
  assign \new_[64066]_  = A199 & ~A166;
  assign \new_[64069]_  = A267 & A200;
  assign \new_[64070]_  = \new_[64069]_  & \new_[64066]_ ;
  assign \new_[64071]_  = \new_[64070]_  & \new_[64063]_ ;
  assign \new_[64075]_  = ~A298 & ~A269;
  assign \new_[64076]_  = ~A268 & \new_[64075]_ ;
  assign \new_[64079]_  = ~A300 & A299;
  assign \new_[64082]_  = ~A302 & ~A301;
  assign \new_[64083]_  = \new_[64082]_  & \new_[64079]_ ;
  assign \new_[64084]_  = \new_[64083]_  & \new_[64076]_ ;
  assign \new_[64088]_  = A167 & A168;
  assign \new_[64089]_  = A169 & \new_[64088]_ ;
  assign \new_[64092]_  = ~A199 & ~A166;
  assign \new_[64095]_  = A201 & A200;
  assign \new_[64096]_  = \new_[64095]_  & \new_[64092]_ ;
  assign \new_[64097]_  = \new_[64096]_  & \new_[64089]_ ;
  assign \new_[64101]_  = A266 & ~A265;
  assign \new_[64102]_  = A202 & \new_[64101]_ ;
  assign \new_[64105]_  = A268 & A267;
  assign \new_[64108]_  = A301 & ~A300;
  assign \new_[64109]_  = \new_[64108]_  & \new_[64105]_ ;
  assign \new_[64110]_  = \new_[64109]_  & \new_[64102]_ ;
  assign \new_[64114]_  = A167 & A168;
  assign \new_[64115]_  = A169 & \new_[64114]_ ;
  assign \new_[64118]_  = ~A199 & ~A166;
  assign \new_[64121]_  = A201 & A200;
  assign \new_[64122]_  = \new_[64121]_  & \new_[64118]_ ;
  assign \new_[64123]_  = \new_[64122]_  & \new_[64115]_ ;
  assign \new_[64127]_  = A266 & ~A265;
  assign \new_[64128]_  = A202 & \new_[64127]_ ;
  assign \new_[64131]_  = A268 & A267;
  assign \new_[64134]_  = A302 & ~A300;
  assign \new_[64135]_  = \new_[64134]_  & \new_[64131]_ ;
  assign \new_[64136]_  = \new_[64135]_  & \new_[64128]_ ;
  assign \new_[64140]_  = A167 & A168;
  assign \new_[64141]_  = A169 & \new_[64140]_ ;
  assign \new_[64144]_  = ~A199 & ~A166;
  assign \new_[64147]_  = A201 & A200;
  assign \new_[64148]_  = \new_[64147]_  & \new_[64144]_ ;
  assign \new_[64149]_  = \new_[64148]_  & \new_[64141]_ ;
  assign \new_[64153]_  = A266 & ~A265;
  assign \new_[64154]_  = A202 & \new_[64153]_ ;
  assign \new_[64157]_  = A268 & A267;
  assign \new_[64160]_  = A299 & A298;
  assign \new_[64161]_  = \new_[64160]_  & \new_[64157]_ ;
  assign \new_[64162]_  = \new_[64161]_  & \new_[64154]_ ;
  assign \new_[64166]_  = A167 & A168;
  assign \new_[64167]_  = A169 & \new_[64166]_ ;
  assign \new_[64170]_  = ~A199 & ~A166;
  assign \new_[64173]_  = A201 & A200;
  assign \new_[64174]_  = \new_[64173]_  & \new_[64170]_ ;
  assign \new_[64175]_  = \new_[64174]_  & \new_[64167]_ ;
  assign \new_[64179]_  = A266 & ~A265;
  assign \new_[64180]_  = A202 & \new_[64179]_ ;
  assign \new_[64183]_  = A268 & A267;
  assign \new_[64186]_  = ~A299 & ~A298;
  assign \new_[64187]_  = \new_[64186]_  & \new_[64183]_ ;
  assign \new_[64188]_  = \new_[64187]_  & \new_[64180]_ ;
  assign \new_[64192]_  = A167 & A168;
  assign \new_[64193]_  = A169 & \new_[64192]_ ;
  assign \new_[64196]_  = ~A199 & ~A166;
  assign \new_[64199]_  = A201 & A200;
  assign \new_[64200]_  = \new_[64199]_  & \new_[64196]_ ;
  assign \new_[64201]_  = \new_[64200]_  & \new_[64193]_ ;
  assign \new_[64205]_  = A266 & ~A265;
  assign \new_[64206]_  = A202 & \new_[64205]_ ;
  assign \new_[64209]_  = A269 & A267;
  assign \new_[64212]_  = A301 & ~A300;
  assign \new_[64213]_  = \new_[64212]_  & \new_[64209]_ ;
  assign \new_[64214]_  = \new_[64213]_  & \new_[64206]_ ;
  assign \new_[64218]_  = A167 & A168;
  assign \new_[64219]_  = A169 & \new_[64218]_ ;
  assign \new_[64222]_  = ~A199 & ~A166;
  assign \new_[64225]_  = A201 & A200;
  assign \new_[64226]_  = \new_[64225]_  & \new_[64222]_ ;
  assign \new_[64227]_  = \new_[64226]_  & \new_[64219]_ ;
  assign \new_[64231]_  = A266 & ~A265;
  assign \new_[64232]_  = A202 & \new_[64231]_ ;
  assign \new_[64235]_  = A269 & A267;
  assign \new_[64238]_  = A302 & ~A300;
  assign \new_[64239]_  = \new_[64238]_  & \new_[64235]_ ;
  assign \new_[64240]_  = \new_[64239]_  & \new_[64232]_ ;
  assign \new_[64244]_  = A167 & A168;
  assign \new_[64245]_  = A169 & \new_[64244]_ ;
  assign \new_[64248]_  = ~A199 & ~A166;
  assign \new_[64251]_  = A201 & A200;
  assign \new_[64252]_  = \new_[64251]_  & \new_[64248]_ ;
  assign \new_[64253]_  = \new_[64252]_  & \new_[64245]_ ;
  assign \new_[64257]_  = A266 & ~A265;
  assign \new_[64258]_  = A202 & \new_[64257]_ ;
  assign \new_[64261]_  = A269 & A267;
  assign \new_[64264]_  = A299 & A298;
  assign \new_[64265]_  = \new_[64264]_  & \new_[64261]_ ;
  assign \new_[64266]_  = \new_[64265]_  & \new_[64258]_ ;
  assign \new_[64270]_  = A167 & A168;
  assign \new_[64271]_  = A169 & \new_[64270]_ ;
  assign \new_[64274]_  = ~A199 & ~A166;
  assign \new_[64277]_  = A201 & A200;
  assign \new_[64278]_  = \new_[64277]_  & \new_[64274]_ ;
  assign \new_[64279]_  = \new_[64278]_  & \new_[64271]_ ;
  assign \new_[64283]_  = A266 & ~A265;
  assign \new_[64284]_  = A202 & \new_[64283]_ ;
  assign \new_[64287]_  = A269 & A267;
  assign \new_[64290]_  = ~A299 & ~A298;
  assign \new_[64291]_  = \new_[64290]_  & \new_[64287]_ ;
  assign \new_[64292]_  = \new_[64291]_  & \new_[64284]_ ;
  assign \new_[64296]_  = A167 & A168;
  assign \new_[64297]_  = A169 & \new_[64296]_ ;
  assign \new_[64300]_  = ~A199 & ~A166;
  assign \new_[64303]_  = A201 & A200;
  assign \new_[64304]_  = \new_[64303]_  & \new_[64300]_ ;
  assign \new_[64305]_  = \new_[64304]_  & \new_[64297]_ ;
  assign \new_[64309]_  = ~A266 & A265;
  assign \new_[64310]_  = A202 & \new_[64309]_ ;
  assign \new_[64313]_  = A268 & A267;
  assign \new_[64316]_  = A301 & ~A300;
  assign \new_[64317]_  = \new_[64316]_  & \new_[64313]_ ;
  assign \new_[64318]_  = \new_[64317]_  & \new_[64310]_ ;
  assign \new_[64322]_  = A167 & A168;
  assign \new_[64323]_  = A169 & \new_[64322]_ ;
  assign \new_[64326]_  = ~A199 & ~A166;
  assign \new_[64329]_  = A201 & A200;
  assign \new_[64330]_  = \new_[64329]_  & \new_[64326]_ ;
  assign \new_[64331]_  = \new_[64330]_  & \new_[64323]_ ;
  assign \new_[64335]_  = ~A266 & A265;
  assign \new_[64336]_  = A202 & \new_[64335]_ ;
  assign \new_[64339]_  = A268 & A267;
  assign \new_[64342]_  = A302 & ~A300;
  assign \new_[64343]_  = \new_[64342]_  & \new_[64339]_ ;
  assign \new_[64344]_  = \new_[64343]_  & \new_[64336]_ ;
  assign \new_[64348]_  = A167 & A168;
  assign \new_[64349]_  = A169 & \new_[64348]_ ;
  assign \new_[64352]_  = ~A199 & ~A166;
  assign \new_[64355]_  = A201 & A200;
  assign \new_[64356]_  = \new_[64355]_  & \new_[64352]_ ;
  assign \new_[64357]_  = \new_[64356]_  & \new_[64349]_ ;
  assign \new_[64361]_  = ~A266 & A265;
  assign \new_[64362]_  = A202 & \new_[64361]_ ;
  assign \new_[64365]_  = A268 & A267;
  assign \new_[64368]_  = A299 & A298;
  assign \new_[64369]_  = \new_[64368]_  & \new_[64365]_ ;
  assign \new_[64370]_  = \new_[64369]_  & \new_[64362]_ ;
  assign \new_[64374]_  = A167 & A168;
  assign \new_[64375]_  = A169 & \new_[64374]_ ;
  assign \new_[64378]_  = ~A199 & ~A166;
  assign \new_[64381]_  = A201 & A200;
  assign \new_[64382]_  = \new_[64381]_  & \new_[64378]_ ;
  assign \new_[64383]_  = \new_[64382]_  & \new_[64375]_ ;
  assign \new_[64387]_  = ~A266 & A265;
  assign \new_[64388]_  = A202 & \new_[64387]_ ;
  assign \new_[64391]_  = A268 & A267;
  assign \new_[64394]_  = ~A299 & ~A298;
  assign \new_[64395]_  = \new_[64394]_  & \new_[64391]_ ;
  assign \new_[64396]_  = \new_[64395]_  & \new_[64388]_ ;
  assign \new_[64400]_  = A167 & A168;
  assign \new_[64401]_  = A169 & \new_[64400]_ ;
  assign \new_[64404]_  = ~A199 & ~A166;
  assign \new_[64407]_  = A201 & A200;
  assign \new_[64408]_  = \new_[64407]_  & \new_[64404]_ ;
  assign \new_[64409]_  = \new_[64408]_  & \new_[64401]_ ;
  assign \new_[64413]_  = ~A266 & A265;
  assign \new_[64414]_  = A202 & \new_[64413]_ ;
  assign \new_[64417]_  = A269 & A267;
  assign \new_[64420]_  = A301 & ~A300;
  assign \new_[64421]_  = \new_[64420]_  & \new_[64417]_ ;
  assign \new_[64422]_  = \new_[64421]_  & \new_[64414]_ ;
  assign \new_[64426]_  = A167 & A168;
  assign \new_[64427]_  = A169 & \new_[64426]_ ;
  assign \new_[64430]_  = ~A199 & ~A166;
  assign \new_[64433]_  = A201 & A200;
  assign \new_[64434]_  = \new_[64433]_  & \new_[64430]_ ;
  assign \new_[64435]_  = \new_[64434]_  & \new_[64427]_ ;
  assign \new_[64439]_  = ~A266 & A265;
  assign \new_[64440]_  = A202 & \new_[64439]_ ;
  assign \new_[64443]_  = A269 & A267;
  assign \new_[64446]_  = A302 & ~A300;
  assign \new_[64447]_  = \new_[64446]_  & \new_[64443]_ ;
  assign \new_[64448]_  = \new_[64447]_  & \new_[64440]_ ;
  assign \new_[64452]_  = A167 & A168;
  assign \new_[64453]_  = A169 & \new_[64452]_ ;
  assign \new_[64456]_  = ~A199 & ~A166;
  assign \new_[64459]_  = A201 & A200;
  assign \new_[64460]_  = \new_[64459]_  & \new_[64456]_ ;
  assign \new_[64461]_  = \new_[64460]_  & \new_[64453]_ ;
  assign \new_[64465]_  = ~A266 & A265;
  assign \new_[64466]_  = A202 & \new_[64465]_ ;
  assign \new_[64469]_  = A269 & A267;
  assign \new_[64472]_  = A299 & A298;
  assign \new_[64473]_  = \new_[64472]_  & \new_[64469]_ ;
  assign \new_[64474]_  = \new_[64473]_  & \new_[64466]_ ;
  assign \new_[64478]_  = A167 & A168;
  assign \new_[64479]_  = A169 & \new_[64478]_ ;
  assign \new_[64482]_  = ~A199 & ~A166;
  assign \new_[64485]_  = A201 & A200;
  assign \new_[64486]_  = \new_[64485]_  & \new_[64482]_ ;
  assign \new_[64487]_  = \new_[64486]_  & \new_[64479]_ ;
  assign \new_[64491]_  = ~A266 & A265;
  assign \new_[64492]_  = A202 & \new_[64491]_ ;
  assign \new_[64495]_  = A269 & A267;
  assign \new_[64498]_  = ~A299 & ~A298;
  assign \new_[64499]_  = \new_[64498]_  & \new_[64495]_ ;
  assign \new_[64500]_  = \new_[64499]_  & \new_[64492]_ ;
  assign \new_[64504]_  = A167 & A168;
  assign \new_[64505]_  = A169 & \new_[64504]_ ;
  assign \new_[64508]_  = ~A199 & ~A166;
  assign \new_[64511]_  = A201 & A200;
  assign \new_[64512]_  = \new_[64511]_  & \new_[64508]_ ;
  assign \new_[64513]_  = \new_[64512]_  & \new_[64505]_ ;
  assign \new_[64517]_  = A266 & ~A265;
  assign \new_[64518]_  = A203 & \new_[64517]_ ;
  assign \new_[64521]_  = A268 & A267;
  assign \new_[64524]_  = A301 & ~A300;
  assign \new_[64525]_  = \new_[64524]_  & \new_[64521]_ ;
  assign \new_[64526]_  = \new_[64525]_  & \new_[64518]_ ;
  assign \new_[64530]_  = A167 & A168;
  assign \new_[64531]_  = A169 & \new_[64530]_ ;
  assign \new_[64534]_  = ~A199 & ~A166;
  assign \new_[64537]_  = A201 & A200;
  assign \new_[64538]_  = \new_[64537]_  & \new_[64534]_ ;
  assign \new_[64539]_  = \new_[64538]_  & \new_[64531]_ ;
  assign \new_[64543]_  = A266 & ~A265;
  assign \new_[64544]_  = A203 & \new_[64543]_ ;
  assign \new_[64547]_  = A268 & A267;
  assign \new_[64550]_  = A302 & ~A300;
  assign \new_[64551]_  = \new_[64550]_  & \new_[64547]_ ;
  assign \new_[64552]_  = \new_[64551]_  & \new_[64544]_ ;
  assign \new_[64556]_  = A167 & A168;
  assign \new_[64557]_  = A169 & \new_[64556]_ ;
  assign \new_[64560]_  = ~A199 & ~A166;
  assign \new_[64563]_  = A201 & A200;
  assign \new_[64564]_  = \new_[64563]_  & \new_[64560]_ ;
  assign \new_[64565]_  = \new_[64564]_  & \new_[64557]_ ;
  assign \new_[64569]_  = A266 & ~A265;
  assign \new_[64570]_  = A203 & \new_[64569]_ ;
  assign \new_[64573]_  = A268 & A267;
  assign \new_[64576]_  = A299 & A298;
  assign \new_[64577]_  = \new_[64576]_  & \new_[64573]_ ;
  assign \new_[64578]_  = \new_[64577]_  & \new_[64570]_ ;
  assign \new_[64582]_  = A167 & A168;
  assign \new_[64583]_  = A169 & \new_[64582]_ ;
  assign \new_[64586]_  = ~A199 & ~A166;
  assign \new_[64589]_  = A201 & A200;
  assign \new_[64590]_  = \new_[64589]_  & \new_[64586]_ ;
  assign \new_[64591]_  = \new_[64590]_  & \new_[64583]_ ;
  assign \new_[64595]_  = A266 & ~A265;
  assign \new_[64596]_  = A203 & \new_[64595]_ ;
  assign \new_[64599]_  = A268 & A267;
  assign \new_[64602]_  = ~A299 & ~A298;
  assign \new_[64603]_  = \new_[64602]_  & \new_[64599]_ ;
  assign \new_[64604]_  = \new_[64603]_  & \new_[64596]_ ;
  assign \new_[64608]_  = A167 & A168;
  assign \new_[64609]_  = A169 & \new_[64608]_ ;
  assign \new_[64612]_  = ~A199 & ~A166;
  assign \new_[64615]_  = A201 & A200;
  assign \new_[64616]_  = \new_[64615]_  & \new_[64612]_ ;
  assign \new_[64617]_  = \new_[64616]_  & \new_[64609]_ ;
  assign \new_[64621]_  = A266 & ~A265;
  assign \new_[64622]_  = A203 & \new_[64621]_ ;
  assign \new_[64625]_  = A269 & A267;
  assign \new_[64628]_  = A301 & ~A300;
  assign \new_[64629]_  = \new_[64628]_  & \new_[64625]_ ;
  assign \new_[64630]_  = \new_[64629]_  & \new_[64622]_ ;
  assign \new_[64634]_  = A167 & A168;
  assign \new_[64635]_  = A169 & \new_[64634]_ ;
  assign \new_[64638]_  = ~A199 & ~A166;
  assign \new_[64641]_  = A201 & A200;
  assign \new_[64642]_  = \new_[64641]_  & \new_[64638]_ ;
  assign \new_[64643]_  = \new_[64642]_  & \new_[64635]_ ;
  assign \new_[64647]_  = A266 & ~A265;
  assign \new_[64648]_  = A203 & \new_[64647]_ ;
  assign \new_[64651]_  = A269 & A267;
  assign \new_[64654]_  = A302 & ~A300;
  assign \new_[64655]_  = \new_[64654]_  & \new_[64651]_ ;
  assign \new_[64656]_  = \new_[64655]_  & \new_[64648]_ ;
  assign \new_[64660]_  = A167 & A168;
  assign \new_[64661]_  = A169 & \new_[64660]_ ;
  assign \new_[64664]_  = ~A199 & ~A166;
  assign \new_[64667]_  = A201 & A200;
  assign \new_[64668]_  = \new_[64667]_  & \new_[64664]_ ;
  assign \new_[64669]_  = \new_[64668]_  & \new_[64661]_ ;
  assign \new_[64673]_  = A266 & ~A265;
  assign \new_[64674]_  = A203 & \new_[64673]_ ;
  assign \new_[64677]_  = A269 & A267;
  assign \new_[64680]_  = A299 & A298;
  assign \new_[64681]_  = \new_[64680]_  & \new_[64677]_ ;
  assign \new_[64682]_  = \new_[64681]_  & \new_[64674]_ ;
  assign \new_[64686]_  = A167 & A168;
  assign \new_[64687]_  = A169 & \new_[64686]_ ;
  assign \new_[64690]_  = ~A199 & ~A166;
  assign \new_[64693]_  = A201 & A200;
  assign \new_[64694]_  = \new_[64693]_  & \new_[64690]_ ;
  assign \new_[64695]_  = \new_[64694]_  & \new_[64687]_ ;
  assign \new_[64699]_  = A266 & ~A265;
  assign \new_[64700]_  = A203 & \new_[64699]_ ;
  assign \new_[64703]_  = A269 & A267;
  assign \new_[64706]_  = ~A299 & ~A298;
  assign \new_[64707]_  = \new_[64706]_  & \new_[64703]_ ;
  assign \new_[64708]_  = \new_[64707]_  & \new_[64700]_ ;
  assign \new_[64712]_  = A167 & A168;
  assign \new_[64713]_  = A169 & \new_[64712]_ ;
  assign \new_[64716]_  = ~A199 & ~A166;
  assign \new_[64719]_  = A201 & A200;
  assign \new_[64720]_  = \new_[64719]_  & \new_[64716]_ ;
  assign \new_[64721]_  = \new_[64720]_  & \new_[64713]_ ;
  assign \new_[64725]_  = ~A266 & A265;
  assign \new_[64726]_  = A203 & \new_[64725]_ ;
  assign \new_[64729]_  = A268 & A267;
  assign \new_[64732]_  = A301 & ~A300;
  assign \new_[64733]_  = \new_[64732]_  & \new_[64729]_ ;
  assign \new_[64734]_  = \new_[64733]_  & \new_[64726]_ ;
  assign \new_[64738]_  = A167 & A168;
  assign \new_[64739]_  = A169 & \new_[64738]_ ;
  assign \new_[64742]_  = ~A199 & ~A166;
  assign \new_[64745]_  = A201 & A200;
  assign \new_[64746]_  = \new_[64745]_  & \new_[64742]_ ;
  assign \new_[64747]_  = \new_[64746]_  & \new_[64739]_ ;
  assign \new_[64751]_  = ~A266 & A265;
  assign \new_[64752]_  = A203 & \new_[64751]_ ;
  assign \new_[64755]_  = A268 & A267;
  assign \new_[64758]_  = A302 & ~A300;
  assign \new_[64759]_  = \new_[64758]_  & \new_[64755]_ ;
  assign \new_[64760]_  = \new_[64759]_  & \new_[64752]_ ;
  assign \new_[64764]_  = A167 & A168;
  assign \new_[64765]_  = A169 & \new_[64764]_ ;
  assign \new_[64768]_  = ~A199 & ~A166;
  assign \new_[64771]_  = A201 & A200;
  assign \new_[64772]_  = \new_[64771]_  & \new_[64768]_ ;
  assign \new_[64773]_  = \new_[64772]_  & \new_[64765]_ ;
  assign \new_[64777]_  = ~A266 & A265;
  assign \new_[64778]_  = A203 & \new_[64777]_ ;
  assign \new_[64781]_  = A268 & A267;
  assign \new_[64784]_  = A299 & A298;
  assign \new_[64785]_  = \new_[64784]_  & \new_[64781]_ ;
  assign \new_[64786]_  = \new_[64785]_  & \new_[64778]_ ;
  assign \new_[64790]_  = A167 & A168;
  assign \new_[64791]_  = A169 & \new_[64790]_ ;
  assign \new_[64794]_  = ~A199 & ~A166;
  assign \new_[64797]_  = A201 & A200;
  assign \new_[64798]_  = \new_[64797]_  & \new_[64794]_ ;
  assign \new_[64799]_  = \new_[64798]_  & \new_[64791]_ ;
  assign \new_[64803]_  = ~A266 & A265;
  assign \new_[64804]_  = A203 & \new_[64803]_ ;
  assign \new_[64807]_  = A268 & A267;
  assign \new_[64810]_  = ~A299 & ~A298;
  assign \new_[64811]_  = \new_[64810]_  & \new_[64807]_ ;
  assign \new_[64812]_  = \new_[64811]_  & \new_[64804]_ ;
  assign \new_[64816]_  = A167 & A168;
  assign \new_[64817]_  = A169 & \new_[64816]_ ;
  assign \new_[64820]_  = ~A199 & ~A166;
  assign \new_[64823]_  = A201 & A200;
  assign \new_[64824]_  = \new_[64823]_  & \new_[64820]_ ;
  assign \new_[64825]_  = \new_[64824]_  & \new_[64817]_ ;
  assign \new_[64829]_  = ~A266 & A265;
  assign \new_[64830]_  = A203 & \new_[64829]_ ;
  assign \new_[64833]_  = A269 & A267;
  assign \new_[64836]_  = A301 & ~A300;
  assign \new_[64837]_  = \new_[64836]_  & \new_[64833]_ ;
  assign \new_[64838]_  = \new_[64837]_  & \new_[64830]_ ;
  assign \new_[64842]_  = A167 & A168;
  assign \new_[64843]_  = A169 & \new_[64842]_ ;
  assign \new_[64846]_  = ~A199 & ~A166;
  assign \new_[64849]_  = A201 & A200;
  assign \new_[64850]_  = \new_[64849]_  & \new_[64846]_ ;
  assign \new_[64851]_  = \new_[64850]_  & \new_[64843]_ ;
  assign \new_[64855]_  = ~A266 & A265;
  assign \new_[64856]_  = A203 & \new_[64855]_ ;
  assign \new_[64859]_  = A269 & A267;
  assign \new_[64862]_  = A302 & ~A300;
  assign \new_[64863]_  = \new_[64862]_  & \new_[64859]_ ;
  assign \new_[64864]_  = \new_[64863]_  & \new_[64856]_ ;
  assign \new_[64868]_  = A167 & A168;
  assign \new_[64869]_  = A169 & \new_[64868]_ ;
  assign \new_[64872]_  = ~A199 & ~A166;
  assign \new_[64875]_  = A201 & A200;
  assign \new_[64876]_  = \new_[64875]_  & \new_[64872]_ ;
  assign \new_[64877]_  = \new_[64876]_  & \new_[64869]_ ;
  assign \new_[64881]_  = ~A266 & A265;
  assign \new_[64882]_  = A203 & \new_[64881]_ ;
  assign \new_[64885]_  = A269 & A267;
  assign \new_[64888]_  = A299 & A298;
  assign \new_[64889]_  = \new_[64888]_  & \new_[64885]_ ;
  assign \new_[64890]_  = \new_[64889]_  & \new_[64882]_ ;
  assign \new_[64894]_  = A167 & A168;
  assign \new_[64895]_  = A169 & \new_[64894]_ ;
  assign \new_[64898]_  = ~A199 & ~A166;
  assign \new_[64901]_  = A201 & A200;
  assign \new_[64902]_  = \new_[64901]_  & \new_[64898]_ ;
  assign \new_[64903]_  = \new_[64902]_  & \new_[64895]_ ;
  assign \new_[64907]_  = ~A266 & A265;
  assign \new_[64908]_  = A203 & \new_[64907]_ ;
  assign \new_[64911]_  = A269 & A267;
  assign \new_[64914]_  = ~A299 & ~A298;
  assign \new_[64915]_  = \new_[64914]_  & \new_[64911]_ ;
  assign \new_[64916]_  = \new_[64915]_  & \new_[64908]_ ;
  assign \new_[64920]_  = A167 & A168;
  assign \new_[64921]_  = A169 & \new_[64920]_ ;
  assign \new_[64924]_  = A199 & ~A166;
  assign \new_[64927]_  = A201 & ~A200;
  assign \new_[64928]_  = \new_[64927]_  & \new_[64924]_ ;
  assign \new_[64929]_  = \new_[64928]_  & \new_[64921]_ ;
  assign \new_[64933]_  = A266 & ~A265;
  assign \new_[64934]_  = A202 & \new_[64933]_ ;
  assign \new_[64937]_  = A268 & A267;
  assign \new_[64940]_  = A301 & ~A300;
  assign \new_[64941]_  = \new_[64940]_  & \new_[64937]_ ;
  assign \new_[64942]_  = \new_[64941]_  & \new_[64934]_ ;
  assign \new_[64946]_  = A167 & A168;
  assign \new_[64947]_  = A169 & \new_[64946]_ ;
  assign \new_[64950]_  = A199 & ~A166;
  assign \new_[64953]_  = A201 & ~A200;
  assign \new_[64954]_  = \new_[64953]_  & \new_[64950]_ ;
  assign \new_[64955]_  = \new_[64954]_  & \new_[64947]_ ;
  assign \new_[64959]_  = A266 & ~A265;
  assign \new_[64960]_  = A202 & \new_[64959]_ ;
  assign \new_[64963]_  = A268 & A267;
  assign \new_[64966]_  = A302 & ~A300;
  assign \new_[64967]_  = \new_[64966]_  & \new_[64963]_ ;
  assign \new_[64968]_  = \new_[64967]_  & \new_[64960]_ ;
  assign \new_[64972]_  = A167 & A168;
  assign \new_[64973]_  = A169 & \new_[64972]_ ;
  assign \new_[64976]_  = A199 & ~A166;
  assign \new_[64979]_  = A201 & ~A200;
  assign \new_[64980]_  = \new_[64979]_  & \new_[64976]_ ;
  assign \new_[64981]_  = \new_[64980]_  & \new_[64973]_ ;
  assign \new_[64985]_  = A266 & ~A265;
  assign \new_[64986]_  = A202 & \new_[64985]_ ;
  assign \new_[64989]_  = A268 & A267;
  assign \new_[64992]_  = A299 & A298;
  assign \new_[64993]_  = \new_[64992]_  & \new_[64989]_ ;
  assign \new_[64994]_  = \new_[64993]_  & \new_[64986]_ ;
  assign \new_[64998]_  = A167 & A168;
  assign \new_[64999]_  = A169 & \new_[64998]_ ;
  assign \new_[65002]_  = A199 & ~A166;
  assign \new_[65005]_  = A201 & ~A200;
  assign \new_[65006]_  = \new_[65005]_  & \new_[65002]_ ;
  assign \new_[65007]_  = \new_[65006]_  & \new_[64999]_ ;
  assign \new_[65011]_  = A266 & ~A265;
  assign \new_[65012]_  = A202 & \new_[65011]_ ;
  assign \new_[65015]_  = A268 & A267;
  assign \new_[65018]_  = ~A299 & ~A298;
  assign \new_[65019]_  = \new_[65018]_  & \new_[65015]_ ;
  assign \new_[65020]_  = \new_[65019]_  & \new_[65012]_ ;
  assign \new_[65024]_  = A167 & A168;
  assign \new_[65025]_  = A169 & \new_[65024]_ ;
  assign \new_[65028]_  = A199 & ~A166;
  assign \new_[65031]_  = A201 & ~A200;
  assign \new_[65032]_  = \new_[65031]_  & \new_[65028]_ ;
  assign \new_[65033]_  = \new_[65032]_  & \new_[65025]_ ;
  assign \new_[65037]_  = A266 & ~A265;
  assign \new_[65038]_  = A202 & \new_[65037]_ ;
  assign \new_[65041]_  = A269 & A267;
  assign \new_[65044]_  = A301 & ~A300;
  assign \new_[65045]_  = \new_[65044]_  & \new_[65041]_ ;
  assign \new_[65046]_  = \new_[65045]_  & \new_[65038]_ ;
  assign \new_[65050]_  = A167 & A168;
  assign \new_[65051]_  = A169 & \new_[65050]_ ;
  assign \new_[65054]_  = A199 & ~A166;
  assign \new_[65057]_  = A201 & ~A200;
  assign \new_[65058]_  = \new_[65057]_  & \new_[65054]_ ;
  assign \new_[65059]_  = \new_[65058]_  & \new_[65051]_ ;
  assign \new_[65063]_  = A266 & ~A265;
  assign \new_[65064]_  = A202 & \new_[65063]_ ;
  assign \new_[65067]_  = A269 & A267;
  assign \new_[65070]_  = A302 & ~A300;
  assign \new_[65071]_  = \new_[65070]_  & \new_[65067]_ ;
  assign \new_[65072]_  = \new_[65071]_  & \new_[65064]_ ;
  assign \new_[65076]_  = A167 & A168;
  assign \new_[65077]_  = A169 & \new_[65076]_ ;
  assign \new_[65080]_  = A199 & ~A166;
  assign \new_[65083]_  = A201 & ~A200;
  assign \new_[65084]_  = \new_[65083]_  & \new_[65080]_ ;
  assign \new_[65085]_  = \new_[65084]_  & \new_[65077]_ ;
  assign \new_[65089]_  = A266 & ~A265;
  assign \new_[65090]_  = A202 & \new_[65089]_ ;
  assign \new_[65093]_  = A269 & A267;
  assign \new_[65096]_  = A299 & A298;
  assign \new_[65097]_  = \new_[65096]_  & \new_[65093]_ ;
  assign \new_[65098]_  = \new_[65097]_  & \new_[65090]_ ;
  assign \new_[65102]_  = A167 & A168;
  assign \new_[65103]_  = A169 & \new_[65102]_ ;
  assign \new_[65106]_  = A199 & ~A166;
  assign \new_[65109]_  = A201 & ~A200;
  assign \new_[65110]_  = \new_[65109]_  & \new_[65106]_ ;
  assign \new_[65111]_  = \new_[65110]_  & \new_[65103]_ ;
  assign \new_[65115]_  = A266 & ~A265;
  assign \new_[65116]_  = A202 & \new_[65115]_ ;
  assign \new_[65119]_  = A269 & A267;
  assign \new_[65122]_  = ~A299 & ~A298;
  assign \new_[65123]_  = \new_[65122]_  & \new_[65119]_ ;
  assign \new_[65124]_  = \new_[65123]_  & \new_[65116]_ ;
  assign \new_[65128]_  = A167 & A168;
  assign \new_[65129]_  = A169 & \new_[65128]_ ;
  assign \new_[65132]_  = A199 & ~A166;
  assign \new_[65135]_  = A201 & ~A200;
  assign \new_[65136]_  = \new_[65135]_  & \new_[65132]_ ;
  assign \new_[65137]_  = \new_[65136]_  & \new_[65129]_ ;
  assign \new_[65141]_  = ~A266 & A265;
  assign \new_[65142]_  = A202 & \new_[65141]_ ;
  assign \new_[65145]_  = A268 & A267;
  assign \new_[65148]_  = A301 & ~A300;
  assign \new_[65149]_  = \new_[65148]_  & \new_[65145]_ ;
  assign \new_[65150]_  = \new_[65149]_  & \new_[65142]_ ;
  assign \new_[65154]_  = A167 & A168;
  assign \new_[65155]_  = A169 & \new_[65154]_ ;
  assign \new_[65158]_  = A199 & ~A166;
  assign \new_[65161]_  = A201 & ~A200;
  assign \new_[65162]_  = \new_[65161]_  & \new_[65158]_ ;
  assign \new_[65163]_  = \new_[65162]_  & \new_[65155]_ ;
  assign \new_[65167]_  = ~A266 & A265;
  assign \new_[65168]_  = A202 & \new_[65167]_ ;
  assign \new_[65171]_  = A268 & A267;
  assign \new_[65174]_  = A302 & ~A300;
  assign \new_[65175]_  = \new_[65174]_  & \new_[65171]_ ;
  assign \new_[65176]_  = \new_[65175]_  & \new_[65168]_ ;
  assign \new_[65180]_  = A167 & A168;
  assign \new_[65181]_  = A169 & \new_[65180]_ ;
  assign \new_[65184]_  = A199 & ~A166;
  assign \new_[65187]_  = A201 & ~A200;
  assign \new_[65188]_  = \new_[65187]_  & \new_[65184]_ ;
  assign \new_[65189]_  = \new_[65188]_  & \new_[65181]_ ;
  assign \new_[65193]_  = ~A266 & A265;
  assign \new_[65194]_  = A202 & \new_[65193]_ ;
  assign \new_[65197]_  = A268 & A267;
  assign \new_[65200]_  = A299 & A298;
  assign \new_[65201]_  = \new_[65200]_  & \new_[65197]_ ;
  assign \new_[65202]_  = \new_[65201]_  & \new_[65194]_ ;
  assign \new_[65206]_  = A167 & A168;
  assign \new_[65207]_  = A169 & \new_[65206]_ ;
  assign \new_[65210]_  = A199 & ~A166;
  assign \new_[65213]_  = A201 & ~A200;
  assign \new_[65214]_  = \new_[65213]_  & \new_[65210]_ ;
  assign \new_[65215]_  = \new_[65214]_  & \new_[65207]_ ;
  assign \new_[65219]_  = ~A266 & A265;
  assign \new_[65220]_  = A202 & \new_[65219]_ ;
  assign \new_[65223]_  = A268 & A267;
  assign \new_[65226]_  = ~A299 & ~A298;
  assign \new_[65227]_  = \new_[65226]_  & \new_[65223]_ ;
  assign \new_[65228]_  = \new_[65227]_  & \new_[65220]_ ;
  assign \new_[65232]_  = A167 & A168;
  assign \new_[65233]_  = A169 & \new_[65232]_ ;
  assign \new_[65236]_  = A199 & ~A166;
  assign \new_[65239]_  = A201 & ~A200;
  assign \new_[65240]_  = \new_[65239]_  & \new_[65236]_ ;
  assign \new_[65241]_  = \new_[65240]_  & \new_[65233]_ ;
  assign \new_[65245]_  = ~A266 & A265;
  assign \new_[65246]_  = A202 & \new_[65245]_ ;
  assign \new_[65249]_  = A269 & A267;
  assign \new_[65252]_  = A301 & ~A300;
  assign \new_[65253]_  = \new_[65252]_  & \new_[65249]_ ;
  assign \new_[65254]_  = \new_[65253]_  & \new_[65246]_ ;
  assign \new_[65258]_  = A167 & A168;
  assign \new_[65259]_  = A169 & \new_[65258]_ ;
  assign \new_[65262]_  = A199 & ~A166;
  assign \new_[65265]_  = A201 & ~A200;
  assign \new_[65266]_  = \new_[65265]_  & \new_[65262]_ ;
  assign \new_[65267]_  = \new_[65266]_  & \new_[65259]_ ;
  assign \new_[65271]_  = ~A266 & A265;
  assign \new_[65272]_  = A202 & \new_[65271]_ ;
  assign \new_[65275]_  = A269 & A267;
  assign \new_[65278]_  = A302 & ~A300;
  assign \new_[65279]_  = \new_[65278]_  & \new_[65275]_ ;
  assign \new_[65280]_  = \new_[65279]_  & \new_[65272]_ ;
  assign \new_[65284]_  = A167 & A168;
  assign \new_[65285]_  = A169 & \new_[65284]_ ;
  assign \new_[65288]_  = A199 & ~A166;
  assign \new_[65291]_  = A201 & ~A200;
  assign \new_[65292]_  = \new_[65291]_  & \new_[65288]_ ;
  assign \new_[65293]_  = \new_[65292]_  & \new_[65285]_ ;
  assign \new_[65297]_  = ~A266 & A265;
  assign \new_[65298]_  = A202 & \new_[65297]_ ;
  assign \new_[65301]_  = A269 & A267;
  assign \new_[65304]_  = A299 & A298;
  assign \new_[65305]_  = \new_[65304]_  & \new_[65301]_ ;
  assign \new_[65306]_  = \new_[65305]_  & \new_[65298]_ ;
  assign \new_[65310]_  = A167 & A168;
  assign \new_[65311]_  = A169 & \new_[65310]_ ;
  assign \new_[65314]_  = A199 & ~A166;
  assign \new_[65317]_  = A201 & ~A200;
  assign \new_[65318]_  = \new_[65317]_  & \new_[65314]_ ;
  assign \new_[65319]_  = \new_[65318]_  & \new_[65311]_ ;
  assign \new_[65323]_  = ~A266 & A265;
  assign \new_[65324]_  = A202 & \new_[65323]_ ;
  assign \new_[65327]_  = A269 & A267;
  assign \new_[65330]_  = ~A299 & ~A298;
  assign \new_[65331]_  = \new_[65330]_  & \new_[65327]_ ;
  assign \new_[65332]_  = \new_[65331]_  & \new_[65324]_ ;
  assign \new_[65336]_  = A167 & A168;
  assign \new_[65337]_  = A169 & \new_[65336]_ ;
  assign \new_[65340]_  = A199 & ~A166;
  assign \new_[65343]_  = A201 & ~A200;
  assign \new_[65344]_  = \new_[65343]_  & \new_[65340]_ ;
  assign \new_[65345]_  = \new_[65344]_  & \new_[65337]_ ;
  assign \new_[65349]_  = A266 & ~A265;
  assign \new_[65350]_  = A203 & \new_[65349]_ ;
  assign \new_[65353]_  = A268 & A267;
  assign \new_[65356]_  = A301 & ~A300;
  assign \new_[65357]_  = \new_[65356]_  & \new_[65353]_ ;
  assign \new_[65358]_  = \new_[65357]_  & \new_[65350]_ ;
  assign \new_[65362]_  = A167 & A168;
  assign \new_[65363]_  = A169 & \new_[65362]_ ;
  assign \new_[65366]_  = A199 & ~A166;
  assign \new_[65369]_  = A201 & ~A200;
  assign \new_[65370]_  = \new_[65369]_  & \new_[65366]_ ;
  assign \new_[65371]_  = \new_[65370]_  & \new_[65363]_ ;
  assign \new_[65375]_  = A266 & ~A265;
  assign \new_[65376]_  = A203 & \new_[65375]_ ;
  assign \new_[65379]_  = A268 & A267;
  assign \new_[65382]_  = A302 & ~A300;
  assign \new_[65383]_  = \new_[65382]_  & \new_[65379]_ ;
  assign \new_[65384]_  = \new_[65383]_  & \new_[65376]_ ;
  assign \new_[65388]_  = A167 & A168;
  assign \new_[65389]_  = A169 & \new_[65388]_ ;
  assign \new_[65392]_  = A199 & ~A166;
  assign \new_[65395]_  = A201 & ~A200;
  assign \new_[65396]_  = \new_[65395]_  & \new_[65392]_ ;
  assign \new_[65397]_  = \new_[65396]_  & \new_[65389]_ ;
  assign \new_[65401]_  = A266 & ~A265;
  assign \new_[65402]_  = A203 & \new_[65401]_ ;
  assign \new_[65405]_  = A268 & A267;
  assign \new_[65408]_  = A299 & A298;
  assign \new_[65409]_  = \new_[65408]_  & \new_[65405]_ ;
  assign \new_[65410]_  = \new_[65409]_  & \new_[65402]_ ;
  assign \new_[65414]_  = A167 & A168;
  assign \new_[65415]_  = A169 & \new_[65414]_ ;
  assign \new_[65418]_  = A199 & ~A166;
  assign \new_[65421]_  = A201 & ~A200;
  assign \new_[65422]_  = \new_[65421]_  & \new_[65418]_ ;
  assign \new_[65423]_  = \new_[65422]_  & \new_[65415]_ ;
  assign \new_[65427]_  = A266 & ~A265;
  assign \new_[65428]_  = A203 & \new_[65427]_ ;
  assign \new_[65431]_  = A268 & A267;
  assign \new_[65434]_  = ~A299 & ~A298;
  assign \new_[65435]_  = \new_[65434]_  & \new_[65431]_ ;
  assign \new_[65436]_  = \new_[65435]_  & \new_[65428]_ ;
  assign \new_[65440]_  = A167 & A168;
  assign \new_[65441]_  = A169 & \new_[65440]_ ;
  assign \new_[65444]_  = A199 & ~A166;
  assign \new_[65447]_  = A201 & ~A200;
  assign \new_[65448]_  = \new_[65447]_  & \new_[65444]_ ;
  assign \new_[65449]_  = \new_[65448]_  & \new_[65441]_ ;
  assign \new_[65453]_  = A266 & ~A265;
  assign \new_[65454]_  = A203 & \new_[65453]_ ;
  assign \new_[65457]_  = A269 & A267;
  assign \new_[65460]_  = A301 & ~A300;
  assign \new_[65461]_  = \new_[65460]_  & \new_[65457]_ ;
  assign \new_[65462]_  = \new_[65461]_  & \new_[65454]_ ;
  assign \new_[65466]_  = A167 & A168;
  assign \new_[65467]_  = A169 & \new_[65466]_ ;
  assign \new_[65470]_  = A199 & ~A166;
  assign \new_[65473]_  = A201 & ~A200;
  assign \new_[65474]_  = \new_[65473]_  & \new_[65470]_ ;
  assign \new_[65475]_  = \new_[65474]_  & \new_[65467]_ ;
  assign \new_[65479]_  = A266 & ~A265;
  assign \new_[65480]_  = A203 & \new_[65479]_ ;
  assign \new_[65483]_  = A269 & A267;
  assign \new_[65486]_  = A302 & ~A300;
  assign \new_[65487]_  = \new_[65486]_  & \new_[65483]_ ;
  assign \new_[65488]_  = \new_[65487]_  & \new_[65480]_ ;
  assign \new_[65492]_  = A167 & A168;
  assign \new_[65493]_  = A169 & \new_[65492]_ ;
  assign \new_[65496]_  = A199 & ~A166;
  assign \new_[65499]_  = A201 & ~A200;
  assign \new_[65500]_  = \new_[65499]_  & \new_[65496]_ ;
  assign \new_[65501]_  = \new_[65500]_  & \new_[65493]_ ;
  assign \new_[65505]_  = A266 & ~A265;
  assign \new_[65506]_  = A203 & \new_[65505]_ ;
  assign \new_[65509]_  = A269 & A267;
  assign \new_[65512]_  = A299 & A298;
  assign \new_[65513]_  = \new_[65512]_  & \new_[65509]_ ;
  assign \new_[65514]_  = \new_[65513]_  & \new_[65506]_ ;
  assign \new_[65518]_  = A167 & A168;
  assign \new_[65519]_  = A169 & \new_[65518]_ ;
  assign \new_[65522]_  = A199 & ~A166;
  assign \new_[65525]_  = A201 & ~A200;
  assign \new_[65526]_  = \new_[65525]_  & \new_[65522]_ ;
  assign \new_[65527]_  = \new_[65526]_  & \new_[65519]_ ;
  assign \new_[65531]_  = A266 & ~A265;
  assign \new_[65532]_  = A203 & \new_[65531]_ ;
  assign \new_[65535]_  = A269 & A267;
  assign \new_[65538]_  = ~A299 & ~A298;
  assign \new_[65539]_  = \new_[65538]_  & \new_[65535]_ ;
  assign \new_[65540]_  = \new_[65539]_  & \new_[65532]_ ;
  assign \new_[65544]_  = A167 & A168;
  assign \new_[65545]_  = A169 & \new_[65544]_ ;
  assign \new_[65548]_  = A199 & ~A166;
  assign \new_[65551]_  = A201 & ~A200;
  assign \new_[65552]_  = \new_[65551]_  & \new_[65548]_ ;
  assign \new_[65553]_  = \new_[65552]_  & \new_[65545]_ ;
  assign \new_[65557]_  = ~A266 & A265;
  assign \new_[65558]_  = A203 & \new_[65557]_ ;
  assign \new_[65561]_  = A268 & A267;
  assign \new_[65564]_  = A301 & ~A300;
  assign \new_[65565]_  = \new_[65564]_  & \new_[65561]_ ;
  assign \new_[65566]_  = \new_[65565]_  & \new_[65558]_ ;
  assign \new_[65570]_  = A167 & A168;
  assign \new_[65571]_  = A169 & \new_[65570]_ ;
  assign \new_[65574]_  = A199 & ~A166;
  assign \new_[65577]_  = A201 & ~A200;
  assign \new_[65578]_  = \new_[65577]_  & \new_[65574]_ ;
  assign \new_[65579]_  = \new_[65578]_  & \new_[65571]_ ;
  assign \new_[65583]_  = ~A266 & A265;
  assign \new_[65584]_  = A203 & \new_[65583]_ ;
  assign \new_[65587]_  = A268 & A267;
  assign \new_[65590]_  = A302 & ~A300;
  assign \new_[65591]_  = \new_[65590]_  & \new_[65587]_ ;
  assign \new_[65592]_  = \new_[65591]_  & \new_[65584]_ ;
  assign \new_[65596]_  = A167 & A168;
  assign \new_[65597]_  = A169 & \new_[65596]_ ;
  assign \new_[65600]_  = A199 & ~A166;
  assign \new_[65603]_  = A201 & ~A200;
  assign \new_[65604]_  = \new_[65603]_  & \new_[65600]_ ;
  assign \new_[65605]_  = \new_[65604]_  & \new_[65597]_ ;
  assign \new_[65609]_  = ~A266 & A265;
  assign \new_[65610]_  = A203 & \new_[65609]_ ;
  assign \new_[65613]_  = A268 & A267;
  assign \new_[65616]_  = A299 & A298;
  assign \new_[65617]_  = \new_[65616]_  & \new_[65613]_ ;
  assign \new_[65618]_  = \new_[65617]_  & \new_[65610]_ ;
  assign \new_[65622]_  = A167 & A168;
  assign \new_[65623]_  = A169 & \new_[65622]_ ;
  assign \new_[65626]_  = A199 & ~A166;
  assign \new_[65629]_  = A201 & ~A200;
  assign \new_[65630]_  = \new_[65629]_  & \new_[65626]_ ;
  assign \new_[65631]_  = \new_[65630]_  & \new_[65623]_ ;
  assign \new_[65635]_  = ~A266 & A265;
  assign \new_[65636]_  = A203 & \new_[65635]_ ;
  assign \new_[65639]_  = A268 & A267;
  assign \new_[65642]_  = ~A299 & ~A298;
  assign \new_[65643]_  = \new_[65642]_  & \new_[65639]_ ;
  assign \new_[65644]_  = \new_[65643]_  & \new_[65636]_ ;
  assign \new_[65648]_  = A167 & A168;
  assign \new_[65649]_  = A169 & \new_[65648]_ ;
  assign \new_[65652]_  = A199 & ~A166;
  assign \new_[65655]_  = A201 & ~A200;
  assign \new_[65656]_  = \new_[65655]_  & \new_[65652]_ ;
  assign \new_[65657]_  = \new_[65656]_  & \new_[65649]_ ;
  assign \new_[65661]_  = ~A266 & A265;
  assign \new_[65662]_  = A203 & \new_[65661]_ ;
  assign \new_[65665]_  = A269 & A267;
  assign \new_[65668]_  = A301 & ~A300;
  assign \new_[65669]_  = \new_[65668]_  & \new_[65665]_ ;
  assign \new_[65670]_  = \new_[65669]_  & \new_[65662]_ ;
  assign \new_[65674]_  = A167 & A168;
  assign \new_[65675]_  = A169 & \new_[65674]_ ;
  assign \new_[65678]_  = A199 & ~A166;
  assign \new_[65681]_  = A201 & ~A200;
  assign \new_[65682]_  = \new_[65681]_  & \new_[65678]_ ;
  assign \new_[65683]_  = \new_[65682]_  & \new_[65675]_ ;
  assign \new_[65687]_  = ~A266 & A265;
  assign \new_[65688]_  = A203 & \new_[65687]_ ;
  assign \new_[65691]_  = A269 & A267;
  assign \new_[65694]_  = A302 & ~A300;
  assign \new_[65695]_  = \new_[65694]_  & \new_[65691]_ ;
  assign \new_[65696]_  = \new_[65695]_  & \new_[65688]_ ;
  assign \new_[65700]_  = A167 & A168;
  assign \new_[65701]_  = A169 & \new_[65700]_ ;
  assign \new_[65704]_  = A199 & ~A166;
  assign \new_[65707]_  = A201 & ~A200;
  assign \new_[65708]_  = \new_[65707]_  & \new_[65704]_ ;
  assign \new_[65709]_  = \new_[65708]_  & \new_[65701]_ ;
  assign \new_[65713]_  = ~A266 & A265;
  assign \new_[65714]_  = A203 & \new_[65713]_ ;
  assign \new_[65717]_  = A269 & A267;
  assign \new_[65720]_  = A299 & A298;
  assign \new_[65721]_  = \new_[65720]_  & \new_[65717]_ ;
  assign \new_[65722]_  = \new_[65721]_  & \new_[65714]_ ;
  assign \new_[65726]_  = A167 & A168;
  assign \new_[65727]_  = A169 & \new_[65726]_ ;
  assign \new_[65730]_  = A199 & ~A166;
  assign \new_[65733]_  = A201 & ~A200;
  assign \new_[65734]_  = \new_[65733]_  & \new_[65730]_ ;
  assign \new_[65735]_  = \new_[65734]_  & \new_[65727]_ ;
  assign \new_[65739]_  = ~A266 & A265;
  assign \new_[65740]_  = A203 & \new_[65739]_ ;
  assign \new_[65743]_  = A269 & A267;
  assign \new_[65746]_  = ~A299 & ~A298;
  assign \new_[65747]_  = \new_[65746]_  & \new_[65743]_ ;
  assign \new_[65748]_  = \new_[65747]_  & \new_[65740]_ ;
  assign \new_[65752]_  = A167 & A168;
  assign \new_[65753]_  = A169 & \new_[65752]_ ;
  assign \new_[65756]_  = ~A199 & ~A166;
  assign \new_[65759]_  = A267 & ~A200;
  assign \new_[65760]_  = \new_[65759]_  & \new_[65756]_ ;
  assign \new_[65761]_  = \new_[65760]_  & \new_[65753]_ ;
  assign \new_[65765]_  = A298 & ~A269;
  assign \new_[65766]_  = ~A268 & \new_[65765]_ ;
  assign \new_[65769]_  = ~A300 & ~A299;
  assign \new_[65772]_  = ~A302 & ~A301;
  assign \new_[65773]_  = \new_[65772]_  & \new_[65769]_ ;
  assign \new_[65774]_  = \new_[65773]_  & \new_[65766]_ ;
  assign \new_[65778]_  = A167 & A168;
  assign \new_[65779]_  = A169 & \new_[65778]_ ;
  assign \new_[65782]_  = ~A199 & ~A166;
  assign \new_[65785]_  = A267 & ~A200;
  assign \new_[65786]_  = \new_[65785]_  & \new_[65782]_ ;
  assign \new_[65787]_  = \new_[65786]_  & \new_[65779]_ ;
  assign \new_[65791]_  = ~A298 & ~A269;
  assign \new_[65792]_  = ~A268 & \new_[65791]_ ;
  assign \new_[65795]_  = ~A300 & A299;
  assign \new_[65798]_  = ~A302 & ~A301;
  assign \new_[65799]_  = \new_[65798]_  & \new_[65795]_ ;
  assign \new_[65800]_  = \new_[65799]_  & \new_[65792]_ ;
  assign \new_[65804]_  = ~A167 & A168;
  assign \new_[65805]_  = A169 & \new_[65804]_ ;
  assign \new_[65808]_  = A201 & A166;
  assign \new_[65811]_  = ~A203 & ~A202;
  assign \new_[65812]_  = \new_[65811]_  & \new_[65808]_ ;
  assign \new_[65813]_  = \new_[65812]_  & \new_[65805]_ ;
  assign \new_[65817]_  = ~A269 & ~A268;
  assign \new_[65818]_  = A267 & \new_[65817]_ ;
  assign \new_[65821]_  = ~A299 & A298;
  assign \new_[65824]_  = A301 & A300;
  assign \new_[65825]_  = \new_[65824]_  & \new_[65821]_ ;
  assign \new_[65826]_  = \new_[65825]_  & \new_[65818]_ ;
  assign \new_[65830]_  = ~A167 & A168;
  assign \new_[65831]_  = A169 & \new_[65830]_ ;
  assign \new_[65834]_  = A201 & A166;
  assign \new_[65837]_  = ~A203 & ~A202;
  assign \new_[65838]_  = \new_[65837]_  & \new_[65834]_ ;
  assign \new_[65839]_  = \new_[65838]_  & \new_[65831]_ ;
  assign \new_[65843]_  = ~A269 & ~A268;
  assign \new_[65844]_  = A267 & \new_[65843]_ ;
  assign \new_[65847]_  = ~A299 & A298;
  assign \new_[65850]_  = A302 & A300;
  assign \new_[65851]_  = \new_[65850]_  & \new_[65847]_ ;
  assign \new_[65852]_  = \new_[65851]_  & \new_[65844]_ ;
  assign \new_[65856]_  = ~A167 & A168;
  assign \new_[65857]_  = A169 & \new_[65856]_ ;
  assign \new_[65860]_  = A201 & A166;
  assign \new_[65863]_  = ~A203 & ~A202;
  assign \new_[65864]_  = \new_[65863]_  & \new_[65860]_ ;
  assign \new_[65865]_  = \new_[65864]_  & \new_[65857]_ ;
  assign \new_[65869]_  = ~A269 & ~A268;
  assign \new_[65870]_  = A267 & \new_[65869]_ ;
  assign \new_[65873]_  = A299 & ~A298;
  assign \new_[65876]_  = A301 & A300;
  assign \new_[65877]_  = \new_[65876]_  & \new_[65873]_ ;
  assign \new_[65878]_  = \new_[65877]_  & \new_[65870]_ ;
  assign \new_[65882]_  = ~A167 & A168;
  assign \new_[65883]_  = A169 & \new_[65882]_ ;
  assign \new_[65886]_  = A201 & A166;
  assign \new_[65889]_  = ~A203 & ~A202;
  assign \new_[65890]_  = \new_[65889]_  & \new_[65886]_ ;
  assign \new_[65891]_  = \new_[65890]_  & \new_[65883]_ ;
  assign \new_[65895]_  = ~A269 & ~A268;
  assign \new_[65896]_  = A267 & \new_[65895]_ ;
  assign \new_[65899]_  = A299 & ~A298;
  assign \new_[65902]_  = A302 & A300;
  assign \new_[65903]_  = \new_[65902]_  & \new_[65899]_ ;
  assign \new_[65904]_  = \new_[65903]_  & \new_[65896]_ ;
  assign \new_[65908]_  = ~A167 & A168;
  assign \new_[65909]_  = A169 & \new_[65908]_ ;
  assign \new_[65912]_  = A201 & A166;
  assign \new_[65915]_  = ~A203 & ~A202;
  assign \new_[65916]_  = \new_[65915]_  & \new_[65912]_ ;
  assign \new_[65917]_  = \new_[65916]_  & \new_[65909]_ ;
  assign \new_[65921]_  = A298 & A268;
  assign \new_[65922]_  = ~A267 & \new_[65921]_ ;
  assign \new_[65925]_  = ~A300 & ~A299;
  assign \new_[65928]_  = ~A302 & ~A301;
  assign \new_[65929]_  = \new_[65928]_  & \new_[65925]_ ;
  assign \new_[65930]_  = \new_[65929]_  & \new_[65922]_ ;
  assign \new_[65934]_  = ~A167 & A168;
  assign \new_[65935]_  = A169 & \new_[65934]_ ;
  assign \new_[65938]_  = A201 & A166;
  assign \new_[65941]_  = ~A203 & ~A202;
  assign \new_[65942]_  = \new_[65941]_  & \new_[65938]_ ;
  assign \new_[65943]_  = \new_[65942]_  & \new_[65935]_ ;
  assign \new_[65947]_  = ~A298 & A268;
  assign \new_[65948]_  = ~A267 & \new_[65947]_ ;
  assign \new_[65951]_  = ~A300 & A299;
  assign \new_[65954]_  = ~A302 & ~A301;
  assign \new_[65955]_  = \new_[65954]_  & \new_[65951]_ ;
  assign \new_[65956]_  = \new_[65955]_  & \new_[65948]_ ;
  assign \new_[65960]_  = ~A167 & A168;
  assign \new_[65961]_  = A169 & \new_[65960]_ ;
  assign \new_[65964]_  = A201 & A166;
  assign \new_[65967]_  = ~A203 & ~A202;
  assign \new_[65968]_  = \new_[65967]_  & \new_[65964]_ ;
  assign \new_[65969]_  = \new_[65968]_  & \new_[65961]_ ;
  assign \new_[65973]_  = A298 & A269;
  assign \new_[65974]_  = ~A267 & \new_[65973]_ ;
  assign \new_[65977]_  = ~A300 & ~A299;
  assign \new_[65980]_  = ~A302 & ~A301;
  assign \new_[65981]_  = \new_[65980]_  & \new_[65977]_ ;
  assign \new_[65982]_  = \new_[65981]_  & \new_[65974]_ ;
  assign \new_[65986]_  = ~A167 & A168;
  assign \new_[65987]_  = A169 & \new_[65986]_ ;
  assign \new_[65990]_  = A201 & A166;
  assign \new_[65993]_  = ~A203 & ~A202;
  assign \new_[65994]_  = \new_[65993]_  & \new_[65990]_ ;
  assign \new_[65995]_  = \new_[65994]_  & \new_[65987]_ ;
  assign \new_[65999]_  = ~A298 & A269;
  assign \new_[66000]_  = ~A267 & \new_[65999]_ ;
  assign \new_[66003]_  = ~A300 & A299;
  assign \new_[66006]_  = ~A302 & ~A301;
  assign \new_[66007]_  = \new_[66006]_  & \new_[66003]_ ;
  assign \new_[66008]_  = \new_[66007]_  & \new_[66000]_ ;
  assign \new_[66012]_  = ~A167 & A168;
  assign \new_[66013]_  = A169 & \new_[66012]_ ;
  assign \new_[66016]_  = A201 & A166;
  assign \new_[66019]_  = ~A203 & ~A202;
  assign \new_[66020]_  = \new_[66019]_  & \new_[66016]_ ;
  assign \new_[66021]_  = \new_[66020]_  & \new_[66013]_ ;
  assign \new_[66025]_  = A298 & A266;
  assign \new_[66026]_  = A265 & \new_[66025]_ ;
  assign \new_[66029]_  = ~A300 & ~A299;
  assign \new_[66032]_  = ~A302 & ~A301;
  assign \new_[66033]_  = \new_[66032]_  & \new_[66029]_ ;
  assign \new_[66034]_  = \new_[66033]_  & \new_[66026]_ ;
  assign \new_[66038]_  = ~A167 & A168;
  assign \new_[66039]_  = A169 & \new_[66038]_ ;
  assign \new_[66042]_  = A201 & A166;
  assign \new_[66045]_  = ~A203 & ~A202;
  assign \new_[66046]_  = \new_[66045]_  & \new_[66042]_ ;
  assign \new_[66047]_  = \new_[66046]_  & \new_[66039]_ ;
  assign \new_[66051]_  = ~A298 & A266;
  assign \new_[66052]_  = A265 & \new_[66051]_ ;
  assign \new_[66055]_  = ~A300 & A299;
  assign \new_[66058]_  = ~A302 & ~A301;
  assign \new_[66059]_  = \new_[66058]_  & \new_[66055]_ ;
  assign \new_[66060]_  = \new_[66059]_  & \new_[66052]_ ;
  assign \new_[66064]_  = ~A167 & A168;
  assign \new_[66065]_  = A169 & \new_[66064]_ ;
  assign \new_[66068]_  = A201 & A166;
  assign \new_[66071]_  = ~A203 & ~A202;
  assign \new_[66072]_  = \new_[66071]_  & \new_[66068]_ ;
  assign \new_[66073]_  = \new_[66072]_  & \new_[66065]_ ;
  assign \new_[66077]_  = A298 & ~A266;
  assign \new_[66078]_  = ~A265 & \new_[66077]_ ;
  assign \new_[66081]_  = ~A300 & ~A299;
  assign \new_[66084]_  = ~A302 & ~A301;
  assign \new_[66085]_  = \new_[66084]_  & \new_[66081]_ ;
  assign \new_[66086]_  = \new_[66085]_  & \new_[66078]_ ;
  assign \new_[66090]_  = ~A167 & A168;
  assign \new_[66091]_  = A169 & \new_[66090]_ ;
  assign \new_[66094]_  = A201 & A166;
  assign \new_[66097]_  = ~A203 & ~A202;
  assign \new_[66098]_  = \new_[66097]_  & \new_[66094]_ ;
  assign \new_[66099]_  = \new_[66098]_  & \new_[66091]_ ;
  assign \new_[66103]_  = ~A298 & ~A266;
  assign \new_[66104]_  = ~A265 & \new_[66103]_ ;
  assign \new_[66107]_  = ~A300 & A299;
  assign \new_[66110]_  = ~A302 & ~A301;
  assign \new_[66111]_  = \new_[66110]_  & \new_[66107]_ ;
  assign \new_[66112]_  = \new_[66111]_  & \new_[66104]_ ;
  assign \new_[66116]_  = ~A167 & A168;
  assign \new_[66117]_  = A169 & \new_[66116]_ ;
  assign \new_[66120]_  = ~A201 & A166;
  assign \new_[66123]_  = A267 & A202;
  assign \new_[66124]_  = \new_[66123]_  & \new_[66120]_ ;
  assign \new_[66125]_  = \new_[66124]_  & \new_[66117]_ ;
  assign \new_[66129]_  = A298 & ~A269;
  assign \new_[66130]_  = ~A268 & \new_[66129]_ ;
  assign \new_[66133]_  = ~A300 & ~A299;
  assign \new_[66136]_  = ~A302 & ~A301;
  assign \new_[66137]_  = \new_[66136]_  & \new_[66133]_ ;
  assign \new_[66138]_  = \new_[66137]_  & \new_[66130]_ ;
  assign \new_[66142]_  = ~A167 & A168;
  assign \new_[66143]_  = A169 & \new_[66142]_ ;
  assign \new_[66146]_  = ~A201 & A166;
  assign \new_[66149]_  = A267 & A202;
  assign \new_[66150]_  = \new_[66149]_  & \new_[66146]_ ;
  assign \new_[66151]_  = \new_[66150]_  & \new_[66143]_ ;
  assign \new_[66155]_  = ~A298 & ~A269;
  assign \new_[66156]_  = ~A268 & \new_[66155]_ ;
  assign \new_[66159]_  = ~A300 & A299;
  assign \new_[66162]_  = ~A302 & ~A301;
  assign \new_[66163]_  = \new_[66162]_  & \new_[66159]_ ;
  assign \new_[66164]_  = \new_[66163]_  & \new_[66156]_ ;
  assign \new_[66168]_  = ~A167 & A168;
  assign \new_[66169]_  = A169 & \new_[66168]_ ;
  assign \new_[66172]_  = ~A201 & A166;
  assign \new_[66175]_  = A267 & A203;
  assign \new_[66176]_  = \new_[66175]_  & \new_[66172]_ ;
  assign \new_[66177]_  = \new_[66176]_  & \new_[66169]_ ;
  assign \new_[66181]_  = A298 & ~A269;
  assign \new_[66182]_  = ~A268 & \new_[66181]_ ;
  assign \new_[66185]_  = ~A300 & ~A299;
  assign \new_[66188]_  = ~A302 & ~A301;
  assign \new_[66189]_  = \new_[66188]_  & \new_[66185]_ ;
  assign \new_[66190]_  = \new_[66189]_  & \new_[66182]_ ;
  assign \new_[66194]_  = ~A167 & A168;
  assign \new_[66195]_  = A169 & \new_[66194]_ ;
  assign \new_[66198]_  = ~A201 & A166;
  assign \new_[66201]_  = A267 & A203;
  assign \new_[66202]_  = \new_[66201]_  & \new_[66198]_ ;
  assign \new_[66203]_  = \new_[66202]_  & \new_[66195]_ ;
  assign \new_[66207]_  = ~A298 & ~A269;
  assign \new_[66208]_  = ~A268 & \new_[66207]_ ;
  assign \new_[66211]_  = ~A300 & A299;
  assign \new_[66214]_  = ~A302 & ~A301;
  assign \new_[66215]_  = \new_[66214]_  & \new_[66211]_ ;
  assign \new_[66216]_  = \new_[66215]_  & \new_[66208]_ ;
  assign \new_[66220]_  = ~A167 & A168;
  assign \new_[66221]_  = A169 & \new_[66220]_ ;
  assign \new_[66224]_  = A199 & A166;
  assign \new_[66227]_  = A267 & A200;
  assign \new_[66228]_  = \new_[66227]_  & \new_[66224]_ ;
  assign \new_[66229]_  = \new_[66228]_  & \new_[66221]_ ;
  assign \new_[66233]_  = A298 & ~A269;
  assign \new_[66234]_  = ~A268 & \new_[66233]_ ;
  assign \new_[66237]_  = ~A300 & ~A299;
  assign \new_[66240]_  = ~A302 & ~A301;
  assign \new_[66241]_  = \new_[66240]_  & \new_[66237]_ ;
  assign \new_[66242]_  = \new_[66241]_  & \new_[66234]_ ;
  assign \new_[66246]_  = ~A167 & A168;
  assign \new_[66247]_  = A169 & \new_[66246]_ ;
  assign \new_[66250]_  = A199 & A166;
  assign \new_[66253]_  = A267 & A200;
  assign \new_[66254]_  = \new_[66253]_  & \new_[66250]_ ;
  assign \new_[66255]_  = \new_[66254]_  & \new_[66247]_ ;
  assign \new_[66259]_  = ~A298 & ~A269;
  assign \new_[66260]_  = ~A268 & \new_[66259]_ ;
  assign \new_[66263]_  = ~A300 & A299;
  assign \new_[66266]_  = ~A302 & ~A301;
  assign \new_[66267]_  = \new_[66266]_  & \new_[66263]_ ;
  assign \new_[66268]_  = \new_[66267]_  & \new_[66260]_ ;
  assign \new_[66272]_  = ~A167 & A168;
  assign \new_[66273]_  = A169 & \new_[66272]_ ;
  assign \new_[66276]_  = ~A199 & A166;
  assign \new_[66279]_  = A201 & A200;
  assign \new_[66280]_  = \new_[66279]_  & \new_[66276]_ ;
  assign \new_[66281]_  = \new_[66280]_  & \new_[66273]_ ;
  assign \new_[66285]_  = A266 & ~A265;
  assign \new_[66286]_  = A202 & \new_[66285]_ ;
  assign \new_[66289]_  = A268 & A267;
  assign \new_[66292]_  = A301 & ~A300;
  assign \new_[66293]_  = \new_[66292]_  & \new_[66289]_ ;
  assign \new_[66294]_  = \new_[66293]_  & \new_[66286]_ ;
  assign \new_[66298]_  = ~A167 & A168;
  assign \new_[66299]_  = A169 & \new_[66298]_ ;
  assign \new_[66302]_  = ~A199 & A166;
  assign \new_[66305]_  = A201 & A200;
  assign \new_[66306]_  = \new_[66305]_  & \new_[66302]_ ;
  assign \new_[66307]_  = \new_[66306]_  & \new_[66299]_ ;
  assign \new_[66311]_  = A266 & ~A265;
  assign \new_[66312]_  = A202 & \new_[66311]_ ;
  assign \new_[66315]_  = A268 & A267;
  assign \new_[66318]_  = A302 & ~A300;
  assign \new_[66319]_  = \new_[66318]_  & \new_[66315]_ ;
  assign \new_[66320]_  = \new_[66319]_  & \new_[66312]_ ;
  assign \new_[66324]_  = ~A167 & A168;
  assign \new_[66325]_  = A169 & \new_[66324]_ ;
  assign \new_[66328]_  = ~A199 & A166;
  assign \new_[66331]_  = A201 & A200;
  assign \new_[66332]_  = \new_[66331]_  & \new_[66328]_ ;
  assign \new_[66333]_  = \new_[66332]_  & \new_[66325]_ ;
  assign \new_[66337]_  = A266 & ~A265;
  assign \new_[66338]_  = A202 & \new_[66337]_ ;
  assign \new_[66341]_  = A268 & A267;
  assign \new_[66344]_  = A299 & A298;
  assign \new_[66345]_  = \new_[66344]_  & \new_[66341]_ ;
  assign \new_[66346]_  = \new_[66345]_  & \new_[66338]_ ;
  assign \new_[66350]_  = ~A167 & A168;
  assign \new_[66351]_  = A169 & \new_[66350]_ ;
  assign \new_[66354]_  = ~A199 & A166;
  assign \new_[66357]_  = A201 & A200;
  assign \new_[66358]_  = \new_[66357]_  & \new_[66354]_ ;
  assign \new_[66359]_  = \new_[66358]_  & \new_[66351]_ ;
  assign \new_[66363]_  = A266 & ~A265;
  assign \new_[66364]_  = A202 & \new_[66363]_ ;
  assign \new_[66367]_  = A268 & A267;
  assign \new_[66370]_  = ~A299 & ~A298;
  assign \new_[66371]_  = \new_[66370]_  & \new_[66367]_ ;
  assign \new_[66372]_  = \new_[66371]_  & \new_[66364]_ ;
  assign \new_[66376]_  = ~A167 & A168;
  assign \new_[66377]_  = A169 & \new_[66376]_ ;
  assign \new_[66380]_  = ~A199 & A166;
  assign \new_[66383]_  = A201 & A200;
  assign \new_[66384]_  = \new_[66383]_  & \new_[66380]_ ;
  assign \new_[66385]_  = \new_[66384]_  & \new_[66377]_ ;
  assign \new_[66389]_  = A266 & ~A265;
  assign \new_[66390]_  = A202 & \new_[66389]_ ;
  assign \new_[66393]_  = A269 & A267;
  assign \new_[66396]_  = A301 & ~A300;
  assign \new_[66397]_  = \new_[66396]_  & \new_[66393]_ ;
  assign \new_[66398]_  = \new_[66397]_  & \new_[66390]_ ;
  assign \new_[66402]_  = ~A167 & A168;
  assign \new_[66403]_  = A169 & \new_[66402]_ ;
  assign \new_[66406]_  = ~A199 & A166;
  assign \new_[66409]_  = A201 & A200;
  assign \new_[66410]_  = \new_[66409]_  & \new_[66406]_ ;
  assign \new_[66411]_  = \new_[66410]_  & \new_[66403]_ ;
  assign \new_[66415]_  = A266 & ~A265;
  assign \new_[66416]_  = A202 & \new_[66415]_ ;
  assign \new_[66419]_  = A269 & A267;
  assign \new_[66422]_  = A302 & ~A300;
  assign \new_[66423]_  = \new_[66422]_  & \new_[66419]_ ;
  assign \new_[66424]_  = \new_[66423]_  & \new_[66416]_ ;
  assign \new_[66428]_  = ~A167 & A168;
  assign \new_[66429]_  = A169 & \new_[66428]_ ;
  assign \new_[66432]_  = ~A199 & A166;
  assign \new_[66435]_  = A201 & A200;
  assign \new_[66436]_  = \new_[66435]_  & \new_[66432]_ ;
  assign \new_[66437]_  = \new_[66436]_  & \new_[66429]_ ;
  assign \new_[66441]_  = A266 & ~A265;
  assign \new_[66442]_  = A202 & \new_[66441]_ ;
  assign \new_[66445]_  = A269 & A267;
  assign \new_[66448]_  = A299 & A298;
  assign \new_[66449]_  = \new_[66448]_  & \new_[66445]_ ;
  assign \new_[66450]_  = \new_[66449]_  & \new_[66442]_ ;
  assign \new_[66454]_  = ~A167 & A168;
  assign \new_[66455]_  = A169 & \new_[66454]_ ;
  assign \new_[66458]_  = ~A199 & A166;
  assign \new_[66461]_  = A201 & A200;
  assign \new_[66462]_  = \new_[66461]_  & \new_[66458]_ ;
  assign \new_[66463]_  = \new_[66462]_  & \new_[66455]_ ;
  assign \new_[66467]_  = A266 & ~A265;
  assign \new_[66468]_  = A202 & \new_[66467]_ ;
  assign \new_[66471]_  = A269 & A267;
  assign \new_[66474]_  = ~A299 & ~A298;
  assign \new_[66475]_  = \new_[66474]_  & \new_[66471]_ ;
  assign \new_[66476]_  = \new_[66475]_  & \new_[66468]_ ;
  assign \new_[66480]_  = ~A167 & A168;
  assign \new_[66481]_  = A169 & \new_[66480]_ ;
  assign \new_[66484]_  = ~A199 & A166;
  assign \new_[66487]_  = A201 & A200;
  assign \new_[66488]_  = \new_[66487]_  & \new_[66484]_ ;
  assign \new_[66489]_  = \new_[66488]_  & \new_[66481]_ ;
  assign \new_[66493]_  = ~A266 & A265;
  assign \new_[66494]_  = A202 & \new_[66493]_ ;
  assign \new_[66497]_  = A268 & A267;
  assign \new_[66500]_  = A301 & ~A300;
  assign \new_[66501]_  = \new_[66500]_  & \new_[66497]_ ;
  assign \new_[66502]_  = \new_[66501]_  & \new_[66494]_ ;
  assign \new_[66506]_  = ~A167 & A168;
  assign \new_[66507]_  = A169 & \new_[66506]_ ;
  assign \new_[66510]_  = ~A199 & A166;
  assign \new_[66513]_  = A201 & A200;
  assign \new_[66514]_  = \new_[66513]_  & \new_[66510]_ ;
  assign \new_[66515]_  = \new_[66514]_  & \new_[66507]_ ;
  assign \new_[66519]_  = ~A266 & A265;
  assign \new_[66520]_  = A202 & \new_[66519]_ ;
  assign \new_[66523]_  = A268 & A267;
  assign \new_[66526]_  = A302 & ~A300;
  assign \new_[66527]_  = \new_[66526]_  & \new_[66523]_ ;
  assign \new_[66528]_  = \new_[66527]_  & \new_[66520]_ ;
  assign \new_[66532]_  = ~A167 & A168;
  assign \new_[66533]_  = A169 & \new_[66532]_ ;
  assign \new_[66536]_  = ~A199 & A166;
  assign \new_[66539]_  = A201 & A200;
  assign \new_[66540]_  = \new_[66539]_  & \new_[66536]_ ;
  assign \new_[66541]_  = \new_[66540]_  & \new_[66533]_ ;
  assign \new_[66545]_  = ~A266 & A265;
  assign \new_[66546]_  = A202 & \new_[66545]_ ;
  assign \new_[66549]_  = A268 & A267;
  assign \new_[66552]_  = A299 & A298;
  assign \new_[66553]_  = \new_[66552]_  & \new_[66549]_ ;
  assign \new_[66554]_  = \new_[66553]_  & \new_[66546]_ ;
  assign \new_[66558]_  = ~A167 & A168;
  assign \new_[66559]_  = A169 & \new_[66558]_ ;
  assign \new_[66562]_  = ~A199 & A166;
  assign \new_[66565]_  = A201 & A200;
  assign \new_[66566]_  = \new_[66565]_  & \new_[66562]_ ;
  assign \new_[66567]_  = \new_[66566]_  & \new_[66559]_ ;
  assign \new_[66571]_  = ~A266 & A265;
  assign \new_[66572]_  = A202 & \new_[66571]_ ;
  assign \new_[66575]_  = A268 & A267;
  assign \new_[66578]_  = ~A299 & ~A298;
  assign \new_[66579]_  = \new_[66578]_  & \new_[66575]_ ;
  assign \new_[66580]_  = \new_[66579]_  & \new_[66572]_ ;
  assign \new_[66584]_  = ~A167 & A168;
  assign \new_[66585]_  = A169 & \new_[66584]_ ;
  assign \new_[66588]_  = ~A199 & A166;
  assign \new_[66591]_  = A201 & A200;
  assign \new_[66592]_  = \new_[66591]_  & \new_[66588]_ ;
  assign \new_[66593]_  = \new_[66592]_  & \new_[66585]_ ;
  assign \new_[66597]_  = ~A266 & A265;
  assign \new_[66598]_  = A202 & \new_[66597]_ ;
  assign \new_[66601]_  = A269 & A267;
  assign \new_[66604]_  = A301 & ~A300;
  assign \new_[66605]_  = \new_[66604]_  & \new_[66601]_ ;
  assign \new_[66606]_  = \new_[66605]_  & \new_[66598]_ ;
  assign \new_[66610]_  = ~A167 & A168;
  assign \new_[66611]_  = A169 & \new_[66610]_ ;
  assign \new_[66614]_  = ~A199 & A166;
  assign \new_[66617]_  = A201 & A200;
  assign \new_[66618]_  = \new_[66617]_  & \new_[66614]_ ;
  assign \new_[66619]_  = \new_[66618]_  & \new_[66611]_ ;
  assign \new_[66623]_  = ~A266 & A265;
  assign \new_[66624]_  = A202 & \new_[66623]_ ;
  assign \new_[66627]_  = A269 & A267;
  assign \new_[66630]_  = A302 & ~A300;
  assign \new_[66631]_  = \new_[66630]_  & \new_[66627]_ ;
  assign \new_[66632]_  = \new_[66631]_  & \new_[66624]_ ;
  assign \new_[66636]_  = ~A167 & A168;
  assign \new_[66637]_  = A169 & \new_[66636]_ ;
  assign \new_[66640]_  = ~A199 & A166;
  assign \new_[66643]_  = A201 & A200;
  assign \new_[66644]_  = \new_[66643]_  & \new_[66640]_ ;
  assign \new_[66645]_  = \new_[66644]_  & \new_[66637]_ ;
  assign \new_[66649]_  = ~A266 & A265;
  assign \new_[66650]_  = A202 & \new_[66649]_ ;
  assign \new_[66653]_  = A269 & A267;
  assign \new_[66656]_  = A299 & A298;
  assign \new_[66657]_  = \new_[66656]_  & \new_[66653]_ ;
  assign \new_[66658]_  = \new_[66657]_  & \new_[66650]_ ;
  assign \new_[66662]_  = ~A167 & A168;
  assign \new_[66663]_  = A169 & \new_[66662]_ ;
  assign \new_[66666]_  = ~A199 & A166;
  assign \new_[66669]_  = A201 & A200;
  assign \new_[66670]_  = \new_[66669]_  & \new_[66666]_ ;
  assign \new_[66671]_  = \new_[66670]_  & \new_[66663]_ ;
  assign \new_[66675]_  = ~A266 & A265;
  assign \new_[66676]_  = A202 & \new_[66675]_ ;
  assign \new_[66679]_  = A269 & A267;
  assign \new_[66682]_  = ~A299 & ~A298;
  assign \new_[66683]_  = \new_[66682]_  & \new_[66679]_ ;
  assign \new_[66684]_  = \new_[66683]_  & \new_[66676]_ ;
  assign \new_[66688]_  = ~A167 & A168;
  assign \new_[66689]_  = A169 & \new_[66688]_ ;
  assign \new_[66692]_  = ~A199 & A166;
  assign \new_[66695]_  = A201 & A200;
  assign \new_[66696]_  = \new_[66695]_  & \new_[66692]_ ;
  assign \new_[66697]_  = \new_[66696]_  & \new_[66689]_ ;
  assign \new_[66701]_  = A266 & ~A265;
  assign \new_[66702]_  = A203 & \new_[66701]_ ;
  assign \new_[66705]_  = A268 & A267;
  assign \new_[66708]_  = A301 & ~A300;
  assign \new_[66709]_  = \new_[66708]_  & \new_[66705]_ ;
  assign \new_[66710]_  = \new_[66709]_  & \new_[66702]_ ;
  assign \new_[66714]_  = ~A167 & A168;
  assign \new_[66715]_  = A169 & \new_[66714]_ ;
  assign \new_[66718]_  = ~A199 & A166;
  assign \new_[66721]_  = A201 & A200;
  assign \new_[66722]_  = \new_[66721]_  & \new_[66718]_ ;
  assign \new_[66723]_  = \new_[66722]_  & \new_[66715]_ ;
  assign \new_[66727]_  = A266 & ~A265;
  assign \new_[66728]_  = A203 & \new_[66727]_ ;
  assign \new_[66731]_  = A268 & A267;
  assign \new_[66734]_  = A302 & ~A300;
  assign \new_[66735]_  = \new_[66734]_  & \new_[66731]_ ;
  assign \new_[66736]_  = \new_[66735]_  & \new_[66728]_ ;
  assign \new_[66740]_  = ~A167 & A168;
  assign \new_[66741]_  = A169 & \new_[66740]_ ;
  assign \new_[66744]_  = ~A199 & A166;
  assign \new_[66747]_  = A201 & A200;
  assign \new_[66748]_  = \new_[66747]_  & \new_[66744]_ ;
  assign \new_[66749]_  = \new_[66748]_  & \new_[66741]_ ;
  assign \new_[66753]_  = A266 & ~A265;
  assign \new_[66754]_  = A203 & \new_[66753]_ ;
  assign \new_[66757]_  = A268 & A267;
  assign \new_[66760]_  = A299 & A298;
  assign \new_[66761]_  = \new_[66760]_  & \new_[66757]_ ;
  assign \new_[66762]_  = \new_[66761]_  & \new_[66754]_ ;
  assign \new_[66766]_  = ~A167 & A168;
  assign \new_[66767]_  = A169 & \new_[66766]_ ;
  assign \new_[66770]_  = ~A199 & A166;
  assign \new_[66773]_  = A201 & A200;
  assign \new_[66774]_  = \new_[66773]_  & \new_[66770]_ ;
  assign \new_[66775]_  = \new_[66774]_  & \new_[66767]_ ;
  assign \new_[66779]_  = A266 & ~A265;
  assign \new_[66780]_  = A203 & \new_[66779]_ ;
  assign \new_[66783]_  = A268 & A267;
  assign \new_[66786]_  = ~A299 & ~A298;
  assign \new_[66787]_  = \new_[66786]_  & \new_[66783]_ ;
  assign \new_[66788]_  = \new_[66787]_  & \new_[66780]_ ;
  assign \new_[66792]_  = ~A167 & A168;
  assign \new_[66793]_  = A169 & \new_[66792]_ ;
  assign \new_[66796]_  = ~A199 & A166;
  assign \new_[66799]_  = A201 & A200;
  assign \new_[66800]_  = \new_[66799]_  & \new_[66796]_ ;
  assign \new_[66801]_  = \new_[66800]_  & \new_[66793]_ ;
  assign \new_[66805]_  = A266 & ~A265;
  assign \new_[66806]_  = A203 & \new_[66805]_ ;
  assign \new_[66809]_  = A269 & A267;
  assign \new_[66812]_  = A301 & ~A300;
  assign \new_[66813]_  = \new_[66812]_  & \new_[66809]_ ;
  assign \new_[66814]_  = \new_[66813]_  & \new_[66806]_ ;
  assign \new_[66818]_  = ~A167 & A168;
  assign \new_[66819]_  = A169 & \new_[66818]_ ;
  assign \new_[66822]_  = ~A199 & A166;
  assign \new_[66825]_  = A201 & A200;
  assign \new_[66826]_  = \new_[66825]_  & \new_[66822]_ ;
  assign \new_[66827]_  = \new_[66826]_  & \new_[66819]_ ;
  assign \new_[66831]_  = A266 & ~A265;
  assign \new_[66832]_  = A203 & \new_[66831]_ ;
  assign \new_[66835]_  = A269 & A267;
  assign \new_[66838]_  = A302 & ~A300;
  assign \new_[66839]_  = \new_[66838]_  & \new_[66835]_ ;
  assign \new_[66840]_  = \new_[66839]_  & \new_[66832]_ ;
  assign \new_[66844]_  = ~A167 & A168;
  assign \new_[66845]_  = A169 & \new_[66844]_ ;
  assign \new_[66848]_  = ~A199 & A166;
  assign \new_[66851]_  = A201 & A200;
  assign \new_[66852]_  = \new_[66851]_  & \new_[66848]_ ;
  assign \new_[66853]_  = \new_[66852]_  & \new_[66845]_ ;
  assign \new_[66857]_  = A266 & ~A265;
  assign \new_[66858]_  = A203 & \new_[66857]_ ;
  assign \new_[66861]_  = A269 & A267;
  assign \new_[66864]_  = A299 & A298;
  assign \new_[66865]_  = \new_[66864]_  & \new_[66861]_ ;
  assign \new_[66866]_  = \new_[66865]_  & \new_[66858]_ ;
  assign \new_[66870]_  = ~A167 & A168;
  assign \new_[66871]_  = A169 & \new_[66870]_ ;
  assign \new_[66874]_  = ~A199 & A166;
  assign \new_[66877]_  = A201 & A200;
  assign \new_[66878]_  = \new_[66877]_  & \new_[66874]_ ;
  assign \new_[66879]_  = \new_[66878]_  & \new_[66871]_ ;
  assign \new_[66883]_  = A266 & ~A265;
  assign \new_[66884]_  = A203 & \new_[66883]_ ;
  assign \new_[66887]_  = A269 & A267;
  assign \new_[66890]_  = ~A299 & ~A298;
  assign \new_[66891]_  = \new_[66890]_  & \new_[66887]_ ;
  assign \new_[66892]_  = \new_[66891]_  & \new_[66884]_ ;
  assign \new_[66896]_  = ~A167 & A168;
  assign \new_[66897]_  = A169 & \new_[66896]_ ;
  assign \new_[66900]_  = ~A199 & A166;
  assign \new_[66903]_  = A201 & A200;
  assign \new_[66904]_  = \new_[66903]_  & \new_[66900]_ ;
  assign \new_[66905]_  = \new_[66904]_  & \new_[66897]_ ;
  assign \new_[66909]_  = ~A266 & A265;
  assign \new_[66910]_  = A203 & \new_[66909]_ ;
  assign \new_[66913]_  = A268 & A267;
  assign \new_[66916]_  = A301 & ~A300;
  assign \new_[66917]_  = \new_[66916]_  & \new_[66913]_ ;
  assign \new_[66918]_  = \new_[66917]_  & \new_[66910]_ ;
  assign \new_[66922]_  = ~A167 & A168;
  assign \new_[66923]_  = A169 & \new_[66922]_ ;
  assign \new_[66926]_  = ~A199 & A166;
  assign \new_[66929]_  = A201 & A200;
  assign \new_[66930]_  = \new_[66929]_  & \new_[66926]_ ;
  assign \new_[66931]_  = \new_[66930]_  & \new_[66923]_ ;
  assign \new_[66935]_  = ~A266 & A265;
  assign \new_[66936]_  = A203 & \new_[66935]_ ;
  assign \new_[66939]_  = A268 & A267;
  assign \new_[66942]_  = A302 & ~A300;
  assign \new_[66943]_  = \new_[66942]_  & \new_[66939]_ ;
  assign \new_[66944]_  = \new_[66943]_  & \new_[66936]_ ;
  assign \new_[66948]_  = ~A167 & A168;
  assign \new_[66949]_  = A169 & \new_[66948]_ ;
  assign \new_[66952]_  = ~A199 & A166;
  assign \new_[66955]_  = A201 & A200;
  assign \new_[66956]_  = \new_[66955]_  & \new_[66952]_ ;
  assign \new_[66957]_  = \new_[66956]_  & \new_[66949]_ ;
  assign \new_[66961]_  = ~A266 & A265;
  assign \new_[66962]_  = A203 & \new_[66961]_ ;
  assign \new_[66965]_  = A268 & A267;
  assign \new_[66968]_  = A299 & A298;
  assign \new_[66969]_  = \new_[66968]_  & \new_[66965]_ ;
  assign \new_[66970]_  = \new_[66969]_  & \new_[66962]_ ;
  assign \new_[66974]_  = ~A167 & A168;
  assign \new_[66975]_  = A169 & \new_[66974]_ ;
  assign \new_[66978]_  = ~A199 & A166;
  assign \new_[66981]_  = A201 & A200;
  assign \new_[66982]_  = \new_[66981]_  & \new_[66978]_ ;
  assign \new_[66983]_  = \new_[66982]_  & \new_[66975]_ ;
  assign \new_[66987]_  = ~A266 & A265;
  assign \new_[66988]_  = A203 & \new_[66987]_ ;
  assign \new_[66991]_  = A268 & A267;
  assign \new_[66994]_  = ~A299 & ~A298;
  assign \new_[66995]_  = \new_[66994]_  & \new_[66991]_ ;
  assign \new_[66996]_  = \new_[66995]_  & \new_[66988]_ ;
  assign \new_[67000]_  = ~A167 & A168;
  assign \new_[67001]_  = A169 & \new_[67000]_ ;
  assign \new_[67004]_  = ~A199 & A166;
  assign \new_[67007]_  = A201 & A200;
  assign \new_[67008]_  = \new_[67007]_  & \new_[67004]_ ;
  assign \new_[67009]_  = \new_[67008]_  & \new_[67001]_ ;
  assign \new_[67013]_  = ~A266 & A265;
  assign \new_[67014]_  = A203 & \new_[67013]_ ;
  assign \new_[67017]_  = A269 & A267;
  assign \new_[67020]_  = A301 & ~A300;
  assign \new_[67021]_  = \new_[67020]_  & \new_[67017]_ ;
  assign \new_[67022]_  = \new_[67021]_  & \new_[67014]_ ;
  assign \new_[67026]_  = ~A167 & A168;
  assign \new_[67027]_  = A169 & \new_[67026]_ ;
  assign \new_[67030]_  = ~A199 & A166;
  assign \new_[67033]_  = A201 & A200;
  assign \new_[67034]_  = \new_[67033]_  & \new_[67030]_ ;
  assign \new_[67035]_  = \new_[67034]_  & \new_[67027]_ ;
  assign \new_[67039]_  = ~A266 & A265;
  assign \new_[67040]_  = A203 & \new_[67039]_ ;
  assign \new_[67043]_  = A269 & A267;
  assign \new_[67046]_  = A302 & ~A300;
  assign \new_[67047]_  = \new_[67046]_  & \new_[67043]_ ;
  assign \new_[67048]_  = \new_[67047]_  & \new_[67040]_ ;
  assign \new_[67052]_  = ~A167 & A168;
  assign \new_[67053]_  = A169 & \new_[67052]_ ;
  assign \new_[67056]_  = ~A199 & A166;
  assign \new_[67059]_  = A201 & A200;
  assign \new_[67060]_  = \new_[67059]_  & \new_[67056]_ ;
  assign \new_[67061]_  = \new_[67060]_  & \new_[67053]_ ;
  assign \new_[67065]_  = ~A266 & A265;
  assign \new_[67066]_  = A203 & \new_[67065]_ ;
  assign \new_[67069]_  = A269 & A267;
  assign \new_[67072]_  = A299 & A298;
  assign \new_[67073]_  = \new_[67072]_  & \new_[67069]_ ;
  assign \new_[67074]_  = \new_[67073]_  & \new_[67066]_ ;
  assign \new_[67078]_  = ~A167 & A168;
  assign \new_[67079]_  = A169 & \new_[67078]_ ;
  assign \new_[67082]_  = ~A199 & A166;
  assign \new_[67085]_  = A201 & A200;
  assign \new_[67086]_  = \new_[67085]_  & \new_[67082]_ ;
  assign \new_[67087]_  = \new_[67086]_  & \new_[67079]_ ;
  assign \new_[67091]_  = ~A266 & A265;
  assign \new_[67092]_  = A203 & \new_[67091]_ ;
  assign \new_[67095]_  = A269 & A267;
  assign \new_[67098]_  = ~A299 & ~A298;
  assign \new_[67099]_  = \new_[67098]_  & \new_[67095]_ ;
  assign \new_[67100]_  = \new_[67099]_  & \new_[67092]_ ;
  assign \new_[67104]_  = ~A167 & A168;
  assign \new_[67105]_  = A169 & \new_[67104]_ ;
  assign \new_[67108]_  = A199 & A166;
  assign \new_[67111]_  = A201 & ~A200;
  assign \new_[67112]_  = \new_[67111]_  & \new_[67108]_ ;
  assign \new_[67113]_  = \new_[67112]_  & \new_[67105]_ ;
  assign \new_[67117]_  = A266 & ~A265;
  assign \new_[67118]_  = A202 & \new_[67117]_ ;
  assign \new_[67121]_  = A268 & A267;
  assign \new_[67124]_  = A301 & ~A300;
  assign \new_[67125]_  = \new_[67124]_  & \new_[67121]_ ;
  assign \new_[67126]_  = \new_[67125]_  & \new_[67118]_ ;
  assign \new_[67130]_  = ~A167 & A168;
  assign \new_[67131]_  = A169 & \new_[67130]_ ;
  assign \new_[67134]_  = A199 & A166;
  assign \new_[67137]_  = A201 & ~A200;
  assign \new_[67138]_  = \new_[67137]_  & \new_[67134]_ ;
  assign \new_[67139]_  = \new_[67138]_  & \new_[67131]_ ;
  assign \new_[67143]_  = A266 & ~A265;
  assign \new_[67144]_  = A202 & \new_[67143]_ ;
  assign \new_[67147]_  = A268 & A267;
  assign \new_[67150]_  = A302 & ~A300;
  assign \new_[67151]_  = \new_[67150]_  & \new_[67147]_ ;
  assign \new_[67152]_  = \new_[67151]_  & \new_[67144]_ ;
  assign \new_[67156]_  = ~A167 & A168;
  assign \new_[67157]_  = A169 & \new_[67156]_ ;
  assign \new_[67160]_  = A199 & A166;
  assign \new_[67163]_  = A201 & ~A200;
  assign \new_[67164]_  = \new_[67163]_  & \new_[67160]_ ;
  assign \new_[67165]_  = \new_[67164]_  & \new_[67157]_ ;
  assign \new_[67169]_  = A266 & ~A265;
  assign \new_[67170]_  = A202 & \new_[67169]_ ;
  assign \new_[67173]_  = A268 & A267;
  assign \new_[67176]_  = A299 & A298;
  assign \new_[67177]_  = \new_[67176]_  & \new_[67173]_ ;
  assign \new_[67178]_  = \new_[67177]_  & \new_[67170]_ ;
  assign \new_[67182]_  = ~A167 & A168;
  assign \new_[67183]_  = A169 & \new_[67182]_ ;
  assign \new_[67186]_  = A199 & A166;
  assign \new_[67189]_  = A201 & ~A200;
  assign \new_[67190]_  = \new_[67189]_  & \new_[67186]_ ;
  assign \new_[67191]_  = \new_[67190]_  & \new_[67183]_ ;
  assign \new_[67195]_  = A266 & ~A265;
  assign \new_[67196]_  = A202 & \new_[67195]_ ;
  assign \new_[67199]_  = A268 & A267;
  assign \new_[67202]_  = ~A299 & ~A298;
  assign \new_[67203]_  = \new_[67202]_  & \new_[67199]_ ;
  assign \new_[67204]_  = \new_[67203]_  & \new_[67196]_ ;
  assign \new_[67208]_  = ~A167 & A168;
  assign \new_[67209]_  = A169 & \new_[67208]_ ;
  assign \new_[67212]_  = A199 & A166;
  assign \new_[67215]_  = A201 & ~A200;
  assign \new_[67216]_  = \new_[67215]_  & \new_[67212]_ ;
  assign \new_[67217]_  = \new_[67216]_  & \new_[67209]_ ;
  assign \new_[67221]_  = A266 & ~A265;
  assign \new_[67222]_  = A202 & \new_[67221]_ ;
  assign \new_[67225]_  = A269 & A267;
  assign \new_[67228]_  = A301 & ~A300;
  assign \new_[67229]_  = \new_[67228]_  & \new_[67225]_ ;
  assign \new_[67230]_  = \new_[67229]_  & \new_[67222]_ ;
  assign \new_[67234]_  = ~A167 & A168;
  assign \new_[67235]_  = A169 & \new_[67234]_ ;
  assign \new_[67238]_  = A199 & A166;
  assign \new_[67241]_  = A201 & ~A200;
  assign \new_[67242]_  = \new_[67241]_  & \new_[67238]_ ;
  assign \new_[67243]_  = \new_[67242]_  & \new_[67235]_ ;
  assign \new_[67247]_  = A266 & ~A265;
  assign \new_[67248]_  = A202 & \new_[67247]_ ;
  assign \new_[67251]_  = A269 & A267;
  assign \new_[67254]_  = A302 & ~A300;
  assign \new_[67255]_  = \new_[67254]_  & \new_[67251]_ ;
  assign \new_[67256]_  = \new_[67255]_  & \new_[67248]_ ;
  assign \new_[67260]_  = ~A167 & A168;
  assign \new_[67261]_  = A169 & \new_[67260]_ ;
  assign \new_[67264]_  = A199 & A166;
  assign \new_[67267]_  = A201 & ~A200;
  assign \new_[67268]_  = \new_[67267]_  & \new_[67264]_ ;
  assign \new_[67269]_  = \new_[67268]_  & \new_[67261]_ ;
  assign \new_[67273]_  = A266 & ~A265;
  assign \new_[67274]_  = A202 & \new_[67273]_ ;
  assign \new_[67277]_  = A269 & A267;
  assign \new_[67280]_  = A299 & A298;
  assign \new_[67281]_  = \new_[67280]_  & \new_[67277]_ ;
  assign \new_[67282]_  = \new_[67281]_  & \new_[67274]_ ;
  assign \new_[67286]_  = ~A167 & A168;
  assign \new_[67287]_  = A169 & \new_[67286]_ ;
  assign \new_[67290]_  = A199 & A166;
  assign \new_[67293]_  = A201 & ~A200;
  assign \new_[67294]_  = \new_[67293]_  & \new_[67290]_ ;
  assign \new_[67295]_  = \new_[67294]_  & \new_[67287]_ ;
  assign \new_[67299]_  = A266 & ~A265;
  assign \new_[67300]_  = A202 & \new_[67299]_ ;
  assign \new_[67303]_  = A269 & A267;
  assign \new_[67306]_  = ~A299 & ~A298;
  assign \new_[67307]_  = \new_[67306]_  & \new_[67303]_ ;
  assign \new_[67308]_  = \new_[67307]_  & \new_[67300]_ ;
  assign \new_[67312]_  = ~A167 & A168;
  assign \new_[67313]_  = A169 & \new_[67312]_ ;
  assign \new_[67316]_  = A199 & A166;
  assign \new_[67319]_  = A201 & ~A200;
  assign \new_[67320]_  = \new_[67319]_  & \new_[67316]_ ;
  assign \new_[67321]_  = \new_[67320]_  & \new_[67313]_ ;
  assign \new_[67325]_  = ~A266 & A265;
  assign \new_[67326]_  = A202 & \new_[67325]_ ;
  assign \new_[67329]_  = A268 & A267;
  assign \new_[67332]_  = A301 & ~A300;
  assign \new_[67333]_  = \new_[67332]_  & \new_[67329]_ ;
  assign \new_[67334]_  = \new_[67333]_  & \new_[67326]_ ;
  assign \new_[67338]_  = ~A167 & A168;
  assign \new_[67339]_  = A169 & \new_[67338]_ ;
  assign \new_[67342]_  = A199 & A166;
  assign \new_[67345]_  = A201 & ~A200;
  assign \new_[67346]_  = \new_[67345]_  & \new_[67342]_ ;
  assign \new_[67347]_  = \new_[67346]_  & \new_[67339]_ ;
  assign \new_[67351]_  = ~A266 & A265;
  assign \new_[67352]_  = A202 & \new_[67351]_ ;
  assign \new_[67355]_  = A268 & A267;
  assign \new_[67358]_  = A302 & ~A300;
  assign \new_[67359]_  = \new_[67358]_  & \new_[67355]_ ;
  assign \new_[67360]_  = \new_[67359]_  & \new_[67352]_ ;
  assign \new_[67364]_  = ~A167 & A168;
  assign \new_[67365]_  = A169 & \new_[67364]_ ;
  assign \new_[67368]_  = A199 & A166;
  assign \new_[67371]_  = A201 & ~A200;
  assign \new_[67372]_  = \new_[67371]_  & \new_[67368]_ ;
  assign \new_[67373]_  = \new_[67372]_  & \new_[67365]_ ;
  assign \new_[67377]_  = ~A266 & A265;
  assign \new_[67378]_  = A202 & \new_[67377]_ ;
  assign \new_[67381]_  = A268 & A267;
  assign \new_[67384]_  = A299 & A298;
  assign \new_[67385]_  = \new_[67384]_  & \new_[67381]_ ;
  assign \new_[67386]_  = \new_[67385]_  & \new_[67378]_ ;
  assign \new_[67390]_  = ~A167 & A168;
  assign \new_[67391]_  = A169 & \new_[67390]_ ;
  assign \new_[67394]_  = A199 & A166;
  assign \new_[67397]_  = A201 & ~A200;
  assign \new_[67398]_  = \new_[67397]_  & \new_[67394]_ ;
  assign \new_[67399]_  = \new_[67398]_  & \new_[67391]_ ;
  assign \new_[67403]_  = ~A266 & A265;
  assign \new_[67404]_  = A202 & \new_[67403]_ ;
  assign \new_[67407]_  = A268 & A267;
  assign \new_[67410]_  = ~A299 & ~A298;
  assign \new_[67411]_  = \new_[67410]_  & \new_[67407]_ ;
  assign \new_[67412]_  = \new_[67411]_  & \new_[67404]_ ;
  assign \new_[67416]_  = ~A167 & A168;
  assign \new_[67417]_  = A169 & \new_[67416]_ ;
  assign \new_[67420]_  = A199 & A166;
  assign \new_[67423]_  = A201 & ~A200;
  assign \new_[67424]_  = \new_[67423]_  & \new_[67420]_ ;
  assign \new_[67425]_  = \new_[67424]_  & \new_[67417]_ ;
  assign \new_[67429]_  = ~A266 & A265;
  assign \new_[67430]_  = A202 & \new_[67429]_ ;
  assign \new_[67433]_  = A269 & A267;
  assign \new_[67436]_  = A301 & ~A300;
  assign \new_[67437]_  = \new_[67436]_  & \new_[67433]_ ;
  assign \new_[67438]_  = \new_[67437]_  & \new_[67430]_ ;
  assign \new_[67442]_  = ~A167 & A168;
  assign \new_[67443]_  = A169 & \new_[67442]_ ;
  assign \new_[67446]_  = A199 & A166;
  assign \new_[67449]_  = A201 & ~A200;
  assign \new_[67450]_  = \new_[67449]_  & \new_[67446]_ ;
  assign \new_[67451]_  = \new_[67450]_  & \new_[67443]_ ;
  assign \new_[67455]_  = ~A266 & A265;
  assign \new_[67456]_  = A202 & \new_[67455]_ ;
  assign \new_[67459]_  = A269 & A267;
  assign \new_[67462]_  = A302 & ~A300;
  assign \new_[67463]_  = \new_[67462]_  & \new_[67459]_ ;
  assign \new_[67464]_  = \new_[67463]_  & \new_[67456]_ ;
  assign \new_[67468]_  = ~A167 & A168;
  assign \new_[67469]_  = A169 & \new_[67468]_ ;
  assign \new_[67472]_  = A199 & A166;
  assign \new_[67475]_  = A201 & ~A200;
  assign \new_[67476]_  = \new_[67475]_  & \new_[67472]_ ;
  assign \new_[67477]_  = \new_[67476]_  & \new_[67469]_ ;
  assign \new_[67481]_  = ~A266 & A265;
  assign \new_[67482]_  = A202 & \new_[67481]_ ;
  assign \new_[67485]_  = A269 & A267;
  assign \new_[67488]_  = A299 & A298;
  assign \new_[67489]_  = \new_[67488]_  & \new_[67485]_ ;
  assign \new_[67490]_  = \new_[67489]_  & \new_[67482]_ ;
  assign \new_[67494]_  = ~A167 & A168;
  assign \new_[67495]_  = A169 & \new_[67494]_ ;
  assign \new_[67498]_  = A199 & A166;
  assign \new_[67501]_  = A201 & ~A200;
  assign \new_[67502]_  = \new_[67501]_  & \new_[67498]_ ;
  assign \new_[67503]_  = \new_[67502]_  & \new_[67495]_ ;
  assign \new_[67507]_  = ~A266 & A265;
  assign \new_[67508]_  = A202 & \new_[67507]_ ;
  assign \new_[67511]_  = A269 & A267;
  assign \new_[67514]_  = ~A299 & ~A298;
  assign \new_[67515]_  = \new_[67514]_  & \new_[67511]_ ;
  assign \new_[67516]_  = \new_[67515]_  & \new_[67508]_ ;
  assign \new_[67520]_  = ~A167 & A168;
  assign \new_[67521]_  = A169 & \new_[67520]_ ;
  assign \new_[67524]_  = A199 & A166;
  assign \new_[67527]_  = A201 & ~A200;
  assign \new_[67528]_  = \new_[67527]_  & \new_[67524]_ ;
  assign \new_[67529]_  = \new_[67528]_  & \new_[67521]_ ;
  assign \new_[67533]_  = A266 & ~A265;
  assign \new_[67534]_  = A203 & \new_[67533]_ ;
  assign \new_[67537]_  = A268 & A267;
  assign \new_[67540]_  = A301 & ~A300;
  assign \new_[67541]_  = \new_[67540]_  & \new_[67537]_ ;
  assign \new_[67542]_  = \new_[67541]_  & \new_[67534]_ ;
  assign \new_[67546]_  = ~A167 & A168;
  assign \new_[67547]_  = A169 & \new_[67546]_ ;
  assign \new_[67550]_  = A199 & A166;
  assign \new_[67553]_  = A201 & ~A200;
  assign \new_[67554]_  = \new_[67553]_  & \new_[67550]_ ;
  assign \new_[67555]_  = \new_[67554]_  & \new_[67547]_ ;
  assign \new_[67559]_  = A266 & ~A265;
  assign \new_[67560]_  = A203 & \new_[67559]_ ;
  assign \new_[67563]_  = A268 & A267;
  assign \new_[67566]_  = A302 & ~A300;
  assign \new_[67567]_  = \new_[67566]_  & \new_[67563]_ ;
  assign \new_[67568]_  = \new_[67567]_  & \new_[67560]_ ;
  assign \new_[67572]_  = ~A167 & A168;
  assign \new_[67573]_  = A169 & \new_[67572]_ ;
  assign \new_[67576]_  = A199 & A166;
  assign \new_[67579]_  = A201 & ~A200;
  assign \new_[67580]_  = \new_[67579]_  & \new_[67576]_ ;
  assign \new_[67581]_  = \new_[67580]_  & \new_[67573]_ ;
  assign \new_[67585]_  = A266 & ~A265;
  assign \new_[67586]_  = A203 & \new_[67585]_ ;
  assign \new_[67589]_  = A268 & A267;
  assign \new_[67592]_  = A299 & A298;
  assign \new_[67593]_  = \new_[67592]_  & \new_[67589]_ ;
  assign \new_[67594]_  = \new_[67593]_  & \new_[67586]_ ;
  assign \new_[67598]_  = ~A167 & A168;
  assign \new_[67599]_  = A169 & \new_[67598]_ ;
  assign \new_[67602]_  = A199 & A166;
  assign \new_[67605]_  = A201 & ~A200;
  assign \new_[67606]_  = \new_[67605]_  & \new_[67602]_ ;
  assign \new_[67607]_  = \new_[67606]_  & \new_[67599]_ ;
  assign \new_[67611]_  = A266 & ~A265;
  assign \new_[67612]_  = A203 & \new_[67611]_ ;
  assign \new_[67615]_  = A268 & A267;
  assign \new_[67618]_  = ~A299 & ~A298;
  assign \new_[67619]_  = \new_[67618]_  & \new_[67615]_ ;
  assign \new_[67620]_  = \new_[67619]_  & \new_[67612]_ ;
  assign \new_[67624]_  = ~A167 & A168;
  assign \new_[67625]_  = A169 & \new_[67624]_ ;
  assign \new_[67628]_  = A199 & A166;
  assign \new_[67631]_  = A201 & ~A200;
  assign \new_[67632]_  = \new_[67631]_  & \new_[67628]_ ;
  assign \new_[67633]_  = \new_[67632]_  & \new_[67625]_ ;
  assign \new_[67637]_  = A266 & ~A265;
  assign \new_[67638]_  = A203 & \new_[67637]_ ;
  assign \new_[67641]_  = A269 & A267;
  assign \new_[67644]_  = A301 & ~A300;
  assign \new_[67645]_  = \new_[67644]_  & \new_[67641]_ ;
  assign \new_[67646]_  = \new_[67645]_  & \new_[67638]_ ;
  assign \new_[67650]_  = ~A167 & A168;
  assign \new_[67651]_  = A169 & \new_[67650]_ ;
  assign \new_[67654]_  = A199 & A166;
  assign \new_[67657]_  = A201 & ~A200;
  assign \new_[67658]_  = \new_[67657]_  & \new_[67654]_ ;
  assign \new_[67659]_  = \new_[67658]_  & \new_[67651]_ ;
  assign \new_[67663]_  = A266 & ~A265;
  assign \new_[67664]_  = A203 & \new_[67663]_ ;
  assign \new_[67667]_  = A269 & A267;
  assign \new_[67670]_  = A302 & ~A300;
  assign \new_[67671]_  = \new_[67670]_  & \new_[67667]_ ;
  assign \new_[67672]_  = \new_[67671]_  & \new_[67664]_ ;
  assign \new_[67676]_  = ~A167 & A168;
  assign \new_[67677]_  = A169 & \new_[67676]_ ;
  assign \new_[67680]_  = A199 & A166;
  assign \new_[67683]_  = A201 & ~A200;
  assign \new_[67684]_  = \new_[67683]_  & \new_[67680]_ ;
  assign \new_[67685]_  = \new_[67684]_  & \new_[67677]_ ;
  assign \new_[67689]_  = A266 & ~A265;
  assign \new_[67690]_  = A203 & \new_[67689]_ ;
  assign \new_[67693]_  = A269 & A267;
  assign \new_[67696]_  = A299 & A298;
  assign \new_[67697]_  = \new_[67696]_  & \new_[67693]_ ;
  assign \new_[67698]_  = \new_[67697]_  & \new_[67690]_ ;
  assign \new_[67702]_  = ~A167 & A168;
  assign \new_[67703]_  = A169 & \new_[67702]_ ;
  assign \new_[67706]_  = A199 & A166;
  assign \new_[67709]_  = A201 & ~A200;
  assign \new_[67710]_  = \new_[67709]_  & \new_[67706]_ ;
  assign \new_[67711]_  = \new_[67710]_  & \new_[67703]_ ;
  assign \new_[67715]_  = A266 & ~A265;
  assign \new_[67716]_  = A203 & \new_[67715]_ ;
  assign \new_[67719]_  = A269 & A267;
  assign \new_[67722]_  = ~A299 & ~A298;
  assign \new_[67723]_  = \new_[67722]_  & \new_[67719]_ ;
  assign \new_[67724]_  = \new_[67723]_  & \new_[67716]_ ;
  assign \new_[67728]_  = ~A167 & A168;
  assign \new_[67729]_  = A169 & \new_[67728]_ ;
  assign \new_[67732]_  = A199 & A166;
  assign \new_[67735]_  = A201 & ~A200;
  assign \new_[67736]_  = \new_[67735]_  & \new_[67732]_ ;
  assign \new_[67737]_  = \new_[67736]_  & \new_[67729]_ ;
  assign \new_[67741]_  = ~A266 & A265;
  assign \new_[67742]_  = A203 & \new_[67741]_ ;
  assign \new_[67745]_  = A268 & A267;
  assign \new_[67748]_  = A301 & ~A300;
  assign \new_[67749]_  = \new_[67748]_  & \new_[67745]_ ;
  assign \new_[67750]_  = \new_[67749]_  & \new_[67742]_ ;
  assign \new_[67754]_  = ~A167 & A168;
  assign \new_[67755]_  = A169 & \new_[67754]_ ;
  assign \new_[67758]_  = A199 & A166;
  assign \new_[67761]_  = A201 & ~A200;
  assign \new_[67762]_  = \new_[67761]_  & \new_[67758]_ ;
  assign \new_[67763]_  = \new_[67762]_  & \new_[67755]_ ;
  assign \new_[67767]_  = ~A266 & A265;
  assign \new_[67768]_  = A203 & \new_[67767]_ ;
  assign \new_[67771]_  = A268 & A267;
  assign \new_[67774]_  = A302 & ~A300;
  assign \new_[67775]_  = \new_[67774]_  & \new_[67771]_ ;
  assign \new_[67776]_  = \new_[67775]_  & \new_[67768]_ ;
  assign \new_[67780]_  = ~A167 & A168;
  assign \new_[67781]_  = A169 & \new_[67780]_ ;
  assign \new_[67784]_  = A199 & A166;
  assign \new_[67787]_  = A201 & ~A200;
  assign \new_[67788]_  = \new_[67787]_  & \new_[67784]_ ;
  assign \new_[67789]_  = \new_[67788]_  & \new_[67781]_ ;
  assign \new_[67793]_  = ~A266 & A265;
  assign \new_[67794]_  = A203 & \new_[67793]_ ;
  assign \new_[67797]_  = A268 & A267;
  assign \new_[67800]_  = A299 & A298;
  assign \new_[67801]_  = \new_[67800]_  & \new_[67797]_ ;
  assign \new_[67802]_  = \new_[67801]_  & \new_[67794]_ ;
  assign \new_[67806]_  = ~A167 & A168;
  assign \new_[67807]_  = A169 & \new_[67806]_ ;
  assign \new_[67810]_  = A199 & A166;
  assign \new_[67813]_  = A201 & ~A200;
  assign \new_[67814]_  = \new_[67813]_  & \new_[67810]_ ;
  assign \new_[67815]_  = \new_[67814]_  & \new_[67807]_ ;
  assign \new_[67819]_  = ~A266 & A265;
  assign \new_[67820]_  = A203 & \new_[67819]_ ;
  assign \new_[67823]_  = A268 & A267;
  assign \new_[67826]_  = ~A299 & ~A298;
  assign \new_[67827]_  = \new_[67826]_  & \new_[67823]_ ;
  assign \new_[67828]_  = \new_[67827]_  & \new_[67820]_ ;
  assign \new_[67832]_  = ~A167 & A168;
  assign \new_[67833]_  = A169 & \new_[67832]_ ;
  assign \new_[67836]_  = A199 & A166;
  assign \new_[67839]_  = A201 & ~A200;
  assign \new_[67840]_  = \new_[67839]_  & \new_[67836]_ ;
  assign \new_[67841]_  = \new_[67840]_  & \new_[67833]_ ;
  assign \new_[67845]_  = ~A266 & A265;
  assign \new_[67846]_  = A203 & \new_[67845]_ ;
  assign \new_[67849]_  = A269 & A267;
  assign \new_[67852]_  = A301 & ~A300;
  assign \new_[67853]_  = \new_[67852]_  & \new_[67849]_ ;
  assign \new_[67854]_  = \new_[67853]_  & \new_[67846]_ ;
  assign \new_[67858]_  = ~A167 & A168;
  assign \new_[67859]_  = A169 & \new_[67858]_ ;
  assign \new_[67862]_  = A199 & A166;
  assign \new_[67865]_  = A201 & ~A200;
  assign \new_[67866]_  = \new_[67865]_  & \new_[67862]_ ;
  assign \new_[67867]_  = \new_[67866]_  & \new_[67859]_ ;
  assign \new_[67871]_  = ~A266 & A265;
  assign \new_[67872]_  = A203 & \new_[67871]_ ;
  assign \new_[67875]_  = A269 & A267;
  assign \new_[67878]_  = A302 & ~A300;
  assign \new_[67879]_  = \new_[67878]_  & \new_[67875]_ ;
  assign \new_[67880]_  = \new_[67879]_  & \new_[67872]_ ;
  assign \new_[67884]_  = ~A167 & A168;
  assign \new_[67885]_  = A169 & \new_[67884]_ ;
  assign \new_[67888]_  = A199 & A166;
  assign \new_[67891]_  = A201 & ~A200;
  assign \new_[67892]_  = \new_[67891]_  & \new_[67888]_ ;
  assign \new_[67893]_  = \new_[67892]_  & \new_[67885]_ ;
  assign \new_[67897]_  = ~A266 & A265;
  assign \new_[67898]_  = A203 & \new_[67897]_ ;
  assign \new_[67901]_  = A269 & A267;
  assign \new_[67904]_  = A299 & A298;
  assign \new_[67905]_  = \new_[67904]_  & \new_[67901]_ ;
  assign \new_[67906]_  = \new_[67905]_  & \new_[67898]_ ;
  assign \new_[67910]_  = ~A167 & A168;
  assign \new_[67911]_  = A169 & \new_[67910]_ ;
  assign \new_[67914]_  = A199 & A166;
  assign \new_[67917]_  = A201 & ~A200;
  assign \new_[67918]_  = \new_[67917]_  & \new_[67914]_ ;
  assign \new_[67919]_  = \new_[67918]_  & \new_[67911]_ ;
  assign \new_[67923]_  = ~A266 & A265;
  assign \new_[67924]_  = A203 & \new_[67923]_ ;
  assign \new_[67927]_  = A269 & A267;
  assign \new_[67930]_  = ~A299 & ~A298;
  assign \new_[67931]_  = \new_[67930]_  & \new_[67927]_ ;
  assign \new_[67932]_  = \new_[67931]_  & \new_[67924]_ ;
  assign \new_[67936]_  = ~A167 & A168;
  assign \new_[67937]_  = A169 & \new_[67936]_ ;
  assign \new_[67940]_  = ~A199 & A166;
  assign \new_[67943]_  = A267 & ~A200;
  assign \new_[67944]_  = \new_[67943]_  & \new_[67940]_ ;
  assign \new_[67945]_  = \new_[67944]_  & \new_[67937]_ ;
  assign \new_[67949]_  = A298 & ~A269;
  assign \new_[67950]_  = ~A268 & \new_[67949]_ ;
  assign \new_[67953]_  = ~A300 & ~A299;
  assign \new_[67956]_  = ~A302 & ~A301;
  assign \new_[67957]_  = \new_[67956]_  & \new_[67953]_ ;
  assign \new_[67958]_  = \new_[67957]_  & \new_[67950]_ ;
  assign \new_[67962]_  = ~A167 & A168;
  assign \new_[67963]_  = A169 & \new_[67962]_ ;
  assign \new_[67966]_  = ~A199 & A166;
  assign \new_[67969]_  = A267 & ~A200;
  assign \new_[67970]_  = \new_[67969]_  & \new_[67966]_ ;
  assign \new_[67971]_  = \new_[67970]_  & \new_[67963]_ ;
  assign \new_[67975]_  = ~A298 & ~A269;
  assign \new_[67976]_  = ~A268 & \new_[67975]_ ;
  assign \new_[67979]_  = ~A300 & A299;
  assign \new_[67982]_  = ~A302 & ~A301;
  assign \new_[67983]_  = \new_[67982]_  & \new_[67979]_ ;
  assign \new_[67984]_  = \new_[67983]_  & \new_[67976]_ ;
  assign \new_[67988]_  = ~A199 & ~A168;
  assign \new_[67989]_  = A169 & \new_[67988]_ ;
  assign \new_[67992]_  = A201 & A200;
  assign \new_[67995]_  = A267 & A202;
  assign \new_[67996]_  = \new_[67995]_  & \new_[67992]_ ;
  assign \new_[67997]_  = \new_[67996]_  & \new_[67989]_ ;
  assign \new_[68001]_  = A298 & ~A269;
  assign \new_[68002]_  = ~A268 & \new_[68001]_ ;
  assign \new_[68005]_  = ~A300 & ~A299;
  assign \new_[68008]_  = ~A302 & ~A301;
  assign \new_[68009]_  = \new_[68008]_  & \new_[68005]_ ;
  assign \new_[68010]_  = \new_[68009]_  & \new_[68002]_ ;
  assign \new_[68014]_  = ~A199 & ~A168;
  assign \new_[68015]_  = A169 & \new_[68014]_ ;
  assign \new_[68018]_  = A201 & A200;
  assign \new_[68021]_  = A267 & A202;
  assign \new_[68022]_  = \new_[68021]_  & \new_[68018]_ ;
  assign \new_[68023]_  = \new_[68022]_  & \new_[68015]_ ;
  assign \new_[68027]_  = ~A298 & ~A269;
  assign \new_[68028]_  = ~A268 & \new_[68027]_ ;
  assign \new_[68031]_  = ~A300 & A299;
  assign \new_[68034]_  = ~A302 & ~A301;
  assign \new_[68035]_  = \new_[68034]_  & \new_[68031]_ ;
  assign \new_[68036]_  = \new_[68035]_  & \new_[68028]_ ;
  assign \new_[68040]_  = ~A199 & ~A168;
  assign \new_[68041]_  = A169 & \new_[68040]_ ;
  assign \new_[68044]_  = A201 & A200;
  assign \new_[68047]_  = A267 & A203;
  assign \new_[68048]_  = \new_[68047]_  & \new_[68044]_ ;
  assign \new_[68049]_  = \new_[68048]_  & \new_[68041]_ ;
  assign \new_[68053]_  = A298 & ~A269;
  assign \new_[68054]_  = ~A268 & \new_[68053]_ ;
  assign \new_[68057]_  = ~A300 & ~A299;
  assign \new_[68060]_  = ~A302 & ~A301;
  assign \new_[68061]_  = \new_[68060]_  & \new_[68057]_ ;
  assign \new_[68062]_  = \new_[68061]_  & \new_[68054]_ ;
  assign \new_[68066]_  = ~A199 & ~A168;
  assign \new_[68067]_  = A169 & \new_[68066]_ ;
  assign \new_[68070]_  = A201 & A200;
  assign \new_[68073]_  = A267 & A203;
  assign \new_[68074]_  = \new_[68073]_  & \new_[68070]_ ;
  assign \new_[68075]_  = \new_[68074]_  & \new_[68067]_ ;
  assign \new_[68079]_  = ~A298 & ~A269;
  assign \new_[68080]_  = ~A268 & \new_[68079]_ ;
  assign \new_[68083]_  = ~A300 & A299;
  assign \new_[68086]_  = ~A302 & ~A301;
  assign \new_[68087]_  = \new_[68086]_  & \new_[68083]_ ;
  assign \new_[68088]_  = \new_[68087]_  & \new_[68080]_ ;
  assign \new_[68092]_  = ~A199 & ~A168;
  assign \new_[68093]_  = A169 & \new_[68092]_ ;
  assign \new_[68096]_  = ~A201 & A200;
  assign \new_[68099]_  = ~A203 & ~A202;
  assign \new_[68100]_  = \new_[68099]_  & \new_[68096]_ ;
  assign \new_[68101]_  = \new_[68100]_  & \new_[68093]_ ;
  assign \new_[68105]_  = ~A269 & ~A268;
  assign \new_[68106]_  = A267 & \new_[68105]_ ;
  assign \new_[68109]_  = ~A299 & A298;
  assign \new_[68112]_  = A301 & A300;
  assign \new_[68113]_  = \new_[68112]_  & \new_[68109]_ ;
  assign \new_[68114]_  = \new_[68113]_  & \new_[68106]_ ;
  assign \new_[68118]_  = ~A199 & ~A168;
  assign \new_[68119]_  = A169 & \new_[68118]_ ;
  assign \new_[68122]_  = ~A201 & A200;
  assign \new_[68125]_  = ~A203 & ~A202;
  assign \new_[68126]_  = \new_[68125]_  & \new_[68122]_ ;
  assign \new_[68127]_  = \new_[68126]_  & \new_[68119]_ ;
  assign \new_[68131]_  = ~A269 & ~A268;
  assign \new_[68132]_  = A267 & \new_[68131]_ ;
  assign \new_[68135]_  = ~A299 & A298;
  assign \new_[68138]_  = A302 & A300;
  assign \new_[68139]_  = \new_[68138]_  & \new_[68135]_ ;
  assign \new_[68140]_  = \new_[68139]_  & \new_[68132]_ ;
  assign \new_[68144]_  = ~A199 & ~A168;
  assign \new_[68145]_  = A169 & \new_[68144]_ ;
  assign \new_[68148]_  = ~A201 & A200;
  assign \new_[68151]_  = ~A203 & ~A202;
  assign \new_[68152]_  = \new_[68151]_  & \new_[68148]_ ;
  assign \new_[68153]_  = \new_[68152]_  & \new_[68145]_ ;
  assign \new_[68157]_  = ~A269 & ~A268;
  assign \new_[68158]_  = A267 & \new_[68157]_ ;
  assign \new_[68161]_  = A299 & ~A298;
  assign \new_[68164]_  = A301 & A300;
  assign \new_[68165]_  = \new_[68164]_  & \new_[68161]_ ;
  assign \new_[68166]_  = \new_[68165]_  & \new_[68158]_ ;
  assign \new_[68170]_  = ~A199 & ~A168;
  assign \new_[68171]_  = A169 & \new_[68170]_ ;
  assign \new_[68174]_  = ~A201 & A200;
  assign \new_[68177]_  = ~A203 & ~A202;
  assign \new_[68178]_  = \new_[68177]_  & \new_[68174]_ ;
  assign \new_[68179]_  = \new_[68178]_  & \new_[68171]_ ;
  assign \new_[68183]_  = ~A269 & ~A268;
  assign \new_[68184]_  = A267 & \new_[68183]_ ;
  assign \new_[68187]_  = A299 & ~A298;
  assign \new_[68190]_  = A302 & A300;
  assign \new_[68191]_  = \new_[68190]_  & \new_[68187]_ ;
  assign \new_[68192]_  = \new_[68191]_  & \new_[68184]_ ;
  assign \new_[68196]_  = ~A199 & ~A168;
  assign \new_[68197]_  = A169 & \new_[68196]_ ;
  assign \new_[68200]_  = ~A201 & A200;
  assign \new_[68203]_  = ~A203 & ~A202;
  assign \new_[68204]_  = \new_[68203]_  & \new_[68200]_ ;
  assign \new_[68205]_  = \new_[68204]_  & \new_[68197]_ ;
  assign \new_[68209]_  = A298 & A268;
  assign \new_[68210]_  = ~A267 & \new_[68209]_ ;
  assign \new_[68213]_  = ~A300 & ~A299;
  assign \new_[68216]_  = ~A302 & ~A301;
  assign \new_[68217]_  = \new_[68216]_  & \new_[68213]_ ;
  assign \new_[68218]_  = \new_[68217]_  & \new_[68210]_ ;
  assign \new_[68222]_  = ~A199 & ~A168;
  assign \new_[68223]_  = A169 & \new_[68222]_ ;
  assign \new_[68226]_  = ~A201 & A200;
  assign \new_[68229]_  = ~A203 & ~A202;
  assign \new_[68230]_  = \new_[68229]_  & \new_[68226]_ ;
  assign \new_[68231]_  = \new_[68230]_  & \new_[68223]_ ;
  assign \new_[68235]_  = ~A298 & A268;
  assign \new_[68236]_  = ~A267 & \new_[68235]_ ;
  assign \new_[68239]_  = ~A300 & A299;
  assign \new_[68242]_  = ~A302 & ~A301;
  assign \new_[68243]_  = \new_[68242]_  & \new_[68239]_ ;
  assign \new_[68244]_  = \new_[68243]_  & \new_[68236]_ ;
  assign \new_[68248]_  = ~A199 & ~A168;
  assign \new_[68249]_  = A169 & \new_[68248]_ ;
  assign \new_[68252]_  = ~A201 & A200;
  assign \new_[68255]_  = ~A203 & ~A202;
  assign \new_[68256]_  = \new_[68255]_  & \new_[68252]_ ;
  assign \new_[68257]_  = \new_[68256]_  & \new_[68249]_ ;
  assign \new_[68261]_  = A298 & A269;
  assign \new_[68262]_  = ~A267 & \new_[68261]_ ;
  assign \new_[68265]_  = ~A300 & ~A299;
  assign \new_[68268]_  = ~A302 & ~A301;
  assign \new_[68269]_  = \new_[68268]_  & \new_[68265]_ ;
  assign \new_[68270]_  = \new_[68269]_  & \new_[68262]_ ;
  assign \new_[68274]_  = ~A199 & ~A168;
  assign \new_[68275]_  = A169 & \new_[68274]_ ;
  assign \new_[68278]_  = ~A201 & A200;
  assign \new_[68281]_  = ~A203 & ~A202;
  assign \new_[68282]_  = \new_[68281]_  & \new_[68278]_ ;
  assign \new_[68283]_  = \new_[68282]_  & \new_[68275]_ ;
  assign \new_[68287]_  = ~A298 & A269;
  assign \new_[68288]_  = ~A267 & \new_[68287]_ ;
  assign \new_[68291]_  = ~A300 & A299;
  assign \new_[68294]_  = ~A302 & ~A301;
  assign \new_[68295]_  = \new_[68294]_  & \new_[68291]_ ;
  assign \new_[68296]_  = \new_[68295]_  & \new_[68288]_ ;
  assign \new_[68300]_  = ~A199 & ~A168;
  assign \new_[68301]_  = A169 & \new_[68300]_ ;
  assign \new_[68304]_  = ~A201 & A200;
  assign \new_[68307]_  = ~A203 & ~A202;
  assign \new_[68308]_  = \new_[68307]_  & \new_[68304]_ ;
  assign \new_[68309]_  = \new_[68308]_  & \new_[68301]_ ;
  assign \new_[68313]_  = A298 & A266;
  assign \new_[68314]_  = A265 & \new_[68313]_ ;
  assign \new_[68317]_  = ~A300 & ~A299;
  assign \new_[68320]_  = ~A302 & ~A301;
  assign \new_[68321]_  = \new_[68320]_  & \new_[68317]_ ;
  assign \new_[68322]_  = \new_[68321]_  & \new_[68314]_ ;
  assign \new_[68326]_  = ~A199 & ~A168;
  assign \new_[68327]_  = A169 & \new_[68326]_ ;
  assign \new_[68330]_  = ~A201 & A200;
  assign \new_[68333]_  = ~A203 & ~A202;
  assign \new_[68334]_  = \new_[68333]_  & \new_[68330]_ ;
  assign \new_[68335]_  = \new_[68334]_  & \new_[68327]_ ;
  assign \new_[68339]_  = ~A298 & A266;
  assign \new_[68340]_  = A265 & \new_[68339]_ ;
  assign \new_[68343]_  = ~A300 & A299;
  assign \new_[68346]_  = ~A302 & ~A301;
  assign \new_[68347]_  = \new_[68346]_  & \new_[68343]_ ;
  assign \new_[68348]_  = \new_[68347]_  & \new_[68340]_ ;
  assign \new_[68352]_  = ~A199 & ~A168;
  assign \new_[68353]_  = A169 & \new_[68352]_ ;
  assign \new_[68356]_  = ~A201 & A200;
  assign \new_[68359]_  = ~A203 & ~A202;
  assign \new_[68360]_  = \new_[68359]_  & \new_[68356]_ ;
  assign \new_[68361]_  = \new_[68360]_  & \new_[68353]_ ;
  assign \new_[68365]_  = A298 & ~A266;
  assign \new_[68366]_  = ~A265 & \new_[68365]_ ;
  assign \new_[68369]_  = ~A300 & ~A299;
  assign \new_[68372]_  = ~A302 & ~A301;
  assign \new_[68373]_  = \new_[68372]_  & \new_[68369]_ ;
  assign \new_[68374]_  = \new_[68373]_  & \new_[68366]_ ;
  assign \new_[68378]_  = ~A199 & ~A168;
  assign \new_[68379]_  = A169 & \new_[68378]_ ;
  assign \new_[68382]_  = ~A201 & A200;
  assign \new_[68385]_  = ~A203 & ~A202;
  assign \new_[68386]_  = \new_[68385]_  & \new_[68382]_ ;
  assign \new_[68387]_  = \new_[68386]_  & \new_[68379]_ ;
  assign \new_[68391]_  = ~A298 & ~A266;
  assign \new_[68392]_  = ~A265 & \new_[68391]_ ;
  assign \new_[68395]_  = ~A300 & A299;
  assign \new_[68398]_  = ~A302 & ~A301;
  assign \new_[68399]_  = \new_[68398]_  & \new_[68395]_ ;
  assign \new_[68400]_  = \new_[68399]_  & \new_[68392]_ ;
  assign \new_[68404]_  = A199 & ~A168;
  assign \new_[68405]_  = A169 & \new_[68404]_ ;
  assign \new_[68408]_  = A201 & ~A200;
  assign \new_[68411]_  = A267 & A202;
  assign \new_[68412]_  = \new_[68411]_  & \new_[68408]_ ;
  assign \new_[68413]_  = \new_[68412]_  & \new_[68405]_ ;
  assign \new_[68417]_  = A298 & ~A269;
  assign \new_[68418]_  = ~A268 & \new_[68417]_ ;
  assign \new_[68421]_  = ~A300 & ~A299;
  assign \new_[68424]_  = ~A302 & ~A301;
  assign \new_[68425]_  = \new_[68424]_  & \new_[68421]_ ;
  assign \new_[68426]_  = \new_[68425]_  & \new_[68418]_ ;
  assign \new_[68430]_  = A199 & ~A168;
  assign \new_[68431]_  = A169 & \new_[68430]_ ;
  assign \new_[68434]_  = A201 & ~A200;
  assign \new_[68437]_  = A267 & A202;
  assign \new_[68438]_  = \new_[68437]_  & \new_[68434]_ ;
  assign \new_[68439]_  = \new_[68438]_  & \new_[68431]_ ;
  assign \new_[68443]_  = ~A298 & ~A269;
  assign \new_[68444]_  = ~A268 & \new_[68443]_ ;
  assign \new_[68447]_  = ~A300 & A299;
  assign \new_[68450]_  = ~A302 & ~A301;
  assign \new_[68451]_  = \new_[68450]_  & \new_[68447]_ ;
  assign \new_[68452]_  = \new_[68451]_  & \new_[68444]_ ;
  assign \new_[68456]_  = A199 & ~A168;
  assign \new_[68457]_  = A169 & \new_[68456]_ ;
  assign \new_[68460]_  = A201 & ~A200;
  assign \new_[68463]_  = A267 & A203;
  assign \new_[68464]_  = \new_[68463]_  & \new_[68460]_ ;
  assign \new_[68465]_  = \new_[68464]_  & \new_[68457]_ ;
  assign \new_[68469]_  = A298 & ~A269;
  assign \new_[68470]_  = ~A268 & \new_[68469]_ ;
  assign \new_[68473]_  = ~A300 & ~A299;
  assign \new_[68476]_  = ~A302 & ~A301;
  assign \new_[68477]_  = \new_[68476]_  & \new_[68473]_ ;
  assign \new_[68478]_  = \new_[68477]_  & \new_[68470]_ ;
  assign \new_[68482]_  = A199 & ~A168;
  assign \new_[68483]_  = A169 & \new_[68482]_ ;
  assign \new_[68486]_  = A201 & ~A200;
  assign \new_[68489]_  = A267 & A203;
  assign \new_[68490]_  = \new_[68489]_  & \new_[68486]_ ;
  assign \new_[68491]_  = \new_[68490]_  & \new_[68483]_ ;
  assign \new_[68495]_  = ~A298 & ~A269;
  assign \new_[68496]_  = ~A268 & \new_[68495]_ ;
  assign \new_[68499]_  = ~A300 & A299;
  assign \new_[68502]_  = ~A302 & ~A301;
  assign \new_[68503]_  = \new_[68502]_  & \new_[68499]_ ;
  assign \new_[68504]_  = \new_[68503]_  & \new_[68496]_ ;
  assign \new_[68508]_  = A199 & ~A168;
  assign \new_[68509]_  = A169 & \new_[68508]_ ;
  assign \new_[68512]_  = ~A201 & ~A200;
  assign \new_[68515]_  = ~A203 & ~A202;
  assign \new_[68516]_  = \new_[68515]_  & \new_[68512]_ ;
  assign \new_[68517]_  = \new_[68516]_  & \new_[68509]_ ;
  assign \new_[68521]_  = ~A269 & ~A268;
  assign \new_[68522]_  = A267 & \new_[68521]_ ;
  assign \new_[68525]_  = ~A299 & A298;
  assign \new_[68528]_  = A301 & A300;
  assign \new_[68529]_  = \new_[68528]_  & \new_[68525]_ ;
  assign \new_[68530]_  = \new_[68529]_  & \new_[68522]_ ;
  assign \new_[68534]_  = A199 & ~A168;
  assign \new_[68535]_  = A169 & \new_[68534]_ ;
  assign \new_[68538]_  = ~A201 & ~A200;
  assign \new_[68541]_  = ~A203 & ~A202;
  assign \new_[68542]_  = \new_[68541]_  & \new_[68538]_ ;
  assign \new_[68543]_  = \new_[68542]_  & \new_[68535]_ ;
  assign \new_[68547]_  = ~A269 & ~A268;
  assign \new_[68548]_  = A267 & \new_[68547]_ ;
  assign \new_[68551]_  = ~A299 & A298;
  assign \new_[68554]_  = A302 & A300;
  assign \new_[68555]_  = \new_[68554]_  & \new_[68551]_ ;
  assign \new_[68556]_  = \new_[68555]_  & \new_[68548]_ ;
  assign \new_[68560]_  = A199 & ~A168;
  assign \new_[68561]_  = A169 & \new_[68560]_ ;
  assign \new_[68564]_  = ~A201 & ~A200;
  assign \new_[68567]_  = ~A203 & ~A202;
  assign \new_[68568]_  = \new_[68567]_  & \new_[68564]_ ;
  assign \new_[68569]_  = \new_[68568]_  & \new_[68561]_ ;
  assign \new_[68573]_  = ~A269 & ~A268;
  assign \new_[68574]_  = A267 & \new_[68573]_ ;
  assign \new_[68577]_  = A299 & ~A298;
  assign \new_[68580]_  = A301 & A300;
  assign \new_[68581]_  = \new_[68580]_  & \new_[68577]_ ;
  assign \new_[68582]_  = \new_[68581]_  & \new_[68574]_ ;
  assign \new_[68586]_  = A199 & ~A168;
  assign \new_[68587]_  = A169 & \new_[68586]_ ;
  assign \new_[68590]_  = ~A201 & ~A200;
  assign \new_[68593]_  = ~A203 & ~A202;
  assign \new_[68594]_  = \new_[68593]_  & \new_[68590]_ ;
  assign \new_[68595]_  = \new_[68594]_  & \new_[68587]_ ;
  assign \new_[68599]_  = ~A269 & ~A268;
  assign \new_[68600]_  = A267 & \new_[68599]_ ;
  assign \new_[68603]_  = A299 & ~A298;
  assign \new_[68606]_  = A302 & A300;
  assign \new_[68607]_  = \new_[68606]_  & \new_[68603]_ ;
  assign \new_[68608]_  = \new_[68607]_  & \new_[68600]_ ;
  assign \new_[68612]_  = A199 & ~A168;
  assign \new_[68613]_  = A169 & \new_[68612]_ ;
  assign \new_[68616]_  = ~A201 & ~A200;
  assign \new_[68619]_  = ~A203 & ~A202;
  assign \new_[68620]_  = \new_[68619]_  & \new_[68616]_ ;
  assign \new_[68621]_  = \new_[68620]_  & \new_[68613]_ ;
  assign \new_[68625]_  = A298 & A268;
  assign \new_[68626]_  = ~A267 & \new_[68625]_ ;
  assign \new_[68629]_  = ~A300 & ~A299;
  assign \new_[68632]_  = ~A302 & ~A301;
  assign \new_[68633]_  = \new_[68632]_  & \new_[68629]_ ;
  assign \new_[68634]_  = \new_[68633]_  & \new_[68626]_ ;
  assign \new_[68638]_  = A199 & ~A168;
  assign \new_[68639]_  = A169 & \new_[68638]_ ;
  assign \new_[68642]_  = ~A201 & ~A200;
  assign \new_[68645]_  = ~A203 & ~A202;
  assign \new_[68646]_  = \new_[68645]_  & \new_[68642]_ ;
  assign \new_[68647]_  = \new_[68646]_  & \new_[68639]_ ;
  assign \new_[68651]_  = ~A298 & A268;
  assign \new_[68652]_  = ~A267 & \new_[68651]_ ;
  assign \new_[68655]_  = ~A300 & A299;
  assign \new_[68658]_  = ~A302 & ~A301;
  assign \new_[68659]_  = \new_[68658]_  & \new_[68655]_ ;
  assign \new_[68660]_  = \new_[68659]_  & \new_[68652]_ ;
  assign \new_[68664]_  = A199 & ~A168;
  assign \new_[68665]_  = A169 & \new_[68664]_ ;
  assign \new_[68668]_  = ~A201 & ~A200;
  assign \new_[68671]_  = ~A203 & ~A202;
  assign \new_[68672]_  = \new_[68671]_  & \new_[68668]_ ;
  assign \new_[68673]_  = \new_[68672]_  & \new_[68665]_ ;
  assign \new_[68677]_  = A298 & A269;
  assign \new_[68678]_  = ~A267 & \new_[68677]_ ;
  assign \new_[68681]_  = ~A300 & ~A299;
  assign \new_[68684]_  = ~A302 & ~A301;
  assign \new_[68685]_  = \new_[68684]_  & \new_[68681]_ ;
  assign \new_[68686]_  = \new_[68685]_  & \new_[68678]_ ;
  assign \new_[68690]_  = A199 & ~A168;
  assign \new_[68691]_  = A169 & \new_[68690]_ ;
  assign \new_[68694]_  = ~A201 & ~A200;
  assign \new_[68697]_  = ~A203 & ~A202;
  assign \new_[68698]_  = \new_[68697]_  & \new_[68694]_ ;
  assign \new_[68699]_  = \new_[68698]_  & \new_[68691]_ ;
  assign \new_[68703]_  = ~A298 & A269;
  assign \new_[68704]_  = ~A267 & \new_[68703]_ ;
  assign \new_[68707]_  = ~A300 & A299;
  assign \new_[68710]_  = ~A302 & ~A301;
  assign \new_[68711]_  = \new_[68710]_  & \new_[68707]_ ;
  assign \new_[68712]_  = \new_[68711]_  & \new_[68704]_ ;
  assign \new_[68716]_  = A199 & ~A168;
  assign \new_[68717]_  = A169 & \new_[68716]_ ;
  assign \new_[68720]_  = ~A201 & ~A200;
  assign \new_[68723]_  = ~A203 & ~A202;
  assign \new_[68724]_  = \new_[68723]_  & \new_[68720]_ ;
  assign \new_[68725]_  = \new_[68724]_  & \new_[68717]_ ;
  assign \new_[68729]_  = A298 & A266;
  assign \new_[68730]_  = A265 & \new_[68729]_ ;
  assign \new_[68733]_  = ~A300 & ~A299;
  assign \new_[68736]_  = ~A302 & ~A301;
  assign \new_[68737]_  = \new_[68736]_  & \new_[68733]_ ;
  assign \new_[68738]_  = \new_[68737]_  & \new_[68730]_ ;
  assign \new_[68742]_  = A199 & ~A168;
  assign \new_[68743]_  = A169 & \new_[68742]_ ;
  assign \new_[68746]_  = ~A201 & ~A200;
  assign \new_[68749]_  = ~A203 & ~A202;
  assign \new_[68750]_  = \new_[68749]_  & \new_[68746]_ ;
  assign \new_[68751]_  = \new_[68750]_  & \new_[68743]_ ;
  assign \new_[68755]_  = ~A298 & A266;
  assign \new_[68756]_  = A265 & \new_[68755]_ ;
  assign \new_[68759]_  = ~A300 & A299;
  assign \new_[68762]_  = ~A302 & ~A301;
  assign \new_[68763]_  = \new_[68762]_  & \new_[68759]_ ;
  assign \new_[68764]_  = \new_[68763]_  & \new_[68756]_ ;
  assign \new_[68768]_  = A199 & ~A168;
  assign \new_[68769]_  = A169 & \new_[68768]_ ;
  assign \new_[68772]_  = ~A201 & ~A200;
  assign \new_[68775]_  = ~A203 & ~A202;
  assign \new_[68776]_  = \new_[68775]_  & \new_[68772]_ ;
  assign \new_[68777]_  = \new_[68776]_  & \new_[68769]_ ;
  assign \new_[68781]_  = A298 & ~A266;
  assign \new_[68782]_  = ~A265 & \new_[68781]_ ;
  assign \new_[68785]_  = ~A300 & ~A299;
  assign \new_[68788]_  = ~A302 & ~A301;
  assign \new_[68789]_  = \new_[68788]_  & \new_[68785]_ ;
  assign \new_[68790]_  = \new_[68789]_  & \new_[68782]_ ;
  assign \new_[68794]_  = A199 & ~A168;
  assign \new_[68795]_  = A169 & \new_[68794]_ ;
  assign \new_[68798]_  = ~A201 & ~A200;
  assign \new_[68801]_  = ~A203 & ~A202;
  assign \new_[68802]_  = \new_[68801]_  & \new_[68798]_ ;
  assign \new_[68803]_  = \new_[68802]_  & \new_[68795]_ ;
  assign \new_[68807]_  = ~A298 & ~A266;
  assign \new_[68808]_  = ~A265 & \new_[68807]_ ;
  assign \new_[68811]_  = ~A300 & A299;
  assign \new_[68814]_  = ~A302 & ~A301;
  assign \new_[68815]_  = \new_[68814]_  & \new_[68811]_ ;
  assign \new_[68816]_  = \new_[68815]_  & \new_[68808]_ ;
  assign \new_[68820]_  = A168 & ~A169;
  assign \new_[68821]_  = A170 & \new_[68820]_ ;
  assign \new_[68824]_  = ~A202 & A201;
  assign \new_[68827]_  = ~A265 & ~A203;
  assign \new_[68828]_  = \new_[68827]_  & \new_[68824]_ ;
  assign \new_[68829]_  = \new_[68828]_  & \new_[68821]_ ;
  assign \new_[68833]_  = ~A268 & ~A267;
  assign \new_[68834]_  = A266 & \new_[68833]_ ;
  assign \new_[68837]_  = A300 & ~A269;
  assign \new_[68840]_  = ~A302 & ~A301;
  assign \new_[68841]_  = \new_[68840]_  & \new_[68837]_ ;
  assign \new_[68842]_  = \new_[68841]_  & \new_[68834]_ ;
  assign \new_[68846]_  = A168 & ~A169;
  assign \new_[68847]_  = A170 & \new_[68846]_ ;
  assign \new_[68850]_  = ~A202 & A201;
  assign \new_[68853]_  = A265 & ~A203;
  assign \new_[68854]_  = \new_[68853]_  & \new_[68850]_ ;
  assign \new_[68855]_  = \new_[68854]_  & \new_[68847]_ ;
  assign \new_[68859]_  = ~A268 & ~A267;
  assign \new_[68860]_  = ~A266 & \new_[68859]_ ;
  assign \new_[68863]_  = A300 & ~A269;
  assign \new_[68866]_  = ~A302 & ~A301;
  assign \new_[68867]_  = \new_[68866]_  & \new_[68863]_ ;
  assign \new_[68868]_  = \new_[68867]_  & \new_[68860]_ ;
  assign \new_[68872]_  = A168 & ~A169;
  assign \new_[68873]_  = A170 & \new_[68872]_ ;
  assign \new_[68876]_  = A200 & ~A199;
  assign \new_[68879]_  = A202 & A201;
  assign \new_[68880]_  = \new_[68879]_  & \new_[68876]_ ;
  assign \new_[68881]_  = \new_[68880]_  & \new_[68873]_ ;
  assign \new_[68885]_  = ~A269 & ~A268;
  assign \new_[68886]_  = A267 & \new_[68885]_ ;
  assign \new_[68889]_  = ~A299 & A298;
  assign \new_[68892]_  = A301 & A300;
  assign \new_[68893]_  = \new_[68892]_  & \new_[68889]_ ;
  assign \new_[68894]_  = \new_[68893]_  & \new_[68886]_ ;
  assign \new_[68898]_  = A168 & ~A169;
  assign \new_[68899]_  = A170 & \new_[68898]_ ;
  assign \new_[68902]_  = A200 & ~A199;
  assign \new_[68905]_  = A202 & A201;
  assign \new_[68906]_  = \new_[68905]_  & \new_[68902]_ ;
  assign \new_[68907]_  = \new_[68906]_  & \new_[68899]_ ;
  assign \new_[68911]_  = ~A269 & ~A268;
  assign \new_[68912]_  = A267 & \new_[68911]_ ;
  assign \new_[68915]_  = ~A299 & A298;
  assign \new_[68918]_  = A302 & A300;
  assign \new_[68919]_  = \new_[68918]_  & \new_[68915]_ ;
  assign \new_[68920]_  = \new_[68919]_  & \new_[68912]_ ;
  assign \new_[68924]_  = A168 & ~A169;
  assign \new_[68925]_  = A170 & \new_[68924]_ ;
  assign \new_[68928]_  = A200 & ~A199;
  assign \new_[68931]_  = A202 & A201;
  assign \new_[68932]_  = \new_[68931]_  & \new_[68928]_ ;
  assign \new_[68933]_  = \new_[68932]_  & \new_[68925]_ ;
  assign \new_[68937]_  = ~A269 & ~A268;
  assign \new_[68938]_  = A267 & \new_[68937]_ ;
  assign \new_[68941]_  = A299 & ~A298;
  assign \new_[68944]_  = A301 & A300;
  assign \new_[68945]_  = \new_[68944]_  & \new_[68941]_ ;
  assign \new_[68946]_  = \new_[68945]_  & \new_[68938]_ ;
  assign \new_[68950]_  = A168 & ~A169;
  assign \new_[68951]_  = A170 & \new_[68950]_ ;
  assign \new_[68954]_  = A200 & ~A199;
  assign \new_[68957]_  = A202 & A201;
  assign \new_[68958]_  = \new_[68957]_  & \new_[68954]_ ;
  assign \new_[68959]_  = \new_[68958]_  & \new_[68951]_ ;
  assign \new_[68963]_  = ~A269 & ~A268;
  assign \new_[68964]_  = A267 & \new_[68963]_ ;
  assign \new_[68967]_  = A299 & ~A298;
  assign \new_[68970]_  = A302 & A300;
  assign \new_[68971]_  = \new_[68970]_  & \new_[68967]_ ;
  assign \new_[68972]_  = \new_[68971]_  & \new_[68964]_ ;
  assign \new_[68976]_  = A168 & ~A169;
  assign \new_[68977]_  = A170 & \new_[68976]_ ;
  assign \new_[68980]_  = A200 & ~A199;
  assign \new_[68983]_  = A202 & A201;
  assign \new_[68984]_  = \new_[68983]_  & \new_[68980]_ ;
  assign \new_[68985]_  = \new_[68984]_  & \new_[68977]_ ;
  assign \new_[68989]_  = A298 & A268;
  assign \new_[68990]_  = ~A267 & \new_[68989]_ ;
  assign \new_[68993]_  = ~A300 & ~A299;
  assign \new_[68996]_  = ~A302 & ~A301;
  assign \new_[68997]_  = \new_[68996]_  & \new_[68993]_ ;
  assign \new_[68998]_  = \new_[68997]_  & \new_[68990]_ ;
  assign \new_[69002]_  = A168 & ~A169;
  assign \new_[69003]_  = A170 & \new_[69002]_ ;
  assign \new_[69006]_  = A200 & ~A199;
  assign \new_[69009]_  = A202 & A201;
  assign \new_[69010]_  = \new_[69009]_  & \new_[69006]_ ;
  assign \new_[69011]_  = \new_[69010]_  & \new_[69003]_ ;
  assign \new_[69015]_  = ~A298 & A268;
  assign \new_[69016]_  = ~A267 & \new_[69015]_ ;
  assign \new_[69019]_  = ~A300 & A299;
  assign \new_[69022]_  = ~A302 & ~A301;
  assign \new_[69023]_  = \new_[69022]_  & \new_[69019]_ ;
  assign \new_[69024]_  = \new_[69023]_  & \new_[69016]_ ;
  assign \new_[69028]_  = A168 & ~A169;
  assign \new_[69029]_  = A170 & \new_[69028]_ ;
  assign \new_[69032]_  = A200 & ~A199;
  assign \new_[69035]_  = A202 & A201;
  assign \new_[69036]_  = \new_[69035]_  & \new_[69032]_ ;
  assign \new_[69037]_  = \new_[69036]_  & \new_[69029]_ ;
  assign \new_[69041]_  = A298 & A269;
  assign \new_[69042]_  = ~A267 & \new_[69041]_ ;
  assign \new_[69045]_  = ~A300 & ~A299;
  assign \new_[69048]_  = ~A302 & ~A301;
  assign \new_[69049]_  = \new_[69048]_  & \new_[69045]_ ;
  assign \new_[69050]_  = \new_[69049]_  & \new_[69042]_ ;
  assign \new_[69054]_  = A168 & ~A169;
  assign \new_[69055]_  = A170 & \new_[69054]_ ;
  assign \new_[69058]_  = A200 & ~A199;
  assign \new_[69061]_  = A202 & A201;
  assign \new_[69062]_  = \new_[69061]_  & \new_[69058]_ ;
  assign \new_[69063]_  = \new_[69062]_  & \new_[69055]_ ;
  assign \new_[69067]_  = ~A298 & A269;
  assign \new_[69068]_  = ~A267 & \new_[69067]_ ;
  assign \new_[69071]_  = ~A300 & A299;
  assign \new_[69074]_  = ~A302 & ~A301;
  assign \new_[69075]_  = \new_[69074]_  & \new_[69071]_ ;
  assign \new_[69076]_  = \new_[69075]_  & \new_[69068]_ ;
  assign \new_[69080]_  = A168 & ~A169;
  assign \new_[69081]_  = A170 & \new_[69080]_ ;
  assign \new_[69084]_  = A200 & ~A199;
  assign \new_[69087]_  = A202 & A201;
  assign \new_[69088]_  = \new_[69087]_  & \new_[69084]_ ;
  assign \new_[69089]_  = \new_[69088]_  & \new_[69081]_ ;
  assign \new_[69093]_  = A298 & A266;
  assign \new_[69094]_  = A265 & \new_[69093]_ ;
  assign \new_[69097]_  = ~A300 & ~A299;
  assign \new_[69100]_  = ~A302 & ~A301;
  assign \new_[69101]_  = \new_[69100]_  & \new_[69097]_ ;
  assign \new_[69102]_  = \new_[69101]_  & \new_[69094]_ ;
  assign \new_[69106]_  = A168 & ~A169;
  assign \new_[69107]_  = A170 & \new_[69106]_ ;
  assign \new_[69110]_  = A200 & ~A199;
  assign \new_[69113]_  = A202 & A201;
  assign \new_[69114]_  = \new_[69113]_  & \new_[69110]_ ;
  assign \new_[69115]_  = \new_[69114]_  & \new_[69107]_ ;
  assign \new_[69119]_  = ~A298 & A266;
  assign \new_[69120]_  = A265 & \new_[69119]_ ;
  assign \new_[69123]_  = ~A300 & A299;
  assign \new_[69126]_  = ~A302 & ~A301;
  assign \new_[69127]_  = \new_[69126]_  & \new_[69123]_ ;
  assign \new_[69128]_  = \new_[69127]_  & \new_[69120]_ ;
  assign \new_[69132]_  = A168 & ~A169;
  assign \new_[69133]_  = A170 & \new_[69132]_ ;
  assign \new_[69136]_  = A200 & ~A199;
  assign \new_[69139]_  = A202 & A201;
  assign \new_[69140]_  = \new_[69139]_  & \new_[69136]_ ;
  assign \new_[69141]_  = \new_[69140]_  & \new_[69133]_ ;
  assign \new_[69145]_  = A298 & ~A266;
  assign \new_[69146]_  = ~A265 & \new_[69145]_ ;
  assign \new_[69149]_  = ~A300 & ~A299;
  assign \new_[69152]_  = ~A302 & ~A301;
  assign \new_[69153]_  = \new_[69152]_  & \new_[69149]_ ;
  assign \new_[69154]_  = \new_[69153]_  & \new_[69146]_ ;
  assign \new_[69158]_  = A168 & ~A169;
  assign \new_[69159]_  = A170 & \new_[69158]_ ;
  assign \new_[69162]_  = A200 & ~A199;
  assign \new_[69165]_  = A202 & A201;
  assign \new_[69166]_  = \new_[69165]_  & \new_[69162]_ ;
  assign \new_[69167]_  = \new_[69166]_  & \new_[69159]_ ;
  assign \new_[69171]_  = ~A298 & ~A266;
  assign \new_[69172]_  = ~A265 & \new_[69171]_ ;
  assign \new_[69175]_  = ~A300 & A299;
  assign \new_[69178]_  = ~A302 & ~A301;
  assign \new_[69179]_  = \new_[69178]_  & \new_[69175]_ ;
  assign \new_[69180]_  = \new_[69179]_  & \new_[69172]_ ;
  assign \new_[69184]_  = A168 & ~A169;
  assign \new_[69185]_  = A170 & \new_[69184]_ ;
  assign \new_[69188]_  = A200 & ~A199;
  assign \new_[69191]_  = A203 & A201;
  assign \new_[69192]_  = \new_[69191]_  & \new_[69188]_ ;
  assign \new_[69193]_  = \new_[69192]_  & \new_[69185]_ ;
  assign \new_[69197]_  = ~A269 & ~A268;
  assign \new_[69198]_  = A267 & \new_[69197]_ ;
  assign \new_[69201]_  = ~A299 & A298;
  assign \new_[69204]_  = A301 & A300;
  assign \new_[69205]_  = \new_[69204]_  & \new_[69201]_ ;
  assign \new_[69206]_  = \new_[69205]_  & \new_[69198]_ ;
  assign \new_[69210]_  = A168 & ~A169;
  assign \new_[69211]_  = A170 & \new_[69210]_ ;
  assign \new_[69214]_  = A200 & ~A199;
  assign \new_[69217]_  = A203 & A201;
  assign \new_[69218]_  = \new_[69217]_  & \new_[69214]_ ;
  assign \new_[69219]_  = \new_[69218]_  & \new_[69211]_ ;
  assign \new_[69223]_  = ~A269 & ~A268;
  assign \new_[69224]_  = A267 & \new_[69223]_ ;
  assign \new_[69227]_  = ~A299 & A298;
  assign \new_[69230]_  = A302 & A300;
  assign \new_[69231]_  = \new_[69230]_  & \new_[69227]_ ;
  assign \new_[69232]_  = \new_[69231]_  & \new_[69224]_ ;
  assign \new_[69236]_  = A168 & ~A169;
  assign \new_[69237]_  = A170 & \new_[69236]_ ;
  assign \new_[69240]_  = A200 & ~A199;
  assign \new_[69243]_  = A203 & A201;
  assign \new_[69244]_  = \new_[69243]_  & \new_[69240]_ ;
  assign \new_[69245]_  = \new_[69244]_  & \new_[69237]_ ;
  assign \new_[69249]_  = ~A269 & ~A268;
  assign \new_[69250]_  = A267 & \new_[69249]_ ;
  assign \new_[69253]_  = A299 & ~A298;
  assign \new_[69256]_  = A301 & A300;
  assign \new_[69257]_  = \new_[69256]_  & \new_[69253]_ ;
  assign \new_[69258]_  = \new_[69257]_  & \new_[69250]_ ;
  assign \new_[69262]_  = A168 & ~A169;
  assign \new_[69263]_  = A170 & \new_[69262]_ ;
  assign \new_[69266]_  = A200 & ~A199;
  assign \new_[69269]_  = A203 & A201;
  assign \new_[69270]_  = \new_[69269]_  & \new_[69266]_ ;
  assign \new_[69271]_  = \new_[69270]_  & \new_[69263]_ ;
  assign \new_[69275]_  = ~A269 & ~A268;
  assign \new_[69276]_  = A267 & \new_[69275]_ ;
  assign \new_[69279]_  = A299 & ~A298;
  assign \new_[69282]_  = A302 & A300;
  assign \new_[69283]_  = \new_[69282]_  & \new_[69279]_ ;
  assign \new_[69284]_  = \new_[69283]_  & \new_[69276]_ ;
  assign \new_[69288]_  = A168 & ~A169;
  assign \new_[69289]_  = A170 & \new_[69288]_ ;
  assign \new_[69292]_  = A200 & ~A199;
  assign \new_[69295]_  = A203 & A201;
  assign \new_[69296]_  = \new_[69295]_  & \new_[69292]_ ;
  assign \new_[69297]_  = \new_[69296]_  & \new_[69289]_ ;
  assign \new_[69301]_  = A298 & A268;
  assign \new_[69302]_  = ~A267 & \new_[69301]_ ;
  assign \new_[69305]_  = ~A300 & ~A299;
  assign \new_[69308]_  = ~A302 & ~A301;
  assign \new_[69309]_  = \new_[69308]_  & \new_[69305]_ ;
  assign \new_[69310]_  = \new_[69309]_  & \new_[69302]_ ;
  assign \new_[69314]_  = A168 & ~A169;
  assign \new_[69315]_  = A170 & \new_[69314]_ ;
  assign \new_[69318]_  = A200 & ~A199;
  assign \new_[69321]_  = A203 & A201;
  assign \new_[69322]_  = \new_[69321]_  & \new_[69318]_ ;
  assign \new_[69323]_  = \new_[69322]_  & \new_[69315]_ ;
  assign \new_[69327]_  = ~A298 & A268;
  assign \new_[69328]_  = ~A267 & \new_[69327]_ ;
  assign \new_[69331]_  = ~A300 & A299;
  assign \new_[69334]_  = ~A302 & ~A301;
  assign \new_[69335]_  = \new_[69334]_  & \new_[69331]_ ;
  assign \new_[69336]_  = \new_[69335]_  & \new_[69328]_ ;
  assign \new_[69340]_  = A168 & ~A169;
  assign \new_[69341]_  = A170 & \new_[69340]_ ;
  assign \new_[69344]_  = A200 & ~A199;
  assign \new_[69347]_  = A203 & A201;
  assign \new_[69348]_  = \new_[69347]_  & \new_[69344]_ ;
  assign \new_[69349]_  = \new_[69348]_  & \new_[69341]_ ;
  assign \new_[69353]_  = A298 & A269;
  assign \new_[69354]_  = ~A267 & \new_[69353]_ ;
  assign \new_[69357]_  = ~A300 & ~A299;
  assign \new_[69360]_  = ~A302 & ~A301;
  assign \new_[69361]_  = \new_[69360]_  & \new_[69357]_ ;
  assign \new_[69362]_  = \new_[69361]_  & \new_[69354]_ ;
  assign \new_[69366]_  = A168 & ~A169;
  assign \new_[69367]_  = A170 & \new_[69366]_ ;
  assign \new_[69370]_  = A200 & ~A199;
  assign \new_[69373]_  = A203 & A201;
  assign \new_[69374]_  = \new_[69373]_  & \new_[69370]_ ;
  assign \new_[69375]_  = \new_[69374]_  & \new_[69367]_ ;
  assign \new_[69379]_  = ~A298 & A269;
  assign \new_[69380]_  = ~A267 & \new_[69379]_ ;
  assign \new_[69383]_  = ~A300 & A299;
  assign \new_[69386]_  = ~A302 & ~A301;
  assign \new_[69387]_  = \new_[69386]_  & \new_[69383]_ ;
  assign \new_[69388]_  = \new_[69387]_  & \new_[69380]_ ;
  assign \new_[69392]_  = A168 & ~A169;
  assign \new_[69393]_  = A170 & \new_[69392]_ ;
  assign \new_[69396]_  = A200 & ~A199;
  assign \new_[69399]_  = A203 & A201;
  assign \new_[69400]_  = \new_[69399]_  & \new_[69396]_ ;
  assign \new_[69401]_  = \new_[69400]_  & \new_[69393]_ ;
  assign \new_[69405]_  = A298 & A266;
  assign \new_[69406]_  = A265 & \new_[69405]_ ;
  assign \new_[69409]_  = ~A300 & ~A299;
  assign \new_[69412]_  = ~A302 & ~A301;
  assign \new_[69413]_  = \new_[69412]_  & \new_[69409]_ ;
  assign \new_[69414]_  = \new_[69413]_  & \new_[69406]_ ;
  assign \new_[69418]_  = A168 & ~A169;
  assign \new_[69419]_  = A170 & \new_[69418]_ ;
  assign \new_[69422]_  = A200 & ~A199;
  assign \new_[69425]_  = A203 & A201;
  assign \new_[69426]_  = \new_[69425]_  & \new_[69422]_ ;
  assign \new_[69427]_  = \new_[69426]_  & \new_[69419]_ ;
  assign \new_[69431]_  = ~A298 & A266;
  assign \new_[69432]_  = A265 & \new_[69431]_ ;
  assign \new_[69435]_  = ~A300 & A299;
  assign \new_[69438]_  = ~A302 & ~A301;
  assign \new_[69439]_  = \new_[69438]_  & \new_[69435]_ ;
  assign \new_[69440]_  = \new_[69439]_  & \new_[69432]_ ;
  assign \new_[69444]_  = A168 & ~A169;
  assign \new_[69445]_  = A170 & \new_[69444]_ ;
  assign \new_[69448]_  = A200 & ~A199;
  assign \new_[69451]_  = A203 & A201;
  assign \new_[69452]_  = \new_[69451]_  & \new_[69448]_ ;
  assign \new_[69453]_  = \new_[69452]_  & \new_[69445]_ ;
  assign \new_[69457]_  = A298 & ~A266;
  assign \new_[69458]_  = ~A265 & \new_[69457]_ ;
  assign \new_[69461]_  = ~A300 & ~A299;
  assign \new_[69464]_  = ~A302 & ~A301;
  assign \new_[69465]_  = \new_[69464]_  & \new_[69461]_ ;
  assign \new_[69466]_  = \new_[69465]_  & \new_[69458]_ ;
  assign \new_[69470]_  = A168 & ~A169;
  assign \new_[69471]_  = A170 & \new_[69470]_ ;
  assign \new_[69474]_  = A200 & ~A199;
  assign \new_[69477]_  = A203 & A201;
  assign \new_[69478]_  = \new_[69477]_  & \new_[69474]_ ;
  assign \new_[69479]_  = \new_[69478]_  & \new_[69471]_ ;
  assign \new_[69483]_  = ~A298 & ~A266;
  assign \new_[69484]_  = ~A265 & \new_[69483]_ ;
  assign \new_[69487]_  = ~A300 & A299;
  assign \new_[69490]_  = ~A302 & ~A301;
  assign \new_[69491]_  = \new_[69490]_  & \new_[69487]_ ;
  assign \new_[69492]_  = \new_[69491]_  & \new_[69484]_ ;
  assign \new_[69496]_  = A168 & ~A169;
  assign \new_[69497]_  = A170 & \new_[69496]_ ;
  assign \new_[69500]_  = A200 & ~A199;
  assign \new_[69503]_  = ~A202 & ~A201;
  assign \new_[69504]_  = \new_[69503]_  & \new_[69500]_ ;
  assign \new_[69505]_  = \new_[69504]_  & \new_[69497]_ ;
  assign \new_[69509]_  = A268 & ~A267;
  assign \new_[69510]_  = ~A203 & \new_[69509]_ ;
  assign \new_[69513]_  = ~A299 & A298;
  assign \new_[69516]_  = A301 & A300;
  assign \new_[69517]_  = \new_[69516]_  & \new_[69513]_ ;
  assign \new_[69518]_  = \new_[69517]_  & \new_[69510]_ ;
  assign \new_[69522]_  = A168 & ~A169;
  assign \new_[69523]_  = A170 & \new_[69522]_ ;
  assign \new_[69526]_  = A200 & ~A199;
  assign \new_[69529]_  = ~A202 & ~A201;
  assign \new_[69530]_  = \new_[69529]_  & \new_[69526]_ ;
  assign \new_[69531]_  = \new_[69530]_  & \new_[69523]_ ;
  assign \new_[69535]_  = A268 & ~A267;
  assign \new_[69536]_  = ~A203 & \new_[69535]_ ;
  assign \new_[69539]_  = ~A299 & A298;
  assign \new_[69542]_  = A302 & A300;
  assign \new_[69543]_  = \new_[69542]_  & \new_[69539]_ ;
  assign \new_[69544]_  = \new_[69543]_  & \new_[69536]_ ;
  assign \new_[69548]_  = A168 & ~A169;
  assign \new_[69549]_  = A170 & \new_[69548]_ ;
  assign \new_[69552]_  = A200 & ~A199;
  assign \new_[69555]_  = ~A202 & ~A201;
  assign \new_[69556]_  = \new_[69555]_  & \new_[69552]_ ;
  assign \new_[69557]_  = \new_[69556]_  & \new_[69549]_ ;
  assign \new_[69561]_  = A268 & ~A267;
  assign \new_[69562]_  = ~A203 & \new_[69561]_ ;
  assign \new_[69565]_  = A299 & ~A298;
  assign \new_[69568]_  = A301 & A300;
  assign \new_[69569]_  = \new_[69568]_  & \new_[69565]_ ;
  assign \new_[69570]_  = \new_[69569]_  & \new_[69562]_ ;
  assign \new_[69574]_  = A168 & ~A169;
  assign \new_[69575]_  = A170 & \new_[69574]_ ;
  assign \new_[69578]_  = A200 & ~A199;
  assign \new_[69581]_  = ~A202 & ~A201;
  assign \new_[69582]_  = \new_[69581]_  & \new_[69578]_ ;
  assign \new_[69583]_  = \new_[69582]_  & \new_[69575]_ ;
  assign \new_[69587]_  = A268 & ~A267;
  assign \new_[69588]_  = ~A203 & \new_[69587]_ ;
  assign \new_[69591]_  = A299 & ~A298;
  assign \new_[69594]_  = A302 & A300;
  assign \new_[69595]_  = \new_[69594]_  & \new_[69591]_ ;
  assign \new_[69596]_  = \new_[69595]_  & \new_[69588]_ ;
  assign \new_[69600]_  = A168 & ~A169;
  assign \new_[69601]_  = A170 & \new_[69600]_ ;
  assign \new_[69604]_  = A200 & ~A199;
  assign \new_[69607]_  = ~A202 & ~A201;
  assign \new_[69608]_  = \new_[69607]_  & \new_[69604]_ ;
  assign \new_[69609]_  = \new_[69608]_  & \new_[69601]_ ;
  assign \new_[69613]_  = A269 & ~A267;
  assign \new_[69614]_  = ~A203 & \new_[69613]_ ;
  assign \new_[69617]_  = ~A299 & A298;
  assign \new_[69620]_  = A301 & A300;
  assign \new_[69621]_  = \new_[69620]_  & \new_[69617]_ ;
  assign \new_[69622]_  = \new_[69621]_  & \new_[69614]_ ;
  assign \new_[69626]_  = A168 & ~A169;
  assign \new_[69627]_  = A170 & \new_[69626]_ ;
  assign \new_[69630]_  = A200 & ~A199;
  assign \new_[69633]_  = ~A202 & ~A201;
  assign \new_[69634]_  = \new_[69633]_  & \new_[69630]_ ;
  assign \new_[69635]_  = \new_[69634]_  & \new_[69627]_ ;
  assign \new_[69639]_  = A269 & ~A267;
  assign \new_[69640]_  = ~A203 & \new_[69639]_ ;
  assign \new_[69643]_  = ~A299 & A298;
  assign \new_[69646]_  = A302 & A300;
  assign \new_[69647]_  = \new_[69646]_  & \new_[69643]_ ;
  assign \new_[69648]_  = \new_[69647]_  & \new_[69640]_ ;
  assign \new_[69652]_  = A168 & ~A169;
  assign \new_[69653]_  = A170 & \new_[69652]_ ;
  assign \new_[69656]_  = A200 & ~A199;
  assign \new_[69659]_  = ~A202 & ~A201;
  assign \new_[69660]_  = \new_[69659]_  & \new_[69656]_ ;
  assign \new_[69661]_  = \new_[69660]_  & \new_[69653]_ ;
  assign \new_[69665]_  = A269 & ~A267;
  assign \new_[69666]_  = ~A203 & \new_[69665]_ ;
  assign \new_[69669]_  = A299 & ~A298;
  assign \new_[69672]_  = A301 & A300;
  assign \new_[69673]_  = \new_[69672]_  & \new_[69669]_ ;
  assign \new_[69674]_  = \new_[69673]_  & \new_[69666]_ ;
  assign \new_[69678]_  = A168 & ~A169;
  assign \new_[69679]_  = A170 & \new_[69678]_ ;
  assign \new_[69682]_  = A200 & ~A199;
  assign \new_[69685]_  = ~A202 & ~A201;
  assign \new_[69686]_  = \new_[69685]_  & \new_[69682]_ ;
  assign \new_[69687]_  = \new_[69686]_  & \new_[69679]_ ;
  assign \new_[69691]_  = A269 & ~A267;
  assign \new_[69692]_  = ~A203 & \new_[69691]_ ;
  assign \new_[69695]_  = A299 & ~A298;
  assign \new_[69698]_  = A302 & A300;
  assign \new_[69699]_  = \new_[69698]_  & \new_[69695]_ ;
  assign \new_[69700]_  = \new_[69699]_  & \new_[69692]_ ;
  assign \new_[69704]_  = A168 & ~A169;
  assign \new_[69705]_  = A170 & \new_[69704]_ ;
  assign \new_[69708]_  = A200 & ~A199;
  assign \new_[69711]_  = ~A202 & ~A201;
  assign \new_[69712]_  = \new_[69711]_  & \new_[69708]_ ;
  assign \new_[69713]_  = \new_[69712]_  & \new_[69705]_ ;
  assign \new_[69717]_  = A266 & A265;
  assign \new_[69718]_  = ~A203 & \new_[69717]_ ;
  assign \new_[69721]_  = ~A299 & A298;
  assign \new_[69724]_  = A301 & A300;
  assign \new_[69725]_  = \new_[69724]_  & \new_[69721]_ ;
  assign \new_[69726]_  = \new_[69725]_  & \new_[69718]_ ;
  assign \new_[69730]_  = A168 & ~A169;
  assign \new_[69731]_  = A170 & \new_[69730]_ ;
  assign \new_[69734]_  = A200 & ~A199;
  assign \new_[69737]_  = ~A202 & ~A201;
  assign \new_[69738]_  = \new_[69737]_  & \new_[69734]_ ;
  assign \new_[69739]_  = \new_[69738]_  & \new_[69731]_ ;
  assign \new_[69743]_  = A266 & A265;
  assign \new_[69744]_  = ~A203 & \new_[69743]_ ;
  assign \new_[69747]_  = ~A299 & A298;
  assign \new_[69750]_  = A302 & A300;
  assign \new_[69751]_  = \new_[69750]_  & \new_[69747]_ ;
  assign \new_[69752]_  = \new_[69751]_  & \new_[69744]_ ;
  assign \new_[69756]_  = A168 & ~A169;
  assign \new_[69757]_  = A170 & \new_[69756]_ ;
  assign \new_[69760]_  = A200 & ~A199;
  assign \new_[69763]_  = ~A202 & ~A201;
  assign \new_[69764]_  = \new_[69763]_  & \new_[69760]_ ;
  assign \new_[69765]_  = \new_[69764]_  & \new_[69757]_ ;
  assign \new_[69769]_  = A266 & A265;
  assign \new_[69770]_  = ~A203 & \new_[69769]_ ;
  assign \new_[69773]_  = A299 & ~A298;
  assign \new_[69776]_  = A301 & A300;
  assign \new_[69777]_  = \new_[69776]_  & \new_[69773]_ ;
  assign \new_[69778]_  = \new_[69777]_  & \new_[69770]_ ;
  assign \new_[69782]_  = A168 & ~A169;
  assign \new_[69783]_  = A170 & \new_[69782]_ ;
  assign \new_[69786]_  = A200 & ~A199;
  assign \new_[69789]_  = ~A202 & ~A201;
  assign \new_[69790]_  = \new_[69789]_  & \new_[69786]_ ;
  assign \new_[69791]_  = \new_[69790]_  & \new_[69783]_ ;
  assign \new_[69795]_  = A266 & A265;
  assign \new_[69796]_  = ~A203 & \new_[69795]_ ;
  assign \new_[69799]_  = A299 & ~A298;
  assign \new_[69802]_  = A302 & A300;
  assign \new_[69803]_  = \new_[69802]_  & \new_[69799]_ ;
  assign \new_[69804]_  = \new_[69803]_  & \new_[69796]_ ;
  assign \new_[69808]_  = A168 & ~A169;
  assign \new_[69809]_  = A170 & \new_[69808]_ ;
  assign \new_[69812]_  = A200 & ~A199;
  assign \new_[69815]_  = ~A202 & ~A201;
  assign \new_[69816]_  = \new_[69815]_  & \new_[69812]_ ;
  assign \new_[69817]_  = \new_[69816]_  & \new_[69809]_ ;
  assign \new_[69821]_  = ~A266 & ~A265;
  assign \new_[69822]_  = ~A203 & \new_[69821]_ ;
  assign \new_[69825]_  = ~A299 & A298;
  assign \new_[69828]_  = A301 & A300;
  assign \new_[69829]_  = \new_[69828]_  & \new_[69825]_ ;
  assign \new_[69830]_  = \new_[69829]_  & \new_[69822]_ ;
  assign \new_[69834]_  = A168 & ~A169;
  assign \new_[69835]_  = A170 & \new_[69834]_ ;
  assign \new_[69838]_  = A200 & ~A199;
  assign \new_[69841]_  = ~A202 & ~A201;
  assign \new_[69842]_  = \new_[69841]_  & \new_[69838]_ ;
  assign \new_[69843]_  = \new_[69842]_  & \new_[69835]_ ;
  assign \new_[69847]_  = ~A266 & ~A265;
  assign \new_[69848]_  = ~A203 & \new_[69847]_ ;
  assign \new_[69851]_  = ~A299 & A298;
  assign \new_[69854]_  = A302 & A300;
  assign \new_[69855]_  = \new_[69854]_  & \new_[69851]_ ;
  assign \new_[69856]_  = \new_[69855]_  & \new_[69848]_ ;
  assign \new_[69860]_  = A168 & ~A169;
  assign \new_[69861]_  = A170 & \new_[69860]_ ;
  assign \new_[69864]_  = A200 & ~A199;
  assign \new_[69867]_  = ~A202 & ~A201;
  assign \new_[69868]_  = \new_[69867]_  & \new_[69864]_ ;
  assign \new_[69869]_  = \new_[69868]_  & \new_[69861]_ ;
  assign \new_[69873]_  = ~A266 & ~A265;
  assign \new_[69874]_  = ~A203 & \new_[69873]_ ;
  assign \new_[69877]_  = A299 & ~A298;
  assign \new_[69880]_  = A301 & A300;
  assign \new_[69881]_  = \new_[69880]_  & \new_[69877]_ ;
  assign \new_[69882]_  = \new_[69881]_  & \new_[69874]_ ;
  assign \new_[69886]_  = A168 & ~A169;
  assign \new_[69887]_  = A170 & \new_[69886]_ ;
  assign \new_[69890]_  = A200 & ~A199;
  assign \new_[69893]_  = ~A202 & ~A201;
  assign \new_[69894]_  = \new_[69893]_  & \new_[69890]_ ;
  assign \new_[69895]_  = \new_[69894]_  & \new_[69887]_ ;
  assign \new_[69899]_  = ~A266 & ~A265;
  assign \new_[69900]_  = ~A203 & \new_[69899]_ ;
  assign \new_[69903]_  = A299 & ~A298;
  assign \new_[69906]_  = A302 & A300;
  assign \new_[69907]_  = \new_[69906]_  & \new_[69903]_ ;
  assign \new_[69908]_  = \new_[69907]_  & \new_[69900]_ ;
  assign \new_[69912]_  = A168 & ~A169;
  assign \new_[69913]_  = A170 & \new_[69912]_ ;
  assign \new_[69916]_  = ~A200 & A199;
  assign \new_[69919]_  = A202 & A201;
  assign \new_[69920]_  = \new_[69919]_  & \new_[69916]_ ;
  assign \new_[69921]_  = \new_[69920]_  & \new_[69913]_ ;
  assign \new_[69925]_  = ~A269 & ~A268;
  assign \new_[69926]_  = A267 & \new_[69925]_ ;
  assign \new_[69929]_  = ~A299 & A298;
  assign \new_[69932]_  = A301 & A300;
  assign \new_[69933]_  = \new_[69932]_  & \new_[69929]_ ;
  assign \new_[69934]_  = \new_[69933]_  & \new_[69926]_ ;
  assign \new_[69938]_  = A168 & ~A169;
  assign \new_[69939]_  = A170 & \new_[69938]_ ;
  assign \new_[69942]_  = ~A200 & A199;
  assign \new_[69945]_  = A202 & A201;
  assign \new_[69946]_  = \new_[69945]_  & \new_[69942]_ ;
  assign \new_[69947]_  = \new_[69946]_  & \new_[69939]_ ;
  assign \new_[69951]_  = ~A269 & ~A268;
  assign \new_[69952]_  = A267 & \new_[69951]_ ;
  assign \new_[69955]_  = ~A299 & A298;
  assign \new_[69958]_  = A302 & A300;
  assign \new_[69959]_  = \new_[69958]_  & \new_[69955]_ ;
  assign \new_[69960]_  = \new_[69959]_  & \new_[69952]_ ;
  assign \new_[69964]_  = A168 & ~A169;
  assign \new_[69965]_  = A170 & \new_[69964]_ ;
  assign \new_[69968]_  = ~A200 & A199;
  assign \new_[69971]_  = A202 & A201;
  assign \new_[69972]_  = \new_[69971]_  & \new_[69968]_ ;
  assign \new_[69973]_  = \new_[69972]_  & \new_[69965]_ ;
  assign \new_[69977]_  = ~A269 & ~A268;
  assign \new_[69978]_  = A267 & \new_[69977]_ ;
  assign \new_[69981]_  = A299 & ~A298;
  assign \new_[69984]_  = A301 & A300;
  assign \new_[69985]_  = \new_[69984]_  & \new_[69981]_ ;
  assign \new_[69986]_  = \new_[69985]_  & \new_[69978]_ ;
  assign \new_[69990]_  = A168 & ~A169;
  assign \new_[69991]_  = A170 & \new_[69990]_ ;
  assign \new_[69994]_  = ~A200 & A199;
  assign \new_[69997]_  = A202 & A201;
  assign \new_[69998]_  = \new_[69997]_  & \new_[69994]_ ;
  assign \new_[69999]_  = \new_[69998]_  & \new_[69991]_ ;
  assign \new_[70003]_  = ~A269 & ~A268;
  assign \new_[70004]_  = A267 & \new_[70003]_ ;
  assign \new_[70007]_  = A299 & ~A298;
  assign \new_[70010]_  = A302 & A300;
  assign \new_[70011]_  = \new_[70010]_  & \new_[70007]_ ;
  assign \new_[70012]_  = \new_[70011]_  & \new_[70004]_ ;
  assign \new_[70016]_  = A168 & ~A169;
  assign \new_[70017]_  = A170 & \new_[70016]_ ;
  assign \new_[70020]_  = ~A200 & A199;
  assign \new_[70023]_  = A202 & A201;
  assign \new_[70024]_  = \new_[70023]_  & \new_[70020]_ ;
  assign \new_[70025]_  = \new_[70024]_  & \new_[70017]_ ;
  assign \new_[70029]_  = A298 & A268;
  assign \new_[70030]_  = ~A267 & \new_[70029]_ ;
  assign \new_[70033]_  = ~A300 & ~A299;
  assign \new_[70036]_  = ~A302 & ~A301;
  assign \new_[70037]_  = \new_[70036]_  & \new_[70033]_ ;
  assign \new_[70038]_  = \new_[70037]_  & \new_[70030]_ ;
  assign \new_[70042]_  = A168 & ~A169;
  assign \new_[70043]_  = A170 & \new_[70042]_ ;
  assign \new_[70046]_  = ~A200 & A199;
  assign \new_[70049]_  = A202 & A201;
  assign \new_[70050]_  = \new_[70049]_  & \new_[70046]_ ;
  assign \new_[70051]_  = \new_[70050]_  & \new_[70043]_ ;
  assign \new_[70055]_  = ~A298 & A268;
  assign \new_[70056]_  = ~A267 & \new_[70055]_ ;
  assign \new_[70059]_  = ~A300 & A299;
  assign \new_[70062]_  = ~A302 & ~A301;
  assign \new_[70063]_  = \new_[70062]_  & \new_[70059]_ ;
  assign \new_[70064]_  = \new_[70063]_  & \new_[70056]_ ;
  assign \new_[70068]_  = A168 & ~A169;
  assign \new_[70069]_  = A170 & \new_[70068]_ ;
  assign \new_[70072]_  = ~A200 & A199;
  assign \new_[70075]_  = A202 & A201;
  assign \new_[70076]_  = \new_[70075]_  & \new_[70072]_ ;
  assign \new_[70077]_  = \new_[70076]_  & \new_[70069]_ ;
  assign \new_[70081]_  = A298 & A269;
  assign \new_[70082]_  = ~A267 & \new_[70081]_ ;
  assign \new_[70085]_  = ~A300 & ~A299;
  assign \new_[70088]_  = ~A302 & ~A301;
  assign \new_[70089]_  = \new_[70088]_  & \new_[70085]_ ;
  assign \new_[70090]_  = \new_[70089]_  & \new_[70082]_ ;
  assign \new_[70094]_  = A168 & ~A169;
  assign \new_[70095]_  = A170 & \new_[70094]_ ;
  assign \new_[70098]_  = ~A200 & A199;
  assign \new_[70101]_  = A202 & A201;
  assign \new_[70102]_  = \new_[70101]_  & \new_[70098]_ ;
  assign \new_[70103]_  = \new_[70102]_  & \new_[70095]_ ;
  assign \new_[70107]_  = ~A298 & A269;
  assign \new_[70108]_  = ~A267 & \new_[70107]_ ;
  assign \new_[70111]_  = ~A300 & A299;
  assign \new_[70114]_  = ~A302 & ~A301;
  assign \new_[70115]_  = \new_[70114]_  & \new_[70111]_ ;
  assign \new_[70116]_  = \new_[70115]_  & \new_[70108]_ ;
  assign \new_[70120]_  = A168 & ~A169;
  assign \new_[70121]_  = A170 & \new_[70120]_ ;
  assign \new_[70124]_  = ~A200 & A199;
  assign \new_[70127]_  = A202 & A201;
  assign \new_[70128]_  = \new_[70127]_  & \new_[70124]_ ;
  assign \new_[70129]_  = \new_[70128]_  & \new_[70121]_ ;
  assign \new_[70133]_  = A298 & A266;
  assign \new_[70134]_  = A265 & \new_[70133]_ ;
  assign \new_[70137]_  = ~A300 & ~A299;
  assign \new_[70140]_  = ~A302 & ~A301;
  assign \new_[70141]_  = \new_[70140]_  & \new_[70137]_ ;
  assign \new_[70142]_  = \new_[70141]_  & \new_[70134]_ ;
  assign \new_[70146]_  = A168 & ~A169;
  assign \new_[70147]_  = A170 & \new_[70146]_ ;
  assign \new_[70150]_  = ~A200 & A199;
  assign \new_[70153]_  = A202 & A201;
  assign \new_[70154]_  = \new_[70153]_  & \new_[70150]_ ;
  assign \new_[70155]_  = \new_[70154]_  & \new_[70147]_ ;
  assign \new_[70159]_  = ~A298 & A266;
  assign \new_[70160]_  = A265 & \new_[70159]_ ;
  assign \new_[70163]_  = ~A300 & A299;
  assign \new_[70166]_  = ~A302 & ~A301;
  assign \new_[70167]_  = \new_[70166]_  & \new_[70163]_ ;
  assign \new_[70168]_  = \new_[70167]_  & \new_[70160]_ ;
  assign \new_[70172]_  = A168 & ~A169;
  assign \new_[70173]_  = A170 & \new_[70172]_ ;
  assign \new_[70176]_  = ~A200 & A199;
  assign \new_[70179]_  = A202 & A201;
  assign \new_[70180]_  = \new_[70179]_  & \new_[70176]_ ;
  assign \new_[70181]_  = \new_[70180]_  & \new_[70173]_ ;
  assign \new_[70185]_  = A298 & ~A266;
  assign \new_[70186]_  = ~A265 & \new_[70185]_ ;
  assign \new_[70189]_  = ~A300 & ~A299;
  assign \new_[70192]_  = ~A302 & ~A301;
  assign \new_[70193]_  = \new_[70192]_  & \new_[70189]_ ;
  assign \new_[70194]_  = \new_[70193]_  & \new_[70186]_ ;
  assign \new_[70198]_  = A168 & ~A169;
  assign \new_[70199]_  = A170 & \new_[70198]_ ;
  assign \new_[70202]_  = ~A200 & A199;
  assign \new_[70205]_  = A202 & A201;
  assign \new_[70206]_  = \new_[70205]_  & \new_[70202]_ ;
  assign \new_[70207]_  = \new_[70206]_  & \new_[70199]_ ;
  assign \new_[70211]_  = ~A298 & ~A266;
  assign \new_[70212]_  = ~A265 & \new_[70211]_ ;
  assign \new_[70215]_  = ~A300 & A299;
  assign \new_[70218]_  = ~A302 & ~A301;
  assign \new_[70219]_  = \new_[70218]_  & \new_[70215]_ ;
  assign \new_[70220]_  = \new_[70219]_  & \new_[70212]_ ;
  assign \new_[70224]_  = A168 & ~A169;
  assign \new_[70225]_  = A170 & \new_[70224]_ ;
  assign \new_[70228]_  = ~A200 & A199;
  assign \new_[70231]_  = A203 & A201;
  assign \new_[70232]_  = \new_[70231]_  & \new_[70228]_ ;
  assign \new_[70233]_  = \new_[70232]_  & \new_[70225]_ ;
  assign \new_[70237]_  = ~A269 & ~A268;
  assign \new_[70238]_  = A267 & \new_[70237]_ ;
  assign \new_[70241]_  = ~A299 & A298;
  assign \new_[70244]_  = A301 & A300;
  assign \new_[70245]_  = \new_[70244]_  & \new_[70241]_ ;
  assign \new_[70246]_  = \new_[70245]_  & \new_[70238]_ ;
  assign \new_[70250]_  = A168 & ~A169;
  assign \new_[70251]_  = A170 & \new_[70250]_ ;
  assign \new_[70254]_  = ~A200 & A199;
  assign \new_[70257]_  = A203 & A201;
  assign \new_[70258]_  = \new_[70257]_  & \new_[70254]_ ;
  assign \new_[70259]_  = \new_[70258]_  & \new_[70251]_ ;
  assign \new_[70263]_  = ~A269 & ~A268;
  assign \new_[70264]_  = A267 & \new_[70263]_ ;
  assign \new_[70267]_  = ~A299 & A298;
  assign \new_[70270]_  = A302 & A300;
  assign \new_[70271]_  = \new_[70270]_  & \new_[70267]_ ;
  assign \new_[70272]_  = \new_[70271]_  & \new_[70264]_ ;
  assign \new_[70276]_  = A168 & ~A169;
  assign \new_[70277]_  = A170 & \new_[70276]_ ;
  assign \new_[70280]_  = ~A200 & A199;
  assign \new_[70283]_  = A203 & A201;
  assign \new_[70284]_  = \new_[70283]_  & \new_[70280]_ ;
  assign \new_[70285]_  = \new_[70284]_  & \new_[70277]_ ;
  assign \new_[70289]_  = ~A269 & ~A268;
  assign \new_[70290]_  = A267 & \new_[70289]_ ;
  assign \new_[70293]_  = A299 & ~A298;
  assign \new_[70296]_  = A301 & A300;
  assign \new_[70297]_  = \new_[70296]_  & \new_[70293]_ ;
  assign \new_[70298]_  = \new_[70297]_  & \new_[70290]_ ;
  assign \new_[70302]_  = A168 & ~A169;
  assign \new_[70303]_  = A170 & \new_[70302]_ ;
  assign \new_[70306]_  = ~A200 & A199;
  assign \new_[70309]_  = A203 & A201;
  assign \new_[70310]_  = \new_[70309]_  & \new_[70306]_ ;
  assign \new_[70311]_  = \new_[70310]_  & \new_[70303]_ ;
  assign \new_[70315]_  = ~A269 & ~A268;
  assign \new_[70316]_  = A267 & \new_[70315]_ ;
  assign \new_[70319]_  = A299 & ~A298;
  assign \new_[70322]_  = A302 & A300;
  assign \new_[70323]_  = \new_[70322]_  & \new_[70319]_ ;
  assign \new_[70324]_  = \new_[70323]_  & \new_[70316]_ ;
  assign \new_[70328]_  = A168 & ~A169;
  assign \new_[70329]_  = A170 & \new_[70328]_ ;
  assign \new_[70332]_  = ~A200 & A199;
  assign \new_[70335]_  = A203 & A201;
  assign \new_[70336]_  = \new_[70335]_  & \new_[70332]_ ;
  assign \new_[70337]_  = \new_[70336]_  & \new_[70329]_ ;
  assign \new_[70341]_  = A298 & A268;
  assign \new_[70342]_  = ~A267 & \new_[70341]_ ;
  assign \new_[70345]_  = ~A300 & ~A299;
  assign \new_[70348]_  = ~A302 & ~A301;
  assign \new_[70349]_  = \new_[70348]_  & \new_[70345]_ ;
  assign \new_[70350]_  = \new_[70349]_  & \new_[70342]_ ;
  assign \new_[70354]_  = A168 & ~A169;
  assign \new_[70355]_  = A170 & \new_[70354]_ ;
  assign \new_[70358]_  = ~A200 & A199;
  assign \new_[70361]_  = A203 & A201;
  assign \new_[70362]_  = \new_[70361]_  & \new_[70358]_ ;
  assign \new_[70363]_  = \new_[70362]_  & \new_[70355]_ ;
  assign \new_[70367]_  = ~A298 & A268;
  assign \new_[70368]_  = ~A267 & \new_[70367]_ ;
  assign \new_[70371]_  = ~A300 & A299;
  assign \new_[70374]_  = ~A302 & ~A301;
  assign \new_[70375]_  = \new_[70374]_  & \new_[70371]_ ;
  assign \new_[70376]_  = \new_[70375]_  & \new_[70368]_ ;
  assign \new_[70380]_  = A168 & ~A169;
  assign \new_[70381]_  = A170 & \new_[70380]_ ;
  assign \new_[70384]_  = ~A200 & A199;
  assign \new_[70387]_  = A203 & A201;
  assign \new_[70388]_  = \new_[70387]_  & \new_[70384]_ ;
  assign \new_[70389]_  = \new_[70388]_  & \new_[70381]_ ;
  assign \new_[70393]_  = A298 & A269;
  assign \new_[70394]_  = ~A267 & \new_[70393]_ ;
  assign \new_[70397]_  = ~A300 & ~A299;
  assign \new_[70400]_  = ~A302 & ~A301;
  assign \new_[70401]_  = \new_[70400]_  & \new_[70397]_ ;
  assign \new_[70402]_  = \new_[70401]_  & \new_[70394]_ ;
  assign \new_[70406]_  = A168 & ~A169;
  assign \new_[70407]_  = A170 & \new_[70406]_ ;
  assign \new_[70410]_  = ~A200 & A199;
  assign \new_[70413]_  = A203 & A201;
  assign \new_[70414]_  = \new_[70413]_  & \new_[70410]_ ;
  assign \new_[70415]_  = \new_[70414]_  & \new_[70407]_ ;
  assign \new_[70419]_  = ~A298 & A269;
  assign \new_[70420]_  = ~A267 & \new_[70419]_ ;
  assign \new_[70423]_  = ~A300 & A299;
  assign \new_[70426]_  = ~A302 & ~A301;
  assign \new_[70427]_  = \new_[70426]_  & \new_[70423]_ ;
  assign \new_[70428]_  = \new_[70427]_  & \new_[70420]_ ;
  assign \new_[70432]_  = A168 & ~A169;
  assign \new_[70433]_  = A170 & \new_[70432]_ ;
  assign \new_[70436]_  = ~A200 & A199;
  assign \new_[70439]_  = A203 & A201;
  assign \new_[70440]_  = \new_[70439]_  & \new_[70436]_ ;
  assign \new_[70441]_  = \new_[70440]_  & \new_[70433]_ ;
  assign \new_[70445]_  = A298 & A266;
  assign \new_[70446]_  = A265 & \new_[70445]_ ;
  assign \new_[70449]_  = ~A300 & ~A299;
  assign \new_[70452]_  = ~A302 & ~A301;
  assign \new_[70453]_  = \new_[70452]_  & \new_[70449]_ ;
  assign \new_[70454]_  = \new_[70453]_  & \new_[70446]_ ;
  assign \new_[70458]_  = A168 & ~A169;
  assign \new_[70459]_  = A170 & \new_[70458]_ ;
  assign \new_[70462]_  = ~A200 & A199;
  assign \new_[70465]_  = A203 & A201;
  assign \new_[70466]_  = \new_[70465]_  & \new_[70462]_ ;
  assign \new_[70467]_  = \new_[70466]_  & \new_[70459]_ ;
  assign \new_[70471]_  = ~A298 & A266;
  assign \new_[70472]_  = A265 & \new_[70471]_ ;
  assign \new_[70475]_  = ~A300 & A299;
  assign \new_[70478]_  = ~A302 & ~A301;
  assign \new_[70479]_  = \new_[70478]_  & \new_[70475]_ ;
  assign \new_[70480]_  = \new_[70479]_  & \new_[70472]_ ;
  assign \new_[70484]_  = A168 & ~A169;
  assign \new_[70485]_  = A170 & \new_[70484]_ ;
  assign \new_[70488]_  = ~A200 & A199;
  assign \new_[70491]_  = A203 & A201;
  assign \new_[70492]_  = \new_[70491]_  & \new_[70488]_ ;
  assign \new_[70493]_  = \new_[70492]_  & \new_[70485]_ ;
  assign \new_[70497]_  = A298 & ~A266;
  assign \new_[70498]_  = ~A265 & \new_[70497]_ ;
  assign \new_[70501]_  = ~A300 & ~A299;
  assign \new_[70504]_  = ~A302 & ~A301;
  assign \new_[70505]_  = \new_[70504]_  & \new_[70501]_ ;
  assign \new_[70506]_  = \new_[70505]_  & \new_[70498]_ ;
  assign \new_[70510]_  = A168 & ~A169;
  assign \new_[70511]_  = A170 & \new_[70510]_ ;
  assign \new_[70514]_  = ~A200 & A199;
  assign \new_[70517]_  = A203 & A201;
  assign \new_[70518]_  = \new_[70517]_  & \new_[70514]_ ;
  assign \new_[70519]_  = \new_[70518]_  & \new_[70511]_ ;
  assign \new_[70523]_  = ~A298 & ~A266;
  assign \new_[70524]_  = ~A265 & \new_[70523]_ ;
  assign \new_[70527]_  = ~A300 & A299;
  assign \new_[70530]_  = ~A302 & ~A301;
  assign \new_[70531]_  = \new_[70530]_  & \new_[70527]_ ;
  assign \new_[70532]_  = \new_[70531]_  & \new_[70524]_ ;
  assign \new_[70536]_  = A168 & ~A169;
  assign \new_[70537]_  = A170 & \new_[70536]_ ;
  assign \new_[70540]_  = ~A200 & A199;
  assign \new_[70543]_  = ~A202 & ~A201;
  assign \new_[70544]_  = \new_[70543]_  & \new_[70540]_ ;
  assign \new_[70545]_  = \new_[70544]_  & \new_[70537]_ ;
  assign \new_[70549]_  = A268 & ~A267;
  assign \new_[70550]_  = ~A203 & \new_[70549]_ ;
  assign \new_[70553]_  = ~A299 & A298;
  assign \new_[70556]_  = A301 & A300;
  assign \new_[70557]_  = \new_[70556]_  & \new_[70553]_ ;
  assign \new_[70558]_  = \new_[70557]_  & \new_[70550]_ ;
  assign \new_[70562]_  = A168 & ~A169;
  assign \new_[70563]_  = A170 & \new_[70562]_ ;
  assign \new_[70566]_  = ~A200 & A199;
  assign \new_[70569]_  = ~A202 & ~A201;
  assign \new_[70570]_  = \new_[70569]_  & \new_[70566]_ ;
  assign \new_[70571]_  = \new_[70570]_  & \new_[70563]_ ;
  assign \new_[70575]_  = A268 & ~A267;
  assign \new_[70576]_  = ~A203 & \new_[70575]_ ;
  assign \new_[70579]_  = ~A299 & A298;
  assign \new_[70582]_  = A302 & A300;
  assign \new_[70583]_  = \new_[70582]_  & \new_[70579]_ ;
  assign \new_[70584]_  = \new_[70583]_  & \new_[70576]_ ;
  assign \new_[70588]_  = A168 & ~A169;
  assign \new_[70589]_  = A170 & \new_[70588]_ ;
  assign \new_[70592]_  = ~A200 & A199;
  assign \new_[70595]_  = ~A202 & ~A201;
  assign \new_[70596]_  = \new_[70595]_  & \new_[70592]_ ;
  assign \new_[70597]_  = \new_[70596]_  & \new_[70589]_ ;
  assign \new_[70601]_  = A268 & ~A267;
  assign \new_[70602]_  = ~A203 & \new_[70601]_ ;
  assign \new_[70605]_  = A299 & ~A298;
  assign \new_[70608]_  = A301 & A300;
  assign \new_[70609]_  = \new_[70608]_  & \new_[70605]_ ;
  assign \new_[70610]_  = \new_[70609]_  & \new_[70602]_ ;
  assign \new_[70614]_  = A168 & ~A169;
  assign \new_[70615]_  = A170 & \new_[70614]_ ;
  assign \new_[70618]_  = ~A200 & A199;
  assign \new_[70621]_  = ~A202 & ~A201;
  assign \new_[70622]_  = \new_[70621]_  & \new_[70618]_ ;
  assign \new_[70623]_  = \new_[70622]_  & \new_[70615]_ ;
  assign \new_[70627]_  = A268 & ~A267;
  assign \new_[70628]_  = ~A203 & \new_[70627]_ ;
  assign \new_[70631]_  = A299 & ~A298;
  assign \new_[70634]_  = A302 & A300;
  assign \new_[70635]_  = \new_[70634]_  & \new_[70631]_ ;
  assign \new_[70636]_  = \new_[70635]_  & \new_[70628]_ ;
  assign \new_[70640]_  = A168 & ~A169;
  assign \new_[70641]_  = A170 & \new_[70640]_ ;
  assign \new_[70644]_  = ~A200 & A199;
  assign \new_[70647]_  = ~A202 & ~A201;
  assign \new_[70648]_  = \new_[70647]_  & \new_[70644]_ ;
  assign \new_[70649]_  = \new_[70648]_  & \new_[70641]_ ;
  assign \new_[70653]_  = A269 & ~A267;
  assign \new_[70654]_  = ~A203 & \new_[70653]_ ;
  assign \new_[70657]_  = ~A299 & A298;
  assign \new_[70660]_  = A301 & A300;
  assign \new_[70661]_  = \new_[70660]_  & \new_[70657]_ ;
  assign \new_[70662]_  = \new_[70661]_  & \new_[70654]_ ;
  assign \new_[70666]_  = A168 & ~A169;
  assign \new_[70667]_  = A170 & \new_[70666]_ ;
  assign \new_[70670]_  = ~A200 & A199;
  assign \new_[70673]_  = ~A202 & ~A201;
  assign \new_[70674]_  = \new_[70673]_  & \new_[70670]_ ;
  assign \new_[70675]_  = \new_[70674]_  & \new_[70667]_ ;
  assign \new_[70679]_  = A269 & ~A267;
  assign \new_[70680]_  = ~A203 & \new_[70679]_ ;
  assign \new_[70683]_  = ~A299 & A298;
  assign \new_[70686]_  = A302 & A300;
  assign \new_[70687]_  = \new_[70686]_  & \new_[70683]_ ;
  assign \new_[70688]_  = \new_[70687]_  & \new_[70680]_ ;
  assign \new_[70692]_  = A168 & ~A169;
  assign \new_[70693]_  = A170 & \new_[70692]_ ;
  assign \new_[70696]_  = ~A200 & A199;
  assign \new_[70699]_  = ~A202 & ~A201;
  assign \new_[70700]_  = \new_[70699]_  & \new_[70696]_ ;
  assign \new_[70701]_  = \new_[70700]_  & \new_[70693]_ ;
  assign \new_[70705]_  = A269 & ~A267;
  assign \new_[70706]_  = ~A203 & \new_[70705]_ ;
  assign \new_[70709]_  = A299 & ~A298;
  assign \new_[70712]_  = A301 & A300;
  assign \new_[70713]_  = \new_[70712]_  & \new_[70709]_ ;
  assign \new_[70714]_  = \new_[70713]_  & \new_[70706]_ ;
  assign \new_[70718]_  = A168 & ~A169;
  assign \new_[70719]_  = A170 & \new_[70718]_ ;
  assign \new_[70722]_  = ~A200 & A199;
  assign \new_[70725]_  = ~A202 & ~A201;
  assign \new_[70726]_  = \new_[70725]_  & \new_[70722]_ ;
  assign \new_[70727]_  = \new_[70726]_  & \new_[70719]_ ;
  assign \new_[70731]_  = A269 & ~A267;
  assign \new_[70732]_  = ~A203 & \new_[70731]_ ;
  assign \new_[70735]_  = A299 & ~A298;
  assign \new_[70738]_  = A302 & A300;
  assign \new_[70739]_  = \new_[70738]_  & \new_[70735]_ ;
  assign \new_[70740]_  = \new_[70739]_  & \new_[70732]_ ;
  assign \new_[70744]_  = A168 & ~A169;
  assign \new_[70745]_  = A170 & \new_[70744]_ ;
  assign \new_[70748]_  = ~A200 & A199;
  assign \new_[70751]_  = ~A202 & ~A201;
  assign \new_[70752]_  = \new_[70751]_  & \new_[70748]_ ;
  assign \new_[70753]_  = \new_[70752]_  & \new_[70745]_ ;
  assign \new_[70757]_  = A266 & A265;
  assign \new_[70758]_  = ~A203 & \new_[70757]_ ;
  assign \new_[70761]_  = ~A299 & A298;
  assign \new_[70764]_  = A301 & A300;
  assign \new_[70765]_  = \new_[70764]_  & \new_[70761]_ ;
  assign \new_[70766]_  = \new_[70765]_  & \new_[70758]_ ;
  assign \new_[70770]_  = A168 & ~A169;
  assign \new_[70771]_  = A170 & \new_[70770]_ ;
  assign \new_[70774]_  = ~A200 & A199;
  assign \new_[70777]_  = ~A202 & ~A201;
  assign \new_[70778]_  = \new_[70777]_  & \new_[70774]_ ;
  assign \new_[70779]_  = \new_[70778]_  & \new_[70771]_ ;
  assign \new_[70783]_  = A266 & A265;
  assign \new_[70784]_  = ~A203 & \new_[70783]_ ;
  assign \new_[70787]_  = ~A299 & A298;
  assign \new_[70790]_  = A302 & A300;
  assign \new_[70791]_  = \new_[70790]_  & \new_[70787]_ ;
  assign \new_[70792]_  = \new_[70791]_  & \new_[70784]_ ;
  assign \new_[70796]_  = A168 & ~A169;
  assign \new_[70797]_  = A170 & \new_[70796]_ ;
  assign \new_[70800]_  = ~A200 & A199;
  assign \new_[70803]_  = ~A202 & ~A201;
  assign \new_[70804]_  = \new_[70803]_  & \new_[70800]_ ;
  assign \new_[70805]_  = \new_[70804]_  & \new_[70797]_ ;
  assign \new_[70809]_  = A266 & A265;
  assign \new_[70810]_  = ~A203 & \new_[70809]_ ;
  assign \new_[70813]_  = A299 & ~A298;
  assign \new_[70816]_  = A301 & A300;
  assign \new_[70817]_  = \new_[70816]_  & \new_[70813]_ ;
  assign \new_[70818]_  = \new_[70817]_  & \new_[70810]_ ;
  assign \new_[70822]_  = A168 & ~A169;
  assign \new_[70823]_  = A170 & \new_[70822]_ ;
  assign \new_[70826]_  = ~A200 & A199;
  assign \new_[70829]_  = ~A202 & ~A201;
  assign \new_[70830]_  = \new_[70829]_  & \new_[70826]_ ;
  assign \new_[70831]_  = \new_[70830]_  & \new_[70823]_ ;
  assign \new_[70835]_  = A266 & A265;
  assign \new_[70836]_  = ~A203 & \new_[70835]_ ;
  assign \new_[70839]_  = A299 & ~A298;
  assign \new_[70842]_  = A302 & A300;
  assign \new_[70843]_  = \new_[70842]_  & \new_[70839]_ ;
  assign \new_[70844]_  = \new_[70843]_  & \new_[70836]_ ;
  assign \new_[70848]_  = A168 & ~A169;
  assign \new_[70849]_  = A170 & \new_[70848]_ ;
  assign \new_[70852]_  = ~A200 & A199;
  assign \new_[70855]_  = ~A202 & ~A201;
  assign \new_[70856]_  = \new_[70855]_  & \new_[70852]_ ;
  assign \new_[70857]_  = \new_[70856]_  & \new_[70849]_ ;
  assign \new_[70861]_  = ~A266 & ~A265;
  assign \new_[70862]_  = ~A203 & \new_[70861]_ ;
  assign \new_[70865]_  = ~A299 & A298;
  assign \new_[70868]_  = A301 & A300;
  assign \new_[70869]_  = \new_[70868]_  & \new_[70865]_ ;
  assign \new_[70870]_  = \new_[70869]_  & \new_[70862]_ ;
  assign \new_[70874]_  = A168 & ~A169;
  assign \new_[70875]_  = A170 & \new_[70874]_ ;
  assign \new_[70878]_  = ~A200 & A199;
  assign \new_[70881]_  = ~A202 & ~A201;
  assign \new_[70882]_  = \new_[70881]_  & \new_[70878]_ ;
  assign \new_[70883]_  = \new_[70882]_  & \new_[70875]_ ;
  assign \new_[70887]_  = ~A266 & ~A265;
  assign \new_[70888]_  = ~A203 & \new_[70887]_ ;
  assign \new_[70891]_  = ~A299 & A298;
  assign \new_[70894]_  = A302 & A300;
  assign \new_[70895]_  = \new_[70894]_  & \new_[70891]_ ;
  assign \new_[70896]_  = \new_[70895]_  & \new_[70888]_ ;
  assign \new_[70900]_  = A168 & ~A169;
  assign \new_[70901]_  = A170 & \new_[70900]_ ;
  assign \new_[70904]_  = ~A200 & A199;
  assign \new_[70907]_  = ~A202 & ~A201;
  assign \new_[70908]_  = \new_[70907]_  & \new_[70904]_ ;
  assign \new_[70909]_  = \new_[70908]_  & \new_[70901]_ ;
  assign \new_[70913]_  = ~A266 & ~A265;
  assign \new_[70914]_  = ~A203 & \new_[70913]_ ;
  assign \new_[70917]_  = A299 & ~A298;
  assign \new_[70920]_  = A301 & A300;
  assign \new_[70921]_  = \new_[70920]_  & \new_[70917]_ ;
  assign \new_[70922]_  = \new_[70921]_  & \new_[70914]_ ;
  assign \new_[70926]_  = A168 & ~A169;
  assign \new_[70927]_  = A170 & \new_[70926]_ ;
  assign \new_[70930]_  = ~A200 & A199;
  assign \new_[70933]_  = ~A202 & ~A201;
  assign \new_[70934]_  = \new_[70933]_  & \new_[70930]_ ;
  assign \new_[70935]_  = \new_[70934]_  & \new_[70927]_ ;
  assign \new_[70939]_  = ~A266 & ~A265;
  assign \new_[70940]_  = ~A203 & \new_[70939]_ ;
  assign \new_[70943]_  = A299 & ~A298;
  assign \new_[70946]_  = A302 & A300;
  assign \new_[70947]_  = \new_[70946]_  & \new_[70943]_ ;
  assign \new_[70948]_  = \new_[70947]_  & \new_[70940]_ ;
  assign \new_[70952]_  = ~A168 & ~A169;
  assign \new_[70953]_  = A170 & \new_[70952]_ ;
  assign \new_[70956]_  = ~A166 & A167;
  assign \new_[70959]_  = ~A202 & A201;
  assign \new_[70960]_  = \new_[70959]_  & \new_[70956]_ ;
  assign \new_[70961]_  = \new_[70960]_  & \new_[70953]_ ;
  assign \new_[70965]_  = A268 & ~A267;
  assign \new_[70966]_  = ~A203 & \new_[70965]_ ;
  assign \new_[70969]_  = ~A299 & A298;
  assign \new_[70972]_  = A301 & A300;
  assign \new_[70973]_  = \new_[70972]_  & \new_[70969]_ ;
  assign \new_[70974]_  = \new_[70973]_  & \new_[70966]_ ;
  assign \new_[70978]_  = ~A168 & ~A169;
  assign \new_[70979]_  = A170 & \new_[70978]_ ;
  assign \new_[70982]_  = ~A166 & A167;
  assign \new_[70985]_  = ~A202 & A201;
  assign \new_[70986]_  = \new_[70985]_  & \new_[70982]_ ;
  assign \new_[70987]_  = \new_[70986]_  & \new_[70979]_ ;
  assign \new_[70991]_  = A268 & ~A267;
  assign \new_[70992]_  = ~A203 & \new_[70991]_ ;
  assign \new_[70995]_  = ~A299 & A298;
  assign \new_[70998]_  = A302 & A300;
  assign \new_[70999]_  = \new_[70998]_  & \new_[70995]_ ;
  assign \new_[71000]_  = \new_[70999]_  & \new_[70992]_ ;
  assign \new_[71004]_  = ~A168 & ~A169;
  assign \new_[71005]_  = A170 & \new_[71004]_ ;
  assign \new_[71008]_  = ~A166 & A167;
  assign \new_[71011]_  = ~A202 & A201;
  assign \new_[71012]_  = \new_[71011]_  & \new_[71008]_ ;
  assign \new_[71013]_  = \new_[71012]_  & \new_[71005]_ ;
  assign \new_[71017]_  = A268 & ~A267;
  assign \new_[71018]_  = ~A203 & \new_[71017]_ ;
  assign \new_[71021]_  = A299 & ~A298;
  assign \new_[71024]_  = A301 & A300;
  assign \new_[71025]_  = \new_[71024]_  & \new_[71021]_ ;
  assign \new_[71026]_  = \new_[71025]_  & \new_[71018]_ ;
  assign \new_[71030]_  = ~A168 & ~A169;
  assign \new_[71031]_  = A170 & \new_[71030]_ ;
  assign \new_[71034]_  = ~A166 & A167;
  assign \new_[71037]_  = ~A202 & A201;
  assign \new_[71038]_  = \new_[71037]_  & \new_[71034]_ ;
  assign \new_[71039]_  = \new_[71038]_  & \new_[71031]_ ;
  assign \new_[71043]_  = A268 & ~A267;
  assign \new_[71044]_  = ~A203 & \new_[71043]_ ;
  assign \new_[71047]_  = A299 & ~A298;
  assign \new_[71050]_  = A302 & A300;
  assign \new_[71051]_  = \new_[71050]_  & \new_[71047]_ ;
  assign \new_[71052]_  = \new_[71051]_  & \new_[71044]_ ;
  assign \new_[71056]_  = ~A168 & ~A169;
  assign \new_[71057]_  = A170 & \new_[71056]_ ;
  assign \new_[71060]_  = ~A166 & A167;
  assign \new_[71063]_  = ~A202 & A201;
  assign \new_[71064]_  = \new_[71063]_  & \new_[71060]_ ;
  assign \new_[71065]_  = \new_[71064]_  & \new_[71057]_ ;
  assign \new_[71069]_  = A269 & ~A267;
  assign \new_[71070]_  = ~A203 & \new_[71069]_ ;
  assign \new_[71073]_  = ~A299 & A298;
  assign \new_[71076]_  = A301 & A300;
  assign \new_[71077]_  = \new_[71076]_  & \new_[71073]_ ;
  assign \new_[71078]_  = \new_[71077]_  & \new_[71070]_ ;
  assign \new_[71082]_  = ~A168 & ~A169;
  assign \new_[71083]_  = A170 & \new_[71082]_ ;
  assign \new_[71086]_  = ~A166 & A167;
  assign \new_[71089]_  = ~A202 & A201;
  assign \new_[71090]_  = \new_[71089]_  & \new_[71086]_ ;
  assign \new_[71091]_  = \new_[71090]_  & \new_[71083]_ ;
  assign \new_[71095]_  = A269 & ~A267;
  assign \new_[71096]_  = ~A203 & \new_[71095]_ ;
  assign \new_[71099]_  = ~A299 & A298;
  assign \new_[71102]_  = A302 & A300;
  assign \new_[71103]_  = \new_[71102]_  & \new_[71099]_ ;
  assign \new_[71104]_  = \new_[71103]_  & \new_[71096]_ ;
  assign \new_[71108]_  = ~A168 & ~A169;
  assign \new_[71109]_  = A170 & \new_[71108]_ ;
  assign \new_[71112]_  = ~A166 & A167;
  assign \new_[71115]_  = ~A202 & A201;
  assign \new_[71116]_  = \new_[71115]_  & \new_[71112]_ ;
  assign \new_[71117]_  = \new_[71116]_  & \new_[71109]_ ;
  assign \new_[71121]_  = A269 & ~A267;
  assign \new_[71122]_  = ~A203 & \new_[71121]_ ;
  assign \new_[71125]_  = A299 & ~A298;
  assign \new_[71128]_  = A301 & A300;
  assign \new_[71129]_  = \new_[71128]_  & \new_[71125]_ ;
  assign \new_[71130]_  = \new_[71129]_  & \new_[71122]_ ;
  assign \new_[71134]_  = ~A168 & ~A169;
  assign \new_[71135]_  = A170 & \new_[71134]_ ;
  assign \new_[71138]_  = ~A166 & A167;
  assign \new_[71141]_  = ~A202 & A201;
  assign \new_[71142]_  = \new_[71141]_  & \new_[71138]_ ;
  assign \new_[71143]_  = \new_[71142]_  & \new_[71135]_ ;
  assign \new_[71147]_  = A269 & ~A267;
  assign \new_[71148]_  = ~A203 & \new_[71147]_ ;
  assign \new_[71151]_  = A299 & ~A298;
  assign \new_[71154]_  = A302 & A300;
  assign \new_[71155]_  = \new_[71154]_  & \new_[71151]_ ;
  assign \new_[71156]_  = \new_[71155]_  & \new_[71148]_ ;
  assign \new_[71160]_  = ~A168 & ~A169;
  assign \new_[71161]_  = A170 & \new_[71160]_ ;
  assign \new_[71164]_  = ~A166 & A167;
  assign \new_[71167]_  = ~A202 & A201;
  assign \new_[71168]_  = \new_[71167]_  & \new_[71164]_ ;
  assign \new_[71169]_  = \new_[71168]_  & \new_[71161]_ ;
  assign \new_[71173]_  = A266 & A265;
  assign \new_[71174]_  = ~A203 & \new_[71173]_ ;
  assign \new_[71177]_  = ~A299 & A298;
  assign \new_[71180]_  = A301 & A300;
  assign \new_[71181]_  = \new_[71180]_  & \new_[71177]_ ;
  assign \new_[71182]_  = \new_[71181]_  & \new_[71174]_ ;
  assign \new_[71186]_  = ~A168 & ~A169;
  assign \new_[71187]_  = A170 & \new_[71186]_ ;
  assign \new_[71190]_  = ~A166 & A167;
  assign \new_[71193]_  = ~A202 & A201;
  assign \new_[71194]_  = \new_[71193]_  & \new_[71190]_ ;
  assign \new_[71195]_  = \new_[71194]_  & \new_[71187]_ ;
  assign \new_[71199]_  = A266 & A265;
  assign \new_[71200]_  = ~A203 & \new_[71199]_ ;
  assign \new_[71203]_  = ~A299 & A298;
  assign \new_[71206]_  = A302 & A300;
  assign \new_[71207]_  = \new_[71206]_  & \new_[71203]_ ;
  assign \new_[71208]_  = \new_[71207]_  & \new_[71200]_ ;
  assign \new_[71212]_  = ~A168 & ~A169;
  assign \new_[71213]_  = A170 & \new_[71212]_ ;
  assign \new_[71216]_  = ~A166 & A167;
  assign \new_[71219]_  = ~A202 & A201;
  assign \new_[71220]_  = \new_[71219]_  & \new_[71216]_ ;
  assign \new_[71221]_  = \new_[71220]_  & \new_[71213]_ ;
  assign \new_[71225]_  = A266 & A265;
  assign \new_[71226]_  = ~A203 & \new_[71225]_ ;
  assign \new_[71229]_  = A299 & ~A298;
  assign \new_[71232]_  = A301 & A300;
  assign \new_[71233]_  = \new_[71232]_  & \new_[71229]_ ;
  assign \new_[71234]_  = \new_[71233]_  & \new_[71226]_ ;
  assign \new_[71238]_  = ~A168 & ~A169;
  assign \new_[71239]_  = A170 & \new_[71238]_ ;
  assign \new_[71242]_  = ~A166 & A167;
  assign \new_[71245]_  = ~A202 & A201;
  assign \new_[71246]_  = \new_[71245]_  & \new_[71242]_ ;
  assign \new_[71247]_  = \new_[71246]_  & \new_[71239]_ ;
  assign \new_[71251]_  = A266 & A265;
  assign \new_[71252]_  = ~A203 & \new_[71251]_ ;
  assign \new_[71255]_  = A299 & ~A298;
  assign \new_[71258]_  = A302 & A300;
  assign \new_[71259]_  = \new_[71258]_  & \new_[71255]_ ;
  assign \new_[71260]_  = \new_[71259]_  & \new_[71252]_ ;
  assign \new_[71264]_  = ~A168 & ~A169;
  assign \new_[71265]_  = A170 & \new_[71264]_ ;
  assign \new_[71268]_  = ~A166 & A167;
  assign \new_[71271]_  = ~A202 & A201;
  assign \new_[71272]_  = \new_[71271]_  & \new_[71268]_ ;
  assign \new_[71273]_  = \new_[71272]_  & \new_[71265]_ ;
  assign \new_[71277]_  = ~A266 & ~A265;
  assign \new_[71278]_  = ~A203 & \new_[71277]_ ;
  assign \new_[71281]_  = ~A299 & A298;
  assign \new_[71284]_  = A301 & A300;
  assign \new_[71285]_  = \new_[71284]_  & \new_[71281]_ ;
  assign \new_[71286]_  = \new_[71285]_  & \new_[71278]_ ;
  assign \new_[71290]_  = ~A168 & ~A169;
  assign \new_[71291]_  = A170 & \new_[71290]_ ;
  assign \new_[71294]_  = ~A166 & A167;
  assign \new_[71297]_  = ~A202 & A201;
  assign \new_[71298]_  = \new_[71297]_  & \new_[71294]_ ;
  assign \new_[71299]_  = \new_[71298]_  & \new_[71291]_ ;
  assign \new_[71303]_  = ~A266 & ~A265;
  assign \new_[71304]_  = ~A203 & \new_[71303]_ ;
  assign \new_[71307]_  = ~A299 & A298;
  assign \new_[71310]_  = A302 & A300;
  assign \new_[71311]_  = \new_[71310]_  & \new_[71307]_ ;
  assign \new_[71312]_  = \new_[71311]_  & \new_[71304]_ ;
  assign \new_[71316]_  = ~A168 & ~A169;
  assign \new_[71317]_  = A170 & \new_[71316]_ ;
  assign \new_[71320]_  = ~A166 & A167;
  assign \new_[71323]_  = ~A202 & A201;
  assign \new_[71324]_  = \new_[71323]_  & \new_[71320]_ ;
  assign \new_[71325]_  = \new_[71324]_  & \new_[71317]_ ;
  assign \new_[71329]_  = ~A266 & ~A265;
  assign \new_[71330]_  = ~A203 & \new_[71329]_ ;
  assign \new_[71333]_  = A299 & ~A298;
  assign \new_[71336]_  = A301 & A300;
  assign \new_[71337]_  = \new_[71336]_  & \new_[71333]_ ;
  assign \new_[71338]_  = \new_[71337]_  & \new_[71330]_ ;
  assign \new_[71342]_  = ~A168 & ~A169;
  assign \new_[71343]_  = A170 & \new_[71342]_ ;
  assign \new_[71346]_  = ~A166 & A167;
  assign \new_[71349]_  = ~A202 & A201;
  assign \new_[71350]_  = \new_[71349]_  & \new_[71346]_ ;
  assign \new_[71351]_  = \new_[71350]_  & \new_[71343]_ ;
  assign \new_[71355]_  = ~A266 & ~A265;
  assign \new_[71356]_  = ~A203 & \new_[71355]_ ;
  assign \new_[71359]_  = A299 & ~A298;
  assign \new_[71362]_  = A302 & A300;
  assign \new_[71363]_  = \new_[71362]_  & \new_[71359]_ ;
  assign \new_[71364]_  = \new_[71363]_  & \new_[71356]_ ;
  assign \new_[71368]_  = ~A168 & ~A169;
  assign \new_[71369]_  = A170 & \new_[71368]_ ;
  assign \new_[71372]_  = ~A166 & A167;
  assign \new_[71375]_  = A202 & ~A201;
  assign \new_[71376]_  = \new_[71375]_  & \new_[71372]_ ;
  assign \new_[71377]_  = \new_[71376]_  & \new_[71369]_ ;
  assign \new_[71381]_  = ~A269 & ~A268;
  assign \new_[71382]_  = A267 & \new_[71381]_ ;
  assign \new_[71385]_  = ~A299 & A298;
  assign \new_[71388]_  = A301 & A300;
  assign \new_[71389]_  = \new_[71388]_  & \new_[71385]_ ;
  assign \new_[71390]_  = \new_[71389]_  & \new_[71382]_ ;
  assign \new_[71394]_  = ~A168 & ~A169;
  assign \new_[71395]_  = A170 & \new_[71394]_ ;
  assign \new_[71398]_  = ~A166 & A167;
  assign \new_[71401]_  = A202 & ~A201;
  assign \new_[71402]_  = \new_[71401]_  & \new_[71398]_ ;
  assign \new_[71403]_  = \new_[71402]_  & \new_[71395]_ ;
  assign \new_[71407]_  = ~A269 & ~A268;
  assign \new_[71408]_  = A267 & \new_[71407]_ ;
  assign \new_[71411]_  = ~A299 & A298;
  assign \new_[71414]_  = A302 & A300;
  assign \new_[71415]_  = \new_[71414]_  & \new_[71411]_ ;
  assign \new_[71416]_  = \new_[71415]_  & \new_[71408]_ ;
  assign \new_[71420]_  = ~A168 & ~A169;
  assign \new_[71421]_  = A170 & \new_[71420]_ ;
  assign \new_[71424]_  = ~A166 & A167;
  assign \new_[71427]_  = A202 & ~A201;
  assign \new_[71428]_  = \new_[71427]_  & \new_[71424]_ ;
  assign \new_[71429]_  = \new_[71428]_  & \new_[71421]_ ;
  assign \new_[71433]_  = ~A269 & ~A268;
  assign \new_[71434]_  = A267 & \new_[71433]_ ;
  assign \new_[71437]_  = A299 & ~A298;
  assign \new_[71440]_  = A301 & A300;
  assign \new_[71441]_  = \new_[71440]_  & \new_[71437]_ ;
  assign \new_[71442]_  = \new_[71441]_  & \new_[71434]_ ;
  assign \new_[71446]_  = ~A168 & ~A169;
  assign \new_[71447]_  = A170 & \new_[71446]_ ;
  assign \new_[71450]_  = ~A166 & A167;
  assign \new_[71453]_  = A202 & ~A201;
  assign \new_[71454]_  = \new_[71453]_  & \new_[71450]_ ;
  assign \new_[71455]_  = \new_[71454]_  & \new_[71447]_ ;
  assign \new_[71459]_  = ~A269 & ~A268;
  assign \new_[71460]_  = A267 & \new_[71459]_ ;
  assign \new_[71463]_  = A299 & ~A298;
  assign \new_[71466]_  = A302 & A300;
  assign \new_[71467]_  = \new_[71466]_  & \new_[71463]_ ;
  assign \new_[71468]_  = \new_[71467]_  & \new_[71460]_ ;
  assign \new_[71472]_  = ~A168 & ~A169;
  assign \new_[71473]_  = A170 & \new_[71472]_ ;
  assign \new_[71476]_  = ~A166 & A167;
  assign \new_[71479]_  = A202 & ~A201;
  assign \new_[71480]_  = \new_[71479]_  & \new_[71476]_ ;
  assign \new_[71481]_  = \new_[71480]_  & \new_[71473]_ ;
  assign \new_[71485]_  = A298 & A268;
  assign \new_[71486]_  = ~A267 & \new_[71485]_ ;
  assign \new_[71489]_  = ~A300 & ~A299;
  assign \new_[71492]_  = ~A302 & ~A301;
  assign \new_[71493]_  = \new_[71492]_  & \new_[71489]_ ;
  assign \new_[71494]_  = \new_[71493]_  & \new_[71486]_ ;
  assign \new_[71498]_  = ~A168 & ~A169;
  assign \new_[71499]_  = A170 & \new_[71498]_ ;
  assign \new_[71502]_  = ~A166 & A167;
  assign \new_[71505]_  = A202 & ~A201;
  assign \new_[71506]_  = \new_[71505]_  & \new_[71502]_ ;
  assign \new_[71507]_  = \new_[71506]_  & \new_[71499]_ ;
  assign \new_[71511]_  = ~A298 & A268;
  assign \new_[71512]_  = ~A267 & \new_[71511]_ ;
  assign \new_[71515]_  = ~A300 & A299;
  assign \new_[71518]_  = ~A302 & ~A301;
  assign \new_[71519]_  = \new_[71518]_  & \new_[71515]_ ;
  assign \new_[71520]_  = \new_[71519]_  & \new_[71512]_ ;
  assign \new_[71524]_  = ~A168 & ~A169;
  assign \new_[71525]_  = A170 & \new_[71524]_ ;
  assign \new_[71528]_  = ~A166 & A167;
  assign \new_[71531]_  = A202 & ~A201;
  assign \new_[71532]_  = \new_[71531]_  & \new_[71528]_ ;
  assign \new_[71533]_  = \new_[71532]_  & \new_[71525]_ ;
  assign \new_[71537]_  = A298 & A269;
  assign \new_[71538]_  = ~A267 & \new_[71537]_ ;
  assign \new_[71541]_  = ~A300 & ~A299;
  assign \new_[71544]_  = ~A302 & ~A301;
  assign \new_[71545]_  = \new_[71544]_  & \new_[71541]_ ;
  assign \new_[71546]_  = \new_[71545]_  & \new_[71538]_ ;
  assign \new_[71550]_  = ~A168 & ~A169;
  assign \new_[71551]_  = A170 & \new_[71550]_ ;
  assign \new_[71554]_  = ~A166 & A167;
  assign \new_[71557]_  = A202 & ~A201;
  assign \new_[71558]_  = \new_[71557]_  & \new_[71554]_ ;
  assign \new_[71559]_  = \new_[71558]_  & \new_[71551]_ ;
  assign \new_[71563]_  = ~A298 & A269;
  assign \new_[71564]_  = ~A267 & \new_[71563]_ ;
  assign \new_[71567]_  = ~A300 & A299;
  assign \new_[71570]_  = ~A302 & ~A301;
  assign \new_[71571]_  = \new_[71570]_  & \new_[71567]_ ;
  assign \new_[71572]_  = \new_[71571]_  & \new_[71564]_ ;
  assign \new_[71576]_  = ~A168 & ~A169;
  assign \new_[71577]_  = A170 & \new_[71576]_ ;
  assign \new_[71580]_  = ~A166 & A167;
  assign \new_[71583]_  = A202 & ~A201;
  assign \new_[71584]_  = \new_[71583]_  & \new_[71580]_ ;
  assign \new_[71585]_  = \new_[71584]_  & \new_[71577]_ ;
  assign \new_[71589]_  = A298 & A266;
  assign \new_[71590]_  = A265 & \new_[71589]_ ;
  assign \new_[71593]_  = ~A300 & ~A299;
  assign \new_[71596]_  = ~A302 & ~A301;
  assign \new_[71597]_  = \new_[71596]_  & \new_[71593]_ ;
  assign \new_[71598]_  = \new_[71597]_  & \new_[71590]_ ;
  assign \new_[71602]_  = ~A168 & ~A169;
  assign \new_[71603]_  = A170 & \new_[71602]_ ;
  assign \new_[71606]_  = ~A166 & A167;
  assign \new_[71609]_  = A202 & ~A201;
  assign \new_[71610]_  = \new_[71609]_  & \new_[71606]_ ;
  assign \new_[71611]_  = \new_[71610]_  & \new_[71603]_ ;
  assign \new_[71615]_  = ~A298 & A266;
  assign \new_[71616]_  = A265 & \new_[71615]_ ;
  assign \new_[71619]_  = ~A300 & A299;
  assign \new_[71622]_  = ~A302 & ~A301;
  assign \new_[71623]_  = \new_[71622]_  & \new_[71619]_ ;
  assign \new_[71624]_  = \new_[71623]_  & \new_[71616]_ ;
  assign \new_[71628]_  = ~A168 & ~A169;
  assign \new_[71629]_  = A170 & \new_[71628]_ ;
  assign \new_[71632]_  = ~A166 & A167;
  assign \new_[71635]_  = A202 & ~A201;
  assign \new_[71636]_  = \new_[71635]_  & \new_[71632]_ ;
  assign \new_[71637]_  = \new_[71636]_  & \new_[71629]_ ;
  assign \new_[71641]_  = A298 & ~A266;
  assign \new_[71642]_  = ~A265 & \new_[71641]_ ;
  assign \new_[71645]_  = ~A300 & ~A299;
  assign \new_[71648]_  = ~A302 & ~A301;
  assign \new_[71649]_  = \new_[71648]_  & \new_[71645]_ ;
  assign \new_[71650]_  = \new_[71649]_  & \new_[71642]_ ;
  assign \new_[71654]_  = ~A168 & ~A169;
  assign \new_[71655]_  = A170 & \new_[71654]_ ;
  assign \new_[71658]_  = ~A166 & A167;
  assign \new_[71661]_  = A202 & ~A201;
  assign \new_[71662]_  = \new_[71661]_  & \new_[71658]_ ;
  assign \new_[71663]_  = \new_[71662]_  & \new_[71655]_ ;
  assign \new_[71667]_  = ~A298 & ~A266;
  assign \new_[71668]_  = ~A265 & \new_[71667]_ ;
  assign \new_[71671]_  = ~A300 & A299;
  assign \new_[71674]_  = ~A302 & ~A301;
  assign \new_[71675]_  = \new_[71674]_  & \new_[71671]_ ;
  assign \new_[71676]_  = \new_[71675]_  & \new_[71668]_ ;
  assign \new_[71680]_  = ~A168 & ~A169;
  assign \new_[71681]_  = A170 & \new_[71680]_ ;
  assign \new_[71684]_  = ~A166 & A167;
  assign \new_[71687]_  = A203 & ~A201;
  assign \new_[71688]_  = \new_[71687]_  & \new_[71684]_ ;
  assign \new_[71689]_  = \new_[71688]_  & \new_[71681]_ ;
  assign \new_[71693]_  = ~A269 & ~A268;
  assign \new_[71694]_  = A267 & \new_[71693]_ ;
  assign \new_[71697]_  = ~A299 & A298;
  assign \new_[71700]_  = A301 & A300;
  assign \new_[71701]_  = \new_[71700]_  & \new_[71697]_ ;
  assign \new_[71702]_  = \new_[71701]_  & \new_[71694]_ ;
  assign \new_[71706]_  = ~A168 & ~A169;
  assign \new_[71707]_  = A170 & \new_[71706]_ ;
  assign \new_[71710]_  = ~A166 & A167;
  assign \new_[71713]_  = A203 & ~A201;
  assign \new_[71714]_  = \new_[71713]_  & \new_[71710]_ ;
  assign \new_[71715]_  = \new_[71714]_  & \new_[71707]_ ;
  assign \new_[71719]_  = ~A269 & ~A268;
  assign \new_[71720]_  = A267 & \new_[71719]_ ;
  assign \new_[71723]_  = ~A299 & A298;
  assign \new_[71726]_  = A302 & A300;
  assign \new_[71727]_  = \new_[71726]_  & \new_[71723]_ ;
  assign \new_[71728]_  = \new_[71727]_  & \new_[71720]_ ;
  assign \new_[71732]_  = ~A168 & ~A169;
  assign \new_[71733]_  = A170 & \new_[71732]_ ;
  assign \new_[71736]_  = ~A166 & A167;
  assign \new_[71739]_  = A203 & ~A201;
  assign \new_[71740]_  = \new_[71739]_  & \new_[71736]_ ;
  assign \new_[71741]_  = \new_[71740]_  & \new_[71733]_ ;
  assign \new_[71745]_  = ~A269 & ~A268;
  assign \new_[71746]_  = A267 & \new_[71745]_ ;
  assign \new_[71749]_  = A299 & ~A298;
  assign \new_[71752]_  = A301 & A300;
  assign \new_[71753]_  = \new_[71752]_  & \new_[71749]_ ;
  assign \new_[71754]_  = \new_[71753]_  & \new_[71746]_ ;
  assign \new_[71758]_  = ~A168 & ~A169;
  assign \new_[71759]_  = A170 & \new_[71758]_ ;
  assign \new_[71762]_  = ~A166 & A167;
  assign \new_[71765]_  = A203 & ~A201;
  assign \new_[71766]_  = \new_[71765]_  & \new_[71762]_ ;
  assign \new_[71767]_  = \new_[71766]_  & \new_[71759]_ ;
  assign \new_[71771]_  = ~A269 & ~A268;
  assign \new_[71772]_  = A267 & \new_[71771]_ ;
  assign \new_[71775]_  = A299 & ~A298;
  assign \new_[71778]_  = A302 & A300;
  assign \new_[71779]_  = \new_[71778]_  & \new_[71775]_ ;
  assign \new_[71780]_  = \new_[71779]_  & \new_[71772]_ ;
  assign \new_[71784]_  = ~A168 & ~A169;
  assign \new_[71785]_  = A170 & \new_[71784]_ ;
  assign \new_[71788]_  = ~A166 & A167;
  assign \new_[71791]_  = A203 & ~A201;
  assign \new_[71792]_  = \new_[71791]_  & \new_[71788]_ ;
  assign \new_[71793]_  = \new_[71792]_  & \new_[71785]_ ;
  assign \new_[71797]_  = A298 & A268;
  assign \new_[71798]_  = ~A267 & \new_[71797]_ ;
  assign \new_[71801]_  = ~A300 & ~A299;
  assign \new_[71804]_  = ~A302 & ~A301;
  assign \new_[71805]_  = \new_[71804]_  & \new_[71801]_ ;
  assign \new_[71806]_  = \new_[71805]_  & \new_[71798]_ ;
  assign \new_[71810]_  = ~A168 & ~A169;
  assign \new_[71811]_  = A170 & \new_[71810]_ ;
  assign \new_[71814]_  = ~A166 & A167;
  assign \new_[71817]_  = A203 & ~A201;
  assign \new_[71818]_  = \new_[71817]_  & \new_[71814]_ ;
  assign \new_[71819]_  = \new_[71818]_  & \new_[71811]_ ;
  assign \new_[71823]_  = ~A298 & A268;
  assign \new_[71824]_  = ~A267 & \new_[71823]_ ;
  assign \new_[71827]_  = ~A300 & A299;
  assign \new_[71830]_  = ~A302 & ~A301;
  assign \new_[71831]_  = \new_[71830]_  & \new_[71827]_ ;
  assign \new_[71832]_  = \new_[71831]_  & \new_[71824]_ ;
  assign \new_[71836]_  = ~A168 & ~A169;
  assign \new_[71837]_  = A170 & \new_[71836]_ ;
  assign \new_[71840]_  = ~A166 & A167;
  assign \new_[71843]_  = A203 & ~A201;
  assign \new_[71844]_  = \new_[71843]_  & \new_[71840]_ ;
  assign \new_[71845]_  = \new_[71844]_  & \new_[71837]_ ;
  assign \new_[71849]_  = A298 & A269;
  assign \new_[71850]_  = ~A267 & \new_[71849]_ ;
  assign \new_[71853]_  = ~A300 & ~A299;
  assign \new_[71856]_  = ~A302 & ~A301;
  assign \new_[71857]_  = \new_[71856]_  & \new_[71853]_ ;
  assign \new_[71858]_  = \new_[71857]_  & \new_[71850]_ ;
  assign \new_[71862]_  = ~A168 & ~A169;
  assign \new_[71863]_  = A170 & \new_[71862]_ ;
  assign \new_[71866]_  = ~A166 & A167;
  assign \new_[71869]_  = A203 & ~A201;
  assign \new_[71870]_  = \new_[71869]_  & \new_[71866]_ ;
  assign \new_[71871]_  = \new_[71870]_  & \new_[71863]_ ;
  assign \new_[71875]_  = ~A298 & A269;
  assign \new_[71876]_  = ~A267 & \new_[71875]_ ;
  assign \new_[71879]_  = ~A300 & A299;
  assign \new_[71882]_  = ~A302 & ~A301;
  assign \new_[71883]_  = \new_[71882]_  & \new_[71879]_ ;
  assign \new_[71884]_  = \new_[71883]_  & \new_[71876]_ ;
  assign \new_[71888]_  = ~A168 & ~A169;
  assign \new_[71889]_  = A170 & \new_[71888]_ ;
  assign \new_[71892]_  = ~A166 & A167;
  assign \new_[71895]_  = A203 & ~A201;
  assign \new_[71896]_  = \new_[71895]_  & \new_[71892]_ ;
  assign \new_[71897]_  = \new_[71896]_  & \new_[71889]_ ;
  assign \new_[71901]_  = A298 & A266;
  assign \new_[71902]_  = A265 & \new_[71901]_ ;
  assign \new_[71905]_  = ~A300 & ~A299;
  assign \new_[71908]_  = ~A302 & ~A301;
  assign \new_[71909]_  = \new_[71908]_  & \new_[71905]_ ;
  assign \new_[71910]_  = \new_[71909]_  & \new_[71902]_ ;
  assign \new_[71914]_  = ~A168 & ~A169;
  assign \new_[71915]_  = A170 & \new_[71914]_ ;
  assign \new_[71918]_  = ~A166 & A167;
  assign \new_[71921]_  = A203 & ~A201;
  assign \new_[71922]_  = \new_[71921]_  & \new_[71918]_ ;
  assign \new_[71923]_  = \new_[71922]_  & \new_[71915]_ ;
  assign \new_[71927]_  = ~A298 & A266;
  assign \new_[71928]_  = A265 & \new_[71927]_ ;
  assign \new_[71931]_  = ~A300 & A299;
  assign \new_[71934]_  = ~A302 & ~A301;
  assign \new_[71935]_  = \new_[71934]_  & \new_[71931]_ ;
  assign \new_[71936]_  = \new_[71935]_  & \new_[71928]_ ;
  assign \new_[71940]_  = ~A168 & ~A169;
  assign \new_[71941]_  = A170 & \new_[71940]_ ;
  assign \new_[71944]_  = ~A166 & A167;
  assign \new_[71947]_  = A203 & ~A201;
  assign \new_[71948]_  = \new_[71947]_  & \new_[71944]_ ;
  assign \new_[71949]_  = \new_[71948]_  & \new_[71941]_ ;
  assign \new_[71953]_  = A298 & ~A266;
  assign \new_[71954]_  = ~A265 & \new_[71953]_ ;
  assign \new_[71957]_  = ~A300 & ~A299;
  assign \new_[71960]_  = ~A302 & ~A301;
  assign \new_[71961]_  = \new_[71960]_  & \new_[71957]_ ;
  assign \new_[71962]_  = \new_[71961]_  & \new_[71954]_ ;
  assign \new_[71966]_  = ~A168 & ~A169;
  assign \new_[71967]_  = A170 & \new_[71966]_ ;
  assign \new_[71970]_  = ~A166 & A167;
  assign \new_[71973]_  = A203 & ~A201;
  assign \new_[71974]_  = \new_[71973]_  & \new_[71970]_ ;
  assign \new_[71975]_  = \new_[71974]_  & \new_[71967]_ ;
  assign \new_[71979]_  = ~A298 & ~A266;
  assign \new_[71980]_  = ~A265 & \new_[71979]_ ;
  assign \new_[71983]_  = ~A300 & A299;
  assign \new_[71986]_  = ~A302 & ~A301;
  assign \new_[71987]_  = \new_[71986]_  & \new_[71983]_ ;
  assign \new_[71988]_  = \new_[71987]_  & \new_[71980]_ ;
  assign \new_[71992]_  = ~A168 & ~A169;
  assign \new_[71993]_  = A170 & \new_[71992]_ ;
  assign \new_[71996]_  = ~A166 & A167;
  assign \new_[71999]_  = A200 & A199;
  assign \new_[72000]_  = \new_[71999]_  & \new_[71996]_ ;
  assign \new_[72001]_  = \new_[72000]_  & \new_[71993]_ ;
  assign \new_[72005]_  = ~A269 & ~A268;
  assign \new_[72006]_  = A267 & \new_[72005]_ ;
  assign \new_[72009]_  = ~A299 & A298;
  assign \new_[72012]_  = A301 & A300;
  assign \new_[72013]_  = \new_[72012]_  & \new_[72009]_ ;
  assign \new_[72014]_  = \new_[72013]_  & \new_[72006]_ ;
  assign \new_[72018]_  = ~A168 & ~A169;
  assign \new_[72019]_  = A170 & \new_[72018]_ ;
  assign \new_[72022]_  = ~A166 & A167;
  assign \new_[72025]_  = A200 & A199;
  assign \new_[72026]_  = \new_[72025]_  & \new_[72022]_ ;
  assign \new_[72027]_  = \new_[72026]_  & \new_[72019]_ ;
  assign \new_[72031]_  = ~A269 & ~A268;
  assign \new_[72032]_  = A267 & \new_[72031]_ ;
  assign \new_[72035]_  = ~A299 & A298;
  assign \new_[72038]_  = A302 & A300;
  assign \new_[72039]_  = \new_[72038]_  & \new_[72035]_ ;
  assign \new_[72040]_  = \new_[72039]_  & \new_[72032]_ ;
  assign \new_[72044]_  = ~A168 & ~A169;
  assign \new_[72045]_  = A170 & \new_[72044]_ ;
  assign \new_[72048]_  = ~A166 & A167;
  assign \new_[72051]_  = A200 & A199;
  assign \new_[72052]_  = \new_[72051]_  & \new_[72048]_ ;
  assign \new_[72053]_  = \new_[72052]_  & \new_[72045]_ ;
  assign \new_[72057]_  = ~A269 & ~A268;
  assign \new_[72058]_  = A267 & \new_[72057]_ ;
  assign \new_[72061]_  = A299 & ~A298;
  assign \new_[72064]_  = A301 & A300;
  assign \new_[72065]_  = \new_[72064]_  & \new_[72061]_ ;
  assign \new_[72066]_  = \new_[72065]_  & \new_[72058]_ ;
  assign \new_[72070]_  = ~A168 & ~A169;
  assign \new_[72071]_  = A170 & \new_[72070]_ ;
  assign \new_[72074]_  = ~A166 & A167;
  assign \new_[72077]_  = A200 & A199;
  assign \new_[72078]_  = \new_[72077]_  & \new_[72074]_ ;
  assign \new_[72079]_  = \new_[72078]_  & \new_[72071]_ ;
  assign \new_[72083]_  = ~A269 & ~A268;
  assign \new_[72084]_  = A267 & \new_[72083]_ ;
  assign \new_[72087]_  = A299 & ~A298;
  assign \new_[72090]_  = A302 & A300;
  assign \new_[72091]_  = \new_[72090]_  & \new_[72087]_ ;
  assign \new_[72092]_  = \new_[72091]_  & \new_[72084]_ ;
  assign \new_[72096]_  = ~A168 & ~A169;
  assign \new_[72097]_  = A170 & \new_[72096]_ ;
  assign \new_[72100]_  = ~A166 & A167;
  assign \new_[72103]_  = A200 & A199;
  assign \new_[72104]_  = \new_[72103]_  & \new_[72100]_ ;
  assign \new_[72105]_  = \new_[72104]_  & \new_[72097]_ ;
  assign \new_[72109]_  = A298 & A268;
  assign \new_[72110]_  = ~A267 & \new_[72109]_ ;
  assign \new_[72113]_  = ~A300 & ~A299;
  assign \new_[72116]_  = ~A302 & ~A301;
  assign \new_[72117]_  = \new_[72116]_  & \new_[72113]_ ;
  assign \new_[72118]_  = \new_[72117]_  & \new_[72110]_ ;
  assign \new_[72122]_  = ~A168 & ~A169;
  assign \new_[72123]_  = A170 & \new_[72122]_ ;
  assign \new_[72126]_  = ~A166 & A167;
  assign \new_[72129]_  = A200 & A199;
  assign \new_[72130]_  = \new_[72129]_  & \new_[72126]_ ;
  assign \new_[72131]_  = \new_[72130]_  & \new_[72123]_ ;
  assign \new_[72135]_  = ~A298 & A268;
  assign \new_[72136]_  = ~A267 & \new_[72135]_ ;
  assign \new_[72139]_  = ~A300 & A299;
  assign \new_[72142]_  = ~A302 & ~A301;
  assign \new_[72143]_  = \new_[72142]_  & \new_[72139]_ ;
  assign \new_[72144]_  = \new_[72143]_  & \new_[72136]_ ;
  assign \new_[72148]_  = ~A168 & ~A169;
  assign \new_[72149]_  = A170 & \new_[72148]_ ;
  assign \new_[72152]_  = ~A166 & A167;
  assign \new_[72155]_  = A200 & A199;
  assign \new_[72156]_  = \new_[72155]_  & \new_[72152]_ ;
  assign \new_[72157]_  = \new_[72156]_  & \new_[72149]_ ;
  assign \new_[72161]_  = A298 & A269;
  assign \new_[72162]_  = ~A267 & \new_[72161]_ ;
  assign \new_[72165]_  = ~A300 & ~A299;
  assign \new_[72168]_  = ~A302 & ~A301;
  assign \new_[72169]_  = \new_[72168]_  & \new_[72165]_ ;
  assign \new_[72170]_  = \new_[72169]_  & \new_[72162]_ ;
  assign \new_[72174]_  = ~A168 & ~A169;
  assign \new_[72175]_  = A170 & \new_[72174]_ ;
  assign \new_[72178]_  = ~A166 & A167;
  assign \new_[72181]_  = A200 & A199;
  assign \new_[72182]_  = \new_[72181]_  & \new_[72178]_ ;
  assign \new_[72183]_  = \new_[72182]_  & \new_[72175]_ ;
  assign \new_[72187]_  = ~A298 & A269;
  assign \new_[72188]_  = ~A267 & \new_[72187]_ ;
  assign \new_[72191]_  = ~A300 & A299;
  assign \new_[72194]_  = ~A302 & ~A301;
  assign \new_[72195]_  = \new_[72194]_  & \new_[72191]_ ;
  assign \new_[72196]_  = \new_[72195]_  & \new_[72188]_ ;
  assign \new_[72200]_  = ~A168 & ~A169;
  assign \new_[72201]_  = A170 & \new_[72200]_ ;
  assign \new_[72204]_  = ~A166 & A167;
  assign \new_[72207]_  = A200 & A199;
  assign \new_[72208]_  = \new_[72207]_  & \new_[72204]_ ;
  assign \new_[72209]_  = \new_[72208]_  & \new_[72201]_ ;
  assign \new_[72213]_  = A298 & A266;
  assign \new_[72214]_  = A265 & \new_[72213]_ ;
  assign \new_[72217]_  = ~A300 & ~A299;
  assign \new_[72220]_  = ~A302 & ~A301;
  assign \new_[72221]_  = \new_[72220]_  & \new_[72217]_ ;
  assign \new_[72222]_  = \new_[72221]_  & \new_[72214]_ ;
  assign \new_[72226]_  = ~A168 & ~A169;
  assign \new_[72227]_  = A170 & \new_[72226]_ ;
  assign \new_[72230]_  = ~A166 & A167;
  assign \new_[72233]_  = A200 & A199;
  assign \new_[72234]_  = \new_[72233]_  & \new_[72230]_ ;
  assign \new_[72235]_  = \new_[72234]_  & \new_[72227]_ ;
  assign \new_[72239]_  = ~A298 & A266;
  assign \new_[72240]_  = A265 & \new_[72239]_ ;
  assign \new_[72243]_  = ~A300 & A299;
  assign \new_[72246]_  = ~A302 & ~A301;
  assign \new_[72247]_  = \new_[72246]_  & \new_[72243]_ ;
  assign \new_[72248]_  = \new_[72247]_  & \new_[72240]_ ;
  assign \new_[72252]_  = ~A168 & ~A169;
  assign \new_[72253]_  = A170 & \new_[72252]_ ;
  assign \new_[72256]_  = ~A166 & A167;
  assign \new_[72259]_  = A200 & A199;
  assign \new_[72260]_  = \new_[72259]_  & \new_[72256]_ ;
  assign \new_[72261]_  = \new_[72260]_  & \new_[72253]_ ;
  assign \new_[72265]_  = A298 & ~A266;
  assign \new_[72266]_  = ~A265 & \new_[72265]_ ;
  assign \new_[72269]_  = ~A300 & ~A299;
  assign \new_[72272]_  = ~A302 & ~A301;
  assign \new_[72273]_  = \new_[72272]_  & \new_[72269]_ ;
  assign \new_[72274]_  = \new_[72273]_  & \new_[72266]_ ;
  assign \new_[72278]_  = ~A168 & ~A169;
  assign \new_[72279]_  = A170 & \new_[72278]_ ;
  assign \new_[72282]_  = ~A166 & A167;
  assign \new_[72285]_  = A200 & A199;
  assign \new_[72286]_  = \new_[72285]_  & \new_[72282]_ ;
  assign \new_[72287]_  = \new_[72286]_  & \new_[72279]_ ;
  assign \new_[72291]_  = ~A298 & ~A266;
  assign \new_[72292]_  = ~A265 & \new_[72291]_ ;
  assign \new_[72295]_  = ~A300 & A299;
  assign \new_[72298]_  = ~A302 & ~A301;
  assign \new_[72299]_  = \new_[72298]_  & \new_[72295]_ ;
  assign \new_[72300]_  = \new_[72299]_  & \new_[72292]_ ;
  assign \new_[72304]_  = ~A168 & ~A169;
  assign \new_[72305]_  = A170 & \new_[72304]_ ;
  assign \new_[72308]_  = ~A166 & A167;
  assign \new_[72311]_  = ~A200 & ~A199;
  assign \new_[72312]_  = \new_[72311]_  & \new_[72308]_ ;
  assign \new_[72313]_  = \new_[72312]_  & \new_[72305]_ ;
  assign \new_[72317]_  = ~A269 & ~A268;
  assign \new_[72318]_  = A267 & \new_[72317]_ ;
  assign \new_[72321]_  = ~A299 & A298;
  assign \new_[72324]_  = A301 & A300;
  assign \new_[72325]_  = \new_[72324]_  & \new_[72321]_ ;
  assign \new_[72326]_  = \new_[72325]_  & \new_[72318]_ ;
  assign \new_[72330]_  = ~A168 & ~A169;
  assign \new_[72331]_  = A170 & \new_[72330]_ ;
  assign \new_[72334]_  = ~A166 & A167;
  assign \new_[72337]_  = ~A200 & ~A199;
  assign \new_[72338]_  = \new_[72337]_  & \new_[72334]_ ;
  assign \new_[72339]_  = \new_[72338]_  & \new_[72331]_ ;
  assign \new_[72343]_  = ~A269 & ~A268;
  assign \new_[72344]_  = A267 & \new_[72343]_ ;
  assign \new_[72347]_  = ~A299 & A298;
  assign \new_[72350]_  = A302 & A300;
  assign \new_[72351]_  = \new_[72350]_  & \new_[72347]_ ;
  assign \new_[72352]_  = \new_[72351]_  & \new_[72344]_ ;
  assign \new_[72356]_  = ~A168 & ~A169;
  assign \new_[72357]_  = A170 & \new_[72356]_ ;
  assign \new_[72360]_  = ~A166 & A167;
  assign \new_[72363]_  = ~A200 & ~A199;
  assign \new_[72364]_  = \new_[72363]_  & \new_[72360]_ ;
  assign \new_[72365]_  = \new_[72364]_  & \new_[72357]_ ;
  assign \new_[72369]_  = ~A269 & ~A268;
  assign \new_[72370]_  = A267 & \new_[72369]_ ;
  assign \new_[72373]_  = A299 & ~A298;
  assign \new_[72376]_  = A301 & A300;
  assign \new_[72377]_  = \new_[72376]_  & \new_[72373]_ ;
  assign \new_[72378]_  = \new_[72377]_  & \new_[72370]_ ;
  assign \new_[72382]_  = ~A168 & ~A169;
  assign \new_[72383]_  = A170 & \new_[72382]_ ;
  assign \new_[72386]_  = ~A166 & A167;
  assign \new_[72389]_  = ~A200 & ~A199;
  assign \new_[72390]_  = \new_[72389]_  & \new_[72386]_ ;
  assign \new_[72391]_  = \new_[72390]_  & \new_[72383]_ ;
  assign \new_[72395]_  = ~A269 & ~A268;
  assign \new_[72396]_  = A267 & \new_[72395]_ ;
  assign \new_[72399]_  = A299 & ~A298;
  assign \new_[72402]_  = A302 & A300;
  assign \new_[72403]_  = \new_[72402]_  & \new_[72399]_ ;
  assign \new_[72404]_  = \new_[72403]_  & \new_[72396]_ ;
  assign \new_[72408]_  = ~A168 & ~A169;
  assign \new_[72409]_  = A170 & \new_[72408]_ ;
  assign \new_[72412]_  = ~A166 & A167;
  assign \new_[72415]_  = ~A200 & ~A199;
  assign \new_[72416]_  = \new_[72415]_  & \new_[72412]_ ;
  assign \new_[72417]_  = \new_[72416]_  & \new_[72409]_ ;
  assign \new_[72421]_  = A298 & A268;
  assign \new_[72422]_  = ~A267 & \new_[72421]_ ;
  assign \new_[72425]_  = ~A300 & ~A299;
  assign \new_[72428]_  = ~A302 & ~A301;
  assign \new_[72429]_  = \new_[72428]_  & \new_[72425]_ ;
  assign \new_[72430]_  = \new_[72429]_  & \new_[72422]_ ;
  assign \new_[72434]_  = ~A168 & ~A169;
  assign \new_[72435]_  = A170 & \new_[72434]_ ;
  assign \new_[72438]_  = ~A166 & A167;
  assign \new_[72441]_  = ~A200 & ~A199;
  assign \new_[72442]_  = \new_[72441]_  & \new_[72438]_ ;
  assign \new_[72443]_  = \new_[72442]_  & \new_[72435]_ ;
  assign \new_[72447]_  = ~A298 & A268;
  assign \new_[72448]_  = ~A267 & \new_[72447]_ ;
  assign \new_[72451]_  = ~A300 & A299;
  assign \new_[72454]_  = ~A302 & ~A301;
  assign \new_[72455]_  = \new_[72454]_  & \new_[72451]_ ;
  assign \new_[72456]_  = \new_[72455]_  & \new_[72448]_ ;
  assign \new_[72460]_  = ~A168 & ~A169;
  assign \new_[72461]_  = A170 & \new_[72460]_ ;
  assign \new_[72464]_  = ~A166 & A167;
  assign \new_[72467]_  = ~A200 & ~A199;
  assign \new_[72468]_  = \new_[72467]_  & \new_[72464]_ ;
  assign \new_[72469]_  = \new_[72468]_  & \new_[72461]_ ;
  assign \new_[72473]_  = A298 & A269;
  assign \new_[72474]_  = ~A267 & \new_[72473]_ ;
  assign \new_[72477]_  = ~A300 & ~A299;
  assign \new_[72480]_  = ~A302 & ~A301;
  assign \new_[72481]_  = \new_[72480]_  & \new_[72477]_ ;
  assign \new_[72482]_  = \new_[72481]_  & \new_[72474]_ ;
  assign \new_[72486]_  = ~A168 & ~A169;
  assign \new_[72487]_  = A170 & \new_[72486]_ ;
  assign \new_[72490]_  = ~A166 & A167;
  assign \new_[72493]_  = ~A200 & ~A199;
  assign \new_[72494]_  = \new_[72493]_  & \new_[72490]_ ;
  assign \new_[72495]_  = \new_[72494]_  & \new_[72487]_ ;
  assign \new_[72499]_  = ~A298 & A269;
  assign \new_[72500]_  = ~A267 & \new_[72499]_ ;
  assign \new_[72503]_  = ~A300 & A299;
  assign \new_[72506]_  = ~A302 & ~A301;
  assign \new_[72507]_  = \new_[72506]_  & \new_[72503]_ ;
  assign \new_[72508]_  = \new_[72507]_  & \new_[72500]_ ;
  assign \new_[72512]_  = ~A168 & ~A169;
  assign \new_[72513]_  = A170 & \new_[72512]_ ;
  assign \new_[72516]_  = ~A166 & A167;
  assign \new_[72519]_  = ~A200 & ~A199;
  assign \new_[72520]_  = \new_[72519]_  & \new_[72516]_ ;
  assign \new_[72521]_  = \new_[72520]_  & \new_[72513]_ ;
  assign \new_[72525]_  = A298 & A266;
  assign \new_[72526]_  = A265 & \new_[72525]_ ;
  assign \new_[72529]_  = ~A300 & ~A299;
  assign \new_[72532]_  = ~A302 & ~A301;
  assign \new_[72533]_  = \new_[72532]_  & \new_[72529]_ ;
  assign \new_[72534]_  = \new_[72533]_  & \new_[72526]_ ;
  assign \new_[72538]_  = ~A168 & ~A169;
  assign \new_[72539]_  = A170 & \new_[72538]_ ;
  assign \new_[72542]_  = ~A166 & A167;
  assign \new_[72545]_  = ~A200 & ~A199;
  assign \new_[72546]_  = \new_[72545]_  & \new_[72542]_ ;
  assign \new_[72547]_  = \new_[72546]_  & \new_[72539]_ ;
  assign \new_[72551]_  = ~A298 & A266;
  assign \new_[72552]_  = A265 & \new_[72551]_ ;
  assign \new_[72555]_  = ~A300 & A299;
  assign \new_[72558]_  = ~A302 & ~A301;
  assign \new_[72559]_  = \new_[72558]_  & \new_[72555]_ ;
  assign \new_[72560]_  = \new_[72559]_  & \new_[72552]_ ;
  assign \new_[72564]_  = ~A168 & ~A169;
  assign \new_[72565]_  = A170 & \new_[72564]_ ;
  assign \new_[72568]_  = ~A166 & A167;
  assign \new_[72571]_  = ~A200 & ~A199;
  assign \new_[72572]_  = \new_[72571]_  & \new_[72568]_ ;
  assign \new_[72573]_  = \new_[72572]_  & \new_[72565]_ ;
  assign \new_[72577]_  = A298 & ~A266;
  assign \new_[72578]_  = ~A265 & \new_[72577]_ ;
  assign \new_[72581]_  = ~A300 & ~A299;
  assign \new_[72584]_  = ~A302 & ~A301;
  assign \new_[72585]_  = \new_[72584]_  & \new_[72581]_ ;
  assign \new_[72586]_  = \new_[72585]_  & \new_[72578]_ ;
  assign \new_[72590]_  = ~A168 & ~A169;
  assign \new_[72591]_  = A170 & \new_[72590]_ ;
  assign \new_[72594]_  = ~A166 & A167;
  assign \new_[72597]_  = ~A200 & ~A199;
  assign \new_[72598]_  = \new_[72597]_  & \new_[72594]_ ;
  assign \new_[72599]_  = \new_[72598]_  & \new_[72591]_ ;
  assign \new_[72603]_  = ~A298 & ~A266;
  assign \new_[72604]_  = ~A265 & \new_[72603]_ ;
  assign \new_[72607]_  = ~A300 & A299;
  assign \new_[72610]_  = ~A302 & ~A301;
  assign \new_[72611]_  = \new_[72610]_  & \new_[72607]_ ;
  assign \new_[72612]_  = \new_[72611]_  & \new_[72604]_ ;
  assign \new_[72616]_  = ~A168 & ~A169;
  assign \new_[72617]_  = A170 & \new_[72616]_ ;
  assign \new_[72620]_  = A166 & ~A167;
  assign \new_[72623]_  = ~A202 & A201;
  assign \new_[72624]_  = \new_[72623]_  & \new_[72620]_ ;
  assign \new_[72625]_  = \new_[72624]_  & \new_[72617]_ ;
  assign \new_[72629]_  = A268 & ~A267;
  assign \new_[72630]_  = ~A203 & \new_[72629]_ ;
  assign \new_[72633]_  = ~A299 & A298;
  assign \new_[72636]_  = A301 & A300;
  assign \new_[72637]_  = \new_[72636]_  & \new_[72633]_ ;
  assign \new_[72638]_  = \new_[72637]_  & \new_[72630]_ ;
  assign \new_[72642]_  = ~A168 & ~A169;
  assign \new_[72643]_  = A170 & \new_[72642]_ ;
  assign \new_[72646]_  = A166 & ~A167;
  assign \new_[72649]_  = ~A202 & A201;
  assign \new_[72650]_  = \new_[72649]_  & \new_[72646]_ ;
  assign \new_[72651]_  = \new_[72650]_  & \new_[72643]_ ;
  assign \new_[72655]_  = A268 & ~A267;
  assign \new_[72656]_  = ~A203 & \new_[72655]_ ;
  assign \new_[72659]_  = ~A299 & A298;
  assign \new_[72662]_  = A302 & A300;
  assign \new_[72663]_  = \new_[72662]_  & \new_[72659]_ ;
  assign \new_[72664]_  = \new_[72663]_  & \new_[72656]_ ;
  assign \new_[72668]_  = ~A168 & ~A169;
  assign \new_[72669]_  = A170 & \new_[72668]_ ;
  assign \new_[72672]_  = A166 & ~A167;
  assign \new_[72675]_  = ~A202 & A201;
  assign \new_[72676]_  = \new_[72675]_  & \new_[72672]_ ;
  assign \new_[72677]_  = \new_[72676]_  & \new_[72669]_ ;
  assign \new_[72681]_  = A268 & ~A267;
  assign \new_[72682]_  = ~A203 & \new_[72681]_ ;
  assign \new_[72685]_  = A299 & ~A298;
  assign \new_[72688]_  = A301 & A300;
  assign \new_[72689]_  = \new_[72688]_  & \new_[72685]_ ;
  assign \new_[72690]_  = \new_[72689]_  & \new_[72682]_ ;
  assign \new_[72694]_  = ~A168 & ~A169;
  assign \new_[72695]_  = A170 & \new_[72694]_ ;
  assign \new_[72698]_  = A166 & ~A167;
  assign \new_[72701]_  = ~A202 & A201;
  assign \new_[72702]_  = \new_[72701]_  & \new_[72698]_ ;
  assign \new_[72703]_  = \new_[72702]_  & \new_[72695]_ ;
  assign \new_[72707]_  = A268 & ~A267;
  assign \new_[72708]_  = ~A203 & \new_[72707]_ ;
  assign \new_[72711]_  = A299 & ~A298;
  assign \new_[72714]_  = A302 & A300;
  assign \new_[72715]_  = \new_[72714]_  & \new_[72711]_ ;
  assign \new_[72716]_  = \new_[72715]_  & \new_[72708]_ ;
  assign \new_[72720]_  = ~A168 & ~A169;
  assign \new_[72721]_  = A170 & \new_[72720]_ ;
  assign \new_[72724]_  = A166 & ~A167;
  assign \new_[72727]_  = ~A202 & A201;
  assign \new_[72728]_  = \new_[72727]_  & \new_[72724]_ ;
  assign \new_[72729]_  = \new_[72728]_  & \new_[72721]_ ;
  assign \new_[72733]_  = A269 & ~A267;
  assign \new_[72734]_  = ~A203 & \new_[72733]_ ;
  assign \new_[72737]_  = ~A299 & A298;
  assign \new_[72740]_  = A301 & A300;
  assign \new_[72741]_  = \new_[72740]_  & \new_[72737]_ ;
  assign \new_[72742]_  = \new_[72741]_  & \new_[72734]_ ;
  assign \new_[72746]_  = ~A168 & ~A169;
  assign \new_[72747]_  = A170 & \new_[72746]_ ;
  assign \new_[72750]_  = A166 & ~A167;
  assign \new_[72753]_  = ~A202 & A201;
  assign \new_[72754]_  = \new_[72753]_  & \new_[72750]_ ;
  assign \new_[72755]_  = \new_[72754]_  & \new_[72747]_ ;
  assign \new_[72759]_  = A269 & ~A267;
  assign \new_[72760]_  = ~A203 & \new_[72759]_ ;
  assign \new_[72763]_  = ~A299 & A298;
  assign \new_[72766]_  = A302 & A300;
  assign \new_[72767]_  = \new_[72766]_  & \new_[72763]_ ;
  assign \new_[72768]_  = \new_[72767]_  & \new_[72760]_ ;
  assign \new_[72772]_  = ~A168 & ~A169;
  assign \new_[72773]_  = A170 & \new_[72772]_ ;
  assign \new_[72776]_  = A166 & ~A167;
  assign \new_[72779]_  = ~A202 & A201;
  assign \new_[72780]_  = \new_[72779]_  & \new_[72776]_ ;
  assign \new_[72781]_  = \new_[72780]_  & \new_[72773]_ ;
  assign \new_[72785]_  = A269 & ~A267;
  assign \new_[72786]_  = ~A203 & \new_[72785]_ ;
  assign \new_[72789]_  = A299 & ~A298;
  assign \new_[72792]_  = A301 & A300;
  assign \new_[72793]_  = \new_[72792]_  & \new_[72789]_ ;
  assign \new_[72794]_  = \new_[72793]_  & \new_[72786]_ ;
  assign \new_[72798]_  = ~A168 & ~A169;
  assign \new_[72799]_  = A170 & \new_[72798]_ ;
  assign \new_[72802]_  = A166 & ~A167;
  assign \new_[72805]_  = ~A202 & A201;
  assign \new_[72806]_  = \new_[72805]_  & \new_[72802]_ ;
  assign \new_[72807]_  = \new_[72806]_  & \new_[72799]_ ;
  assign \new_[72811]_  = A269 & ~A267;
  assign \new_[72812]_  = ~A203 & \new_[72811]_ ;
  assign \new_[72815]_  = A299 & ~A298;
  assign \new_[72818]_  = A302 & A300;
  assign \new_[72819]_  = \new_[72818]_  & \new_[72815]_ ;
  assign \new_[72820]_  = \new_[72819]_  & \new_[72812]_ ;
  assign \new_[72824]_  = ~A168 & ~A169;
  assign \new_[72825]_  = A170 & \new_[72824]_ ;
  assign \new_[72828]_  = A166 & ~A167;
  assign \new_[72831]_  = ~A202 & A201;
  assign \new_[72832]_  = \new_[72831]_  & \new_[72828]_ ;
  assign \new_[72833]_  = \new_[72832]_  & \new_[72825]_ ;
  assign \new_[72837]_  = A266 & A265;
  assign \new_[72838]_  = ~A203 & \new_[72837]_ ;
  assign \new_[72841]_  = ~A299 & A298;
  assign \new_[72844]_  = A301 & A300;
  assign \new_[72845]_  = \new_[72844]_  & \new_[72841]_ ;
  assign \new_[72846]_  = \new_[72845]_  & \new_[72838]_ ;
  assign \new_[72850]_  = ~A168 & ~A169;
  assign \new_[72851]_  = A170 & \new_[72850]_ ;
  assign \new_[72854]_  = A166 & ~A167;
  assign \new_[72857]_  = ~A202 & A201;
  assign \new_[72858]_  = \new_[72857]_  & \new_[72854]_ ;
  assign \new_[72859]_  = \new_[72858]_  & \new_[72851]_ ;
  assign \new_[72863]_  = A266 & A265;
  assign \new_[72864]_  = ~A203 & \new_[72863]_ ;
  assign \new_[72867]_  = ~A299 & A298;
  assign \new_[72870]_  = A302 & A300;
  assign \new_[72871]_  = \new_[72870]_  & \new_[72867]_ ;
  assign \new_[72872]_  = \new_[72871]_  & \new_[72864]_ ;
  assign \new_[72876]_  = ~A168 & ~A169;
  assign \new_[72877]_  = A170 & \new_[72876]_ ;
  assign \new_[72880]_  = A166 & ~A167;
  assign \new_[72883]_  = ~A202 & A201;
  assign \new_[72884]_  = \new_[72883]_  & \new_[72880]_ ;
  assign \new_[72885]_  = \new_[72884]_  & \new_[72877]_ ;
  assign \new_[72889]_  = A266 & A265;
  assign \new_[72890]_  = ~A203 & \new_[72889]_ ;
  assign \new_[72893]_  = A299 & ~A298;
  assign \new_[72896]_  = A301 & A300;
  assign \new_[72897]_  = \new_[72896]_  & \new_[72893]_ ;
  assign \new_[72898]_  = \new_[72897]_  & \new_[72890]_ ;
  assign \new_[72902]_  = ~A168 & ~A169;
  assign \new_[72903]_  = A170 & \new_[72902]_ ;
  assign \new_[72906]_  = A166 & ~A167;
  assign \new_[72909]_  = ~A202 & A201;
  assign \new_[72910]_  = \new_[72909]_  & \new_[72906]_ ;
  assign \new_[72911]_  = \new_[72910]_  & \new_[72903]_ ;
  assign \new_[72915]_  = A266 & A265;
  assign \new_[72916]_  = ~A203 & \new_[72915]_ ;
  assign \new_[72919]_  = A299 & ~A298;
  assign \new_[72922]_  = A302 & A300;
  assign \new_[72923]_  = \new_[72922]_  & \new_[72919]_ ;
  assign \new_[72924]_  = \new_[72923]_  & \new_[72916]_ ;
  assign \new_[72928]_  = ~A168 & ~A169;
  assign \new_[72929]_  = A170 & \new_[72928]_ ;
  assign \new_[72932]_  = A166 & ~A167;
  assign \new_[72935]_  = ~A202 & A201;
  assign \new_[72936]_  = \new_[72935]_  & \new_[72932]_ ;
  assign \new_[72937]_  = \new_[72936]_  & \new_[72929]_ ;
  assign \new_[72941]_  = ~A266 & ~A265;
  assign \new_[72942]_  = ~A203 & \new_[72941]_ ;
  assign \new_[72945]_  = ~A299 & A298;
  assign \new_[72948]_  = A301 & A300;
  assign \new_[72949]_  = \new_[72948]_  & \new_[72945]_ ;
  assign \new_[72950]_  = \new_[72949]_  & \new_[72942]_ ;
  assign \new_[72954]_  = ~A168 & ~A169;
  assign \new_[72955]_  = A170 & \new_[72954]_ ;
  assign \new_[72958]_  = A166 & ~A167;
  assign \new_[72961]_  = ~A202 & A201;
  assign \new_[72962]_  = \new_[72961]_  & \new_[72958]_ ;
  assign \new_[72963]_  = \new_[72962]_  & \new_[72955]_ ;
  assign \new_[72967]_  = ~A266 & ~A265;
  assign \new_[72968]_  = ~A203 & \new_[72967]_ ;
  assign \new_[72971]_  = ~A299 & A298;
  assign \new_[72974]_  = A302 & A300;
  assign \new_[72975]_  = \new_[72974]_  & \new_[72971]_ ;
  assign \new_[72976]_  = \new_[72975]_  & \new_[72968]_ ;
  assign \new_[72980]_  = ~A168 & ~A169;
  assign \new_[72981]_  = A170 & \new_[72980]_ ;
  assign \new_[72984]_  = A166 & ~A167;
  assign \new_[72987]_  = ~A202 & A201;
  assign \new_[72988]_  = \new_[72987]_  & \new_[72984]_ ;
  assign \new_[72989]_  = \new_[72988]_  & \new_[72981]_ ;
  assign \new_[72993]_  = ~A266 & ~A265;
  assign \new_[72994]_  = ~A203 & \new_[72993]_ ;
  assign \new_[72997]_  = A299 & ~A298;
  assign \new_[73000]_  = A301 & A300;
  assign \new_[73001]_  = \new_[73000]_  & \new_[72997]_ ;
  assign \new_[73002]_  = \new_[73001]_  & \new_[72994]_ ;
  assign \new_[73006]_  = ~A168 & ~A169;
  assign \new_[73007]_  = A170 & \new_[73006]_ ;
  assign \new_[73010]_  = A166 & ~A167;
  assign \new_[73013]_  = ~A202 & A201;
  assign \new_[73014]_  = \new_[73013]_  & \new_[73010]_ ;
  assign \new_[73015]_  = \new_[73014]_  & \new_[73007]_ ;
  assign \new_[73019]_  = ~A266 & ~A265;
  assign \new_[73020]_  = ~A203 & \new_[73019]_ ;
  assign \new_[73023]_  = A299 & ~A298;
  assign \new_[73026]_  = A302 & A300;
  assign \new_[73027]_  = \new_[73026]_  & \new_[73023]_ ;
  assign \new_[73028]_  = \new_[73027]_  & \new_[73020]_ ;
  assign \new_[73032]_  = ~A168 & ~A169;
  assign \new_[73033]_  = A170 & \new_[73032]_ ;
  assign \new_[73036]_  = A166 & ~A167;
  assign \new_[73039]_  = A202 & ~A201;
  assign \new_[73040]_  = \new_[73039]_  & \new_[73036]_ ;
  assign \new_[73041]_  = \new_[73040]_  & \new_[73033]_ ;
  assign \new_[73045]_  = ~A269 & ~A268;
  assign \new_[73046]_  = A267 & \new_[73045]_ ;
  assign \new_[73049]_  = ~A299 & A298;
  assign \new_[73052]_  = A301 & A300;
  assign \new_[73053]_  = \new_[73052]_  & \new_[73049]_ ;
  assign \new_[73054]_  = \new_[73053]_  & \new_[73046]_ ;
  assign \new_[73058]_  = ~A168 & ~A169;
  assign \new_[73059]_  = A170 & \new_[73058]_ ;
  assign \new_[73062]_  = A166 & ~A167;
  assign \new_[73065]_  = A202 & ~A201;
  assign \new_[73066]_  = \new_[73065]_  & \new_[73062]_ ;
  assign \new_[73067]_  = \new_[73066]_  & \new_[73059]_ ;
  assign \new_[73071]_  = ~A269 & ~A268;
  assign \new_[73072]_  = A267 & \new_[73071]_ ;
  assign \new_[73075]_  = ~A299 & A298;
  assign \new_[73078]_  = A302 & A300;
  assign \new_[73079]_  = \new_[73078]_  & \new_[73075]_ ;
  assign \new_[73080]_  = \new_[73079]_  & \new_[73072]_ ;
  assign \new_[73084]_  = ~A168 & ~A169;
  assign \new_[73085]_  = A170 & \new_[73084]_ ;
  assign \new_[73088]_  = A166 & ~A167;
  assign \new_[73091]_  = A202 & ~A201;
  assign \new_[73092]_  = \new_[73091]_  & \new_[73088]_ ;
  assign \new_[73093]_  = \new_[73092]_  & \new_[73085]_ ;
  assign \new_[73097]_  = ~A269 & ~A268;
  assign \new_[73098]_  = A267 & \new_[73097]_ ;
  assign \new_[73101]_  = A299 & ~A298;
  assign \new_[73104]_  = A301 & A300;
  assign \new_[73105]_  = \new_[73104]_  & \new_[73101]_ ;
  assign \new_[73106]_  = \new_[73105]_  & \new_[73098]_ ;
  assign \new_[73110]_  = ~A168 & ~A169;
  assign \new_[73111]_  = A170 & \new_[73110]_ ;
  assign \new_[73114]_  = A166 & ~A167;
  assign \new_[73117]_  = A202 & ~A201;
  assign \new_[73118]_  = \new_[73117]_  & \new_[73114]_ ;
  assign \new_[73119]_  = \new_[73118]_  & \new_[73111]_ ;
  assign \new_[73123]_  = ~A269 & ~A268;
  assign \new_[73124]_  = A267 & \new_[73123]_ ;
  assign \new_[73127]_  = A299 & ~A298;
  assign \new_[73130]_  = A302 & A300;
  assign \new_[73131]_  = \new_[73130]_  & \new_[73127]_ ;
  assign \new_[73132]_  = \new_[73131]_  & \new_[73124]_ ;
  assign \new_[73136]_  = ~A168 & ~A169;
  assign \new_[73137]_  = A170 & \new_[73136]_ ;
  assign \new_[73140]_  = A166 & ~A167;
  assign \new_[73143]_  = A202 & ~A201;
  assign \new_[73144]_  = \new_[73143]_  & \new_[73140]_ ;
  assign \new_[73145]_  = \new_[73144]_  & \new_[73137]_ ;
  assign \new_[73149]_  = A298 & A268;
  assign \new_[73150]_  = ~A267 & \new_[73149]_ ;
  assign \new_[73153]_  = ~A300 & ~A299;
  assign \new_[73156]_  = ~A302 & ~A301;
  assign \new_[73157]_  = \new_[73156]_  & \new_[73153]_ ;
  assign \new_[73158]_  = \new_[73157]_  & \new_[73150]_ ;
  assign \new_[73162]_  = ~A168 & ~A169;
  assign \new_[73163]_  = A170 & \new_[73162]_ ;
  assign \new_[73166]_  = A166 & ~A167;
  assign \new_[73169]_  = A202 & ~A201;
  assign \new_[73170]_  = \new_[73169]_  & \new_[73166]_ ;
  assign \new_[73171]_  = \new_[73170]_  & \new_[73163]_ ;
  assign \new_[73175]_  = ~A298 & A268;
  assign \new_[73176]_  = ~A267 & \new_[73175]_ ;
  assign \new_[73179]_  = ~A300 & A299;
  assign \new_[73182]_  = ~A302 & ~A301;
  assign \new_[73183]_  = \new_[73182]_  & \new_[73179]_ ;
  assign \new_[73184]_  = \new_[73183]_  & \new_[73176]_ ;
  assign \new_[73188]_  = ~A168 & ~A169;
  assign \new_[73189]_  = A170 & \new_[73188]_ ;
  assign \new_[73192]_  = A166 & ~A167;
  assign \new_[73195]_  = A202 & ~A201;
  assign \new_[73196]_  = \new_[73195]_  & \new_[73192]_ ;
  assign \new_[73197]_  = \new_[73196]_  & \new_[73189]_ ;
  assign \new_[73201]_  = A298 & A269;
  assign \new_[73202]_  = ~A267 & \new_[73201]_ ;
  assign \new_[73205]_  = ~A300 & ~A299;
  assign \new_[73208]_  = ~A302 & ~A301;
  assign \new_[73209]_  = \new_[73208]_  & \new_[73205]_ ;
  assign \new_[73210]_  = \new_[73209]_  & \new_[73202]_ ;
  assign \new_[73214]_  = ~A168 & ~A169;
  assign \new_[73215]_  = A170 & \new_[73214]_ ;
  assign \new_[73218]_  = A166 & ~A167;
  assign \new_[73221]_  = A202 & ~A201;
  assign \new_[73222]_  = \new_[73221]_  & \new_[73218]_ ;
  assign \new_[73223]_  = \new_[73222]_  & \new_[73215]_ ;
  assign \new_[73227]_  = ~A298 & A269;
  assign \new_[73228]_  = ~A267 & \new_[73227]_ ;
  assign \new_[73231]_  = ~A300 & A299;
  assign \new_[73234]_  = ~A302 & ~A301;
  assign \new_[73235]_  = \new_[73234]_  & \new_[73231]_ ;
  assign \new_[73236]_  = \new_[73235]_  & \new_[73228]_ ;
  assign \new_[73240]_  = ~A168 & ~A169;
  assign \new_[73241]_  = A170 & \new_[73240]_ ;
  assign \new_[73244]_  = A166 & ~A167;
  assign \new_[73247]_  = A202 & ~A201;
  assign \new_[73248]_  = \new_[73247]_  & \new_[73244]_ ;
  assign \new_[73249]_  = \new_[73248]_  & \new_[73241]_ ;
  assign \new_[73253]_  = A298 & A266;
  assign \new_[73254]_  = A265 & \new_[73253]_ ;
  assign \new_[73257]_  = ~A300 & ~A299;
  assign \new_[73260]_  = ~A302 & ~A301;
  assign \new_[73261]_  = \new_[73260]_  & \new_[73257]_ ;
  assign \new_[73262]_  = \new_[73261]_  & \new_[73254]_ ;
  assign \new_[73266]_  = ~A168 & ~A169;
  assign \new_[73267]_  = A170 & \new_[73266]_ ;
  assign \new_[73270]_  = A166 & ~A167;
  assign \new_[73273]_  = A202 & ~A201;
  assign \new_[73274]_  = \new_[73273]_  & \new_[73270]_ ;
  assign \new_[73275]_  = \new_[73274]_  & \new_[73267]_ ;
  assign \new_[73279]_  = ~A298 & A266;
  assign \new_[73280]_  = A265 & \new_[73279]_ ;
  assign \new_[73283]_  = ~A300 & A299;
  assign \new_[73286]_  = ~A302 & ~A301;
  assign \new_[73287]_  = \new_[73286]_  & \new_[73283]_ ;
  assign \new_[73288]_  = \new_[73287]_  & \new_[73280]_ ;
  assign \new_[73292]_  = ~A168 & ~A169;
  assign \new_[73293]_  = A170 & \new_[73292]_ ;
  assign \new_[73296]_  = A166 & ~A167;
  assign \new_[73299]_  = A202 & ~A201;
  assign \new_[73300]_  = \new_[73299]_  & \new_[73296]_ ;
  assign \new_[73301]_  = \new_[73300]_  & \new_[73293]_ ;
  assign \new_[73305]_  = A298 & ~A266;
  assign \new_[73306]_  = ~A265 & \new_[73305]_ ;
  assign \new_[73309]_  = ~A300 & ~A299;
  assign \new_[73312]_  = ~A302 & ~A301;
  assign \new_[73313]_  = \new_[73312]_  & \new_[73309]_ ;
  assign \new_[73314]_  = \new_[73313]_  & \new_[73306]_ ;
  assign \new_[73318]_  = ~A168 & ~A169;
  assign \new_[73319]_  = A170 & \new_[73318]_ ;
  assign \new_[73322]_  = A166 & ~A167;
  assign \new_[73325]_  = A202 & ~A201;
  assign \new_[73326]_  = \new_[73325]_  & \new_[73322]_ ;
  assign \new_[73327]_  = \new_[73326]_  & \new_[73319]_ ;
  assign \new_[73331]_  = ~A298 & ~A266;
  assign \new_[73332]_  = ~A265 & \new_[73331]_ ;
  assign \new_[73335]_  = ~A300 & A299;
  assign \new_[73338]_  = ~A302 & ~A301;
  assign \new_[73339]_  = \new_[73338]_  & \new_[73335]_ ;
  assign \new_[73340]_  = \new_[73339]_  & \new_[73332]_ ;
  assign \new_[73344]_  = ~A168 & ~A169;
  assign \new_[73345]_  = A170 & \new_[73344]_ ;
  assign \new_[73348]_  = A166 & ~A167;
  assign \new_[73351]_  = A203 & ~A201;
  assign \new_[73352]_  = \new_[73351]_  & \new_[73348]_ ;
  assign \new_[73353]_  = \new_[73352]_  & \new_[73345]_ ;
  assign \new_[73357]_  = ~A269 & ~A268;
  assign \new_[73358]_  = A267 & \new_[73357]_ ;
  assign \new_[73361]_  = ~A299 & A298;
  assign \new_[73364]_  = A301 & A300;
  assign \new_[73365]_  = \new_[73364]_  & \new_[73361]_ ;
  assign \new_[73366]_  = \new_[73365]_  & \new_[73358]_ ;
  assign \new_[73370]_  = ~A168 & ~A169;
  assign \new_[73371]_  = A170 & \new_[73370]_ ;
  assign \new_[73374]_  = A166 & ~A167;
  assign \new_[73377]_  = A203 & ~A201;
  assign \new_[73378]_  = \new_[73377]_  & \new_[73374]_ ;
  assign \new_[73379]_  = \new_[73378]_  & \new_[73371]_ ;
  assign \new_[73383]_  = ~A269 & ~A268;
  assign \new_[73384]_  = A267 & \new_[73383]_ ;
  assign \new_[73387]_  = ~A299 & A298;
  assign \new_[73390]_  = A302 & A300;
  assign \new_[73391]_  = \new_[73390]_  & \new_[73387]_ ;
  assign \new_[73392]_  = \new_[73391]_  & \new_[73384]_ ;
  assign \new_[73396]_  = ~A168 & ~A169;
  assign \new_[73397]_  = A170 & \new_[73396]_ ;
  assign \new_[73400]_  = A166 & ~A167;
  assign \new_[73403]_  = A203 & ~A201;
  assign \new_[73404]_  = \new_[73403]_  & \new_[73400]_ ;
  assign \new_[73405]_  = \new_[73404]_  & \new_[73397]_ ;
  assign \new_[73409]_  = ~A269 & ~A268;
  assign \new_[73410]_  = A267 & \new_[73409]_ ;
  assign \new_[73413]_  = A299 & ~A298;
  assign \new_[73416]_  = A301 & A300;
  assign \new_[73417]_  = \new_[73416]_  & \new_[73413]_ ;
  assign \new_[73418]_  = \new_[73417]_  & \new_[73410]_ ;
  assign \new_[73422]_  = ~A168 & ~A169;
  assign \new_[73423]_  = A170 & \new_[73422]_ ;
  assign \new_[73426]_  = A166 & ~A167;
  assign \new_[73429]_  = A203 & ~A201;
  assign \new_[73430]_  = \new_[73429]_  & \new_[73426]_ ;
  assign \new_[73431]_  = \new_[73430]_  & \new_[73423]_ ;
  assign \new_[73435]_  = ~A269 & ~A268;
  assign \new_[73436]_  = A267 & \new_[73435]_ ;
  assign \new_[73439]_  = A299 & ~A298;
  assign \new_[73442]_  = A302 & A300;
  assign \new_[73443]_  = \new_[73442]_  & \new_[73439]_ ;
  assign \new_[73444]_  = \new_[73443]_  & \new_[73436]_ ;
  assign \new_[73448]_  = ~A168 & ~A169;
  assign \new_[73449]_  = A170 & \new_[73448]_ ;
  assign \new_[73452]_  = A166 & ~A167;
  assign \new_[73455]_  = A203 & ~A201;
  assign \new_[73456]_  = \new_[73455]_  & \new_[73452]_ ;
  assign \new_[73457]_  = \new_[73456]_  & \new_[73449]_ ;
  assign \new_[73461]_  = A298 & A268;
  assign \new_[73462]_  = ~A267 & \new_[73461]_ ;
  assign \new_[73465]_  = ~A300 & ~A299;
  assign \new_[73468]_  = ~A302 & ~A301;
  assign \new_[73469]_  = \new_[73468]_  & \new_[73465]_ ;
  assign \new_[73470]_  = \new_[73469]_  & \new_[73462]_ ;
  assign \new_[73474]_  = ~A168 & ~A169;
  assign \new_[73475]_  = A170 & \new_[73474]_ ;
  assign \new_[73478]_  = A166 & ~A167;
  assign \new_[73481]_  = A203 & ~A201;
  assign \new_[73482]_  = \new_[73481]_  & \new_[73478]_ ;
  assign \new_[73483]_  = \new_[73482]_  & \new_[73475]_ ;
  assign \new_[73487]_  = ~A298 & A268;
  assign \new_[73488]_  = ~A267 & \new_[73487]_ ;
  assign \new_[73491]_  = ~A300 & A299;
  assign \new_[73494]_  = ~A302 & ~A301;
  assign \new_[73495]_  = \new_[73494]_  & \new_[73491]_ ;
  assign \new_[73496]_  = \new_[73495]_  & \new_[73488]_ ;
  assign \new_[73500]_  = ~A168 & ~A169;
  assign \new_[73501]_  = A170 & \new_[73500]_ ;
  assign \new_[73504]_  = A166 & ~A167;
  assign \new_[73507]_  = A203 & ~A201;
  assign \new_[73508]_  = \new_[73507]_  & \new_[73504]_ ;
  assign \new_[73509]_  = \new_[73508]_  & \new_[73501]_ ;
  assign \new_[73513]_  = A298 & A269;
  assign \new_[73514]_  = ~A267 & \new_[73513]_ ;
  assign \new_[73517]_  = ~A300 & ~A299;
  assign \new_[73520]_  = ~A302 & ~A301;
  assign \new_[73521]_  = \new_[73520]_  & \new_[73517]_ ;
  assign \new_[73522]_  = \new_[73521]_  & \new_[73514]_ ;
  assign \new_[73526]_  = ~A168 & ~A169;
  assign \new_[73527]_  = A170 & \new_[73526]_ ;
  assign \new_[73530]_  = A166 & ~A167;
  assign \new_[73533]_  = A203 & ~A201;
  assign \new_[73534]_  = \new_[73533]_  & \new_[73530]_ ;
  assign \new_[73535]_  = \new_[73534]_  & \new_[73527]_ ;
  assign \new_[73539]_  = ~A298 & A269;
  assign \new_[73540]_  = ~A267 & \new_[73539]_ ;
  assign \new_[73543]_  = ~A300 & A299;
  assign \new_[73546]_  = ~A302 & ~A301;
  assign \new_[73547]_  = \new_[73546]_  & \new_[73543]_ ;
  assign \new_[73548]_  = \new_[73547]_  & \new_[73540]_ ;
  assign \new_[73552]_  = ~A168 & ~A169;
  assign \new_[73553]_  = A170 & \new_[73552]_ ;
  assign \new_[73556]_  = A166 & ~A167;
  assign \new_[73559]_  = A203 & ~A201;
  assign \new_[73560]_  = \new_[73559]_  & \new_[73556]_ ;
  assign \new_[73561]_  = \new_[73560]_  & \new_[73553]_ ;
  assign \new_[73565]_  = A298 & A266;
  assign \new_[73566]_  = A265 & \new_[73565]_ ;
  assign \new_[73569]_  = ~A300 & ~A299;
  assign \new_[73572]_  = ~A302 & ~A301;
  assign \new_[73573]_  = \new_[73572]_  & \new_[73569]_ ;
  assign \new_[73574]_  = \new_[73573]_  & \new_[73566]_ ;
  assign \new_[73578]_  = ~A168 & ~A169;
  assign \new_[73579]_  = A170 & \new_[73578]_ ;
  assign \new_[73582]_  = A166 & ~A167;
  assign \new_[73585]_  = A203 & ~A201;
  assign \new_[73586]_  = \new_[73585]_  & \new_[73582]_ ;
  assign \new_[73587]_  = \new_[73586]_  & \new_[73579]_ ;
  assign \new_[73591]_  = ~A298 & A266;
  assign \new_[73592]_  = A265 & \new_[73591]_ ;
  assign \new_[73595]_  = ~A300 & A299;
  assign \new_[73598]_  = ~A302 & ~A301;
  assign \new_[73599]_  = \new_[73598]_  & \new_[73595]_ ;
  assign \new_[73600]_  = \new_[73599]_  & \new_[73592]_ ;
  assign \new_[73604]_  = ~A168 & ~A169;
  assign \new_[73605]_  = A170 & \new_[73604]_ ;
  assign \new_[73608]_  = A166 & ~A167;
  assign \new_[73611]_  = A203 & ~A201;
  assign \new_[73612]_  = \new_[73611]_  & \new_[73608]_ ;
  assign \new_[73613]_  = \new_[73612]_  & \new_[73605]_ ;
  assign \new_[73617]_  = A298 & ~A266;
  assign \new_[73618]_  = ~A265 & \new_[73617]_ ;
  assign \new_[73621]_  = ~A300 & ~A299;
  assign \new_[73624]_  = ~A302 & ~A301;
  assign \new_[73625]_  = \new_[73624]_  & \new_[73621]_ ;
  assign \new_[73626]_  = \new_[73625]_  & \new_[73618]_ ;
  assign \new_[73630]_  = ~A168 & ~A169;
  assign \new_[73631]_  = A170 & \new_[73630]_ ;
  assign \new_[73634]_  = A166 & ~A167;
  assign \new_[73637]_  = A203 & ~A201;
  assign \new_[73638]_  = \new_[73637]_  & \new_[73634]_ ;
  assign \new_[73639]_  = \new_[73638]_  & \new_[73631]_ ;
  assign \new_[73643]_  = ~A298 & ~A266;
  assign \new_[73644]_  = ~A265 & \new_[73643]_ ;
  assign \new_[73647]_  = ~A300 & A299;
  assign \new_[73650]_  = ~A302 & ~A301;
  assign \new_[73651]_  = \new_[73650]_  & \new_[73647]_ ;
  assign \new_[73652]_  = \new_[73651]_  & \new_[73644]_ ;
  assign \new_[73656]_  = ~A168 & ~A169;
  assign \new_[73657]_  = A170 & \new_[73656]_ ;
  assign \new_[73660]_  = A166 & ~A167;
  assign \new_[73663]_  = A200 & A199;
  assign \new_[73664]_  = \new_[73663]_  & \new_[73660]_ ;
  assign \new_[73665]_  = \new_[73664]_  & \new_[73657]_ ;
  assign \new_[73669]_  = ~A269 & ~A268;
  assign \new_[73670]_  = A267 & \new_[73669]_ ;
  assign \new_[73673]_  = ~A299 & A298;
  assign \new_[73676]_  = A301 & A300;
  assign \new_[73677]_  = \new_[73676]_  & \new_[73673]_ ;
  assign \new_[73678]_  = \new_[73677]_  & \new_[73670]_ ;
  assign \new_[73682]_  = ~A168 & ~A169;
  assign \new_[73683]_  = A170 & \new_[73682]_ ;
  assign \new_[73686]_  = A166 & ~A167;
  assign \new_[73689]_  = A200 & A199;
  assign \new_[73690]_  = \new_[73689]_  & \new_[73686]_ ;
  assign \new_[73691]_  = \new_[73690]_  & \new_[73683]_ ;
  assign \new_[73695]_  = ~A269 & ~A268;
  assign \new_[73696]_  = A267 & \new_[73695]_ ;
  assign \new_[73699]_  = ~A299 & A298;
  assign \new_[73702]_  = A302 & A300;
  assign \new_[73703]_  = \new_[73702]_  & \new_[73699]_ ;
  assign \new_[73704]_  = \new_[73703]_  & \new_[73696]_ ;
  assign \new_[73708]_  = ~A168 & ~A169;
  assign \new_[73709]_  = A170 & \new_[73708]_ ;
  assign \new_[73712]_  = A166 & ~A167;
  assign \new_[73715]_  = A200 & A199;
  assign \new_[73716]_  = \new_[73715]_  & \new_[73712]_ ;
  assign \new_[73717]_  = \new_[73716]_  & \new_[73709]_ ;
  assign \new_[73721]_  = ~A269 & ~A268;
  assign \new_[73722]_  = A267 & \new_[73721]_ ;
  assign \new_[73725]_  = A299 & ~A298;
  assign \new_[73728]_  = A301 & A300;
  assign \new_[73729]_  = \new_[73728]_  & \new_[73725]_ ;
  assign \new_[73730]_  = \new_[73729]_  & \new_[73722]_ ;
  assign \new_[73734]_  = ~A168 & ~A169;
  assign \new_[73735]_  = A170 & \new_[73734]_ ;
  assign \new_[73738]_  = A166 & ~A167;
  assign \new_[73741]_  = A200 & A199;
  assign \new_[73742]_  = \new_[73741]_  & \new_[73738]_ ;
  assign \new_[73743]_  = \new_[73742]_  & \new_[73735]_ ;
  assign \new_[73747]_  = ~A269 & ~A268;
  assign \new_[73748]_  = A267 & \new_[73747]_ ;
  assign \new_[73751]_  = A299 & ~A298;
  assign \new_[73754]_  = A302 & A300;
  assign \new_[73755]_  = \new_[73754]_  & \new_[73751]_ ;
  assign \new_[73756]_  = \new_[73755]_  & \new_[73748]_ ;
  assign \new_[73760]_  = ~A168 & ~A169;
  assign \new_[73761]_  = A170 & \new_[73760]_ ;
  assign \new_[73764]_  = A166 & ~A167;
  assign \new_[73767]_  = A200 & A199;
  assign \new_[73768]_  = \new_[73767]_  & \new_[73764]_ ;
  assign \new_[73769]_  = \new_[73768]_  & \new_[73761]_ ;
  assign \new_[73773]_  = A298 & A268;
  assign \new_[73774]_  = ~A267 & \new_[73773]_ ;
  assign \new_[73777]_  = ~A300 & ~A299;
  assign \new_[73780]_  = ~A302 & ~A301;
  assign \new_[73781]_  = \new_[73780]_  & \new_[73777]_ ;
  assign \new_[73782]_  = \new_[73781]_  & \new_[73774]_ ;
  assign \new_[73786]_  = ~A168 & ~A169;
  assign \new_[73787]_  = A170 & \new_[73786]_ ;
  assign \new_[73790]_  = A166 & ~A167;
  assign \new_[73793]_  = A200 & A199;
  assign \new_[73794]_  = \new_[73793]_  & \new_[73790]_ ;
  assign \new_[73795]_  = \new_[73794]_  & \new_[73787]_ ;
  assign \new_[73799]_  = ~A298 & A268;
  assign \new_[73800]_  = ~A267 & \new_[73799]_ ;
  assign \new_[73803]_  = ~A300 & A299;
  assign \new_[73806]_  = ~A302 & ~A301;
  assign \new_[73807]_  = \new_[73806]_  & \new_[73803]_ ;
  assign \new_[73808]_  = \new_[73807]_  & \new_[73800]_ ;
  assign \new_[73812]_  = ~A168 & ~A169;
  assign \new_[73813]_  = A170 & \new_[73812]_ ;
  assign \new_[73816]_  = A166 & ~A167;
  assign \new_[73819]_  = A200 & A199;
  assign \new_[73820]_  = \new_[73819]_  & \new_[73816]_ ;
  assign \new_[73821]_  = \new_[73820]_  & \new_[73813]_ ;
  assign \new_[73825]_  = A298 & A269;
  assign \new_[73826]_  = ~A267 & \new_[73825]_ ;
  assign \new_[73829]_  = ~A300 & ~A299;
  assign \new_[73832]_  = ~A302 & ~A301;
  assign \new_[73833]_  = \new_[73832]_  & \new_[73829]_ ;
  assign \new_[73834]_  = \new_[73833]_  & \new_[73826]_ ;
  assign \new_[73838]_  = ~A168 & ~A169;
  assign \new_[73839]_  = A170 & \new_[73838]_ ;
  assign \new_[73842]_  = A166 & ~A167;
  assign \new_[73845]_  = A200 & A199;
  assign \new_[73846]_  = \new_[73845]_  & \new_[73842]_ ;
  assign \new_[73847]_  = \new_[73846]_  & \new_[73839]_ ;
  assign \new_[73851]_  = ~A298 & A269;
  assign \new_[73852]_  = ~A267 & \new_[73851]_ ;
  assign \new_[73855]_  = ~A300 & A299;
  assign \new_[73858]_  = ~A302 & ~A301;
  assign \new_[73859]_  = \new_[73858]_  & \new_[73855]_ ;
  assign \new_[73860]_  = \new_[73859]_  & \new_[73852]_ ;
  assign \new_[73864]_  = ~A168 & ~A169;
  assign \new_[73865]_  = A170 & \new_[73864]_ ;
  assign \new_[73868]_  = A166 & ~A167;
  assign \new_[73871]_  = A200 & A199;
  assign \new_[73872]_  = \new_[73871]_  & \new_[73868]_ ;
  assign \new_[73873]_  = \new_[73872]_  & \new_[73865]_ ;
  assign \new_[73877]_  = A298 & A266;
  assign \new_[73878]_  = A265 & \new_[73877]_ ;
  assign \new_[73881]_  = ~A300 & ~A299;
  assign \new_[73884]_  = ~A302 & ~A301;
  assign \new_[73885]_  = \new_[73884]_  & \new_[73881]_ ;
  assign \new_[73886]_  = \new_[73885]_  & \new_[73878]_ ;
  assign \new_[73890]_  = ~A168 & ~A169;
  assign \new_[73891]_  = A170 & \new_[73890]_ ;
  assign \new_[73894]_  = A166 & ~A167;
  assign \new_[73897]_  = A200 & A199;
  assign \new_[73898]_  = \new_[73897]_  & \new_[73894]_ ;
  assign \new_[73899]_  = \new_[73898]_  & \new_[73891]_ ;
  assign \new_[73903]_  = ~A298 & A266;
  assign \new_[73904]_  = A265 & \new_[73903]_ ;
  assign \new_[73907]_  = ~A300 & A299;
  assign \new_[73910]_  = ~A302 & ~A301;
  assign \new_[73911]_  = \new_[73910]_  & \new_[73907]_ ;
  assign \new_[73912]_  = \new_[73911]_  & \new_[73904]_ ;
  assign \new_[73916]_  = ~A168 & ~A169;
  assign \new_[73917]_  = A170 & \new_[73916]_ ;
  assign \new_[73920]_  = A166 & ~A167;
  assign \new_[73923]_  = A200 & A199;
  assign \new_[73924]_  = \new_[73923]_  & \new_[73920]_ ;
  assign \new_[73925]_  = \new_[73924]_  & \new_[73917]_ ;
  assign \new_[73929]_  = A298 & ~A266;
  assign \new_[73930]_  = ~A265 & \new_[73929]_ ;
  assign \new_[73933]_  = ~A300 & ~A299;
  assign \new_[73936]_  = ~A302 & ~A301;
  assign \new_[73937]_  = \new_[73936]_  & \new_[73933]_ ;
  assign \new_[73938]_  = \new_[73937]_  & \new_[73930]_ ;
  assign \new_[73942]_  = ~A168 & ~A169;
  assign \new_[73943]_  = A170 & \new_[73942]_ ;
  assign \new_[73946]_  = A166 & ~A167;
  assign \new_[73949]_  = A200 & A199;
  assign \new_[73950]_  = \new_[73949]_  & \new_[73946]_ ;
  assign \new_[73951]_  = \new_[73950]_  & \new_[73943]_ ;
  assign \new_[73955]_  = ~A298 & ~A266;
  assign \new_[73956]_  = ~A265 & \new_[73955]_ ;
  assign \new_[73959]_  = ~A300 & A299;
  assign \new_[73962]_  = ~A302 & ~A301;
  assign \new_[73963]_  = \new_[73962]_  & \new_[73959]_ ;
  assign \new_[73964]_  = \new_[73963]_  & \new_[73956]_ ;
  assign \new_[73968]_  = ~A168 & ~A169;
  assign \new_[73969]_  = A170 & \new_[73968]_ ;
  assign \new_[73972]_  = A166 & ~A167;
  assign \new_[73975]_  = ~A200 & ~A199;
  assign \new_[73976]_  = \new_[73975]_  & \new_[73972]_ ;
  assign \new_[73977]_  = \new_[73976]_  & \new_[73969]_ ;
  assign \new_[73981]_  = ~A269 & ~A268;
  assign \new_[73982]_  = A267 & \new_[73981]_ ;
  assign \new_[73985]_  = ~A299 & A298;
  assign \new_[73988]_  = A301 & A300;
  assign \new_[73989]_  = \new_[73988]_  & \new_[73985]_ ;
  assign \new_[73990]_  = \new_[73989]_  & \new_[73982]_ ;
  assign \new_[73994]_  = ~A168 & ~A169;
  assign \new_[73995]_  = A170 & \new_[73994]_ ;
  assign \new_[73998]_  = A166 & ~A167;
  assign \new_[74001]_  = ~A200 & ~A199;
  assign \new_[74002]_  = \new_[74001]_  & \new_[73998]_ ;
  assign \new_[74003]_  = \new_[74002]_  & \new_[73995]_ ;
  assign \new_[74007]_  = ~A269 & ~A268;
  assign \new_[74008]_  = A267 & \new_[74007]_ ;
  assign \new_[74011]_  = ~A299 & A298;
  assign \new_[74014]_  = A302 & A300;
  assign \new_[74015]_  = \new_[74014]_  & \new_[74011]_ ;
  assign \new_[74016]_  = \new_[74015]_  & \new_[74008]_ ;
  assign \new_[74020]_  = ~A168 & ~A169;
  assign \new_[74021]_  = A170 & \new_[74020]_ ;
  assign \new_[74024]_  = A166 & ~A167;
  assign \new_[74027]_  = ~A200 & ~A199;
  assign \new_[74028]_  = \new_[74027]_  & \new_[74024]_ ;
  assign \new_[74029]_  = \new_[74028]_  & \new_[74021]_ ;
  assign \new_[74033]_  = ~A269 & ~A268;
  assign \new_[74034]_  = A267 & \new_[74033]_ ;
  assign \new_[74037]_  = A299 & ~A298;
  assign \new_[74040]_  = A301 & A300;
  assign \new_[74041]_  = \new_[74040]_  & \new_[74037]_ ;
  assign \new_[74042]_  = \new_[74041]_  & \new_[74034]_ ;
  assign \new_[74046]_  = ~A168 & ~A169;
  assign \new_[74047]_  = A170 & \new_[74046]_ ;
  assign \new_[74050]_  = A166 & ~A167;
  assign \new_[74053]_  = ~A200 & ~A199;
  assign \new_[74054]_  = \new_[74053]_  & \new_[74050]_ ;
  assign \new_[74055]_  = \new_[74054]_  & \new_[74047]_ ;
  assign \new_[74059]_  = ~A269 & ~A268;
  assign \new_[74060]_  = A267 & \new_[74059]_ ;
  assign \new_[74063]_  = A299 & ~A298;
  assign \new_[74066]_  = A302 & A300;
  assign \new_[74067]_  = \new_[74066]_  & \new_[74063]_ ;
  assign \new_[74068]_  = \new_[74067]_  & \new_[74060]_ ;
  assign \new_[74072]_  = ~A168 & ~A169;
  assign \new_[74073]_  = A170 & \new_[74072]_ ;
  assign \new_[74076]_  = A166 & ~A167;
  assign \new_[74079]_  = ~A200 & ~A199;
  assign \new_[74080]_  = \new_[74079]_  & \new_[74076]_ ;
  assign \new_[74081]_  = \new_[74080]_  & \new_[74073]_ ;
  assign \new_[74085]_  = A298 & A268;
  assign \new_[74086]_  = ~A267 & \new_[74085]_ ;
  assign \new_[74089]_  = ~A300 & ~A299;
  assign \new_[74092]_  = ~A302 & ~A301;
  assign \new_[74093]_  = \new_[74092]_  & \new_[74089]_ ;
  assign \new_[74094]_  = \new_[74093]_  & \new_[74086]_ ;
  assign \new_[74098]_  = ~A168 & ~A169;
  assign \new_[74099]_  = A170 & \new_[74098]_ ;
  assign \new_[74102]_  = A166 & ~A167;
  assign \new_[74105]_  = ~A200 & ~A199;
  assign \new_[74106]_  = \new_[74105]_  & \new_[74102]_ ;
  assign \new_[74107]_  = \new_[74106]_  & \new_[74099]_ ;
  assign \new_[74111]_  = ~A298 & A268;
  assign \new_[74112]_  = ~A267 & \new_[74111]_ ;
  assign \new_[74115]_  = ~A300 & A299;
  assign \new_[74118]_  = ~A302 & ~A301;
  assign \new_[74119]_  = \new_[74118]_  & \new_[74115]_ ;
  assign \new_[74120]_  = \new_[74119]_  & \new_[74112]_ ;
  assign \new_[74124]_  = ~A168 & ~A169;
  assign \new_[74125]_  = A170 & \new_[74124]_ ;
  assign \new_[74128]_  = A166 & ~A167;
  assign \new_[74131]_  = ~A200 & ~A199;
  assign \new_[74132]_  = \new_[74131]_  & \new_[74128]_ ;
  assign \new_[74133]_  = \new_[74132]_  & \new_[74125]_ ;
  assign \new_[74137]_  = A298 & A269;
  assign \new_[74138]_  = ~A267 & \new_[74137]_ ;
  assign \new_[74141]_  = ~A300 & ~A299;
  assign \new_[74144]_  = ~A302 & ~A301;
  assign \new_[74145]_  = \new_[74144]_  & \new_[74141]_ ;
  assign \new_[74146]_  = \new_[74145]_  & \new_[74138]_ ;
  assign \new_[74150]_  = ~A168 & ~A169;
  assign \new_[74151]_  = A170 & \new_[74150]_ ;
  assign \new_[74154]_  = A166 & ~A167;
  assign \new_[74157]_  = ~A200 & ~A199;
  assign \new_[74158]_  = \new_[74157]_  & \new_[74154]_ ;
  assign \new_[74159]_  = \new_[74158]_  & \new_[74151]_ ;
  assign \new_[74163]_  = ~A298 & A269;
  assign \new_[74164]_  = ~A267 & \new_[74163]_ ;
  assign \new_[74167]_  = ~A300 & A299;
  assign \new_[74170]_  = ~A302 & ~A301;
  assign \new_[74171]_  = \new_[74170]_  & \new_[74167]_ ;
  assign \new_[74172]_  = \new_[74171]_  & \new_[74164]_ ;
  assign \new_[74176]_  = ~A168 & ~A169;
  assign \new_[74177]_  = A170 & \new_[74176]_ ;
  assign \new_[74180]_  = A166 & ~A167;
  assign \new_[74183]_  = ~A200 & ~A199;
  assign \new_[74184]_  = \new_[74183]_  & \new_[74180]_ ;
  assign \new_[74185]_  = \new_[74184]_  & \new_[74177]_ ;
  assign \new_[74189]_  = A298 & A266;
  assign \new_[74190]_  = A265 & \new_[74189]_ ;
  assign \new_[74193]_  = ~A300 & ~A299;
  assign \new_[74196]_  = ~A302 & ~A301;
  assign \new_[74197]_  = \new_[74196]_  & \new_[74193]_ ;
  assign \new_[74198]_  = \new_[74197]_  & \new_[74190]_ ;
  assign \new_[74202]_  = ~A168 & ~A169;
  assign \new_[74203]_  = A170 & \new_[74202]_ ;
  assign \new_[74206]_  = A166 & ~A167;
  assign \new_[74209]_  = ~A200 & ~A199;
  assign \new_[74210]_  = \new_[74209]_  & \new_[74206]_ ;
  assign \new_[74211]_  = \new_[74210]_  & \new_[74203]_ ;
  assign \new_[74215]_  = ~A298 & A266;
  assign \new_[74216]_  = A265 & \new_[74215]_ ;
  assign \new_[74219]_  = ~A300 & A299;
  assign \new_[74222]_  = ~A302 & ~A301;
  assign \new_[74223]_  = \new_[74222]_  & \new_[74219]_ ;
  assign \new_[74224]_  = \new_[74223]_  & \new_[74216]_ ;
  assign \new_[74228]_  = ~A168 & ~A169;
  assign \new_[74229]_  = A170 & \new_[74228]_ ;
  assign \new_[74232]_  = A166 & ~A167;
  assign \new_[74235]_  = ~A200 & ~A199;
  assign \new_[74236]_  = \new_[74235]_  & \new_[74232]_ ;
  assign \new_[74237]_  = \new_[74236]_  & \new_[74229]_ ;
  assign \new_[74241]_  = A298 & ~A266;
  assign \new_[74242]_  = ~A265 & \new_[74241]_ ;
  assign \new_[74245]_  = ~A300 & ~A299;
  assign \new_[74248]_  = ~A302 & ~A301;
  assign \new_[74249]_  = \new_[74248]_  & \new_[74245]_ ;
  assign \new_[74250]_  = \new_[74249]_  & \new_[74242]_ ;
  assign \new_[74254]_  = ~A168 & ~A169;
  assign \new_[74255]_  = A170 & \new_[74254]_ ;
  assign \new_[74258]_  = A166 & ~A167;
  assign \new_[74261]_  = ~A200 & ~A199;
  assign \new_[74262]_  = \new_[74261]_  & \new_[74258]_ ;
  assign \new_[74263]_  = \new_[74262]_  & \new_[74255]_ ;
  assign \new_[74267]_  = ~A298 & ~A266;
  assign \new_[74268]_  = ~A265 & \new_[74267]_ ;
  assign \new_[74271]_  = ~A300 & A299;
  assign \new_[74274]_  = ~A302 & ~A301;
  assign \new_[74275]_  = \new_[74274]_  & \new_[74271]_ ;
  assign \new_[74276]_  = \new_[74275]_  & \new_[74268]_ ;
  assign \new_[74280]_  = ~A199 & A166;
  assign \new_[74281]_  = A167 & \new_[74280]_ ;
  assign \new_[74284]_  = ~A201 & A200;
  assign \new_[74287]_  = ~A203 & ~A202;
  assign \new_[74288]_  = \new_[74287]_  & \new_[74284]_ ;
  assign \new_[74289]_  = \new_[74288]_  & \new_[74281]_ ;
  assign \new_[74292]_  = ~A268 & A267;
  assign \new_[74295]_  = A298 & ~A269;
  assign \new_[74296]_  = \new_[74295]_  & \new_[74292]_ ;
  assign \new_[74299]_  = ~A300 & ~A299;
  assign \new_[74302]_  = ~A302 & ~A301;
  assign \new_[74303]_  = \new_[74302]_  & \new_[74299]_ ;
  assign \new_[74304]_  = \new_[74303]_  & \new_[74296]_ ;
  assign \new_[74308]_  = ~A199 & A166;
  assign \new_[74309]_  = A167 & \new_[74308]_ ;
  assign \new_[74312]_  = ~A201 & A200;
  assign \new_[74315]_  = ~A203 & ~A202;
  assign \new_[74316]_  = \new_[74315]_  & \new_[74312]_ ;
  assign \new_[74317]_  = \new_[74316]_  & \new_[74309]_ ;
  assign \new_[74320]_  = ~A268 & A267;
  assign \new_[74323]_  = ~A298 & ~A269;
  assign \new_[74324]_  = \new_[74323]_  & \new_[74320]_ ;
  assign \new_[74327]_  = ~A300 & A299;
  assign \new_[74330]_  = ~A302 & ~A301;
  assign \new_[74331]_  = \new_[74330]_  & \new_[74327]_ ;
  assign \new_[74332]_  = \new_[74331]_  & \new_[74324]_ ;
  assign \new_[74336]_  = A199 & A166;
  assign \new_[74337]_  = A167 & \new_[74336]_ ;
  assign \new_[74340]_  = ~A201 & ~A200;
  assign \new_[74343]_  = ~A203 & ~A202;
  assign \new_[74344]_  = \new_[74343]_  & \new_[74340]_ ;
  assign \new_[74345]_  = \new_[74344]_  & \new_[74337]_ ;
  assign \new_[74348]_  = ~A268 & A267;
  assign \new_[74351]_  = A298 & ~A269;
  assign \new_[74352]_  = \new_[74351]_  & \new_[74348]_ ;
  assign \new_[74355]_  = ~A300 & ~A299;
  assign \new_[74358]_  = ~A302 & ~A301;
  assign \new_[74359]_  = \new_[74358]_  & \new_[74355]_ ;
  assign \new_[74360]_  = \new_[74359]_  & \new_[74352]_ ;
  assign \new_[74364]_  = A199 & A166;
  assign \new_[74365]_  = A167 & \new_[74364]_ ;
  assign \new_[74368]_  = ~A201 & ~A200;
  assign \new_[74371]_  = ~A203 & ~A202;
  assign \new_[74372]_  = \new_[74371]_  & \new_[74368]_ ;
  assign \new_[74373]_  = \new_[74372]_  & \new_[74365]_ ;
  assign \new_[74376]_  = ~A268 & A267;
  assign \new_[74379]_  = ~A298 & ~A269;
  assign \new_[74380]_  = \new_[74379]_  & \new_[74376]_ ;
  assign \new_[74383]_  = ~A300 & A299;
  assign \new_[74386]_  = ~A302 & ~A301;
  assign \new_[74387]_  = \new_[74386]_  & \new_[74383]_ ;
  assign \new_[74388]_  = \new_[74387]_  & \new_[74380]_ ;
  assign \new_[74392]_  = ~A199 & ~A166;
  assign \new_[74393]_  = ~A167 & \new_[74392]_ ;
  assign \new_[74396]_  = ~A201 & A200;
  assign \new_[74399]_  = ~A203 & ~A202;
  assign \new_[74400]_  = \new_[74399]_  & \new_[74396]_ ;
  assign \new_[74401]_  = \new_[74400]_  & \new_[74393]_ ;
  assign \new_[74404]_  = ~A268 & A267;
  assign \new_[74407]_  = A298 & ~A269;
  assign \new_[74408]_  = \new_[74407]_  & \new_[74404]_ ;
  assign \new_[74411]_  = ~A300 & ~A299;
  assign \new_[74414]_  = ~A302 & ~A301;
  assign \new_[74415]_  = \new_[74414]_  & \new_[74411]_ ;
  assign \new_[74416]_  = \new_[74415]_  & \new_[74408]_ ;
  assign \new_[74420]_  = ~A199 & ~A166;
  assign \new_[74421]_  = ~A167 & \new_[74420]_ ;
  assign \new_[74424]_  = ~A201 & A200;
  assign \new_[74427]_  = ~A203 & ~A202;
  assign \new_[74428]_  = \new_[74427]_  & \new_[74424]_ ;
  assign \new_[74429]_  = \new_[74428]_  & \new_[74421]_ ;
  assign \new_[74432]_  = ~A268 & A267;
  assign \new_[74435]_  = ~A298 & ~A269;
  assign \new_[74436]_  = \new_[74435]_  & \new_[74432]_ ;
  assign \new_[74439]_  = ~A300 & A299;
  assign \new_[74442]_  = ~A302 & ~A301;
  assign \new_[74443]_  = \new_[74442]_  & \new_[74439]_ ;
  assign \new_[74444]_  = \new_[74443]_  & \new_[74436]_ ;
  assign \new_[74448]_  = A199 & ~A166;
  assign \new_[74449]_  = ~A167 & \new_[74448]_ ;
  assign \new_[74452]_  = ~A201 & ~A200;
  assign \new_[74455]_  = ~A203 & ~A202;
  assign \new_[74456]_  = \new_[74455]_  & \new_[74452]_ ;
  assign \new_[74457]_  = \new_[74456]_  & \new_[74449]_ ;
  assign \new_[74460]_  = ~A268 & A267;
  assign \new_[74463]_  = A298 & ~A269;
  assign \new_[74464]_  = \new_[74463]_  & \new_[74460]_ ;
  assign \new_[74467]_  = ~A300 & ~A299;
  assign \new_[74470]_  = ~A302 & ~A301;
  assign \new_[74471]_  = \new_[74470]_  & \new_[74467]_ ;
  assign \new_[74472]_  = \new_[74471]_  & \new_[74464]_ ;
  assign \new_[74476]_  = A199 & ~A166;
  assign \new_[74477]_  = ~A167 & \new_[74476]_ ;
  assign \new_[74480]_  = ~A201 & ~A200;
  assign \new_[74483]_  = ~A203 & ~A202;
  assign \new_[74484]_  = \new_[74483]_  & \new_[74480]_ ;
  assign \new_[74485]_  = \new_[74484]_  & \new_[74477]_ ;
  assign \new_[74488]_  = ~A268 & A267;
  assign \new_[74491]_  = ~A298 & ~A269;
  assign \new_[74492]_  = \new_[74491]_  & \new_[74488]_ ;
  assign \new_[74495]_  = ~A300 & A299;
  assign \new_[74498]_  = ~A302 & ~A301;
  assign \new_[74499]_  = \new_[74498]_  & \new_[74495]_ ;
  assign \new_[74500]_  = \new_[74499]_  & \new_[74492]_ ;
  assign \new_[74504]_  = A167 & A168;
  assign \new_[74505]_  = ~A170 & \new_[74504]_ ;
  assign \new_[74508]_  = A201 & ~A166;
  assign \new_[74511]_  = ~A203 & ~A202;
  assign \new_[74512]_  = \new_[74511]_  & \new_[74508]_ ;
  assign \new_[74513]_  = \new_[74512]_  & \new_[74505]_ ;
  assign \new_[74516]_  = ~A268 & A267;
  assign \new_[74519]_  = A298 & ~A269;
  assign \new_[74520]_  = \new_[74519]_  & \new_[74516]_ ;
  assign \new_[74523]_  = ~A300 & ~A299;
  assign \new_[74526]_  = ~A302 & ~A301;
  assign \new_[74527]_  = \new_[74526]_  & \new_[74523]_ ;
  assign \new_[74528]_  = \new_[74527]_  & \new_[74520]_ ;
  assign \new_[74532]_  = A167 & A168;
  assign \new_[74533]_  = ~A170 & \new_[74532]_ ;
  assign \new_[74536]_  = A201 & ~A166;
  assign \new_[74539]_  = ~A203 & ~A202;
  assign \new_[74540]_  = \new_[74539]_  & \new_[74536]_ ;
  assign \new_[74541]_  = \new_[74540]_  & \new_[74533]_ ;
  assign \new_[74544]_  = ~A268 & A267;
  assign \new_[74547]_  = ~A298 & ~A269;
  assign \new_[74548]_  = \new_[74547]_  & \new_[74544]_ ;
  assign \new_[74551]_  = ~A300 & A299;
  assign \new_[74554]_  = ~A302 & ~A301;
  assign \new_[74555]_  = \new_[74554]_  & \new_[74551]_ ;
  assign \new_[74556]_  = \new_[74555]_  & \new_[74548]_ ;
  assign \new_[74560]_  = A167 & A168;
  assign \new_[74561]_  = ~A170 & \new_[74560]_ ;
  assign \new_[74564]_  = ~A199 & ~A166;
  assign \new_[74567]_  = A201 & A200;
  assign \new_[74568]_  = \new_[74567]_  & \new_[74564]_ ;
  assign \new_[74569]_  = \new_[74568]_  & \new_[74561]_ ;
  assign \new_[74572]_  = ~A265 & A202;
  assign \new_[74575]_  = A267 & A266;
  assign \new_[74576]_  = \new_[74575]_  & \new_[74572]_ ;
  assign \new_[74579]_  = A300 & A268;
  assign \new_[74582]_  = ~A302 & ~A301;
  assign \new_[74583]_  = \new_[74582]_  & \new_[74579]_ ;
  assign \new_[74584]_  = \new_[74583]_  & \new_[74576]_ ;
  assign \new_[74588]_  = A167 & A168;
  assign \new_[74589]_  = ~A170 & \new_[74588]_ ;
  assign \new_[74592]_  = ~A199 & ~A166;
  assign \new_[74595]_  = A201 & A200;
  assign \new_[74596]_  = \new_[74595]_  & \new_[74592]_ ;
  assign \new_[74597]_  = \new_[74596]_  & \new_[74589]_ ;
  assign \new_[74600]_  = ~A265 & A202;
  assign \new_[74603]_  = A267 & A266;
  assign \new_[74604]_  = \new_[74603]_  & \new_[74600]_ ;
  assign \new_[74607]_  = A300 & A269;
  assign \new_[74610]_  = ~A302 & ~A301;
  assign \new_[74611]_  = \new_[74610]_  & \new_[74607]_ ;
  assign \new_[74612]_  = \new_[74611]_  & \new_[74604]_ ;
  assign \new_[74616]_  = A167 & A168;
  assign \new_[74617]_  = ~A170 & \new_[74616]_ ;
  assign \new_[74620]_  = ~A199 & ~A166;
  assign \new_[74623]_  = A201 & A200;
  assign \new_[74624]_  = \new_[74623]_  & \new_[74620]_ ;
  assign \new_[74625]_  = \new_[74624]_  & \new_[74617]_ ;
  assign \new_[74628]_  = ~A265 & A202;
  assign \new_[74631]_  = ~A267 & A266;
  assign \new_[74632]_  = \new_[74631]_  & \new_[74628]_ ;
  assign \new_[74635]_  = ~A269 & ~A268;
  assign \new_[74638]_  = A301 & ~A300;
  assign \new_[74639]_  = \new_[74638]_  & \new_[74635]_ ;
  assign \new_[74640]_  = \new_[74639]_  & \new_[74632]_ ;
  assign \new_[74644]_  = A167 & A168;
  assign \new_[74645]_  = ~A170 & \new_[74644]_ ;
  assign \new_[74648]_  = ~A199 & ~A166;
  assign \new_[74651]_  = A201 & A200;
  assign \new_[74652]_  = \new_[74651]_  & \new_[74648]_ ;
  assign \new_[74653]_  = \new_[74652]_  & \new_[74645]_ ;
  assign \new_[74656]_  = ~A265 & A202;
  assign \new_[74659]_  = ~A267 & A266;
  assign \new_[74660]_  = \new_[74659]_  & \new_[74656]_ ;
  assign \new_[74663]_  = ~A269 & ~A268;
  assign \new_[74666]_  = A302 & ~A300;
  assign \new_[74667]_  = \new_[74666]_  & \new_[74663]_ ;
  assign \new_[74668]_  = \new_[74667]_  & \new_[74660]_ ;
  assign \new_[74672]_  = A167 & A168;
  assign \new_[74673]_  = ~A170 & \new_[74672]_ ;
  assign \new_[74676]_  = ~A199 & ~A166;
  assign \new_[74679]_  = A201 & A200;
  assign \new_[74680]_  = \new_[74679]_  & \new_[74676]_ ;
  assign \new_[74681]_  = \new_[74680]_  & \new_[74673]_ ;
  assign \new_[74684]_  = ~A265 & A202;
  assign \new_[74687]_  = ~A267 & A266;
  assign \new_[74688]_  = \new_[74687]_  & \new_[74684]_ ;
  assign \new_[74691]_  = ~A269 & ~A268;
  assign \new_[74694]_  = A299 & A298;
  assign \new_[74695]_  = \new_[74694]_  & \new_[74691]_ ;
  assign \new_[74696]_  = \new_[74695]_  & \new_[74688]_ ;
  assign \new_[74700]_  = A167 & A168;
  assign \new_[74701]_  = ~A170 & \new_[74700]_ ;
  assign \new_[74704]_  = ~A199 & ~A166;
  assign \new_[74707]_  = A201 & A200;
  assign \new_[74708]_  = \new_[74707]_  & \new_[74704]_ ;
  assign \new_[74709]_  = \new_[74708]_  & \new_[74701]_ ;
  assign \new_[74712]_  = ~A265 & A202;
  assign \new_[74715]_  = ~A267 & A266;
  assign \new_[74716]_  = \new_[74715]_  & \new_[74712]_ ;
  assign \new_[74719]_  = ~A269 & ~A268;
  assign \new_[74722]_  = ~A299 & ~A298;
  assign \new_[74723]_  = \new_[74722]_  & \new_[74719]_ ;
  assign \new_[74724]_  = \new_[74723]_  & \new_[74716]_ ;
  assign \new_[74728]_  = A167 & A168;
  assign \new_[74729]_  = ~A170 & \new_[74728]_ ;
  assign \new_[74732]_  = ~A199 & ~A166;
  assign \new_[74735]_  = A201 & A200;
  assign \new_[74736]_  = \new_[74735]_  & \new_[74732]_ ;
  assign \new_[74737]_  = \new_[74736]_  & \new_[74729]_ ;
  assign \new_[74740]_  = A265 & A202;
  assign \new_[74743]_  = A267 & ~A266;
  assign \new_[74744]_  = \new_[74743]_  & \new_[74740]_ ;
  assign \new_[74747]_  = A300 & A268;
  assign \new_[74750]_  = ~A302 & ~A301;
  assign \new_[74751]_  = \new_[74750]_  & \new_[74747]_ ;
  assign \new_[74752]_  = \new_[74751]_  & \new_[74744]_ ;
  assign \new_[74756]_  = A167 & A168;
  assign \new_[74757]_  = ~A170 & \new_[74756]_ ;
  assign \new_[74760]_  = ~A199 & ~A166;
  assign \new_[74763]_  = A201 & A200;
  assign \new_[74764]_  = \new_[74763]_  & \new_[74760]_ ;
  assign \new_[74765]_  = \new_[74764]_  & \new_[74757]_ ;
  assign \new_[74768]_  = A265 & A202;
  assign \new_[74771]_  = A267 & ~A266;
  assign \new_[74772]_  = \new_[74771]_  & \new_[74768]_ ;
  assign \new_[74775]_  = A300 & A269;
  assign \new_[74778]_  = ~A302 & ~A301;
  assign \new_[74779]_  = \new_[74778]_  & \new_[74775]_ ;
  assign \new_[74780]_  = \new_[74779]_  & \new_[74772]_ ;
  assign \new_[74784]_  = A167 & A168;
  assign \new_[74785]_  = ~A170 & \new_[74784]_ ;
  assign \new_[74788]_  = ~A199 & ~A166;
  assign \new_[74791]_  = A201 & A200;
  assign \new_[74792]_  = \new_[74791]_  & \new_[74788]_ ;
  assign \new_[74793]_  = \new_[74792]_  & \new_[74785]_ ;
  assign \new_[74796]_  = A265 & A202;
  assign \new_[74799]_  = ~A267 & ~A266;
  assign \new_[74800]_  = \new_[74799]_  & \new_[74796]_ ;
  assign \new_[74803]_  = ~A269 & ~A268;
  assign \new_[74806]_  = A301 & ~A300;
  assign \new_[74807]_  = \new_[74806]_  & \new_[74803]_ ;
  assign \new_[74808]_  = \new_[74807]_  & \new_[74800]_ ;
  assign \new_[74812]_  = A167 & A168;
  assign \new_[74813]_  = ~A170 & \new_[74812]_ ;
  assign \new_[74816]_  = ~A199 & ~A166;
  assign \new_[74819]_  = A201 & A200;
  assign \new_[74820]_  = \new_[74819]_  & \new_[74816]_ ;
  assign \new_[74821]_  = \new_[74820]_  & \new_[74813]_ ;
  assign \new_[74824]_  = A265 & A202;
  assign \new_[74827]_  = ~A267 & ~A266;
  assign \new_[74828]_  = \new_[74827]_  & \new_[74824]_ ;
  assign \new_[74831]_  = ~A269 & ~A268;
  assign \new_[74834]_  = A302 & ~A300;
  assign \new_[74835]_  = \new_[74834]_  & \new_[74831]_ ;
  assign \new_[74836]_  = \new_[74835]_  & \new_[74828]_ ;
  assign \new_[74840]_  = A167 & A168;
  assign \new_[74841]_  = ~A170 & \new_[74840]_ ;
  assign \new_[74844]_  = ~A199 & ~A166;
  assign \new_[74847]_  = A201 & A200;
  assign \new_[74848]_  = \new_[74847]_  & \new_[74844]_ ;
  assign \new_[74849]_  = \new_[74848]_  & \new_[74841]_ ;
  assign \new_[74852]_  = A265 & A202;
  assign \new_[74855]_  = ~A267 & ~A266;
  assign \new_[74856]_  = \new_[74855]_  & \new_[74852]_ ;
  assign \new_[74859]_  = ~A269 & ~A268;
  assign \new_[74862]_  = A299 & A298;
  assign \new_[74863]_  = \new_[74862]_  & \new_[74859]_ ;
  assign \new_[74864]_  = \new_[74863]_  & \new_[74856]_ ;
  assign \new_[74868]_  = A167 & A168;
  assign \new_[74869]_  = ~A170 & \new_[74868]_ ;
  assign \new_[74872]_  = ~A199 & ~A166;
  assign \new_[74875]_  = A201 & A200;
  assign \new_[74876]_  = \new_[74875]_  & \new_[74872]_ ;
  assign \new_[74877]_  = \new_[74876]_  & \new_[74869]_ ;
  assign \new_[74880]_  = A265 & A202;
  assign \new_[74883]_  = ~A267 & ~A266;
  assign \new_[74884]_  = \new_[74883]_  & \new_[74880]_ ;
  assign \new_[74887]_  = ~A269 & ~A268;
  assign \new_[74890]_  = ~A299 & ~A298;
  assign \new_[74891]_  = \new_[74890]_  & \new_[74887]_ ;
  assign \new_[74892]_  = \new_[74891]_  & \new_[74884]_ ;
  assign \new_[74896]_  = A167 & A168;
  assign \new_[74897]_  = ~A170 & \new_[74896]_ ;
  assign \new_[74900]_  = ~A199 & ~A166;
  assign \new_[74903]_  = A201 & A200;
  assign \new_[74904]_  = \new_[74903]_  & \new_[74900]_ ;
  assign \new_[74905]_  = \new_[74904]_  & \new_[74897]_ ;
  assign \new_[74908]_  = ~A265 & A203;
  assign \new_[74911]_  = A267 & A266;
  assign \new_[74912]_  = \new_[74911]_  & \new_[74908]_ ;
  assign \new_[74915]_  = A300 & A268;
  assign \new_[74918]_  = ~A302 & ~A301;
  assign \new_[74919]_  = \new_[74918]_  & \new_[74915]_ ;
  assign \new_[74920]_  = \new_[74919]_  & \new_[74912]_ ;
  assign \new_[74924]_  = A167 & A168;
  assign \new_[74925]_  = ~A170 & \new_[74924]_ ;
  assign \new_[74928]_  = ~A199 & ~A166;
  assign \new_[74931]_  = A201 & A200;
  assign \new_[74932]_  = \new_[74931]_  & \new_[74928]_ ;
  assign \new_[74933]_  = \new_[74932]_  & \new_[74925]_ ;
  assign \new_[74936]_  = ~A265 & A203;
  assign \new_[74939]_  = A267 & A266;
  assign \new_[74940]_  = \new_[74939]_  & \new_[74936]_ ;
  assign \new_[74943]_  = A300 & A269;
  assign \new_[74946]_  = ~A302 & ~A301;
  assign \new_[74947]_  = \new_[74946]_  & \new_[74943]_ ;
  assign \new_[74948]_  = \new_[74947]_  & \new_[74940]_ ;
  assign \new_[74952]_  = A167 & A168;
  assign \new_[74953]_  = ~A170 & \new_[74952]_ ;
  assign \new_[74956]_  = ~A199 & ~A166;
  assign \new_[74959]_  = A201 & A200;
  assign \new_[74960]_  = \new_[74959]_  & \new_[74956]_ ;
  assign \new_[74961]_  = \new_[74960]_  & \new_[74953]_ ;
  assign \new_[74964]_  = ~A265 & A203;
  assign \new_[74967]_  = ~A267 & A266;
  assign \new_[74968]_  = \new_[74967]_  & \new_[74964]_ ;
  assign \new_[74971]_  = ~A269 & ~A268;
  assign \new_[74974]_  = A301 & ~A300;
  assign \new_[74975]_  = \new_[74974]_  & \new_[74971]_ ;
  assign \new_[74976]_  = \new_[74975]_  & \new_[74968]_ ;
  assign \new_[74980]_  = A167 & A168;
  assign \new_[74981]_  = ~A170 & \new_[74980]_ ;
  assign \new_[74984]_  = ~A199 & ~A166;
  assign \new_[74987]_  = A201 & A200;
  assign \new_[74988]_  = \new_[74987]_  & \new_[74984]_ ;
  assign \new_[74989]_  = \new_[74988]_  & \new_[74981]_ ;
  assign \new_[74992]_  = ~A265 & A203;
  assign \new_[74995]_  = ~A267 & A266;
  assign \new_[74996]_  = \new_[74995]_  & \new_[74992]_ ;
  assign \new_[74999]_  = ~A269 & ~A268;
  assign \new_[75002]_  = A302 & ~A300;
  assign \new_[75003]_  = \new_[75002]_  & \new_[74999]_ ;
  assign \new_[75004]_  = \new_[75003]_  & \new_[74996]_ ;
  assign \new_[75008]_  = A167 & A168;
  assign \new_[75009]_  = ~A170 & \new_[75008]_ ;
  assign \new_[75012]_  = ~A199 & ~A166;
  assign \new_[75015]_  = A201 & A200;
  assign \new_[75016]_  = \new_[75015]_  & \new_[75012]_ ;
  assign \new_[75017]_  = \new_[75016]_  & \new_[75009]_ ;
  assign \new_[75020]_  = ~A265 & A203;
  assign \new_[75023]_  = ~A267 & A266;
  assign \new_[75024]_  = \new_[75023]_  & \new_[75020]_ ;
  assign \new_[75027]_  = ~A269 & ~A268;
  assign \new_[75030]_  = A299 & A298;
  assign \new_[75031]_  = \new_[75030]_  & \new_[75027]_ ;
  assign \new_[75032]_  = \new_[75031]_  & \new_[75024]_ ;
  assign \new_[75036]_  = A167 & A168;
  assign \new_[75037]_  = ~A170 & \new_[75036]_ ;
  assign \new_[75040]_  = ~A199 & ~A166;
  assign \new_[75043]_  = A201 & A200;
  assign \new_[75044]_  = \new_[75043]_  & \new_[75040]_ ;
  assign \new_[75045]_  = \new_[75044]_  & \new_[75037]_ ;
  assign \new_[75048]_  = ~A265 & A203;
  assign \new_[75051]_  = ~A267 & A266;
  assign \new_[75052]_  = \new_[75051]_  & \new_[75048]_ ;
  assign \new_[75055]_  = ~A269 & ~A268;
  assign \new_[75058]_  = ~A299 & ~A298;
  assign \new_[75059]_  = \new_[75058]_  & \new_[75055]_ ;
  assign \new_[75060]_  = \new_[75059]_  & \new_[75052]_ ;
  assign \new_[75064]_  = A167 & A168;
  assign \new_[75065]_  = ~A170 & \new_[75064]_ ;
  assign \new_[75068]_  = ~A199 & ~A166;
  assign \new_[75071]_  = A201 & A200;
  assign \new_[75072]_  = \new_[75071]_  & \new_[75068]_ ;
  assign \new_[75073]_  = \new_[75072]_  & \new_[75065]_ ;
  assign \new_[75076]_  = A265 & A203;
  assign \new_[75079]_  = A267 & ~A266;
  assign \new_[75080]_  = \new_[75079]_  & \new_[75076]_ ;
  assign \new_[75083]_  = A300 & A268;
  assign \new_[75086]_  = ~A302 & ~A301;
  assign \new_[75087]_  = \new_[75086]_  & \new_[75083]_ ;
  assign \new_[75088]_  = \new_[75087]_  & \new_[75080]_ ;
  assign \new_[75092]_  = A167 & A168;
  assign \new_[75093]_  = ~A170 & \new_[75092]_ ;
  assign \new_[75096]_  = ~A199 & ~A166;
  assign \new_[75099]_  = A201 & A200;
  assign \new_[75100]_  = \new_[75099]_  & \new_[75096]_ ;
  assign \new_[75101]_  = \new_[75100]_  & \new_[75093]_ ;
  assign \new_[75104]_  = A265 & A203;
  assign \new_[75107]_  = A267 & ~A266;
  assign \new_[75108]_  = \new_[75107]_  & \new_[75104]_ ;
  assign \new_[75111]_  = A300 & A269;
  assign \new_[75114]_  = ~A302 & ~A301;
  assign \new_[75115]_  = \new_[75114]_  & \new_[75111]_ ;
  assign \new_[75116]_  = \new_[75115]_  & \new_[75108]_ ;
  assign \new_[75120]_  = A167 & A168;
  assign \new_[75121]_  = ~A170 & \new_[75120]_ ;
  assign \new_[75124]_  = ~A199 & ~A166;
  assign \new_[75127]_  = A201 & A200;
  assign \new_[75128]_  = \new_[75127]_  & \new_[75124]_ ;
  assign \new_[75129]_  = \new_[75128]_  & \new_[75121]_ ;
  assign \new_[75132]_  = A265 & A203;
  assign \new_[75135]_  = ~A267 & ~A266;
  assign \new_[75136]_  = \new_[75135]_  & \new_[75132]_ ;
  assign \new_[75139]_  = ~A269 & ~A268;
  assign \new_[75142]_  = A301 & ~A300;
  assign \new_[75143]_  = \new_[75142]_  & \new_[75139]_ ;
  assign \new_[75144]_  = \new_[75143]_  & \new_[75136]_ ;
  assign \new_[75148]_  = A167 & A168;
  assign \new_[75149]_  = ~A170 & \new_[75148]_ ;
  assign \new_[75152]_  = ~A199 & ~A166;
  assign \new_[75155]_  = A201 & A200;
  assign \new_[75156]_  = \new_[75155]_  & \new_[75152]_ ;
  assign \new_[75157]_  = \new_[75156]_  & \new_[75149]_ ;
  assign \new_[75160]_  = A265 & A203;
  assign \new_[75163]_  = ~A267 & ~A266;
  assign \new_[75164]_  = \new_[75163]_  & \new_[75160]_ ;
  assign \new_[75167]_  = ~A269 & ~A268;
  assign \new_[75170]_  = A302 & ~A300;
  assign \new_[75171]_  = \new_[75170]_  & \new_[75167]_ ;
  assign \new_[75172]_  = \new_[75171]_  & \new_[75164]_ ;
  assign \new_[75176]_  = A167 & A168;
  assign \new_[75177]_  = ~A170 & \new_[75176]_ ;
  assign \new_[75180]_  = ~A199 & ~A166;
  assign \new_[75183]_  = A201 & A200;
  assign \new_[75184]_  = \new_[75183]_  & \new_[75180]_ ;
  assign \new_[75185]_  = \new_[75184]_  & \new_[75177]_ ;
  assign \new_[75188]_  = A265 & A203;
  assign \new_[75191]_  = ~A267 & ~A266;
  assign \new_[75192]_  = \new_[75191]_  & \new_[75188]_ ;
  assign \new_[75195]_  = ~A269 & ~A268;
  assign \new_[75198]_  = A299 & A298;
  assign \new_[75199]_  = \new_[75198]_  & \new_[75195]_ ;
  assign \new_[75200]_  = \new_[75199]_  & \new_[75192]_ ;
  assign \new_[75204]_  = A167 & A168;
  assign \new_[75205]_  = ~A170 & \new_[75204]_ ;
  assign \new_[75208]_  = ~A199 & ~A166;
  assign \new_[75211]_  = A201 & A200;
  assign \new_[75212]_  = \new_[75211]_  & \new_[75208]_ ;
  assign \new_[75213]_  = \new_[75212]_  & \new_[75205]_ ;
  assign \new_[75216]_  = A265 & A203;
  assign \new_[75219]_  = ~A267 & ~A266;
  assign \new_[75220]_  = \new_[75219]_  & \new_[75216]_ ;
  assign \new_[75223]_  = ~A269 & ~A268;
  assign \new_[75226]_  = ~A299 & ~A298;
  assign \new_[75227]_  = \new_[75226]_  & \new_[75223]_ ;
  assign \new_[75228]_  = \new_[75227]_  & \new_[75220]_ ;
  assign \new_[75232]_  = A167 & A168;
  assign \new_[75233]_  = ~A170 & \new_[75232]_ ;
  assign \new_[75236]_  = ~A199 & ~A166;
  assign \new_[75239]_  = ~A201 & A200;
  assign \new_[75240]_  = \new_[75239]_  & \new_[75236]_ ;
  assign \new_[75241]_  = \new_[75240]_  & \new_[75233]_ ;
  assign \new_[75244]_  = ~A203 & ~A202;
  assign \new_[75247]_  = A266 & ~A265;
  assign \new_[75248]_  = \new_[75247]_  & \new_[75244]_ ;
  assign \new_[75251]_  = A268 & A267;
  assign \new_[75254]_  = A301 & ~A300;
  assign \new_[75255]_  = \new_[75254]_  & \new_[75251]_ ;
  assign \new_[75256]_  = \new_[75255]_  & \new_[75248]_ ;
  assign \new_[75260]_  = A167 & A168;
  assign \new_[75261]_  = ~A170 & \new_[75260]_ ;
  assign \new_[75264]_  = ~A199 & ~A166;
  assign \new_[75267]_  = ~A201 & A200;
  assign \new_[75268]_  = \new_[75267]_  & \new_[75264]_ ;
  assign \new_[75269]_  = \new_[75268]_  & \new_[75261]_ ;
  assign \new_[75272]_  = ~A203 & ~A202;
  assign \new_[75275]_  = A266 & ~A265;
  assign \new_[75276]_  = \new_[75275]_  & \new_[75272]_ ;
  assign \new_[75279]_  = A268 & A267;
  assign \new_[75282]_  = A302 & ~A300;
  assign \new_[75283]_  = \new_[75282]_  & \new_[75279]_ ;
  assign \new_[75284]_  = \new_[75283]_  & \new_[75276]_ ;
  assign \new_[75288]_  = A167 & A168;
  assign \new_[75289]_  = ~A170 & \new_[75288]_ ;
  assign \new_[75292]_  = ~A199 & ~A166;
  assign \new_[75295]_  = ~A201 & A200;
  assign \new_[75296]_  = \new_[75295]_  & \new_[75292]_ ;
  assign \new_[75297]_  = \new_[75296]_  & \new_[75289]_ ;
  assign \new_[75300]_  = ~A203 & ~A202;
  assign \new_[75303]_  = A266 & ~A265;
  assign \new_[75304]_  = \new_[75303]_  & \new_[75300]_ ;
  assign \new_[75307]_  = A268 & A267;
  assign \new_[75310]_  = A299 & A298;
  assign \new_[75311]_  = \new_[75310]_  & \new_[75307]_ ;
  assign \new_[75312]_  = \new_[75311]_  & \new_[75304]_ ;
  assign \new_[75316]_  = A167 & A168;
  assign \new_[75317]_  = ~A170 & \new_[75316]_ ;
  assign \new_[75320]_  = ~A199 & ~A166;
  assign \new_[75323]_  = ~A201 & A200;
  assign \new_[75324]_  = \new_[75323]_  & \new_[75320]_ ;
  assign \new_[75325]_  = \new_[75324]_  & \new_[75317]_ ;
  assign \new_[75328]_  = ~A203 & ~A202;
  assign \new_[75331]_  = A266 & ~A265;
  assign \new_[75332]_  = \new_[75331]_  & \new_[75328]_ ;
  assign \new_[75335]_  = A268 & A267;
  assign \new_[75338]_  = ~A299 & ~A298;
  assign \new_[75339]_  = \new_[75338]_  & \new_[75335]_ ;
  assign \new_[75340]_  = \new_[75339]_  & \new_[75332]_ ;
  assign \new_[75344]_  = A167 & A168;
  assign \new_[75345]_  = ~A170 & \new_[75344]_ ;
  assign \new_[75348]_  = ~A199 & ~A166;
  assign \new_[75351]_  = ~A201 & A200;
  assign \new_[75352]_  = \new_[75351]_  & \new_[75348]_ ;
  assign \new_[75353]_  = \new_[75352]_  & \new_[75345]_ ;
  assign \new_[75356]_  = ~A203 & ~A202;
  assign \new_[75359]_  = A266 & ~A265;
  assign \new_[75360]_  = \new_[75359]_  & \new_[75356]_ ;
  assign \new_[75363]_  = A269 & A267;
  assign \new_[75366]_  = A301 & ~A300;
  assign \new_[75367]_  = \new_[75366]_  & \new_[75363]_ ;
  assign \new_[75368]_  = \new_[75367]_  & \new_[75360]_ ;
  assign \new_[75372]_  = A167 & A168;
  assign \new_[75373]_  = ~A170 & \new_[75372]_ ;
  assign \new_[75376]_  = ~A199 & ~A166;
  assign \new_[75379]_  = ~A201 & A200;
  assign \new_[75380]_  = \new_[75379]_  & \new_[75376]_ ;
  assign \new_[75381]_  = \new_[75380]_  & \new_[75373]_ ;
  assign \new_[75384]_  = ~A203 & ~A202;
  assign \new_[75387]_  = A266 & ~A265;
  assign \new_[75388]_  = \new_[75387]_  & \new_[75384]_ ;
  assign \new_[75391]_  = A269 & A267;
  assign \new_[75394]_  = A302 & ~A300;
  assign \new_[75395]_  = \new_[75394]_  & \new_[75391]_ ;
  assign \new_[75396]_  = \new_[75395]_  & \new_[75388]_ ;
  assign \new_[75400]_  = A167 & A168;
  assign \new_[75401]_  = ~A170 & \new_[75400]_ ;
  assign \new_[75404]_  = ~A199 & ~A166;
  assign \new_[75407]_  = ~A201 & A200;
  assign \new_[75408]_  = \new_[75407]_  & \new_[75404]_ ;
  assign \new_[75409]_  = \new_[75408]_  & \new_[75401]_ ;
  assign \new_[75412]_  = ~A203 & ~A202;
  assign \new_[75415]_  = A266 & ~A265;
  assign \new_[75416]_  = \new_[75415]_  & \new_[75412]_ ;
  assign \new_[75419]_  = A269 & A267;
  assign \new_[75422]_  = A299 & A298;
  assign \new_[75423]_  = \new_[75422]_  & \new_[75419]_ ;
  assign \new_[75424]_  = \new_[75423]_  & \new_[75416]_ ;
  assign \new_[75428]_  = A167 & A168;
  assign \new_[75429]_  = ~A170 & \new_[75428]_ ;
  assign \new_[75432]_  = ~A199 & ~A166;
  assign \new_[75435]_  = ~A201 & A200;
  assign \new_[75436]_  = \new_[75435]_  & \new_[75432]_ ;
  assign \new_[75437]_  = \new_[75436]_  & \new_[75429]_ ;
  assign \new_[75440]_  = ~A203 & ~A202;
  assign \new_[75443]_  = A266 & ~A265;
  assign \new_[75444]_  = \new_[75443]_  & \new_[75440]_ ;
  assign \new_[75447]_  = A269 & A267;
  assign \new_[75450]_  = ~A299 & ~A298;
  assign \new_[75451]_  = \new_[75450]_  & \new_[75447]_ ;
  assign \new_[75452]_  = \new_[75451]_  & \new_[75444]_ ;
  assign \new_[75456]_  = A167 & A168;
  assign \new_[75457]_  = ~A170 & \new_[75456]_ ;
  assign \new_[75460]_  = ~A199 & ~A166;
  assign \new_[75463]_  = ~A201 & A200;
  assign \new_[75464]_  = \new_[75463]_  & \new_[75460]_ ;
  assign \new_[75465]_  = \new_[75464]_  & \new_[75457]_ ;
  assign \new_[75468]_  = ~A203 & ~A202;
  assign \new_[75471]_  = ~A266 & A265;
  assign \new_[75472]_  = \new_[75471]_  & \new_[75468]_ ;
  assign \new_[75475]_  = A268 & A267;
  assign \new_[75478]_  = A301 & ~A300;
  assign \new_[75479]_  = \new_[75478]_  & \new_[75475]_ ;
  assign \new_[75480]_  = \new_[75479]_  & \new_[75472]_ ;
  assign \new_[75484]_  = A167 & A168;
  assign \new_[75485]_  = ~A170 & \new_[75484]_ ;
  assign \new_[75488]_  = ~A199 & ~A166;
  assign \new_[75491]_  = ~A201 & A200;
  assign \new_[75492]_  = \new_[75491]_  & \new_[75488]_ ;
  assign \new_[75493]_  = \new_[75492]_  & \new_[75485]_ ;
  assign \new_[75496]_  = ~A203 & ~A202;
  assign \new_[75499]_  = ~A266 & A265;
  assign \new_[75500]_  = \new_[75499]_  & \new_[75496]_ ;
  assign \new_[75503]_  = A268 & A267;
  assign \new_[75506]_  = A302 & ~A300;
  assign \new_[75507]_  = \new_[75506]_  & \new_[75503]_ ;
  assign \new_[75508]_  = \new_[75507]_  & \new_[75500]_ ;
  assign \new_[75512]_  = A167 & A168;
  assign \new_[75513]_  = ~A170 & \new_[75512]_ ;
  assign \new_[75516]_  = ~A199 & ~A166;
  assign \new_[75519]_  = ~A201 & A200;
  assign \new_[75520]_  = \new_[75519]_  & \new_[75516]_ ;
  assign \new_[75521]_  = \new_[75520]_  & \new_[75513]_ ;
  assign \new_[75524]_  = ~A203 & ~A202;
  assign \new_[75527]_  = ~A266 & A265;
  assign \new_[75528]_  = \new_[75527]_  & \new_[75524]_ ;
  assign \new_[75531]_  = A268 & A267;
  assign \new_[75534]_  = A299 & A298;
  assign \new_[75535]_  = \new_[75534]_  & \new_[75531]_ ;
  assign \new_[75536]_  = \new_[75535]_  & \new_[75528]_ ;
  assign \new_[75540]_  = A167 & A168;
  assign \new_[75541]_  = ~A170 & \new_[75540]_ ;
  assign \new_[75544]_  = ~A199 & ~A166;
  assign \new_[75547]_  = ~A201 & A200;
  assign \new_[75548]_  = \new_[75547]_  & \new_[75544]_ ;
  assign \new_[75549]_  = \new_[75548]_  & \new_[75541]_ ;
  assign \new_[75552]_  = ~A203 & ~A202;
  assign \new_[75555]_  = ~A266 & A265;
  assign \new_[75556]_  = \new_[75555]_  & \new_[75552]_ ;
  assign \new_[75559]_  = A268 & A267;
  assign \new_[75562]_  = ~A299 & ~A298;
  assign \new_[75563]_  = \new_[75562]_  & \new_[75559]_ ;
  assign \new_[75564]_  = \new_[75563]_  & \new_[75556]_ ;
  assign \new_[75568]_  = A167 & A168;
  assign \new_[75569]_  = ~A170 & \new_[75568]_ ;
  assign \new_[75572]_  = ~A199 & ~A166;
  assign \new_[75575]_  = ~A201 & A200;
  assign \new_[75576]_  = \new_[75575]_  & \new_[75572]_ ;
  assign \new_[75577]_  = \new_[75576]_  & \new_[75569]_ ;
  assign \new_[75580]_  = ~A203 & ~A202;
  assign \new_[75583]_  = ~A266 & A265;
  assign \new_[75584]_  = \new_[75583]_  & \new_[75580]_ ;
  assign \new_[75587]_  = A269 & A267;
  assign \new_[75590]_  = A301 & ~A300;
  assign \new_[75591]_  = \new_[75590]_  & \new_[75587]_ ;
  assign \new_[75592]_  = \new_[75591]_  & \new_[75584]_ ;
  assign \new_[75596]_  = A167 & A168;
  assign \new_[75597]_  = ~A170 & \new_[75596]_ ;
  assign \new_[75600]_  = ~A199 & ~A166;
  assign \new_[75603]_  = ~A201 & A200;
  assign \new_[75604]_  = \new_[75603]_  & \new_[75600]_ ;
  assign \new_[75605]_  = \new_[75604]_  & \new_[75597]_ ;
  assign \new_[75608]_  = ~A203 & ~A202;
  assign \new_[75611]_  = ~A266 & A265;
  assign \new_[75612]_  = \new_[75611]_  & \new_[75608]_ ;
  assign \new_[75615]_  = A269 & A267;
  assign \new_[75618]_  = A302 & ~A300;
  assign \new_[75619]_  = \new_[75618]_  & \new_[75615]_ ;
  assign \new_[75620]_  = \new_[75619]_  & \new_[75612]_ ;
  assign \new_[75624]_  = A167 & A168;
  assign \new_[75625]_  = ~A170 & \new_[75624]_ ;
  assign \new_[75628]_  = ~A199 & ~A166;
  assign \new_[75631]_  = ~A201 & A200;
  assign \new_[75632]_  = \new_[75631]_  & \new_[75628]_ ;
  assign \new_[75633]_  = \new_[75632]_  & \new_[75625]_ ;
  assign \new_[75636]_  = ~A203 & ~A202;
  assign \new_[75639]_  = ~A266 & A265;
  assign \new_[75640]_  = \new_[75639]_  & \new_[75636]_ ;
  assign \new_[75643]_  = A269 & A267;
  assign \new_[75646]_  = A299 & A298;
  assign \new_[75647]_  = \new_[75646]_  & \new_[75643]_ ;
  assign \new_[75648]_  = \new_[75647]_  & \new_[75640]_ ;
  assign \new_[75652]_  = A167 & A168;
  assign \new_[75653]_  = ~A170 & \new_[75652]_ ;
  assign \new_[75656]_  = ~A199 & ~A166;
  assign \new_[75659]_  = ~A201 & A200;
  assign \new_[75660]_  = \new_[75659]_  & \new_[75656]_ ;
  assign \new_[75661]_  = \new_[75660]_  & \new_[75653]_ ;
  assign \new_[75664]_  = ~A203 & ~A202;
  assign \new_[75667]_  = ~A266 & A265;
  assign \new_[75668]_  = \new_[75667]_  & \new_[75664]_ ;
  assign \new_[75671]_  = A269 & A267;
  assign \new_[75674]_  = ~A299 & ~A298;
  assign \new_[75675]_  = \new_[75674]_  & \new_[75671]_ ;
  assign \new_[75676]_  = \new_[75675]_  & \new_[75668]_ ;
  assign \new_[75680]_  = A167 & A168;
  assign \new_[75681]_  = ~A170 & \new_[75680]_ ;
  assign \new_[75684]_  = A199 & ~A166;
  assign \new_[75687]_  = A201 & ~A200;
  assign \new_[75688]_  = \new_[75687]_  & \new_[75684]_ ;
  assign \new_[75689]_  = \new_[75688]_  & \new_[75681]_ ;
  assign \new_[75692]_  = ~A265 & A202;
  assign \new_[75695]_  = A267 & A266;
  assign \new_[75696]_  = \new_[75695]_  & \new_[75692]_ ;
  assign \new_[75699]_  = A300 & A268;
  assign \new_[75702]_  = ~A302 & ~A301;
  assign \new_[75703]_  = \new_[75702]_  & \new_[75699]_ ;
  assign \new_[75704]_  = \new_[75703]_  & \new_[75696]_ ;
  assign \new_[75708]_  = A167 & A168;
  assign \new_[75709]_  = ~A170 & \new_[75708]_ ;
  assign \new_[75712]_  = A199 & ~A166;
  assign \new_[75715]_  = A201 & ~A200;
  assign \new_[75716]_  = \new_[75715]_  & \new_[75712]_ ;
  assign \new_[75717]_  = \new_[75716]_  & \new_[75709]_ ;
  assign \new_[75720]_  = ~A265 & A202;
  assign \new_[75723]_  = A267 & A266;
  assign \new_[75724]_  = \new_[75723]_  & \new_[75720]_ ;
  assign \new_[75727]_  = A300 & A269;
  assign \new_[75730]_  = ~A302 & ~A301;
  assign \new_[75731]_  = \new_[75730]_  & \new_[75727]_ ;
  assign \new_[75732]_  = \new_[75731]_  & \new_[75724]_ ;
  assign \new_[75736]_  = A167 & A168;
  assign \new_[75737]_  = ~A170 & \new_[75736]_ ;
  assign \new_[75740]_  = A199 & ~A166;
  assign \new_[75743]_  = A201 & ~A200;
  assign \new_[75744]_  = \new_[75743]_  & \new_[75740]_ ;
  assign \new_[75745]_  = \new_[75744]_  & \new_[75737]_ ;
  assign \new_[75748]_  = ~A265 & A202;
  assign \new_[75751]_  = ~A267 & A266;
  assign \new_[75752]_  = \new_[75751]_  & \new_[75748]_ ;
  assign \new_[75755]_  = ~A269 & ~A268;
  assign \new_[75758]_  = A301 & ~A300;
  assign \new_[75759]_  = \new_[75758]_  & \new_[75755]_ ;
  assign \new_[75760]_  = \new_[75759]_  & \new_[75752]_ ;
  assign \new_[75764]_  = A167 & A168;
  assign \new_[75765]_  = ~A170 & \new_[75764]_ ;
  assign \new_[75768]_  = A199 & ~A166;
  assign \new_[75771]_  = A201 & ~A200;
  assign \new_[75772]_  = \new_[75771]_  & \new_[75768]_ ;
  assign \new_[75773]_  = \new_[75772]_  & \new_[75765]_ ;
  assign \new_[75776]_  = ~A265 & A202;
  assign \new_[75779]_  = ~A267 & A266;
  assign \new_[75780]_  = \new_[75779]_  & \new_[75776]_ ;
  assign \new_[75783]_  = ~A269 & ~A268;
  assign \new_[75786]_  = A302 & ~A300;
  assign \new_[75787]_  = \new_[75786]_  & \new_[75783]_ ;
  assign \new_[75788]_  = \new_[75787]_  & \new_[75780]_ ;
  assign \new_[75792]_  = A167 & A168;
  assign \new_[75793]_  = ~A170 & \new_[75792]_ ;
  assign \new_[75796]_  = A199 & ~A166;
  assign \new_[75799]_  = A201 & ~A200;
  assign \new_[75800]_  = \new_[75799]_  & \new_[75796]_ ;
  assign \new_[75801]_  = \new_[75800]_  & \new_[75793]_ ;
  assign \new_[75804]_  = ~A265 & A202;
  assign \new_[75807]_  = ~A267 & A266;
  assign \new_[75808]_  = \new_[75807]_  & \new_[75804]_ ;
  assign \new_[75811]_  = ~A269 & ~A268;
  assign \new_[75814]_  = A299 & A298;
  assign \new_[75815]_  = \new_[75814]_  & \new_[75811]_ ;
  assign \new_[75816]_  = \new_[75815]_  & \new_[75808]_ ;
  assign \new_[75820]_  = A167 & A168;
  assign \new_[75821]_  = ~A170 & \new_[75820]_ ;
  assign \new_[75824]_  = A199 & ~A166;
  assign \new_[75827]_  = A201 & ~A200;
  assign \new_[75828]_  = \new_[75827]_  & \new_[75824]_ ;
  assign \new_[75829]_  = \new_[75828]_  & \new_[75821]_ ;
  assign \new_[75832]_  = ~A265 & A202;
  assign \new_[75835]_  = ~A267 & A266;
  assign \new_[75836]_  = \new_[75835]_  & \new_[75832]_ ;
  assign \new_[75839]_  = ~A269 & ~A268;
  assign \new_[75842]_  = ~A299 & ~A298;
  assign \new_[75843]_  = \new_[75842]_  & \new_[75839]_ ;
  assign \new_[75844]_  = \new_[75843]_  & \new_[75836]_ ;
  assign \new_[75848]_  = A167 & A168;
  assign \new_[75849]_  = ~A170 & \new_[75848]_ ;
  assign \new_[75852]_  = A199 & ~A166;
  assign \new_[75855]_  = A201 & ~A200;
  assign \new_[75856]_  = \new_[75855]_  & \new_[75852]_ ;
  assign \new_[75857]_  = \new_[75856]_  & \new_[75849]_ ;
  assign \new_[75860]_  = A265 & A202;
  assign \new_[75863]_  = A267 & ~A266;
  assign \new_[75864]_  = \new_[75863]_  & \new_[75860]_ ;
  assign \new_[75867]_  = A300 & A268;
  assign \new_[75870]_  = ~A302 & ~A301;
  assign \new_[75871]_  = \new_[75870]_  & \new_[75867]_ ;
  assign \new_[75872]_  = \new_[75871]_  & \new_[75864]_ ;
  assign \new_[75876]_  = A167 & A168;
  assign \new_[75877]_  = ~A170 & \new_[75876]_ ;
  assign \new_[75880]_  = A199 & ~A166;
  assign \new_[75883]_  = A201 & ~A200;
  assign \new_[75884]_  = \new_[75883]_  & \new_[75880]_ ;
  assign \new_[75885]_  = \new_[75884]_  & \new_[75877]_ ;
  assign \new_[75888]_  = A265 & A202;
  assign \new_[75891]_  = A267 & ~A266;
  assign \new_[75892]_  = \new_[75891]_  & \new_[75888]_ ;
  assign \new_[75895]_  = A300 & A269;
  assign \new_[75898]_  = ~A302 & ~A301;
  assign \new_[75899]_  = \new_[75898]_  & \new_[75895]_ ;
  assign \new_[75900]_  = \new_[75899]_  & \new_[75892]_ ;
  assign \new_[75904]_  = A167 & A168;
  assign \new_[75905]_  = ~A170 & \new_[75904]_ ;
  assign \new_[75908]_  = A199 & ~A166;
  assign \new_[75911]_  = A201 & ~A200;
  assign \new_[75912]_  = \new_[75911]_  & \new_[75908]_ ;
  assign \new_[75913]_  = \new_[75912]_  & \new_[75905]_ ;
  assign \new_[75916]_  = A265 & A202;
  assign \new_[75919]_  = ~A267 & ~A266;
  assign \new_[75920]_  = \new_[75919]_  & \new_[75916]_ ;
  assign \new_[75923]_  = ~A269 & ~A268;
  assign \new_[75926]_  = A301 & ~A300;
  assign \new_[75927]_  = \new_[75926]_  & \new_[75923]_ ;
  assign \new_[75928]_  = \new_[75927]_  & \new_[75920]_ ;
  assign \new_[75932]_  = A167 & A168;
  assign \new_[75933]_  = ~A170 & \new_[75932]_ ;
  assign \new_[75936]_  = A199 & ~A166;
  assign \new_[75939]_  = A201 & ~A200;
  assign \new_[75940]_  = \new_[75939]_  & \new_[75936]_ ;
  assign \new_[75941]_  = \new_[75940]_  & \new_[75933]_ ;
  assign \new_[75944]_  = A265 & A202;
  assign \new_[75947]_  = ~A267 & ~A266;
  assign \new_[75948]_  = \new_[75947]_  & \new_[75944]_ ;
  assign \new_[75951]_  = ~A269 & ~A268;
  assign \new_[75954]_  = A302 & ~A300;
  assign \new_[75955]_  = \new_[75954]_  & \new_[75951]_ ;
  assign \new_[75956]_  = \new_[75955]_  & \new_[75948]_ ;
  assign \new_[75960]_  = A167 & A168;
  assign \new_[75961]_  = ~A170 & \new_[75960]_ ;
  assign \new_[75964]_  = A199 & ~A166;
  assign \new_[75967]_  = A201 & ~A200;
  assign \new_[75968]_  = \new_[75967]_  & \new_[75964]_ ;
  assign \new_[75969]_  = \new_[75968]_  & \new_[75961]_ ;
  assign \new_[75972]_  = A265 & A202;
  assign \new_[75975]_  = ~A267 & ~A266;
  assign \new_[75976]_  = \new_[75975]_  & \new_[75972]_ ;
  assign \new_[75979]_  = ~A269 & ~A268;
  assign \new_[75982]_  = A299 & A298;
  assign \new_[75983]_  = \new_[75982]_  & \new_[75979]_ ;
  assign \new_[75984]_  = \new_[75983]_  & \new_[75976]_ ;
  assign \new_[75988]_  = A167 & A168;
  assign \new_[75989]_  = ~A170 & \new_[75988]_ ;
  assign \new_[75992]_  = A199 & ~A166;
  assign \new_[75995]_  = A201 & ~A200;
  assign \new_[75996]_  = \new_[75995]_  & \new_[75992]_ ;
  assign \new_[75997]_  = \new_[75996]_  & \new_[75989]_ ;
  assign \new_[76000]_  = A265 & A202;
  assign \new_[76003]_  = ~A267 & ~A266;
  assign \new_[76004]_  = \new_[76003]_  & \new_[76000]_ ;
  assign \new_[76007]_  = ~A269 & ~A268;
  assign \new_[76010]_  = ~A299 & ~A298;
  assign \new_[76011]_  = \new_[76010]_  & \new_[76007]_ ;
  assign \new_[76012]_  = \new_[76011]_  & \new_[76004]_ ;
  assign \new_[76016]_  = A167 & A168;
  assign \new_[76017]_  = ~A170 & \new_[76016]_ ;
  assign \new_[76020]_  = A199 & ~A166;
  assign \new_[76023]_  = A201 & ~A200;
  assign \new_[76024]_  = \new_[76023]_  & \new_[76020]_ ;
  assign \new_[76025]_  = \new_[76024]_  & \new_[76017]_ ;
  assign \new_[76028]_  = ~A265 & A203;
  assign \new_[76031]_  = A267 & A266;
  assign \new_[76032]_  = \new_[76031]_  & \new_[76028]_ ;
  assign \new_[76035]_  = A300 & A268;
  assign \new_[76038]_  = ~A302 & ~A301;
  assign \new_[76039]_  = \new_[76038]_  & \new_[76035]_ ;
  assign \new_[76040]_  = \new_[76039]_  & \new_[76032]_ ;
  assign \new_[76044]_  = A167 & A168;
  assign \new_[76045]_  = ~A170 & \new_[76044]_ ;
  assign \new_[76048]_  = A199 & ~A166;
  assign \new_[76051]_  = A201 & ~A200;
  assign \new_[76052]_  = \new_[76051]_  & \new_[76048]_ ;
  assign \new_[76053]_  = \new_[76052]_  & \new_[76045]_ ;
  assign \new_[76056]_  = ~A265 & A203;
  assign \new_[76059]_  = A267 & A266;
  assign \new_[76060]_  = \new_[76059]_  & \new_[76056]_ ;
  assign \new_[76063]_  = A300 & A269;
  assign \new_[76066]_  = ~A302 & ~A301;
  assign \new_[76067]_  = \new_[76066]_  & \new_[76063]_ ;
  assign \new_[76068]_  = \new_[76067]_  & \new_[76060]_ ;
  assign \new_[76072]_  = A167 & A168;
  assign \new_[76073]_  = ~A170 & \new_[76072]_ ;
  assign \new_[76076]_  = A199 & ~A166;
  assign \new_[76079]_  = A201 & ~A200;
  assign \new_[76080]_  = \new_[76079]_  & \new_[76076]_ ;
  assign \new_[76081]_  = \new_[76080]_  & \new_[76073]_ ;
  assign \new_[76084]_  = ~A265 & A203;
  assign \new_[76087]_  = ~A267 & A266;
  assign \new_[76088]_  = \new_[76087]_  & \new_[76084]_ ;
  assign \new_[76091]_  = ~A269 & ~A268;
  assign \new_[76094]_  = A301 & ~A300;
  assign \new_[76095]_  = \new_[76094]_  & \new_[76091]_ ;
  assign \new_[76096]_  = \new_[76095]_  & \new_[76088]_ ;
  assign \new_[76100]_  = A167 & A168;
  assign \new_[76101]_  = ~A170 & \new_[76100]_ ;
  assign \new_[76104]_  = A199 & ~A166;
  assign \new_[76107]_  = A201 & ~A200;
  assign \new_[76108]_  = \new_[76107]_  & \new_[76104]_ ;
  assign \new_[76109]_  = \new_[76108]_  & \new_[76101]_ ;
  assign \new_[76112]_  = ~A265 & A203;
  assign \new_[76115]_  = ~A267 & A266;
  assign \new_[76116]_  = \new_[76115]_  & \new_[76112]_ ;
  assign \new_[76119]_  = ~A269 & ~A268;
  assign \new_[76122]_  = A302 & ~A300;
  assign \new_[76123]_  = \new_[76122]_  & \new_[76119]_ ;
  assign \new_[76124]_  = \new_[76123]_  & \new_[76116]_ ;
  assign \new_[76128]_  = A167 & A168;
  assign \new_[76129]_  = ~A170 & \new_[76128]_ ;
  assign \new_[76132]_  = A199 & ~A166;
  assign \new_[76135]_  = A201 & ~A200;
  assign \new_[76136]_  = \new_[76135]_  & \new_[76132]_ ;
  assign \new_[76137]_  = \new_[76136]_  & \new_[76129]_ ;
  assign \new_[76140]_  = ~A265 & A203;
  assign \new_[76143]_  = ~A267 & A266;
  assign \new_[76144]_  = \new_[76143]_  & \new_[76140]_ ;
  assign \new_[76147]_  = ~A269 & ~A268;
  assign \new_[76150]_  = A299 & A298;
  assign \new_[76151]_  = \new_[76150]_  & \new_[76147]_ ;
  assign \new_[76152]_  = \new_[76151]_  & \new_[76144]_ ;
  assign \new_[76156]_  = A167 & A168;
  assign \new_[76157]_  = ~A170 & \new_[76156]_ ;
  assign \new_[76160]_  = A199 & ~A166;
  assign \new_[76163]_  = A201 & ~A200;
  assign \new_[76164]_  = \new_[76163]_  & \new_[76160]_ ;
  assign \new_[76165]_  = \new_[76164]_  & \new_[76157]_ ;
  assign \new_[76168]_  = ~A265 & A203;
  assign \new_[76171]_  = ~A267 & A266;
  assign \new_[76172]_  = \new_[76171]_  & \new_[76168]_ ;
  assign \new_[76175]_  = ~A269 & ~A268;
  assign \new_[76178]_  = ~A299 & ~A298;
  assign \new_[76179]_  = \new_[76178]_  & \new_[76175]_ ;
  assign \new_[76180]_  = \new_[76179]_  & \new_[76172]_ ;
  assign \new_[76184]_  = A167 & A168;
  assign \new_[76185]_  = ~A170 & \new_[76184]_ ;
  assign \new_[76188]_  = A199 & ~A166;
  assign \new_[76191]_  = A201 & ~A200;
  assign \new_[76192]_  = \new_[76191]_  & \new_[76188]_ ;
  assign \new_[76193]_  = \new_[76192]_  & \new_[76185]_ ;
  assign \new_[76196]_  = A265 & A203;
  assign \new_[76199]_  = A267 & ~A266;
  assign \new_[76200]_  = \new_[76199]_  & \new_[76196]_ ;
  assign \new_[76203]_  = A300 & A268;
  assign \new_[76206]_  = ~A302 & ~A301;
  assign \new_[76207]_  = \new_[76206]_  & \new_[76203]_ ;
  assign \new_[76208]_  = \new_[76207]_  & \new_[76200]_ ;
  assign \new_[76212]_  = A167 & A168;
  assign \new_[76213]_  = ~A170 & \new_[76212]_ ;
  assign \new_[76216]_  = A199 & ~A166;
  assign \new_[76219]_  = A201 & ~A200;
  assign \new_[76220]_  = \new_[76219]_  & \new_[76216]_ ;
  assign \new_[76221]_  = \new_[76220]_  & \new_[76213]_ ;
  assign \new_[76224]_  = A265 & A203;
  assign \new_[76227]_  = A267 & ~A266;
  assign \new_[76228]_  = \new_[76227]_  & \new_[76224]_ ;
  assign \new_[76231]_  = A300 & A269;
  assign \new_[76234]_  = ~A302 & ~A301;
  assign \new_[76235]_  = \new_[76234]_  & \new_[76231]_ ;
  assign \new_[76236]_  = \new_[76235]_  & \new_[76228]_ ;
  assign \new_[76240]_  = A167 & A168;
  assign \new_[76241]_  = ~A170 & \new_[76240]_ ;
  assign \new_[76244]_  = A199 & ~A166;
  assign \new_[76247]_  = A201 & ~A200;
  assign \new_[76248]_  = \new_[76247]_  & \new_[76244]_ ;
  assign \new_[76249]_  = \new_[76248]_  & \new_[76241]_ ;
  assign \new_[76252]_  = A265 & A203;
  assign \new_[76255]_  = ~A267 & ~A266;
  assign \new_[76256]_  = \new_[76255]_  & \new_[76252]_ ;
  assign \new_[76259]_  = ~A269 & ~A268;
  assign \new_[76262]_  = A301 & ~A300;
  assign \new_[76263]_  = \new_[76262]_  & \new_[76259]_ ;
  assign \new_[76264]_  = \new_[76263]_  & \new_[76256]_ ;
  assign \new_[76268]_  = A167 & A168;
  assign \new_[76269]_  = ~A170 & \new_[76268]_ ;
  assign \new_[76272]_  = A199 & ~A166;
  assign \new_[76275]_  = A201 & ~A200;
  assign \new_[76276]_  = \new_[76275]_  & \new_[76272]_ ;
  assign \new_[76277]_  = \new_[76276]_  & \new_[76269]_ ;
  assign \new_[76280]_  = A265 & A203;
  assign \new_[76283]_  = ~A267 & ~A266;
  assign \new_[76284]_  = \new_[76283]_  & \new_[76280]_ ;
  assign \new_[76287]_  = ~A269 & ~A268;
  assign \new_[76290]_  = A302 & ~A300;
  assign \new_[76291]_  = \new_[76290]_  & \new_[76287]_ ;
  assign \new_[76292]_  = \new_[76291]_  & \new_[76284]_ ;
  assign \new_[76296]_  = A167 & A168;
  assign \new_[76297]_  = ~A170 & \new_[76296]_ ;
  assign \new_[76300]_  = A199 & ~A166;
  assign \new_[76303]_  = A201 & ~A200;
  assign \new_[76304]_  = \new_[76303]_  & \new_[76300]_ ;
  assign \new_[76305]_  = \new_[76304]_  & \new_[76297]_ ;
  assign \new_[76308]_  = A265 & A203;
  assign \new_[76311]_  = ~A267 & ~A266;
  assign \new_[76312]_  = \new_[76311]_  & \new_[76308]_ ;
  assign \new_[76315]_  = ~A269 & ~A268;
  assign \new_[76318]_  = A299 & A298;
  assign \new_[76319]_  = \new_[76318]_  & \new_[76315]_ ;
  assign \new_[76320]_  = \new_[76319]_  & \new_[76312]_ ;
  assign \new_[76324]_  = A167 & A168;
  assign \new_[76325]_  = ~A170 & \new_[76324]_ ;
  assign \new_[76328]_  = A199 & ~A166;
  assign \new_[76331]_  = A201 & ~A200;
  assign \new_[76332]_  = \new_[76331]_  & \new_[76328]_ ;
  assign \new_[76333]_  = \new_[76332]_  & \new_[76325]_ ;
  assign \new_[76336]_  = A265 & A203;
  assign \new_[76339]_  = ~A267 & ~A266;
  assign \new_[76340]_  = \new_[76339]_  & \new_[76336]_ ;
  assign \new_[76343]_  = ~A269 & ~A268;
  assign \new_[76346]_  = ~A299 & ~A298;
  assign \new_[76347]_  = \new_[76346]_  & \new_[76343]_ ;
  assign \new_[76348]_  = \new_[76347]_  & \new_[76340]_ ;
  assign \new_[76352]_  = A167 & A168;
  assign \new_[76353]_  = ~A170 & \new_[76352]_ ;
  assign \new_[76356]_  = A199 & ~A166;
  assign \new_[76359]_  = ~A201 & ~A200;
  assign \new_[76360]_  = \new_[76359]_  & \new_[76356]_ ;
  assign \new_[76361]_  = \new_[76360]_  & \new_[76353]_ ;
  assign \new_[76364]_  = ~A203 & ~A202;
  assign \new_[76367]_  = A266 & ~A265;
  assign \new_[76368]_  = \new_[76367]_  & \new_[76364]_ ;
  assign \new_[76371]_  = A268 & A267;
  assign \new_[76374]_  = A301 & ~A300;
  assign \new_[76375]_  = \new_[76374]_  & \new_[76371]_ ;
  assign \new_[76376]_  = \new_[76375]_  & \new_[76368]_ ;
  assign \new_[76380]_  = A167 & A168;
  assign \new_[76381]_  = ~A170 & \new_[76380]_ ;
  assign \new_[76384]_  = A199 & ~A166;
  assign \new_[76387]_  = ~A201 & ~A200;
  assign \new_[76388]_  = \new_[76387]_  & \new_[76384]_ ;
  assign \new_[76389]_  = \new_[76388]_  & \new_[76381]_ ;
  assign \new_[76392]_  = ~A203 & ~A202;
  assign \new_[76395]_  = A266 & ~A265;
  assign \new_[76396]_  = \new_[76395]_  & \new_[76392]_ ;
  assign \new_[76399]_  = A268 & A267;
  assign \new_[76402]_  = A302 & ~A300;
  assign \new_[76403]_  = \new_[76402]_  & \new_[76399]_ ;
  assign \new_[76404]_  = \new_[76403]_  & \new_[76396]_ ;
  assign \new_[76408]_  = A167 & A168;
  assign \new_[76409]_  = ~A170 & \new_[76408]_ ;
  assign \new_[76412]_  = A199 & ~A166;
  assign \new_[76415]_  = ~A201 & ~A200;
  assign \new_[76416]_  = \new_[76415]_  & \new_[76412]_ ;
  assign \new_[76417]_  = \new_[76416]_  & \new_[76409]_ ;
  assign \new_[76420]_  = ~A203 & ~A202;
  assign \new_[76423]_  = A266 & ~A265;
  assign \new_[76424]_  = \new_[76423]_  & \new_[76420]_ ;
  assign \new_[76427]_  = A268 & A267;
  assign \new_[76430]_  = A299 & A298;
  assign \new_[76431]_  = \new_[76430]_  & \new_[76427]_ ;
  assign \new_[76432]_  = \new_[76431]_  & \new_[76424]_ ;
  assign \new_[76436]_  = A167 & A168;
  assign \new_[76437]_  = ~A170 & \new_[76436]_ ;
  assign \new_[76440]_  = A199 & ~A166;
  assign \new_[76443]_  = ~A201 & ~A200;
  assign \new_[76444]_  = \new_[76443]_  & \new_[76440]_ ;
  assign \new_[76445]_  = \new_[76444]_  & \new_[76437]_ ;
  assign \new_[76448]_  = ~A203 & ~A202;
  assign \new_[76451]_  = A266 & ~A265;
  assign \new_[76452]_  = \new_[76451]_  & \new_[76448]_ ;
  assign \new_[76455]_  = A268 & A267;
  assign \new_[76458]_  = ~A299 & ~A298;
  assign \new_[76459]_  = \new_[76458]_  & \new_[76455]_ ;
  assign \new_[76460]_  = \new_[76459]_  & \new_[76452]_ ;
  assign \new_[76464]_  = A167 & A168;
  assign \new_[76465]_  = ~A170 & \new_[76464]_ ;
  assign \new_[76468]_  = A199 & ~A166;
  assign \new_[76471]_  = ~A201 & ~A200;
  assign \new_[76472]_  = \new_[76471]_  & \new_[76468]_ ;
  assign \new_[76473]_  = \new_[76472]_  & \new_[76465]_ ;
  assign \new_[76476]_  = ~A203 & ~A202;
  assign \new_[76479]_  = A266 & ~A265;
  assign \new_[76480]_  = \new_[76479]_  & \new_[76476]_ ;
  assign \new_[76483]_  = A269 & A267;
  assign \new_[76486]_  = A301 & ~A300;
  assign \new_[76487]_  = \new_[76486]_  & \new_[76483]_ ;
  assign \new_[76488]_  = \new_[76487]_  & \new_[76480]_ ;
  assign \new_[76492]_  = A167 & A168;
  assign \new_[76493]_  = ~A170 & \new_[76492]_ ;
  assign \new_[76496]_  = A199 & ~A166;
  assign \new_[76499]_  = ~A201 & ~A200;
  assign \new_[76500]_  = \new_[76499]_  & \new_[76496]_ ;
  assign \new_[76501]_  = \new_[76500]_  & \new_[76493]_ ;
  assign \new_[76504]_  = ~A203 & ~A202;
  assign \new_[76507]_  = A266 & ~A265;
  assign \new_[76508]_  = \new_[76507]_  & \new_[76504]_ ;
  assign \new_[76511]_  = A269 & A267;
  assign \new_[76514]_  = A302 & ~A300;
  assign \new_[76515]_  = \new_[76514]_  & \new_[76511]_ ;
  assign \new_[76516]_  = \new_[76515]_  & \new_[76508]_ ;
  assign \new_[76520]_  = A167 & A168;
  assign \new_[76521]_  = ~A170 & \new_[76520]_ ;
  assign \new_[76524]_  = A199 & ~A166;
  assign \new_[76527]_  = ~A201 & ~A200;
  assign \new_[76528]_  = \new_[76527]_  & \new_[76524]_ ;
  assign \new_[76529]_  = \new_[76528]_  & \new_[76521]_ ;
  assign \new_[76532]_  = ~A203 & ~A202;
  assign \new_[76535]_  = A266 & ~A265;
  assign \new_[76536]_  = \new_[76535]_  & \new_[76532]_ ;
  assign \new_[76539]_  = A269 & A267;
  assign \new_[76542]_  = A299 & A298;
  assign \new_[76543]_  = \new_[76542]_  & \new_[76539]_ ;
  assign \new_[76544]_  = \new_[76543]_  & \new_[76536]_ ;
  assign \new_[76548]_  = A167 & A168;
  assign \new_[76549]_  = ~A170 & \new_[76548]_ ;
  assign \new_[76552]_  = A199 & ~A166;
  assign \new_[76555]_  = ~A201 & ~A200;
  assign \new_[76556]_  = \new_[76555]_  & \new_[76552]_ ;
  assign \new_[76557]_  = \new_[76556]_  & \new_[76549]_ ;
  assign \new_[76560]_  = ~A203 & ~A202;
  assign \new_[76563]_  = A266 & ~A265;
  assign \new_[76564]_  = \new_[76563]_  & \new_[76560]_ ;
  assign \new_[76567]_  = A269 & A267;
  assign \new_[76570]_  = ~A299 & ~A298;
  assign \new_[76571]_  = \new_[76570]_  & \new_[76567]_ ;
  assign \new_[76572]_  = \new_[76571]_  & \new_[76564]_ ;
  assign \new_[76576]_  = A167 & A168;
  assign \new_[76577]_  = ~A170 & \new_[76576]_ ;
  assign \new_[76580]_  = A199 & ~A166;
  assign \new_[76583]_  = ~A201 & ~A200;
  assign \new_[76584]_  = \new_[76583]_  & \new_[76580]_ ;
  assign \new_[76585]_  = \new_[76584]_  & \new_[76577]_ ;
  assign \new_[76588]_  = ~A203 & ~A202;
  assign \new_[76591]_  = ~A266 & A265;
  assign \new_[76592]_  = \new_[76591]_  & \new_[76588]_ ;
  assign \new_[76595]_  = A268 & A267;
  assign \new_[76598]_  = A301 & ~A300;
  assign \new_[76599]_  = \new_[76598]_  & \new_[76595]_ ;
  assign \new_[76600]_  = \new_[76599]_  & \new_[76592]_ ;
  assign \new_[76604]_  = A167 & A168;
  assign \new_[76605]_  = ~A170 & \new_[76604]_ ;
  assign \new_[76608]_  = A199 & ~A166;
  assign \new_[76611]_  = ~A201 & ~A200;
  assign \new_[76612]_  = \new_[76611]_  & \new_[76608]_ ;
  assign \new_[76613]_  = \new_[76612]_  & \new_[76605]_ ;
  assign \new_[76616]_  = ~A203 & ~A202;
  assign \new_[76619]_  = ~A266 & A265;
  assign \new_[76620]_  = \new_[76619]_  & \new_[76616]_ ;
  assign \new_[76623]_  = A268 & A267;
  assign \new_[76626]_  = A302 & ~A300;
  assign \new_[76627]_  = \new_[76626]_  & \new_[76623]_ ;
  assign \new_[76628]_  = \new_[76627]_  & \new_[76620]_ ;
  assign \new_[76632]_  = A167 & A168;
  assign \new_[76633]_  = ~A170 & \new_[76632]_ ;
  assign \new_[76636]_  = A199 & ~A166;
  assign \new_[76639]_  = ~A201 & ~A200;
  assign \new_[76640]_  = \new_[76639]_  & \new_[76636]_ ;
  assign \new_[76641]_  = \new_[76640]_  & \new_[76633]_ ;
  assign \new_[76644]_  = ~A203 & ~A202;
  assign \new_[76647]_  = ~A266 & A265;
  assign \new_[76648]_  = \new_[76647]_  & \new_[76644]_ ;
  assign \new_[76651]_  = A268 & A267;
  assign \new_[76654]_  = A299 & A298;
  assign \new_[76655]_  = \new_[76654]_  & \new_[76651]_ ;
  assign \new_[76656]_  = \new_[76655]_  & \new_[76648]_ ;
  assign \new_[76660]_  = A167 & A168;
  assign \new_[76661]_  = ~A170 & \new_[76660]_ ;
  assign \new_[76664]_  = A199 & ~A166;
  assign \new_[76667]_  = ~A201 & ~A200;
  assign \new_[76668]_  = \new_[76667]_  & \new_[76664]_ ;
  assign \new_[76669]_  = \new_[76668]_  & \new_[76661]_ ;
  assign \new_[76672]_  = ~A203 & ~A202;
  assign \new_[76675]_  = ~A266 & A265;
  assign \new_[76676]_  = \new_[76675]_  & \new_[76672]_ ;
  assign \new_[76679]_  = A268 & A267;
  assign \new_[76682]_  = ~A299 & ~A298;
  assign \new_[76683]_  = \new_[76682]_  & \new_[76679]_ ;
  assign \new_[76684]_  = \new_[76683]_  & \new_[76676]_ ;
  assign \new_[76688]_  = A167 & A168;
  assign \new_[76689]_  = ~A170 & \new_[76688]_ ;
  assign \new_[76692]_  = A199 & ~A166;
  assign \new_[76695]_  = ~A201 & ~A200;
  assign \new_[76696]_  = \new_[76695]_  & \new_[76692]_ ;
  assign \new_[76697]_  = \new_[76696]_  & \new_[76689]_ ;
  assign \new_[76700]_  = ~A203 & ~A202;
  assign \new_[76703]_  = ~A266 & A265;
  assign \new_[76704]_  = \new_[76703]_  & \new_[76700]_ ;
  assign \new_[76707]_  = A269 & A267;
  assign \new_[76710]_  = A301 & ~A300;
  assign \new_[76711]_  = \new_[76710]_  & \new_[76707]_ ;
  assign \new_[76712]_  = \new_[76711]_  & \new_[76704]_ ;
  assign \new_[76716]_  = A167 & A168;
  assign \new_[76717]_  = ~A170 & \new_[76716]_ ;
  assign \new_[76720]_  = A199 & ~A166;
  assign \new_[76723]_  = ~A201 & ~A200;
  assign \new_[76724]_  = \new_[76723]_  & \new_[76720]_ ;
  assign \new_[76725]_  = \new_[76724]_  & \new_[76717]_ ;
  assign \new_[76728]_  = ~A203 & ~A202;
  assign \new_[76731]_  = ~A266 & A265;
  assign \new_[76732]_  = \new_[76731]_  & \new_[76728]_ ;
  assign \new_[76735]_  = A269 & A267;
  assign \new_[76738]_  = A302 & ~A300;
  assign \new_[76739]_  = \new_[76738]_  & \new_[76735]_ ;
  assign \new_[76740]_  = \new_[76739]_  & \new_[76732]_ ;
  assign \new_[76744]_  = A167 & A168;
  assign \new_[76745]_  = ~A170 & \new_[76744]_ ;
  assign \new_[76748]_  = A199 & ~A166;
  assign \new_[76751]_  = ~A201 & ~A200;
  assign \new_[76752]_  = \new_[76751]_  & \new_[76748]_ ;
  assign \new_[76753]_  = \new_[76752]_  & \new_[76745]_ ;
  assign \new_[76756]_  = ~A203 & ~A202;
  assign \new_[76759]_  = ~A266 & A265;
  assign \new_[76760]_  = \new_[76759]_  & \new_[76756]_ ;
  assign \new_[76763]_  = A269 & A267;
  assign \new_[76766]_  = A299 & A298;
  assign \new_[76767]_  = \new_[76766]_  & \new_[76763]_ ;
  assign \new_[76768]_  = \new_[76767]_  & \new_[76760]_ ;
  assign \new_[76772]_  = A167 & A168;
  assign \new_[76773]_  = ~A170 & \new_[76772]_ ;
  assign \new_[76776]_  = A199 & ~A166;
  assign \new_[76779]_  = ~A201 & ~A200;
  assign \new_[76780]_  = \new_[76779]_  & \new_[76776]_ ;
  assign \new_[76781]_  = \new_[76780]_  & \new_[76773]_ ;
  assign \new_[76784]_  = ~A203 & ~A202;
  assign \new_[76787]_  = ~A266 & A265;
  assign \new_[76788]_  = \new_[76787]_  & \new_[76784]_ ;
  assign \new_[76791]_  = A269 & A267;
  assign \new_[76794]_  = ~A299 & ~A298;
  assign \new_[76795]_  = \new_[76794]_  & \new_[76791]_ ;
  assign \new_[76796]_  = \new_[76795]_  & \new_[76788]_ ;
  assign \new_[76800]_  = ~A167 & A168;
  assign \new_[76801]_  = ~A170 & \new_[76800]_ ;
  assign \new_[76804]_  = A201 & A166;
  assign \new_[76807]_  = ~A203 & ~A202;
  assign \new_[76808]_  = \new_[76807]_  & \new_[76804]_ ;
  assign \new_[76809]_  = \new_[76808]_  & \new_[76801]_ ;
  assign \new_[76812]_  = ~A268 & A267;
  assign \new_[76815]_  = A298 & ~A269;
  assign \new_[76816]_  = \new_[76815]_  & \new_[76812]_ ;
  assign \new_[76819]_  = ~A300 & ~A299;
  assign \new_[76822]_  = ~A302 & ~A301;
  assign \new_[76823]_  = \new_[76822]_  & \new_[76819]_ ;
  assign \new_[76824]_  = \new_[76823]_  & \new_[76816]_ ;
  assign \new_[76828]_  = ~A167 & A168;
  assign \new_[76829]_  = ~A170 & \new_[76828]_ ;
  assign \new_[76832]_  = A201 & A166;
  assign \new_[76835]_  = ~A203 & ~A202;
  assign \new_[76836]_  = \new_[76835]_  & \new_[76832]_ ;
  assign \new_[76837]_  = \new_[76836]_  & \new_[76829]_ ;
  assign \new_[76840]_  = ~A268 & A267;
  assign \new_[76843]_  = ~A298 & ~A269;
  assign \new_[76844]_  = \new_[76843]_  & \new_[76840]_ ;
  assign \new_[76847]_  = ~A300 & A299;
  assign \new_[76850]_  = ~A302 & ~A301;
  assign \new_[76851]_  = \new_[76850]_  & \new_[76847]_ ;
  assign \new_[76852]_  = \new_[76851]_  & \new_[76844]_ ;
  assign \new_[76856]_  = ~A167 & A168;
  assign \new_[76857]_  = ~A170 & \new_[76856]_ ;
  assign \new_[76860]_  = ~A199 & A166;
  assign \new_[76863]_  = A201 & A200;
  assign \new_[76864]_  = \new_[76863]_  & \new_[76860]_ ;
  assign \new_[76865]_  = \new_[76864]_  & \new_[76857]_ ;
  assign \new_[76868]_  = ~A265 & A202;
  assign \new_[76871]_  = A267 & A266;
  assign \new_[76872]_  = \new_[76871]_  & \new_[76868]_ ;
  assign \new_[76875]_  = A300 & A268;
  assign \new_[76878]_  = ~A302 & ~A301;
  assign \new_[76879]_  = \new_[76878]_  & \new_[76875]_ ;
  assign \new_[76880]_  = \new_[76879]_  & \new_[76872]_ ;
  assign \new_[76884]_  = ~A167 & A168;
  assign \new_[76885]_  = ~A170 & \new_[76884]_ ;
  assign \new_[76888]_  = ~A199 & A166;
  assign \new_[76891]_  = A201 & A200;
  assign \new_[76892]_  = \new_[76891]_  & \new_[76888]_ ;
  assign \new_[76893]_  = \new_[76892]_  & \new_[76885]_ ;
  assign \new_[76896]_  = ~A265 & A202;
  assign \new_[76899]_  = A267 & A266;
  assign \new_[76900]_  = \new_[76899]_  & \new_[76896]_ ;
  assign \new_[76903]_  = A300 & A269;
  assign \new_[76906]_  = ~A302 & ~A301;
  assign \new_[76907]_  = \new_[76906]_  & \new_[76903]_ ;
  assign \new_[76908]_  = \new_[76907]_  & \new_[76900]_ ;
  assign \new_[76912]_  = ~A167 & A168;
  assign \new_[76913]_  = ~A170 & \new_[76912]_ ;
  assign \new_[76916]_  = ~A199 & A166;
  assign \new_[76919]_  = A201 & A200;
  assign \new_[76920]_  = \new_[76919]_  & \new_[76916]_ ;
  assign \new_[76921]_  = \new_[76920]_  & \new_[76913]_ ;
  assign \new_[76924]_  = ~A265 & A202;
  assign \new_[76927]_  = ~A267 & A266;
  assign \new_[76928]_  = \new_[76927]_  & \new_[76924]_ ;
  assign \new_[76931]_  = ~A269 & ~A268;
  assign \new_[76934]_  = A301 & ~A300;
  assign \new_[76935]_  = \new_[76934]_  & \new_[76931]_ ;
  assign \new_[76936]_  = \new_[76935]_  & \new_[76928]_ ;
  assign \new_[76940]_  = ~A167 & A168;
  assign \new_[76941]_  = ~A170 & \new_[76940]_ ;
  assign \new_[76944]_  = ~A199 & A166;
  assign \new_[76947]_  = A201 & A200;
  assign \new_[76948]_  = \new_[76947]_  & \new_[76944]_ ;
  assign \new_[76949]_  = \new_[76948]_  & \new_[76941]_ ;
  assign \new_[76952]_  = ~A265 & A202;
  assign \new_[76955]_  = ~A267 & A266;
  assign \new_[76956]_  = \new_[76955]_  & \new_[76952]_ ;
  assign \new_[76959]_  = ~A269 & ~A268;
  assign \new_[76962]_  = A302 & ~A300;
  assign \new_[76963]_  = \new_[76962]_  & \new_[76959]_ ;
  assign \new_[76964]_  = \new_[76963]_  & \new_[76956]_ ;
  assign \new_[76968]_  = ~A167 & A168;
  assign \new_[76969]_  = ~A170 & \new_[76968]_ ;
  assign \new_[76972]_  = ~A199 & A166;
  assign \new_[76975]_  = A201 & A200;
  assign \new_[76976]_  = \new_[76975]_  & \new_[76972]_ ;
  assign \new_[76977]_  = \new_[76976]_  & \new_[76969]_ ;
  assign \new_[76980]_  = ~A265 & A202;
  assign \new_[76983]_  = ~A267 & A266;
  assign \new_[76984]_  = \new_[76983]_  & \new_[76980]_ ;
  assign \new_[76987]_  = ~A269 & ~A268;
  assign \new_[76990]_  = A299 & A298;
  assign \new_[76991]_  = \new_[76990]_  & \new_[76987]_ ;
  assign \new_[76992]_  = \new_[76991]_  & \new_[76984]_ ;
  assign \new_[76996]_  = ~A167 & A168;
  assign \new_[76997]_  = ~A170 & \new_[76996]_ ;
  assign \new_[77000]_  = ~A199 & A166;
  assign \new_[77003]_  = A201 & A200;
  assign \new_[77004]_  = \new_[77003]_  & \new_[77000]_ ;
  assign \new_[77005]_  = \new_[77004]_  & \new_[76997]_ ;
  assign \new_[77008]_  = ~A265 & A202;
  assign \new_[77011]_  = ~A267 & A266;
  assign \new_[77012]_  = \new_[77011]_  & \new_[77008]_ ;
  assign \new_[77015]_  = ~A269 & ~A268;
  assign \new_[77018]_  = ~A299 & ~A298;
  assign \new_[77019]_  = \new_[77018]_  & \new_[77015]_ ;
  assign \new_[77020]_  = \new_[77019]_  & \new_[77012]_ ;
  assign \new_[77024]_  = ~A167 & A168;
  assign \new_[77025]_  = ~A170 & \new_[77024]_ ;
  assign \new_[77028]_  = ~A199 & A166;
  assign \new_[77031]_  = A201 & A200;
  assign \new_[77032]_  = \new_[77031]_  & \new_[77028]_ ;
  assign \new_[77033]_  = \new_[77032]_  & \new_[77025]_ ;
  assign \new_[77036]_  = A265 & A202;
  assign \new_[77039]_  = A267 & ~A266;
  assign \new_[77040]_  = \new_[77039]_  & \new_[77036]_ ;
  assign \new_[77043]_  = A300 & A268;
  assign \new_[77046]_  = ~A302 & ~A301;
  assign \new_[77047]_  = \new_[77046]_  & \new_[77043]_ ;
  assign \new_[77048]_  = \new_[77047]_  & \new_[77040]_ ;
  assign \new_[77052]_  = ~A167 & A168;
  assign \new_[77053]_  = ~A170 & \new_[77052]_ ;
  assign \new_[77056]_  = ~A199 & A166;
  assign \new_[77059]_  = A201 & A200;
  assign \new_[77060]_  = \new_[77059]_  & \new_[77056]_ ;
  assign \new_[77061]_  = \new_[77060]_  & \new_[77053]_ ;
  assign \new_[77064]_  = A265 & A202;
  assign \new_[77067]_  = A267 & ~A266;
  assign \new_[77068]_  = \new_[77067]_  & \new_[77064]_ ;
  assign \new_[77071]_  = A300 & A269;
  assign \new_[77074]_  = ~A302 & ~A301;
  assign \new_[77075]_  = \new_[77074]_  & \new_[77071]_ ;
  assign \new_[77076]_  = \new_[77075]_  & \new_[77068]_ ;
  assign \new_[77080]_  = ~A167 & A168;
  assign \new_[77081]_  = ~A170 & \new_[77080]_ ;
  assign \new_[77084]_  = ~A199 & A166;
  assign \new_[77087]_  = A201 & A200;
  assign \new_[77088]_  = \new_[77087]_  & \new_[77084]_ ;
  assign \new_[77089]_  = \new_[77088]_  & \new_[77081]_ ;
  assign \new_[77092]_  = A265 & A202;
  assign \new_[77095]_  = ~A267 & ~A266;
  assign \new_[77096]_  = \new_[77095]_  & \new_[77092]_ ;
  assign \new_[77099]_  = ~A269 & ~A268;
  assign \new_[77102]_  = A301 & ~A300;
  assign \new_[77103]_  = \new_[77102]_  & \new_[77099]_ ;
  assign \new_[77104]_  = \new_[77103]_  & \new_[77096]_ ;
  assign \new_[77108]_  = ~A167 & A168;
  assign \new_[77109]_  = ~A170 & \new_[77108]_ ;
  assign \new_[77112]_  = ~A199 & A166;
  assign \new_[77115]_  = A201 & A200;
  assign \new_[77116]_  = \new_[77115]_  & \new_[77112]_ ;
  assign \new_[77117]_  = \new_[77116]_  & \new_[77109]_ ;
  assign \new_[77120]_  = A265 & A202;
  assign \new_[77123]_  = ~A267 & ~A266;
  assign \new_[77124]_  = \new_[77123]_  & \new_[77120]_ ;
  assign \new_[77127]_  = ~A269 & ~A268;
  assign \new_[77130]_  = A302 & ~A300;
  assign \new_[77131]_  = \new_[77130]_  & \new_[77127]_ ;
  assign \new_[77132]_  = \new_[77131]_  & \new_[77124]_ ;
  assign \new_[77136]_  = ~A167 & A168;
  assign \new_[77137]_  = ~A170 & \new_[77136]_ ;
  assign \new_[77140]_  = ~A199 & A166;
  assign \new_[77143]_  = A201 & A200;
  assign \new_[77144]_  = \new_[77143]_  & \new_[77140]_ ;
  assign \new_[77145]_  = \new_[77144]_  & \new_[77137]_ ;
  assign \new_[77148]_  = A265 & A202;
  assign \new_[77151]_  = ~A267 & ~A266;
  assign \new_[77152]_  = \new_[77151]_  & \new_[77148]_ ;
  assign \new_[77155]_  = ~A269 & ~A268;
  assign \new_[77158]_  = A299 & A298;
  assign \new_[77159]_  = \new_[77158]_  & \new_[77155]_ ;
  assign \new_[77160]_  = \new_[77159]_  & \new_[77152]_ ;
  assign \new_[77164]_  = ~A167 & A168;
  assign \new_[77165]_  = ~A170 & \new_[77164]_ ;
  assign \new_[77168]_  = ~A199 & A166;
  assign \new_[77171]_  = A201 & A200;
  assign \new_[77172]_  = \new_[77171]_  & \new_[77168]_ ;
  assign \new_[77173]_  = \new_[77172]_  & \new_[77165]_ ;
  assign \new_[77176]_  = A265 & A202;
  assign \new_[77179]_  = ~A267 & ~A266;
  assign \new_[77180]_  = \new_[77179]_  & \new_[77176]_ ;
  assign \new_[77183]_  = ~A269 & ~A268;
  assign \new_[77186]_  = ~A299 & ~A298;
  assign \new_[77187]_  = \new_[77186]_  & \new_[77183]_ ;
  assign \new_[77188]_  = \new_[77187]_  & \new_[77180]_ ;
  assign \new_[77192]_  = ~A167 & A168;
  assign \new_[77193]_  = ~A170 & \new_[77192]_ ;
  assign \new_[77196]_  = ~A199 & A166;
  assign \new_[77199]_  = A201 & A200;
  assign \new_[77200]_  = \new_[77199]_  & \new_[77196]_ ;
  assign \new_[77201]_  = \new_[77200]_  & \new_[77193]_ ;
  assign \new_[77204]_  = ~A265 & A203;
  assign \new_[77207]_  = A267 & A266;
  assign \new_[77208]_  = \new_[77207]_  & \new_[77204]_ ;
  assign \new_[77211]_  = A300 & A268;
  assign \new_[77214]_  = ~A302 & ~A301;
  assign \new_[77215]_  = \new_[77214]_  & \new_[77211]_ ;
  assign \new_[77216]_  = \new_[77215]_  & \new_[77208]_ ;
  assign \new_[77220]_  = ~A167 & A168;
  assign \new_[77221]_  = ~A170 & \new_[77220]_ ;
  assign \new_[77224]_  = ~A199 & A166;
  assign \new_[77227]_  = A201 & A200;
  assign \new_[77228]_  = \new_[77227]_  & \new_[77224]_ ;
  assign \new_[77229]_  = \new_[77228]_  & \new_[77221]_ ;
  assign \new_[77232]_  = ~A265 & A203;
  assign \new_[77235]_  = A267 & A266;
  assign \new_[77236]_  = \new_[77235]_  & \new_[77232]_ ;
  assign \new_[77239]_  = A300 & A269;
  assign \new_[77242]_  = ~A302 & ~A301;
  assign \new_[77243]_  = \new_[77242]_  & \new_[77239]_ ;
  assign \new_[77244]_  = \new_[77243]_  & \new_[77236]_ ;
  assign \new_[77248]_  = ~A167 & A168;
  assign \new_[77249]_  = ~A170 & \new_[77248]_ ;
  assign \new_[77252]_  = ~A199 & A166;
  assign \new_[77255]_  = A201 & A200;
  assign \new_[77256]_  = \new_[77255]_  & \new_[77252]_ ;
  assign \new_[77257]_  = \new_[77256]_  & \new_[77249]_ ;
  assign \new_[77260]_  = ~A265 & A203;
  assign \new_[77263]_  = ~A267 & A266;
  assign \new_[77264]_  = \new_[77263]_  & \new_[77260]_ ;
  assign \new_[77267]_  = ~A269 & ~A268;
  assign \new_[77270]_  = A301 & ~A300;
  assign \new_[77271]_  = \new_[77270]_  & \new_[77267]_ ;
  assign \new_[77272]_  = \new_[77271]_  & \new_[77264]_ ;
  assign \new_[77276]_  = ~A167 & A168;
  assign \new_[77277]_  = ~A170 & \new_[77276]_ ;
  assign \new_[77280]_  = ~A199 & A166;
  assign \new_[77283]_  = A201 & A200;
  assign \new_[77284]_  = \new_[77283]_  & \new_[77280]_ ;
  assign \new_[77285]_  = \new_[77284]_  & \new_[77277]_ ;
  assign \new_[77288]_  = ~A265 & A203;
  assign \new_[77291]_  = ~A267 & A266;
  assign \new_[77292]_  = \new_[77291]_  & \new_[77288]_ ;
  assign \new_[77295]_  = ~A269 & ~A268;
  assign \new_[77298]_  = A302 & ~A300;
  assign \new_[77299]_  = \new_[77298]_  & \new_[77295]_ ;
  assign \new_[77300]_  = \new_[77299]_  & \new_[77292]_ ;
  assign \new_[77304]_  = ~A167 & A168;
  assign \new_[77305]_  = ~A170 & \new_[77304]_ ;
  assign \new_[77308]_  = ~A199 & A166;
  assign \new_[77311]_  = A201 & A200;
  assign \new_[77312]_  = \new_[77311]_  & \new_[77308]_ ;
  assign \new_[77313]_  = \new_[77312]_  & \new_[77305]_ ;
  assign \new_[77316]_  = ~A265 & A203;
  assign \new_[77319]_  = ~A267 & A266;
  assign \new_[77320]_  = \new_[77319]_  & \new_[77316]_ ;
  assign \new_[77323]_  = ~A269 & ~A268;
  assign \new_[77326]_  = A299 & A298;
  assign \new_[77327]_  = \new_[77326]_  & \new_[77323]_ ;
  assign \new_[77328]_  = \new_[77327]_  & \new_[77320]_ ;
  assign \new_[77332]_  = ~A167 & A168;
  assign \new_[77333]_  = ~A170 & \new_[77332]_ ;
  assign \new_[77336]_  = ~A199 & A166;
  assign \new_[77339]_  = A201 & A200;
  assign \new_[77340]_  = \new_[77339]_  & \new_[77336]_ ;
  assign \new_[77341]_  = \new_[77340]_  & \new_[77333]_ ;
  assign \new_[77344]_  = ~A265 & A203;
  assign \new_[77347]_  = ~A267 & A266;
  assign \new_[77348]_  = \new_[77347]_  & \new_[77344]_ ;
  assign \new_[77351]_  = ~A269 & ~A268;
  assign \new_[77354]_  = ~A299 & ~A298;
  assign \new_[77355]_  = \new_[77354]_  & \new_[77351]_ ;
  assign \new_[77356]_  = \new_[77355]_  & \new_[77348]_ ;
  assign \new_[77360]_  = ~A167 & A168;
  assign \new_[77361]_  = ~A170 & \new_[77360]_ ;
  assign \new_[77364]_  = ~A199 & A166;
  assign \new_[77367]_  = A201 & A200;
  assign \new_[77368]_  = \new_[77367]_  & \new_[77364]_ ;
  assign \new_[77369]_  = \new_[77368]_  & \new_[77361]_ ;
  assign \new_[77372]_  = A265 & A203;
  assign \new_[77375]_  = A267 & ~A266;
  assign \new_[77376]_  = \new_[77375]_  & \new_[77372]_ ;
  assign \new_[77379]_  = A300 & A268;
  assign \new_[77382]_  = ~A302 & ~A301;
  assign \new_[77383]_  = \new_[77382]_  & \new_[77379]_ ;
  assign \new_[77384]_  = \new_[77383]_  & \new_[77376]_ ;
  assign \new_[77388]_  = ~A167 & A168;
  assign \new_[77389]_  = ~A170 & \new_[77388]_ ;
  assign \new_[77392]_  = ~A199 & A166;
  assign \new_[77395]_  = A201 & A200;
  assign \new_[77396]_  = \new_[77395]_  & \new_[77392]_ ;
  assign \new_[77397]_  = \new_[77396]_  & \new_[77389]_ ;
  assign \new_[77400]_  = A265 & A203;
  assign \new_[77403]_  = A267 & ~A266;
  assign \new_[77404]_  = \new_[77403]_  & \new_[77400]_ ;
  assign \new_[77407]_  = A300 & A269;
  assign \new_[77410]_  = ~A302 & ~A301;
  assign \new_[77411]_  = \new_[77410]_  & \new_[77407]_ ;
  assign \new_[77412]_  = \new_[77411]_  & \new_[77404]_ ;
  assign \new_[77416]_  = ~A167 & A168;
  assign \new_[77417]_  = ~A170 & \new_[77416]_ ;
  assign \new_[77420]_  = ~A199 & A166;
  assign \new_[77423]_  = A201 & A200;
  assign \new_[77424]_  = \new_[77423]_  & \new_[77420]_ ;
  assign \new_[77425]_  = \new_[77424]_  & \new_[77417]_ ;
  assign \new_[77428]_  = A265 & A203;
  assign \new_[77431]_  = ~A267 & ~A266;
  assign \new_[77432]_  = \new_[77431]_  & \new_[77428]_ ;
  assign \new_[77435]_  = ~A269 & ~A268;
  assign \new_[77438]_  = A301 & ~A300;
  assign \new_[77439]_  = \new_[77438]_  & \new_[77435]_ ;
  assign \new_[77440]_  = \new_[77439]_  & \new_[77432]_ ;
  assign \new_[77444]_  = ~A167 & A168;
  assign \new_[77445]_  = ~A170 & \new_[77444]_ ;
  assign \new_[77448]_  = ~A199 & A166;
  assign \new_[77451]_  = A201 & A200;
  assign \new_[77452]_  = \new_[77451]_  & \new_[77448]_ ;
  assign \new_[77453]_  = \new_[77452]_  & \new_[77445]_ ;
  assign \new_[77456]_  = A265 & A203;
  assign \new_[77459]_  = ~A267 & ~A266;
  assign \new_[77460]_  = \new_[77459]_  & \new_[77456]_ ;
  assign \new_[77463]_  = ~A269 & ~A268;
  assign \new_[77466]_  = A302 & ~A300;
  assign \new_[77467]_  = \new_[77466]_  & \new_[77463]_ ;
  assign \new_[77468]_  = \new_[77467]_  & \new_[77460]_ ;
  assign \new_[77472]_  = ~A167 & A168;
  assign \new_[77473]_  = ~A170 & \new_[77472]_ ;
  assign \new_[77476]_  = ~A199 & A166;
  assign \new_[77479]_  = A201 & A200;
  assign \new_[77480]_  = \new_[77479]_  & \new_[77476]_ ;
  assign \new_[77481]_  = \new_[77480]_  & \new_[77473]_ ;
  assign \new_[77484]_  = A265 & A203;
  assign \new_[77487]_  = ~A267 & ~A266;
  assign \new_[77488]_  = \new_[77487]_  & \new_[77484]_ ;
  assign \new_[77491]_  = ~A269 & ~A268;
  assign \new_[77494]_  = A299 & A298;
  assign \new_[77495]_  = \new_[77494]_  & \new_[77491]_ ;
  assign \new_[77496]_  = \new_[77495]_  & \new_[77488]_ ;
  assign \new_[77500]_  = ~A167 & A168;
  assign \new_[77501]_  = ~A170 & \new_[77500]_ ;
  assign \new_[77504]_  = ~A199 & A166;
  assign \new_[77507]_  = A201 & A200;
  assign \new_[77508]_  = \new_[77507]_  & \new_[77504]_ ;
  assign \new_[77509]_  = \new_[77508]_  & \new_[77501]_ ;
  assign \new_[77512]_  = A265 & A203;
  assign \new_[77515]_  = ~A267 & ~A266;
  assign \new_[77516]_  = \new_[77515]_  & \new_[77512]_ ;
  assign \new_[77519]_  = ~A269 & ~A268;
  assign \new_[77522]_  = ~A299 & ~A298;
  assign \new_[77523]_  = \new_[77522]_  & \new_[77519]_ ;
  assign \new_[77524]_  = \new_[77523]_  & \new_[77516]_ ;
  assign \new_[77528]_  = ~A167 & A168;
  assign \new_[77529]_  = ~A170 & \new_[77528]_ ;
  assign \new_[77532]_  = ~A199 & A166;
  assign \new_[77535]_  = ~A201 & A200;
  assign \new_[77536]_  = \new_[77535]_  & \new_[77532]_ ;
  assign \new_[77537]_  = \new_[77536]_  & \new_[77529]_ ;
  assign \new_[77540]_  = ~A203 & ~A202;
  assign \new_[77543]_  = A266 & ~A265;
  assign \new_[77544]_  = \new_[77543]_  & \new_[77540]_ ;
  assign \new_[77547]_  = A268 & A267;
  assign \new_[77550]_  = A301 & ~A300;
  assign \new_[77551]_  = \new_[77550]_  & \new_[77547]_ ;
  assign \new_[77552]_  = \new_[77551]_  & \new_[77544]_ ;
  assign \new_[77556]_  = ~A167 & A168;
  assign \new_[77557]_  = ~A170 & \new_[77556]_ ;
  assign \new_[77560]_  = ~A199 & A166;
  assign \new_[77563]_  = ~A201 & A200;
  assign \new_[77564]_  = \new_[77563]_  & \new_[77560]_ ;
  assign \new_[77565]_  = \new_[77564]_  & \new_[77557]_ ;
  assign \new_[77568]_  = ~A203 & ~A202;
  assign \new_[77571]_  = A266 & ~A265;
  assign \new_[77572]_  = \new_[77571]_  & \new_[77568]_ ;
  assign \new_[77575]_  = A268 & A267;
  assign \new_[77578]_  = A302 & ~A300;
  assign \new_[77579]_  = \new_[77578]_  & \new_[77575]_ ;
  assign \new_[77580]_  = \new_[77579]_  & \new_[77572]_ ;
  assign \new_[77584]_  = ~A167 & A168;
  assign \new_[77585]_  = ~A170 & \new_[77584]_ ;
  assign \new_[77588]_  = ~A199 & A166;
  assign \new_[77591]_  = ~A201 & A200;
  assign \new_[77592]_  = \new_[77591]_  & \new_[77588]_ ;
  assign \new_[77593]_  = \new_[77592]_  & \new_[77585]_ ;
  assign \new_[77596]_  = ~A203 & ~A202;
  assign \new_[77599]_  = A266 & ~A265;
  assign \new_[77600]_  = \new_[77599]_  & \new_[77596]_ ;
  assign \new_[77603]_  = A268 & A267;
  assign \new_[77606]_  = A299 & A298;
  assign \new_[77607]_  = \new_[77606]_  & \new_[77603]_ ;
  assign \new_[77608]_  = \new_[77607]_  & \new_[77600]_ ;
  assign \new_[77612]_  = ~A167 & A168;
  assign \new_[77613]_  = ~A170 & \new_[77612]_ ;
  assign \new_[77616]_  = ~A199 & A166;
  assign \new_[77619]_  = ~A201 & A200;
  assign \new_[77620]_  = \new_[77619]_  & \new_[77616]_ ;
  assign \new_[77621]_  = \new_[77620]_  & \new_[77613]_ ;
  assign \new_[77624]_  = ~A203 & ~A202;
  assign \new_[77627]_  = A266 & ~A265;
  assign \new_[77628]_  = \new_[77627]_  & \new_[77624]_ ;
  assign \new_[77631]_  = A268 & A267;
  assign \new_[77634]_  = ~A299 & ~A298;
  assign \new_[77635]_  = \new_[77634]_  & \new_[77631]_ ;
  assign \new_[77636]_  = \new_[77635]_  & \new_[77628]_ ;
  assign \new_[77640]_  = ~A167 & A168;
  assign \new_[77641]_  = ~A170 & \new_[77640]_ ;
  assign \new_[77644]_  = ~A199 & A166;
  assign \new_[77647]_  = ~A201 & A200;
  assign \new_[77648]_  = \new_[77647]_  & \new_[77644]_ ;
  assign \new_[77649]_  = \new_[77648]_  & \new_[77641]_ ;
  assign \new_[77652]_  = ~A203 & ~A202;
  assign \new_[77655]_  = A266 & ~A265;
  assign \new_[77656]_  = \new_[77655]_  & \new_[77652]_ ;
  assign \new_[77659]_  = A269 & A267;
  assign \new_[77662]_  = A301 & ~A300;
  assign \new_[77663]_  = \new_[77662]_  & \new_[77659]_ ;
  assign \new_[77664]_  = \new_[77663]_  & \new_[77656]_ ;
  assign \new_[77668]_  = ~A167 & A168;
  assign \new_[77669]_  = ~A170 & \new_[77668]_ ;
  assign \new_[77672]_  = ~A199 & A166;
  assign \new_[77675]_  = ~A201 & A200;
  assign \new_[77676]_  = \new_[77675]_  & \new_[77672]_ ;
  assign \new_[77677]_  = \new_[77676]_  & \new_[77669]_ ;
  assign \new_[77680]_  = ~A203 & ~A202;
  assign \new_[77683]_  = A266 & ~A265;
  assign \new_[77684]_  = \new_[77683]_  & \new_[77680]_ ;
  assign \new_[77687]_  = A269 & A267;
  assign \new_[77690]_  = A302 & ~A300;
  assign \new_[77691]_  = \new_[77690]_  & \new_[77687]_ ;
  assign \new_[77692]_  = \new_[77691]_  & \new_[77684]_ ;
  assign \new_[77696]_  = ~A167 & A168;
  assign \new_[77697]_  = ~A170 & \new_[77696]_ ;
  assign \new_[77700]_  = ~A199 & A166;
  assign \new_[77703]_  = ~A201 & A200;
  assign \new_[77704]_  = \new_[77703]_  & \new_[77700]_ ;
  assign \new_[77705]_  = \new_[77704]_  & \new_[77697]_ ;
  assign \new_[77708]_  = ~A203 & ~A202;
  assign \new_[77711]_  = A266 & ~A265;
  assign \new_[77712]_  = \new_[77711]_  & \new_[77708]_ ;
  assign \new_[77715]_  = A269 & A267;
  assign \new_[77718]_  = A299 & A298;
  assign \new_[77719]_  = \new_[77718]_  & \new_[77715]_ ;
  assign \new_[77720]_  = \new_[77719]_  & \new_[77712]_ ;
  assign \new_[77724]_  = ~A167 & A168;
  assign \new_[77725]_  = ~A170 & \new_[77724]_ ;
  assign \new_[77728]_  = ~A199 & A166;
  assign \new_[77731]_  = ~A201 & A200;
  assign \new_[77732]_  = \new_[77731]_  & \new_[77728]_ ;
  assign \new_[77733]_  = \new_[77732]_  & \new_[77725]_ ;
  assign \new_[77736]_  = ~A203 & ~A202;
  assign \new_[77739]_  = A266 & ~A265;
  assign \new_[77740]_  = \new_[77739]_  & \new_[77736]_ ;
  assign \new_[77743]_  = A269 & A267;
  assign \new_[77746]_  = ~A299 & ~A298;
  assign \new_[77747]_  = \new_[77746]_  & \new_[77743]_ ;
  assign \new_[77748]_  = \new_[77747]_  & \new_[77740]_ ;
  assign \new_[77752]_  = ~A167 & A168;
  assign \new_[77753]_  = ~A170 & \new_[77752]_ ;
  assign \new_[77756]_  = ~A199 & A166;
  assign \new_[77759]_  = ~A201 & A200;
  assign \new_[77760]_  = \new_[77759]_  & \new_[77756]_ ;
  assign \new_[77761]_  = \new_[77760]_  & \new_[77753]_ ;
  assign \new_[77764]_  = ~A203 & ~A202;
  assign \new_[77767]_  = ~A266 & A265;
  assign \new_[77768]_  = \new_[77767]_  & \new_[77764]_ ;
  assign \new_[77771]_  = A268 & A267;
  assign \new_[77774]_  = A301 & ~A300;
  assign \new_[77775]_  = \new_[77774]_  & \new_[77771]_ ;
  assign \new_[77776]_  = \new_[77775]_  & \new_[77768]_ ;
  assign \new_[77780]_  = ~A167 & A168;
  assign \new_[77781]_  = ~A170 & \new_[77780]_ ;
  assign \new_[77784]_  = ~A199 & A166;
  assign \new_[77787]_  = ~A201 & A200;
  assign \new_[77788]_  = \new_[77787]_  & \new_[77784]_ ;
  assign \new_[77789]_  = \new_[77788]_  & \new_[77781]_ ;
  assign \new_[77792]_  = ~A203 & ~A202;
  assign \new_[77795]_  = ~A266 & A265;
  assign \new_[77796]_  = \new_[77795]_  & \new_[77792]_ ;
  assign \new_[77799]_  = A268 & A267;
  assign \new_[77802]_  = A302 & ~A300;
  assign \new_[77803]_  = \new_[77802]_  & \new_[77799]_ ;
  assign \new_[77804]_  = \new_[77803]_  & \new_[77796]_ ;
  assign \new_[77808]_  = ~A167 & A168;
  assign \new_[77809]_  = ~A170 & \new_[77808]_ ;
  assign \new_[77812]_  = ~A199 & A166;
  assign \new_[77815]_  = ~A201 & A200;
  assign \new_[77816]_  = \new_[77815]_  & \new_[77812]_ ;
  assign \new_[77817]_  = \new_[77816]_  & \new_[77809]_ ;
  assign \new_[77820]_  = ~A203 & ~A202;
  assign \new_[77823]_  = ~A266 & A265;
  assign \new_[77824]_  = \new_[77823]_  & \new_[77820]_ ;
  assign \new_[77827]_  = A268 & A267;
  assign \new_[77830]_  = A299 & A298;
  assign \new_[77831]_  = \new_[77830]_  & \new_[77827]_ ;
  assign \new_[77832]_  = \new_[77831]_  & \new_[77824]_ ;
  assign \new_[77836]_  = ~A167 & A168;
  assign \new_[77837]_  = ~A170 & \new_[77836]_ ;
  assign \new_[77840]_  = ~A199 & A166;
  assign \new_[77843]_  = ~A201 & A200;
  assign \new_[77844]_  = \new_[77843]_  & \new_[77840]_ ;
  assign \new_[77845]_  = \new_[77844]_  & \new_[77837]_ ;
  assign \new_[77848]_  = ~A203 & ~A202;
  assign \new_[77851]_  = ~A266 & A265;
  assign \new_[77852]_  = \new_[77851]_  & \new_[77848]_ ;
  assign \new_[77855]_  = A268 & A267;
  assign \new_[77858]_  = ~A299 & ~A298;
  assign \new_[77859]_  = \new_[77858]_  & \new_[77855]_ ;
  assign \new_[77860]_  = \new_[77859]_  & \new_[77852]_ ;
  assign \new_[77864]_  = ~A167 & A168;
  assign \new_[77865]_  = ~A170 & \new_[77864]_ ;
  assign \new_[77868]_  = ~A199 & A166;
  assign \new_[77871]_  = ~A201 & A200;
  assign \new_[77872]_  = \new_[77871]_  & \new_[77868]_ ;
  assign \new_[77873]_  = \new_[77872]_  & \new_[77865]_ ;
  assign \new_[77876]_  = ~A203 & ~A202;
  assign \new_[77879]_  = ~A266 & A265;
  assign \new_[77880]_  = \new_[77879]_  & \new_[77876]_ ;
  assign \new_[77883]_  = A269 & A267;
  assign \new_[77886]_  = A301 & ~A300;
  assign \new_[77887]_  = \new_[77886]_  & \new_[77883]_ ;
  assign \new_[77888]_  = \new_[77887]_  & \new_[77880]_ ;
  assign \new_[77892]_  = ~A167 & A168;
  assign \new_[77893]_  = ~A170 & \new_[77892]_ ;
  assign \new_[77896]_  = ~A199 & A166;
  assign \new_[77899]_  = ~A201 & A200;
  assign \new_[77900]_  = \new_[77899]_  & \new_[77896]_ ;
  assign \new_[77901]_  = \new_[77900]_  & \new_[77893]_ ;
  assign \new_[77904]_  = ~A203 & ~A202;
  assign \new_[77907]_  = ~A266 & A265;
  assign \new_[77908]_  = \new_[77907]_  & \new_[77904]_ ;
  assign \new_[77911]_  = A269 & A267;
  assign \new_[77914]_  = A302 & ~A300;
  assign \new_[77915]_  = \new_[77914]_  & \new_[77911]_ ;
  assign \new_[77916]_  = \new_[77915]_  & \new_[77908]_ ;
  assign \new_[77920]_  = ~A167 & A168;
  assign \new_[77921]_  = ~A170 & \new_[77920]_ ;
  assign \new_[77924]_  = ~A199 & A166;
  assign \new_[77927]_  = ~A201 & A200;
  assign \new_[77928]_  = \new_[77927]_  & \new_[77924]_ ;
  assign \new_[77929]_  = \new_[77928]_  & \new_[77921]_ ;
  assign \new_[77932]_  = ~A203 & ~A202;
  assign \new_[77935]_  = ~A266 & A265;
  assign \new_[77936]_  = \new_[77935]_  & \new_[77932]_ ;
  assign \new_[77939]_  = A269 & A267;
  assign \new_[77942]_  = A299 & A298;
  assign \new_[77943]_  = \new_[77942]_  & \new_[77939]_ ;
  assign \new_[77944]_  = \new_[77943]_  & \new_[77936]_ ;
  assign \new_[77948]_  = ~A167 & A168;
  assign \new_[77949]_  = ~A170 & \new_[77948]_ ;
  assign \new_[77952]_  = ~A199 & A166;
  assign \new_[77955]_  = ~A201 & A200;
  assign \new_[77956]_  = \new_[77955]_  & \new_[77952]_ ;
  assign \new_[77957]_  = \new_[77956]_  & \new_[77949]_ ;
  assign \new_[77960]_  = ~A203 & ~A202;
  assign \new_[77963]_  = ~A266 & A265;
  assign \new_[77964]_  = \new_[77963]_  & \new_[77960]_ ;
  assign \new_[77967]_  = A269 & A267;
  assign \new_[77970]_  = ~A299 & ~A298;
  assign \new_[77971]_  = \new_[77970]_  & \new_[77967]_ ;
  assign \new_[77972]_  = \new_[77971]_  & \new_[77964]_ ;
  assign \new_[77976]_  = ~A167 & A168;
  assign \new_[77977]_  = ~A170 & \new_[77976]_ ;
  assign \new_[77980]_  = A199 & A166;
  assign \new_[77983]_  = A201 & ~A200;
  assign \new_[77984]_  = \new_[77983]_  & \new_[77980]_ ;
  assign \new_[77985]_  = \new_[77984]_  & \new_[77977]_ ;
  assign \new_[77988]_  = ~A265 & A202;
  assign \new_[77991]_  = A267 & A266;
  assign \new_[77992]_  = \new_[77991]_  & \new_[77988]_ ;
  assign \new_[77995]_  = A300 & A268;
  assign \new_[77998]_  = ~A302 & ~A301;
  assign \new_[77999]_  = \new_[77998]_  & \new_[77995]_ ;
  assign \new_[78000]_  = \new_[77999]_  & \new_[77992]_ ;
  assign \new_[78004]_  = ~A167 & A168;
  assign \new_[78005]_  = ~A170 & \new_[78004]_ ;
  assign \new_[78008]_  = A199 & A166;
  assign \new_[78011]_  = A201 & ~A200;
  assign \new_[78012]_  = \new_[78011]_  & \new_[78008]_ ;
  assign \new_[78013]_  = \new_[78012]_  & \new_[78005]_ ;
  assign \new_[78016]_  = ~A265 & A202;
  assign \new_[78019]_  = A267 & A266;
  assign \new_[78020]_  = \new_[78019]_  & \new_[78016]_ ;
  assign \new_[78023]_  = A300 & A269;
  assign \new_[78026]_  = ~A302 & ~A301;
  assign \new_[78027]_  = \new_[78026]_  & \new_[78023]_ ;
  assign \new_[78028]_  = \new_[78027]_  & \new_[78020]_ ;
  assign \new_[78032]_  = ~A167 & A168;
  assign \new_[78033]_  = ~A170 & \new_[78032]_ ;
  assign \new_[78036]_  = A199 & A166;
  assign \new_[78039]_  = A201 & ~A200;
  assign \new_[78040]_  = \new_[78039]_  & \new_[78036]_ ;
  assign \new_[78041]_  = \new_[78040]_  & \new_[78033]_ ;
  assign \new_[78044]_  = ~A265 & A202;
  assign \new_[78047]_  = ~A267 & A266;
  assign \new_[78048]_  = \new_[78047]_  & \new_[78044]_ ;
  assign \new_[78051]_  = ~A269 & ~A268;
  assign \new_[78054]_  = A301 & ~A300;
  assign \new_[78055]_  = \new_[78054]_  & \new_[78051]_ ;
  assign \new_[78056]_  = \new_[78055]_  & \new_[78048]_ ;
  assign \new_[78060]_  = ~A167 & A168;
  assign \new_[78061]_  = ~A170 & \new_[78060]_ ;
  assign \new_[78064]_  = A199 & A166;
  assign \new_[78067]_  = A201 & ~A200;
  assign \new_[78068]_  = \new_[78067]_  & \new_[78064]_ ;
  assign \new_[78069]_  = \new_[78068]_  & \new_[78061]_ ;
  assign \new_[78072]_  = ~A265 & A202;
  assign \new_[78075]_  = ~A267 & A266;
  assign \new_[78076]_  = \new_[78075]_  & \new_[78072]_ ;
  assign \new_[78079]_  = ~A269 & ~A268;
  assign \new_[78082]_  = A302 & ~A300;
  assign \new_[78083]_  = \new_[78082]_  & \new_[78079]_ ;
  assign \new_[78084]_  = \new_[78083]_  & \new_[78076]_ ;
  assign \new_[78088]_  = ~A167 & A168;
  assign \new_[78089]_  = ~A170 & \new_[78088]_ ;
  assign \new_[78092]_  = A199 & A166;
  assign \new_[78095]_  = A201 & ~A200;
  assign \new_[78096]_  = \new_[78095]_  & \new_[78092]_ ;
  assign \new_[78097]_  = \new_[78096]_  & \new_[78089]_ ;
  assign \new_[78100]_  = ~A265 & A202;
  assign \new_[78103]_  = ~A267 & A266;
  assign \new_[78104]_  = \new_[78103]_  & \new_[78100]_ ;
  assign \new_[78107]_  = ~A269 & ~A268;
  assign \new_[78110]_  = A299 & A298;
  assign \new_[78111]_  = \new_[78110]_  & \new_[78107]_ ;
  assign \new_[78112]_  = \new_[78111]_  & \new_[78104]_ ;
  assign \new_[78116]_  = ~A167 & A168;
  assign \new_[78117]_  = ~A170 & \new_[78116]_ ;
  assign \new_[78120]_  = A199 & A166;
  assign \new_[78123]_  = A201 & ~A200;
  assign \new_[78124]_  = \new_[78123]_  & \new_[78120]_ ;
  assign \new_[78125]_  = \new_[78124]_  & \new_[78117]_ ;
  assign \new_[78128]_  = ~A265 & A202;
  assign \new_[78131]_  = ~A267 & A266;
  assign \new_[78132]_  = \new_[78131]_  & \new_[78128]_ ;
  assign \new_[78135]_  = ~A269 & ~A268;
  assign \new_[78138]_  = ~A299 & ~A298;
  assign \new_[78139]_  = \new_[78138]_  & \new_[78135]_ ;
  assign \new_[78140]_  = \new_[78139]_  & \new_[78132]_ ;
  assign \new_[78144]_  = ~A167 & A168;
  assign \new_[78145]_  = ~A170 & \new_[78144]_ ;
  assign \new_[78148]_  = A199 & A166;
  assign \new_[78151]_  = A201 & ~A200;
  assign \new_[78152]_  = \new_[78151]_  & \new_[78148]_ ;
  assign \new_[78153]_  = \new_[78152]_  & \new_[78145]_ ;
  assign \new_[78156]_  = A265 & A202;
  assign \new_[78159]_  = A267 & ~A266;
  assign \new_[78160]_  = \new_[78159]_  & \new_[78156]_ ;
  assign \new_[78163]_  = A300 & A268;
  assign \new_[78166]_  = ~A302 & ~A301;
  assign \new_[78167]_  = \new_[78166]_  & \new_[78163]_ ;
  assign \new_[78168]_  = \new_[78167]_  & \new_[78160]_ ;
  assign \new_[78172]_  = ~A167 & A168;
  assign \new_[78173]_  = ~A170 & \new_[78172]_ ;
  assign \new_[78176]_  = A199 & A166;
  assign \new_[78179]_  = A201 & ~A200;
  assign \new_[78180]_  = \new_[78179]_  & \new_[78176]_ ;
  assign \new_[78181]_  = \new_[78180]_  & \new_[78173]_ ;
  assign \new_[78184]_  = A265 & A202;
  assign \new_[78187]_  = A267 & ~A266;
  assign \new_[78188]_  = \new_[78187]_  & \new_[78184]_ ;
  assign \new_[78191]_  = A300 & A269;
  assign \new_[78194]_  = ~A302 & ~A301;
  assign \new_[78195]_  = \new_[78194]_  & \new_[78191]_ ;
  assign \new_[78196]_  = \new_[78195]_  & \new_[78188]_ ;
  assign \new_[78200]_  = ~A167 & A168;
  assign \new_[78201]_  = ~A170 & \new_[78200]_ ;
  assign \new_[78204]_  = A199 & A166;
  assign \new_[78207]_  = A201 & ~A200;
  assign \new_[78208]_  = \new_[78207]_  & \new_[78204]_ ;
  assign \new_[78209]_  = \new_[78208]_  & \new_[78201]_ ;
  assign \new_[78212]_  = A265 & A202;
  assign \new_[78215]_  = ~A267 & ~A266;
  assign \new_[78216]_  = \new_[78215]_  & \new_[78212]_ ;
  assign \new_[78219]_  = ~A269 & ~A268;
  assign \new_[78222]_  = A301 & ~A300;
  assign \new_[78223]_  = \new_[78222]_  & \new_[78219]_ ;
  assign \new_[78224]_  = \new_[78223]_  & \new_[78216]_ ;
  assign \new_[78228]_  = ~A167 & A168;
  assign \new_[78229]_  = ~A170 & \new_[78228]_ ;
  assign \new_[78232]_  = A199 & A166;
  assign \new_[78235]_  = A201 & ~A200;
  assign \new_[78236]_  = \new_[78235]_  & \new_[78232]_ ;
  assign \new_[78237]_  = \new_[78236]_  & \new_[78229]_ ;
  assign \new_[78240]_  = A265 & A202;
  assign \new_[78243]_  = ~A267 & ~A266;
  assign \new_[78244]_  = \new_[78243]_  & \new_[78240]_ ;
  assign \new_[78247]_  = ~A269 & ~A268;
  assign \new_[78250]_  = A302 & ~A300;
  assign \new_[78251]_  = \new_[78250]_  & \new_[78247]_ ;
  assign \new_[78252]_  = \new_[78251]_  & \new_[78244]_ ;
  assign \new_[78256]_  = ~A167 & A168;
  assign \new_[78257]_  = ~A170 & \new_[78256]_ ;
  assign \new_[78260]_  = A199 & A166;
  assign \new_[78263]_  = A201 & ~A200;
  assign \new_[78264]_  = \new_[78263]_  & \new_[78260]_ ;
  assign \new_[78265]_  = \new_[78264]_  & \new_[78257]_ ;
  assign \new_[78268]_  = A265 & A202;
  assign \new_[78271]_  = ~A267 & ~A266;
  assign \new_[78272]_  = \new_[78271]_  & \new_[78268]_ ;
  assign \new_[78275]_  = ~A269 & ~A268;
  assign \new_[78278]_  = A299 & A298;
  assign \new_[78279]_  = \new_[78278]_  & \new_[78275]_ ;
  assign \new_[78280]_  = \new_[78279]_  & \new_[78272]_ ;
  assign \new_[78284]_  = ~A167 & A168;
  assign \new_[78285]_  = ~A170 & \new_[78284]_ ;
  assign \new_[78288]_  = A199 & A166;
  assign \new_[78291]_  = A201 & ~A200;
  assign \new_[78292]_  = \new_[78291]_  & \new_[78288]_ ;
  assign \new_[78293]_  = \new_[78292]_  & \new_[78285]_ ;
  assign \new_[78296]_  = A265 & A202;
  assign \new_[78299]_  = ~A267 & ~A266;
  assign \new_[78300]_  = \new_[78299]_  & \new_[78296]_ ;
  assign \new_[78303]_  = ~A269 & ~A268;
  assign \new_[78306]_  = ~A299 & ~A298;
  assign \new_[78307]_  = \new_[78306]_  & \new_[78303]_ ;
  assign \new_[78308]_  = \new_[78307]_  & \new_[78300]_ ;
  assign \new_[78312]_  = ~A167 & A168;
  assign \new_[78313]_  = ~A170 & \new_[78312]_ ;
  assign \new_[78316]_  = A199 & A166;
  assign \new_[78319]_  = A201 & ~A200;
  assign \new_[78320]_  = \new_[78319]_  & \new_[78316]_ ;
  assign \new_[78321]_  = \new_[78320]_  & \new_[78313]_ ;
  assign \new_[78324]_  = ~A265 & A203;
  assign \new_[78327]_  = A267 & A266;
  assign \new_[78328]_  = \new_[78327]_  & \new_[78324]_ ;
  assign \new_[78331]_  = A300 & A268;
  assign \new_[78334]_  = ~A302 & ~A301;
  assign \new_[78335]_  = \new_[78334]_  & \new_[78331]_ ;
  assign \new_[78336]_  = \new_[78335]_  & \new_[78328]_ ;
  assign \new_[78340]_  = ~A167 & A168;
  assign \new_[78341]_  = ~A170 & \new_[78340]_ ;
  assign \new_[78344]_  = A199 & A166;
  assign \new_[78347]_  = A201 & ~A200;
  assign \new_[78348]_  = \new_[78347]_  & \new_[78344]_ ;
  assign \new_[78349]_  = \new_[78348]_  & \new_[78341]_ ;
  assign \new_[78352]_  = ~A265 & A203;
  assign \new_[78355]_  = A267 & A266;
  assign \new_[78356]_  = \new_[78355]_  & \new_[78352]_ ;
  assign \new_[78359]_  = A300 & A269;
  assign \new_[78362]_  = ~A302 & ~A301;
  assign \new_[78363]_  = \new_[78362]_  & \new_[78359]_ ;
  assign \new_[78364]_  = \new_[78363]_  & \new_[78356]_ ;
  assign \new_[78368]_  = ~A167 & A168;
  assign \new_[78369]_  = ~A170 & \new_[78368]_ ;
  assign \new_[78372]_  = A199 & A166;
  assign \new_[78375]_  = A201 & ~A200;
  assign \new_[78376]_  = \new_[78375]_  & \new_[78372]_ ;
  assign \new_[78377]_  = \new_[78376]_  & \new_[78369]_ ;
  assign \new_[78380]_  = ~A265 & A203;
  assign \new_[78383]_  = ~A267 & A266;
  assign \new_[78384]_  = \new_[78383]_  & \new_[78380]_ ;
  assign \new_[78387]_  = ~A269 & ~A268;
  assign \new_[78390]_  = A301 & ~A300;
  assign \new_[78391]_  = \new_[78390]_  & \new_[78387]_ ;
  assign \new_[78392]_  = \new_[78391]_  & \new_[78384]_ ;
  assign \new_[78396]_  = ~A167 & A168;
  assign \new_[78397]_  = ~A170 & \new_[78396]_ ;
  assign \new_[78400]_  = A199 & A166;
  assign \new_[78403]_  = A201 & ~A200;
  assign \new_[78404]_  = \new_[78403]_  & \new_[78400]_ ;
  assign \new_[78405]_  = \new_[78404]_  & \new_[78397]_ ;
  assign \new_[78408]_  = ~A265 & A203;
  assign \new_[78411]_  = ~A267 & A266;
  assign \new_[78412]_  = \new_[78411]_  & \new_[78408]_ ;
  assign \new_[78415]_  = ~A269 & ~A268;
  assign \new_[78418]_  = A302 & ~A300;
  assign \new_[78419]_  = \new_[78418]_  & \new_[78415]_ ;
  assign \new_[78420]_  = \new_[78419]_  & \new_[78412]_ ;
  assign \new_[78424]_  = ~A167 & A168;
  assign \new_[78425]_  = ~A170 & \new_[78424]_ ;
  assign \new_[78428]_  = A199 & A166;
  assign \new_[78431]_  = A201 & ~A200;
  assign \new_[78432]_  = \new_[78431]_  & \new_[78428]_ ;
  assign \new_[78433]_  = \new_[78432]_  & \new_[78425]_ ;
  assign \new_[78436]_  = ~A265 & A203;
  assign \new_[78439]_  = ~A267 & A266;
  assign \new_[78440]_  = \new_[78439]_  & \new_[78436]_ ;
  assign \new_[78443]_  = ~A269 & ~A268;
  assign \new_[78446]_  = A299 & A298;
  assign \new_[78447]_  = \new_[78446]_  & \new_[78443]_ ;
  assign \new_[78448]_  = \new_[78447]_  & \new_[78440]_ ;
  assign \new_[78452]_  = ~A167 & A168;
  assign \new_[78453]_  = ~A170 & \new_[78452]_ ;
  assign \new_[78456]_  = A199 & A166;
  assign \new_[78459]_  = A201 & ~A200;
  assign \new_[78460]_  = \new_[78459]_  & \new_[78456]_ ;
  assign \new_[78461]_  = \new_[78460]_  & \new_[78453]_ ;
  assign \new_[78464]_  = ~A265 & A203;
  assign \new_[78467]_  = ~A267 & A266;
  assign \new_[78468]_  = \new_[78467]_  & \new_[78464]_ ;
  assign \new_[78471]_  = ~A269 & ~A268;
  assign \new_[78474]_  = ~A299 & ~A298;
  assign \new_[78475]_  = \new_[78474]_  & \new_[78471]_ ;
  assign \new_[78476]_  = \new_[78475]_  & \new_[78468]_ ;
  assign \new_[78480]_  = ~A167 & A168;
  assign \new_[78481]_  = ~A170 & \new_[78480]_ ;
  assign \new_[78484]_  = A199 & A166;
  assign \new_[78487]_  = A201 & ~A200;
  assign \new_[78488]_  = \new_[78487]_  & \new_[78484]_ ;
  assign \new_[78489]_  = \new_[78488]_  & \new_[78481]_ ;
  assign \new_[78492]_  = A265 & A203;
  assign \new_[78495]_  = A267 & ~A266;
  assign \new_[78496]_  = \new_[78495]_  & \new_[78492]_ ;
  assign \new_[78499]_  = A300 & A268;
  assign \new_[78502]_  = ~A302 & ~A301;
  assign \new_[78503]_  = \new_[78502]_  & \new_[78499]_ ;
  assign \new_[78504]_  = \new_[78503]_  & \new_[78496]_ ;
  assign \new_[78508]_  = ~A167 & A168;
  assign \new_[78509]_  = ~A170 & \new_[78508]_ ;
  assign \new_[78512]_  = A199 & A166;
  assign \new_[78515]_  = A201 & ~A200;
  assign \new_[78516]_  = \new_[78515]_  & \new_[78512]_ ;
  assign \new_[78517]_  = \new_[78516]_  & \new_[78509]_ ;
  assign \new_[78520]_  = A265 & A203;
  assign \new_[78523]_  = A267 & ~A266;
  assign \new_[78524]_  = \new_[78523]_  & \new_[78520]_ ;
  assign \new_[78527]_  = A300 & A269;
  assign \new_[78530]_  = ~A302 & ~A301;
  assign \new_[78531]_  = \new_[78530]_  & \new_[78527]_ ;
  assign \new_[78532]_  = \new_[78531]_  & \new_[78524]_ ;
  assign \new_[78536]_  = ~A167 & A168;
  assign \new_[78537]_  = ~A170 & \new_[78536]_ ;
  assign \new_[78540]_  = A199 & A166;
  assign \new_[78543]_  = A201 & ~A200;
  assign \new_[78544]_  = \new_[78543]_  & \new_[78540]_ ;
  assign \new_[78545]_  = \new_[78544]_  & \new_[78537]_ ;
  assign \new_[78548]_  = A265 & A203;
  assign \new_[78551]_  = ~A267 & ~A266;
  assign \new_[78552]_  = \new_[78551]_  & \new_[78548]_ ;
  assign \new_[78555]_  = ~A269 & ~A268;
  assign \new_[78558]_  = A301 & ~A300;
  assign \new_[78559]_  = \new_[78558]_  & \new_[78555]_ ;
  assign \new_[78560]_  = \new_[78559]_  & \new_[78552]_ ;
  assign \new_[78564]_  = ~A167 & A168;
  assign \new_[78565]_  = ~A170 & \new_[78564]_ ;
  assign \new_[78568]_  = A199 & A166;
  assign \new_[78571]_  = A201 & ~A200;
  assign \new_[78572]_  = \new_[78571]_  & \new_[78568]_ ;
  assign \new_[78573]_  = \new_[78572]_  & \new_[78565]_ ;
  assign \new_[78576]_  = A265 & A203;
  assign \new_[78579]_  = ~A267 & ~A266;
  assign \new_[78580]_  = \new_[78579]_  & \new_[78576]_ ;
  assign \new_[78583]_  = ~A269 & ~A268;
  assign \new_[78586]_  = A302 & ~A300;
  assign \new_[78587]_  = \new_[78586]_  & \new_[78583]_ ;
  assign \new_[78588]_  = \new_[78587]_  & \new_[78580]_ ;
  assign \new_[78592]_  = ~A167 & A168;
  assign \new_[78593]_  = ~A170 & \new_[78592]_ ;
  assign \new_[78596]_  = A199 & A166;
  assign \new_[78599]_  = A201 & ~A200;
  assign \new_[78600]_  = \new_[78599]_  & \new_[78596]_ ;
  assign \new_[78601]_  = \new_[78600]_  & \new_[78593]_ ;
  assign \new_[78604]_  = A265 & A203;
  assign \new_[78607]_  = ~A267 & ~A266;
  assign \new_[78608]_  = \new_[78607]_  & \new_[78604]_ ;
  assign \new_[78611]_  = ~A269 & ~A268;
  assign \new_[78614]_  = A299 & A298;
  assign \new_[78615]_  = \new_[78614]_  & \new_[78611]_ ;
  assign \new_[78616]_  = \new_[78615]_  & \new_[78608]_ ;
  assign \new_[78620]_  = ~A167 & A168;
  assign \new_[78621]_  = ~A170 & \new_[78620]_ ;
  assign \new_[78624]_  = A199 & A166;
  assign \new_[78627]_  = A201 & ~A200;
  assign \new_[78628]_  = \new_[78627]_  & \new_[78624]_ ;
  assign \new_[78629]_  = \new_[78628]_  & \new_[78621]_ ;
  assign \new_[78632]_  = A265 & A203;
  assign \new_[78635]_  = ~A267 & ~A266;
  assign \new_[78636]_  = \new_[78635]_  & \new_[78632]_ ;
  assign \new_[78639]_  = ~A269 & ~A268;
  assign \new_[78642]_  = ~A299 & ~A298;
  assign \new_[78643]_  = \new_[78642]_  & \new_[78639]_ ;
  assign \new_[78644]_  = \new_[78643]_  & \new_[78636]_ ;
  assign \new_[78648]_  = ~A167 & A168;
  assign \new_[78649]_  = ~A170 & \new_[78648]_ ;
  assign \new_[78652]_  = A199 & A166;
  assign \new_[78655]_  = ~A201 & ~A200;
  assign \new_[78656]_  = \new_[78655]_  & \new_[78652]_ ;
  assign \new_[78657]_  = \new_[78656]_  & \new_[78649]_ ;
  assign \new_[78660]_  = ~A203 & ~A202;
  assign \new_[78663]_  = A266 & ~A265;
  assign \new_[78664]_  = \new_[78663]_  & \new_[78660]_ ;
  assign \new_[78667]_  = A268 & A267;
  assign \new_[78670]_  = A301 & ~A300;
  assign \new_[78671]_  = \new_[78670]_  & \new_[78667]_ ;
  assign \new_[78672]_  = \new_[78671]_  & \new_[78664]_ ;
  assign \new_[78676]_  = ~A167 & A168;
  assign \new_[78677]_  = ~A170 & \new_[78676]_ ;
  assign \new_[78680]_  = A199 & A166;
  assign \new_[78683]_  = ~A201 & ~A200;
  assign \new_[78684]_  = \new_[78683]_  & \new_[78680]_ ;
  assign \new_[78685]_  = \new_[78684]_  & \new_[78677]_ ;
  assign \new_[78688]_  = ~A203 & ~A202;
  assign \new_[78691]_  = A266 & ~A265;
  assign \new_[78692]_  = \new_[78691]_  & \new_[78688]_ ;
  assign \new_[78695]_  = A268 & A267;
  assign \new_[78698]_  = A302 & ~A300;
  assign \new_[78699]_  = \new_[78698]_  & \new_[78695]_ ;
  assign \new_[78700]_  = \new_[78699]_  & \new_[78692]_ ;
  assign \new_[78704]_  = ~A167 & A168;
  assign \new_[78705]_  = ~A170 & \new_[78704]_ ;
  assign \new_[78708]_  = A199 & A166;
  assign \new_[78711]_  = ~A201 & ~A200;
  assign \new_[78712]_  = \new_[78711]_  & \new_[78708]_ ;
  assign \new_[78713]_  = \new_[78712]_  & \new_[78705]_ ;
  assign \new_[78716]_  = ~A203 & ~A202;
  assign \new_[78719]_  = A266 & ~A265;
  assign \new_[78720]_  = \new_[78719]_  & \new_[78716]_ ;
  assign \new_[78723]_  = A268 & A267;
  assign \new_[78726]_  = A299 & A298;
  assign \new_[78727]_  = \new_[78726]_  & \new_[78723]_ ;
  assign \new_[78728]_  = \new_[78727]_  & \new_[78720]_ ;
  assign \new_[78732]_  = ~A167 & A168;
  assign \new_[78733]_  = ~A170 & \new_[78732]_ ;
  assign \new_[78736]_  = A199 & A166;
  assign \new_[78739]_  = ~A201 & ~A200;
  assign \new_[78740]_  = \new_[78739]_  & \new_[78736]_ ;
  assign \new_[78741]_  = \new_[78740]_  & \new_[78733]_ ;
  assign \new_[78744]_  = ~A203 & ~A202;
  assign \new_[78747]_  = A266 & ~A265;
  assign \new_[78748]_  = \new_[78747]_  & \new_[78744]_ ;
  assign \new_[78751]_  = A268 & A267;
  assign \new_[78754]_  = ~A299 & ~A298;
  assign \new_[78755]_  = \new_[78754]_  & \new_[78751]_ ;
  assign \new_[78756]_  = \new_[78755]_  & \new_[78748]_ ;
  assign \new_[78760]_  = ~A167 & A168;
  assign \new_[78761]_  = ~A170 & \new_[78760]_ ;
  assign \new_[78764]_  = A199 & A166;
  assign \new_[78767]_  = ~A201 & ~A200;
  assign \new_[78768]_  = \new_[78767]_  & \new_[78764]_ ;
  assign \new_[78769]_  = \new_[78768]_  & \new_[78761]_ ;
  assign \new_[78772]_  = ~A203 & ~A202;
  assign \new_[78775]_  = A266 & ~A265;
  assign \new_[78776]_  = \new_[78775]_  & \new_[78772]_ ;
  assign \new_[78779]_  = A269 & A267;
  assign \new_[78782]_  = A301 & ~A300;
  assign \new_[78783]_  = \new_[78782]_  & \new_[78779]_ ;
  assign \new_[78784]_  = \new_[78783]_  & \new_[78776]_ ;
  assign \new_[78788]_  = ~A167 & A168;
  assign \new_[78789]_  = ~A170 & \new_[78788]_ ;
  assign \new_[78792]_  = A199 & A166;
  assign \new_[78795]_  = ~A201 & ~A200;
  assign \new_[78796]_  = \new_[78795]_  & \new_[78792]_ ;
  assign \new_[78797]_  = \new_[78796]_  & \new_[78789]_ ;
  assign \new_[78800]_  = ~A203 & ~A202;
  assign \new_[78803]_  = A266 & ~A265;
  assign \new_[78804]_  = \new_[78803]_  & \new_[78800]_ ;
  assign \new_[78807]_  = A269 & A267;
  assign \new_[78810]_  = A302 & ~A300;
  assign \new_[78811]_  = \new_[78810]_  & \new_[78807]_ ;
  assign \new_[78812]_  = \new_[78811]_  & \new_[78804]_ ;
  assign \new_[78816]_  = ~A167 & A168;
  assign \new_[78817]_  = ~A170 & \new_[78816]_ ;
  assign \new_[78820]_  = A199 & A166;
  assign \new_[78823]_  = ~A201 & ~A200;
  assign \new_[78824]_  = \new_[78823]_  & \new_[78820]_ ;
  assign \new_[78825]_  = \new_[78824]_  & \new_[78817]_ ;
  assign \new_[78828]_  = ~A203 & ~A202;
  assign \new_[78831]_  = A266 & ~A265;
  assign \new_[78832]_  = \new_[78831]_  & \new_[78828]_ ;
  assign \new_[78835]_  = A269 & A267;
  assign \new_[78838]_  = A299 & A298;
  assign \new_[78839]_  = \new_[78838]_  & \new_[78835]_ ;
  assign \new_[78840]_  = \new_[78839]_  & \new_[78832]_ ;
  assign \new_[78844]_  = ~A167 & A168;
  assign \new_[78845]_  = ~A170 & \new_[78844]_ ;
  assign \new_[78848]_  = A199 & A166;
  assign \new_[78851]_  = ~A201 & ~A200;
  assign \new_[78852]_  = \new_[78851]_  & \new_[78848]_ ;
  assign \new_[78853]_  = \new_[78852]_  & \new_[78845]_ ;
  assign \new_[78856]_  = ~A203 & ~A202;
  assign \new_[78859]_  = A266 & ~A265;
  assign \new_[78860]_  = \new_[78859]_  & \new_[78856]_ ;
  assign \new_[78863]_  = A269 & A267;
  assign \new_[78866]_  = ~A299 & ~A298;
  assign \new_[78867]_  = \new_[78866]_  & \new_[78863]_ ;
  assign \new_[78868]_  = \new_[78867]_  & \new_[78860]_ ;
  assign \new_[78872]_  = ~A167 & A168;
  assign \new_[78873]_  = ~A170 & \new_[78872]_ ;
  assign \new_[78876]_  = A199 & A166;
  assign \new_[78879]_  = ~A201 & ~A200;
  assign \new_[78880]_  = \new_[78879]_  & \new_[78876]_ ;
  assign \new_[78881]_  = \new_[78880]_  & \new_[78873]_ ;
  assign \new_[78884]_  = ~A203 & ~A202;
  assign \new_[78887]_  = ~A266 & A265;
  assign \new_[78888]_  = \new_[78887]_  & \new_[78884]_ ;
  assign \new_[78891]_  = A268 & A267;
  assign \new_[78894]_  = A301 & ~A300;
  assign \new_[78895]_  = \new_[78894]_  & \new_[78891]_ ;
  assign \new_[78896]_  = \new_[78895]_  & \new_[78888]_ ;
  assign \new_[78900]_  = ~A167 & A168;
  assign \new_[78901]_  = ~A170 & \new_[78900]_ ;
  assign \new_[78904]_  = A199 & A166;
  assign \new_[78907]_  = ~A201 & ~A200;
  assign \new_[78908]_  = \new_[78907]_  & \new_[78904]_ ;
  assign \new_[78909]_  = \new_[78908]_  & \new_[78901]_ ;
  assign \new_[78912]_  = ~A203 & ~A202;
  assign \new_[78915]_  = ~A266 & A265;
  assign \new_[78916]_  = \new_[78915]_  & \new_[78912]_ ;
  assign \new_[78919]_  = A268 & A267;
  assign \new_[78922]_  = A302 & ~A300;
  assign \new_[78923]_  = \new_[78922]_  & \new_[78919]_ ;
  assign \new_[78924]_  = \new_[78923]_  & \new_[78916]_ ;
  assign \new_[78928]_  = ~A167 & A168;
  assign \new_[78929]_  = ~A170 & \new_[78928]_ ;
  assign \new_[78932]_  = A199 & A166;
  assign \new_[78935]_  = ~A201 & ~A200;
  assign \new_[78936]_  = \new_[78935]_  & \new_[78932]_ ;
  assign \new_[78937]_  = \new_[78936]_  & \new_[78929]_ ;
  assign \new_[78940]_  = ~A203 & ~A202;
  assign \new_[78943]_  = ~A266 & A265;
  assign \new_[78944]_  = \new_[78943]_  & \new_[78940]_ ;
  assign \new_[78947]_  = A268 & A267;
  assign \new_[78950]_  = A299 & A298;
  assign \new_[78951]_  = \new_[78950]_  & \new_[78947]_ ;
  assign \new_[78952]_  = \new_[78951]_  & \new_[78944]_ ;
  assign \new_[78956]_  = ~A167 & A168;
  assign \new_[78957]_  = ~A170 & \new_[78956]_ ;
  assign \new_[78960]_  = A199 & A166;
  assign \new_[78963]_  = ~A201 & ~A200;
  assign \new_[78964]_  = \new_[78963]_  & \new_[78960]_ ;
  assign \new_[78965]_  = \new_[78964]_  & \new_[78957]_ ;
  assign \new_[78968]_  = ~A203 & ~A202;
  assign \new_[78971]_  = ~A266 & A265;
  assign \new_[78972]_  = \new_[78971]_  & \new_[78968]_ ;
  assign \new_[78975]_  = A268 & A267;
  assign \new_[78978]_  = ~A299 & ~A298;
  assign \new_[78979]_  = \new_[78978]_  & \new_[78975]_ ;
  assign \new_[78980]_  = \new_[78979]_  & \new_[78972]_ ;
  assign \new_[78984]_  = ~A167 & A168;
  assign \new_[78985]_  = ~A170 & \new_[78984]_ ;
  assign \new_[78988]_  = A199 & A166;
  assign \new_[78991]_  = ~A201 & ~A200;
  assign \new_[78992]_  = \new_[78991]_  & \new_[78988]_ ;
  assign \new_[78993]_  = \new_[78992]_  & \new_[78985]_ ;
  assign \new_[78996]_  = ~A203 & ~A202;
  assign \new_[78999]_  = ~A266 & A265;
  assign \new_[79000]_  = \new_[78999]_  & \new_[78996]_ ;
  assign \new_[79003]_  = A269 & A267;
  assign \new_[79006]_  = A301 & ~A300;
  assign \new_[79007]_  = \new_[79006]_  & \new_[79003]_ ;
  assign \new_[79008]_  = \new_[79007]_  & \new_[79000]_ ;
  assign \new_[79012]_  = ~A167 & A168;
  assign \new_[79013]_  = ~A170 & \new_[79012]_ ;
  assign \new_[79016]_  = A199 & A166;
  assign \new_[79019]_  = ~A201 & ~A200;
  assign \new_[79020]_  = \new_[79019]_  & \new_[79016]_ ;
  assign \new_[79021]_  = \new_[79020]_  & \new_[79013]_ ;
  assign \new_[79024]_  = ~A203 & ~A202;
  assign \new_[79027]_  = ~A266 & A265;
  assign \new_[79028]_  = \new_[79027]_  & \new_[79024]_ ;
  assign \new_[79031]_  = A269 & A267;
  assign \new_[79034]_  = A302 & ~A300;
  assign \new_[79035]_  = \new_[79034]_  & \new_[79031]_ ;
  assign \new_[79036]_  = \new_[79035]_  & \new_[79028]_ ;
  assign \new_[79040]_  = ~A167 & A168;
  assign \new_[79041]_  = ~A170 & \new_[79040]_ ;
  assign \new_[79044]_  = A199 & A166;
  assign \new_[79047]_  = ~A201 & ~A200;
  assign \new_[79048]_  = \new_[79047]_  & \new_[79044]_ ;
  assign \new_[79049]_  = \new_[79048]_  & \new_[79041]_ ;
  assign \new_[79052]_  = ~A203 & ~A202;
  assign \new_[79055]_  = ~A266 & A265;
  assign \new_[79056]_  = \new_[79055]_  & \new_[79052]_ ;
  assign \new_[79059]_  = A269 & A267;
  assign \new_[79062]_  = A299 & A298;
  assign \new_[79063]_  = \new_[79062]_  & \new_[79059]_ ;
  assign \new_[79064]_  = \new_[79063]_  & \new_[79056]_ ;
  assign \new_[79068]_  = ~A167 & A168;
  assign \new_[79069]_  = ~A170 & \new_[79068]_ ;
  assign \new_[79072]_  = A199 & A166;
  assign \new_[79075]_  = ~A201 & ~A200;
  assign \new_[79076]_  = \new_[79075]_  & \new_[79072]_ ;
  assign \new_[79077]_  = \new_[79076]_  & \new_[79069]_ ;
  assign \new_[79080]_  = ~A203 & ~A202;
  assign \new_[79083]_  = ~A266 & A265;
  assign \new_[79084]_  = \new_[79083]_  & \new_[79080]_ ;
  assign \new_[79087]_  = A269 & A267;
  assign \new_[79090]_  = ~A299 & ~A298;
  assign \new_[79091]_  = \new_[79090]_  & \new_[79087]_ ;
  assign \new_[79092]_  = \new_[79091]_  & \new_[79084]_ ;
  assign \new_[79096]_  = ~A199 & ~A168;
  assign \new_[79097]_  = ~A170 & \new_[79096]_ ;
  assign \new_[79100]_  = ~A201 & A200;
  assign \new_[79103]_  = ~A203 & ~A202;
  assign \new_[79104]_  = \new_[79103]_  & \new_[79100]_ ;
  assign \new_[79105]_  = \new_[79104]_  & \new_[79097]_ ;
  assign \new_[79108]_  = ~A268 & A267;
  assign \new_[79111]_  = A298 & ~A269;
  assign \new_[79112]_  = \new_[79111]_  & \new_[79108]_ ;
  assign \new_[79115]_  = ~A300 & ~A299;
  assign \new_[79118]_  = ~A302 & ~A301;
  assign \new_[79119]_  = \new_[79118]_  & \new_[79115]_ ;
  assign \new_[79120]_  = \new_[79119]_  & \new_[79112]_ ;
  assign \new_[79124]_  = ~A199 & ~A168;
  assign \new_[79125]_  = ~A170 & \new_[79124]_ ;
  assign \new_[79128]_  = ~A201 & A200;
  assign \new_[79131]_  = ~A203 & ~A202;
  assign \new_[79132]_  = \new_[79131]_  & \new_[79128]_ ;
  assign \new_[79133]_  = \new_[79132]_  & \new_[79125]_ ;
  assign \new_[79136]_  = ~A268 & A267;
  assign \new_[79139]_  = ~A298 & ~A269;
  assign \new_[79140]_  = \new_[79139]_  & \new_[79136]_ ;
  assign \new_[79143]_  = ~A300 & A299;
  assign \new_[79146]_  = ~A302 & ~A301;
  assign \new_[79147]_  = \new_[79146]_  & \new_[79143]_ ;
  assign \new_[79148]_  = \new_[79147]_  & \new_[79140]_ ;
  assign \new_[79152]_  = A199 & ~A168;
  assign \new_[79153]_  = ~A170 & \new_[79152]_ ;
  assign \new_[79156]_  = ~A201 & ~A200;
  assign \new_[79159]_  = ~A203 & ~A202;
  assign \new_[79160]_  = \new_[79159]_  & \new_[79156]_ ;
  assign \new_[79161]_  = \new_[79160]_  & \new_[79153]_ ;
  assign \new_[79164]_  = ~A268 & A267;
  assign \new_[79167]_  = A298 & ~A269;
  assign \new_[79168]_  = \new_[79167]_  & \new_[79164]_ ;
  assign \new_[79171]_  = ~A300 & ~A299;
  assign \new_[79174]_  = ~A302 & ~A301;
  assign \new_[79175]_  = \new_[79174]_  & \new_[79171]_ ;
  assign \new_[79176]_  = \new_[79175]_  & \new_[79168]_ ;
  assign \new_[79180]_  = A199 & ~A168;
  assign \new_[79181]_  = ~A170 & \new_[79180]_ ;
  assign \new_[79184]_  = ~A201 & ~A200;
  assign \new_[79187]_  = ~A203 & ~A202;
  assign \new_[79188]_  = \new_[79187]_  & \new_[79184]_ ;
  assign \new_[79189]_  = \new_[79188]_  & \new_[79181]_ ;
  assign \new_[79192]_  = ~A268 & A267;
  assign \new_[79195]_  = ~A298 & ~A269;
  assign \new_[79196]_  = \new_[79195]_  & \new_[79192]_ ;
  assign \new_[79199]_  = ~A300 & A299;
  assign \new_[79202]_  = ~A302 & ~A301;
  assign \new_[79203]_  = \new_[79202]_  & \new_[79199]_ ;
  assign \new_[79204]_  = \new_[79203]_  & \new_[79196]_ ;
  assign \new_[79208]_  = A167 & A168;
  assign \new_[79209]_  = A169 & \new_[79208]_ ;
  assign \new_[79212]_  = A201 & ~A166;
  assign \new_[79215]_  = ~A203 & ~A202;
  assign \new_[79216]_  = \new_[79215]_  & \new_[79212]_ ;
  assign \new_[79217]_  = \new_[79216]_  & \new_[79209]_ ;
  assign \new_[79220]_  = ~A268 & A267;
  assign \new_[79223]_  = A298 & ~A269;
  assign \new_[79224]_  = \new_[79223]_  & \new_[79220]_ ;
  assign \new_[79227]_  = ~A300 & ~A299;
  assign \new_[79230]_  = ~A302 & ~A301;
  assign \new_[79231]_  = \new_[79230]_  & \new_[79227]_ ;
  assign \new_[79232]_  = \new_[79231]_  & \new_[79224]_ ;
  assign \new_[79236]_  = A167 & A168;
  assign \new_[79237]_  = A169 & \new_[79236]_ ;
  assign \new_[79240]_  = A201 & ~A166;
  assign \new_[79243]_  = ~A203 & ~A202;
  assign \new_[79244]_  = \new_[79243]_  & \new_[79240]_ ;
  assign \new_[79245]_  = \new_[79244]_  & \new_[79237]_ ;
  assign \new_[79248]_  = ~A268 & A267;
  assign \new_[79251]_  = ~A298 & ~A269;
  assign \new_[79252]_  = \new_[79251]_  & \new_[79248]_ ;
  assign \new_[79255]_  = ~A300 & A299;
  assign \new_[79258]_  = ~A302 & ~A301;
  assign \new_[79259]_  = \new_[79258]_  & \new_[79255]_ ;
  assign \new_[79260]_  = \new_[79259]_  & \new_[79252]_ ;
  assign \new_[79264]_  = A167 & A168;
  assign \new_[79265]_  = A169 & \new_[79264]_ ;
  assign \new_[79268]_  = ~A199 & ~A166;
  assign \new_[79271]_  = A201 & A200;
  assign \new_[79272]_  = \new_[79271]_  & \new_[79268]_ ;
  assign \new_[79273]_  = \new_[79272]_  & \new_[79265]_ ;
  assign \new_[79276]_  = ~A265 & A202;
  assign \new_[79279]_  = A267 & A266;
  assign \new_[79280]_  = \new_[79279]_  & \new_[79276]_ ;
  assign \new_[79283]_  = A300 & A268;
  assign \new_[79286]_  = ~A302 & ~A301;
  assign \new_[79287]_  = \new_[79286]_  & \new_[79283]_ ;
  assign \new_[79288]_  = \new_[79287]_  & \new_[79280]_ ;
  assign \new_[79292]_  = A167 & A168;
  assign \new_[79293]_  = A169 & \new_[79292]_ ;
  assign \new_[79296]_  = ~A199 & ~A166;
  assign \new_[79299]_  = A201 & A200;
  assign \new_[79300]_  = \new_[79299]_  & \new_[79296]_ ;
  assign \new_[79301]_  = \new_[79300]_  & \new_[79293]_ ;
  assign \new_[79304]_  = ~A265 & A202;
  assign \new_[79307]_  = A267 & A266;
  assign \new_[79308]_  = \new_[79307]_  & \new_[79304]_ ;
  assign \new_[79311]_  = A300 & A269;
  assign \new_[79314]_  = ~A302 & ~A301;
  assign \new_[79315]_  = \new_[79314]_  & \new_[79311]_ ;
  assign \new_[79316]_  = \new_[79315]_  & \new_[79308]_ ;
  assign \new_[79320]_  = A167 & A168;
  assign \new_[79321]_  = A169 & \new_[79320]_ ;
  assign \new_[79324]_  = ~A199 & ~A166;
  assign \new_[79327]_  = A201 & A200;
  assign \new_[79328]_  = \new_[79327]_  & \new_[79324]_ ;
  assign \new_[79329]_  = \new_[79328]_  & \new_[79321]_ ;
  assign \new_[79332]_  = ~A265 & A202;
  assign \new_[79335]_  = ~A267 & A266;
  assign \new_[79336]_  = \new_[79335]_  & \new_[79332]_ ;
  assign \new_[79339]_  = ~A269 & ~A268;
  assign \new_[79342]_  = A301 & ~A300;
  assign \new_[79343]_  = \new_[79342]_  & \new_[79339]_ ;
  assign \new_[79344]_  = \new_[79343]_  & \new_[79336]_ ;
  assign \new_[79348]_  = A167 & A168;
  assign \new_[79349]_  = A169 & \new_[79348]_ ;
  assign \new_[79352]_  = ~A199 & ~A166;
  assign \new_[79355]_  = A201 & A200;
  assign \new_[79356]_  = \new_[79355]_  & \new_[79352]_ ;
  assign \new_[79357]_  = \new_[79356]_  & \new_[79349]_ ;
  assign \new_[79360]_  = ~A265 & A202;
  assign \new_[79363]_  = ~A267 & A266;
  assign \new_[79364]_  = \new_[79363]_  & \new_[79360]_ ;
  assign \new_[79367]_  = ~A269 & ~A268;
  assign \new_[79370]_  = A302 & ~A300;
  assign \new_[79371]_  = \new_[79370]_  & \new_[79367]_ ;
  assign \new_[79372]_  = \new_[79371]_  & \new_[79364]_ ;
  assign \new_[79376]_  = A167 & A168;
  assign \new_[79377]_  = A169 & \new_[79376]_ ;
  assign \new_[79380]_  = ~A199 & ~A166;
  assign \new_[79383]_  = A201 & A200;
  assign \new_[79384]_  = \new_[79383]_  & \new_[79380]_ ;
  assign \new_[79385]_  = \new_[79384]_  & \new_[79377]_ ;
  assign \new_[79388]_  = ~A265 & A202;
  assign \new_[79391]_  = ~A267 & A266;
  assign \new_[79392]_  = \new_[79391]_  & \new_[79388]_ ;
  assign \new_[79395]_  = ~A269 & ~A268;
  assign \new_[79398]_  = A299 & A298;
  assign \new_[79399]_  = \new_[79398]_  & \new_[79395]_ ;
  assign \new_[79400]_  = \new_[79399]_  & \new_[79392]_ ;
  assign \new_[79404]_  = A167 & A168;
  assign \new_[79405]_  = A169 & \new_[79404]_ ;
  assign \new_[79408]_  = ~A199 & ~A166;
  assign \new_[79411]_  = A201 & A200;
  assign \new_[79412]_  = \new_[79411]_  & \new_[79408]_ ;
  assign \new_[79413]_  = \new_[79412]_  & \new_[79405]_ ;
  assign \new_[79416]_  = ~A265 & A202;
  assign \new_[79419]_  = ~A267 & A266;
  assign \new_[79420]_  = \new_[79419]_  & \new_[79416]_ ;
  assign \new_[79423]_  = ~A269 & ~A268;
  assign \new_[79426]_  = ~A299 & ~A298;
  assign \new_[79427]_  = \new_[79426]_  & \new_[79423]_ ;
  assign \new_[79428]_  = \new_[79427]_  & \new_[79420]_ ;
  assign \new_[79432]_  = A167 & A168;
  assign \new_[79433]_  = A169 & \new_[79432]_ ;
  assign \new_[79436]_  = ~A199 & ~A166;
  assign \new_[79439]_  = A201 & A200;
  assign \new_[79440]_  = \new_[79439]_  & \new_[79436]_ ;
  assign \new_[79441]_  = \new_[79440]_  & \new_[79433]_ ;
  assign \new_[79444]_  = A265 & A202;
  assign \new_[79447]_  = A267 & ~A266;
  assign \new_[79448]_  = \new_[79447]_  & \new_[79444]_ ;
  assign \new_[79451]_  = A300 & A268;
  assign \new_[79454]_  = ~A302 & ~A301;
  assign \new_[79455]_  = \new_[79454]_  & \new_[79451]_ ;
  assign \new_[79456]_  = \new_[79455]_  & \new_[79448]_ ;
  assign \new_[79460]_  = A167 & A168;
  assign \new_[79461]_  = A169 & \new_[79460]_ ;
  assign \new_[79464]_  = ~A199 & ~A166;
  assign \new_[79467]_  = A201 & A200;
  assign \new_[79468]_  = \new_[79467]_  & \new_[79464]_ ;
  assign \new_[79469]_  = \new_[79468]_  & \new_[79461]_ ;
  assign \new_[79472]_  = A265 & A202;
  assign \new_[79475]_  = A267 & ~A266;
  assign \new_[79476]_  = \new_[79475]_  & \new_[79472]_ ;
  assign \new_[79479]_  = A300 & A269;
  assign \new_[79482]_  = ~A302 & ~A301;
  assign \new_[79483]_  = \new_[79482]_  & \new_[79479]_ ;
  assign \new_[79484]_  = \new_[79483]_  & \new_[79476]_ ;
  assign \new_[79488]_  = A167 & A168;
  assign \new_[79489]_  = A169 & \new_[79488]_ ;
  assign \new_[79492]_  = ~A199 & ~A166;
  assign \new_[79495]_  = A201 & A200;
  assign \new_[79496]_  = \new_[79495]_  & \new_[79492]_ ;
  assign \new_[79497]_  = \new_[79496]_  & \new_[79489]_ ;
  assign \new_[79500]_  = A265 & A202;
  assign \new_[79503]_  = ~A267 & ~A266;
  assign \new_[79504]_  = \new_[79503]_  & \new_[79500]_ ;
  assign \new_[79507]_  = ~A269 & ~A268;
  assign \new_[79510]_  = A301 & ~A300;
  assign \new_[79511]_  = \new_[79510]_  & \new_[79507]_ ;
  assign \new_[79512]_  = \new_[79511]_  & \new_[79504]_ ;
  assign \new_[79516]_  = A167 & A168;
  assign \new_[79517]_  = A169 & \new_[79516]_ ;
  assign \new_[79520]_  = ~A199 & ~A166;
  assign \new_[79523]_  = A201 & A200;
  assign \new_[79524]_  = \new_[79523]_  & \new_[79520]_ ;
  assign \new_[79525]_  = \new_[79524]_  & \new_[79517]_ ;
  assign \new_[79528]_  = A265 & A202;
  assign \new_[79531]_  = ~A267 & ~A266;
  assign \new_[79532]_  = \new_[79531]_  & \new_[79528]_ ;
  assign \new_[79535]_  = ~A269 & ~A268;
  assign \new_[79538]_  = A302 & ~A300;
  assign \new_[79539]_  = \new_[79538]_  & \new_[79535]_ ;
  assign \new_[79540]_  = \new_[79539]_  & \new_[79532]_ ;
  assign \new_[79544]_  = A167 & A168;
  assign \new_[79545]_  = A169 & \new_[79544]_ ;
  assign \new_[79548]_  = ~A199 & ~A166;
  assign \new_[79551]_  = A201 & A200;
  assign \new_[79552]_  = \new_[79551]_  & \new_[79548]_ ;
  assign \new_[79553]_  = \new_[79552]_  & \new_[79545]_ ;
  assign \new_[79556]_  = A265 & A202;
  assign \new_[79559]_  = ~A267 & ~A266;
  assign \new_[79560]_  = \new_[79559]_  & \new_[79556]_ ;
  assign \new_[79563]_  = ~A269 & ~A268;
  assign \new_[79566]_  = A299 & A298;
  assign \new_[79567]_  = \new_[79566]_  & \new_[79563]_ ;
  assign \new_[79568]_  = \new_[79567]_  & \new_[79560]_ ;
  assign \new_[79572]_  = A167 & A168;
  assign \new_[79573]_  = A169 & \new_[79572]_ ;
  assign \new_[79576]_  = ~A199 & ~A166;
  assign \new_[79579]_  = A201 & A200;
  assign \new_[79580]_  = \new_[79579]_  & \new_[79576]_ ;
  assign \new_[79581]_  = \new_[79580]_  & \new_[79573]_ ;
  assign \new_[79584]_  = A265 & A202;
  assign \new_[79587]_  = ~A267 & ~A266;
  assign \new_[79588]_  = \new_[79587]_  & \new_[79584]_ ;
  assign \new_[79591]_  = ~A269 & ~A268;
  assign \new_[79594]_  = ~A299 & ~A298;
  assign \new_[79595]_  = \new_[79594]_  & \new_[79591]_ ;
  assign \new_[79596]_  = \new_[79595]_  & \new_[79588]_ ;
  assign \new_[79600]_  = A167 & A168;
  assign \new_[79601]_  = A169 & \new_[79600]_ ;
  assign \new_[79604]_  = ~A199 & ~A166;
  assign \new_[79607]_  = A201 & A200;
  assign \new_[79608]_  = \new_[79607]_  & \new_[79604]_ ;
  assign \new_[79609]_  = \new_[79608]_  & \new_[79601]_ ;
  assign \new_[79612]_  = ~A265 & A203;
  assign \new_[79615]_  = A267 & A266;
  assign \new_[79616]_  = \new_[79615]_  & \new_[79612]_ ;
  assign \new_[79619]_  = A300 & A268;
  assign \new_[79622]_  = ~A302 & ~A301;
  assign \new_[79623]_  = \new_[79622]_  & \new_[79619]_ ;
  assign \new_[79624]_  = \new_[79623]_  & \new_[79616]_ ;
  assign \new_[79628]_  = A167 & A168;
  assign \new_[79629]_  = A169 & \new_[79628]_ ;
  assign \new_[79632]_  = ~A199 & ~A166;
  assign \new_[79635]_  = A201 & A200;
  assign \new_[79636]_  = \new_[79635]_  & \new_[79632]_ ;
  assign \new_[79637]_  = \new_[79636]_  & \new_[79629]_ ;
  assign \new_[79640]_  = ~A265 & A203;
  assign \new_[79643]_  = A267 & A266;
  assign \new_[79644]_  = \new_[79643]_  & \new_[79640]_ ;
  assign \new_[79647]_  = A300 & A269;
  assign \new_[79650]_  = ~A302 & ~A301;
  assign \new_[79651]_  = \new_[79650]_  & \new_[79647]_ ;
  assign \new_[79652]_  = \new_[79651]_  & \new_[79644]_ ;
  assign \new_[79656]_  = A167 & A168;
  assign \new_[79657]_  = A169 & \new_[79656]_ ;
  assign \new_[79660]_  = ~A199 & ~A166;
  assign \new_[79663]_  = A201 & A200;
  assign \new_[79664]_  = \new_[79663]_  & \new_[79660]_ ;
  assign \new_[79665]_  = \new_[79664]_  & \new_[79657]_ ;
  assign \new_[79668]_  = ~A265 & A203;
  assign \new_[79671]_  = ~A267 & A266;
  assign \new_[79672]_  = \new_[79671]_  & \new_[79668]_ ;
  assign \new_[79675]_  = ~A269 & ~A268;
  assign \new_[79678]_  = A301 & ~A300;
  assign \new_[79679]_  = \new_[79678]_  & \new_[79675]_ ;
  assign \new_[79680]_  = \new_[79679]_  & \new_[79672]_ ;
  assign \new_[79684]_  = A167 & A168;
  assign \new_[79685]_  = A169 & \new_[79684]_ ;
  assign \new_[79688]_  = ~A199 & ~A166;
  assign \new_[79691]_  = A201 & A200;
  assign \new_[79692]_  = \new_[79691]_  & \new_[79688]_ ;
  assign \new_[79693]_  = \new_[79692]_  & \new_[79685]_ ;
  assign \new_[79696]_  = ~A265 & A203;
  assign \new_[79699]_  = ~A267 & A266;
  assign \new_[79700]_  = \new_[79699]_  & \new_[79696]_ ;
  assign \new_[79703]_  = ~A269 & ~A268;
  assign \new_[79706]_  = A302 & ~A300;
  assign \new_[79707]_  = \new_[79706]_  & \new_[79703]_ ;
  assign \new_[79708]_  = \new_[79707]_  & \new_[79700]_ ;
  assign \new_[79712]_  = A167 & A168;
  assign \new_[79713]_  = A169 & \new_[79712]_ ;
  assign \new_[79716]_  = ~A199 & ~A166;
  assign \new_[79719]_  = A201 & A200;
  assign \new_[79720]_  = \new_[79719]_  & \new_[79716]_ ;
  assign \new_[79721]_  = \new_[79720]_  & \new_[79713]_ ;
  assign \new_[79724]_  = ~A265 & A203;
  assign \new_[79727]_  = ~A267 & A266;
  assign \new_[79728]_  = \new_[79727]_  & \new_[79724]_ ;
  assign \new_[79731]_  = ~A269 & ~A268;
  assign \new_[79734]_  = A299 & A298;
  assign \new_[79735]_  = \new_[79734]_  & \new_[79731]_ ;
  assign \new_[79736]_  = \new_[79735]_  & \new_[79728]_ ;
  assign \new_[79740]_  = A167 & A168;
  assign \new_[79741]_  = A169 & \new_[79740]_ ;
  assign \new_[79744]_  = ~A199 & ~A166;
  assign \new_[79747]_  = A201 & A200;
  assign \new_[79748]_  = \new_[79747]_  & \new_[79744]_ ;
  assign \new_[79749]_  = \new_[79748]_  & \new_[79741]_ ;
  assign \new_[79752]_  = ~A265 & A203;
  assign \new_[79755]_  = ~A267 & A266;
  assign \new_[79756]_  = \new_[79755]_  & \new_[79752]_ ;
  assign \new_[79759]_  = ~A269 & ~A268;
  assign \new_[79762]_  = ~A299 & ~A298;
  assign \new_[79763]_  = \new_[79762]_  & \new_[79759]_ ;
  assign \new_[79764]_  = \new_[79763]_  & \new_[79756]_ ;
  assign \new_[79768]_  = A167 & A168;
  assign \new_[79769]_  = A169 & \new_[79768]_ ;
  assign \new_[79772]_  = ~A199 & ~A166;
  assign \new_[79775]_  = A201 & A200;
  assign \new_[79776]_  = \new_[79775]_  & \new_[79772]_ ;
  assign \new_[79777]_  = \new_[79776]_  & \new_[79769]_ ;
  assign \new_[79780]_  = A265 & A203;
  assign \new_[79783]_  = A267 & ~A266;
  assign \new_[79784]_  = \new_[79783]_  & \new_[79780]_ ;
  assign \new_[79787]_  = A300 & A268;
  assign \new_[79790]_  = ~A302 & ~A301;
  assign \new_[79791]_  = \new_[79790]_  & \new_[79787]_ ;
  assign \new_[79792]_  = \new_[79791]_  & \new_[79784]_ ;
  assign \new_[79796]_  = A167 & A168;
  assign \new_[79797]_  = A169 & \new_[79796]_ ;
  assign \new_[79800]_  = ~A199 & ~A166;
  assign \new_[79803]_  = A201 & A200;
  assign \new_[79804]_  = \new_[79803]_  & \new_[79800]_ ;
  assign \new_[79805]_  = \new_[79804]_  & \new_[79797]_ ;
  assign \new_[79808]_  = A265 & A203;
  assign \new_[79811]_  = A267 & ~A266;
  assign \new_[79812]_  = \new_[79811]_  & \new_[79808]_ ;
  assign \new_[79815]_  = A300 & A269;
  assign \new_[79818]_  = ~A302 & ~A301;
  assign \new_[79819]_  = \new_[79818]_  & \new_[79815]_ ;
  assign \new_[79820]_  = \new_[79819]_  & \new_[79812]_ ;
  assign \new_[79824]_  = A167 & A168;
  assign \new_[79825]_  = A169 & \new_[79824]_ ;
  assign \new_[79828]_  = ~A199 & ~A166;
  assign \new_[79831]_  = A201 & A200;
  assign \new_[79832]_  = \new_[79831]_  & \new_[79828]_ ;
  assign \new_[79833]_  = \new_[79832]_  & \new_[79825]_ ;
  assign \new_[79836]_  = A265 & A203;
  assign \new_[79839]_  = ~A267 & ~A266;
  assign \new_[79840]_  = \new_[79839]_  & \new_[79836]_ ;
  assign \new_[79843]_  = ~A269 & ~A268;
  assign \new_[79846]_  = A301 & ~A300;
  assign \new_[79847]_  = \new_[79846]_  & \new_[79843]_ ;
  assign \new_[79848]_  = \new_[79847]_  & \new_[79840]_ ;
  assign \new_[79852]_  = A167 & A168;
  assign \new_[79853]_  = A169 & \new_[79852]_ ;
  assign \new_[79856]_  = ~A199 & ~A166;
  assign \new_[79859]_  = A201 & A200;
  assign \new_[79860]_  = \new_[79859]_  & \new_[79856]_ ;
  assign \new_[79861]_  = \new_[79860]_  & \new_[79853]_ ;
  assign \new_[79864]_  = A265 & A203;
  assign \new_[79867]_  = ~A267 & ~A266;
  assign \new_[79868]_  = \new_[79867]_  & \new_[79864]_ ;
  assign \new_[79871]_  = ~A269 & ~A268;
  assign \new_[79874]_  = A302 & ~A300;
  assign \new_[79875]_  = \new_[79874]_  & \new_[79871]_ ;
  assign \new_[79876]_  = \new_[79875]_  & \new_[79868]_ ;
  assign \new_[79880]_  = A167 & A168;
  assign \new_[79881]_  = A169 & \new_[79880]_ ;
  assign \new_[79884]_  = ~A199 & ~A166;
  assign \new_[79887]_  = A201 & A200;
  assign \new_[79888]_  = \new_[79887]_  & \new_[79884]_ ;
  assign \new_[79889]_  = \new_[79888]_  & \new_[79881]_ ;
  assign \new_[79892]_  = A265 & A203;
  assign \new_[79895]_  = ~A267 & ~A266;
  assign \new_[79896]_  = \new_[79895]_  & \new_[79892]_ ;
  assign \new_[79899]_  = ~A269 & ~A268;
  assign \new_[79902]_  = A299 & A298;
  assign \new_[79903]_  = \new_[79902]_  & \new_[79899]_ ;
  assign \new_[79904]_  = \new_[79903]_  & \new_[79896]_ ;
  assign \new_[79908]_  = A167 & A168;
  assign \new_[79909]_  = A169 & \new_[79908]_ ;
  assign \new_[79912]_  = ~A199 & ~A166;
  assign \new_[79915]_  = A201 & A200;
  assign \new_[79916]_  = \new_[79915]_  & \new_[79912]_ ;
  assign \new_[79917]_  = \new_[79916]_  & \new_[79909]_ ;
  assign \new_[79920]_  = A265 & A203;
  assign \new_[79923]_  = ~A267 & ~A266;
  assign \new_[79924]_  = \new_[79923]_  & \new_[79920]_ ;
  assign \new_[79927]_  = ~A269 & ~A268;
  assign \new_[79930]_  = ~A299 & ~A298;
  assign \new_[79931]_  = \new_[79930]_  & \new_[79927]_ ;
  assign \new_[79932]_  = \new_[79931]_  & \new_[79924]_ ;
  assign \new_[79936]_  = A167 & A168;
  assign \new_[79937]_  = A169 & \new_[79936]_ ;
  assign \new_[79940]_  = ~A199 & ~A166;
  assign \new_[79943]_  = ~A201 & A200;
  assign \new_[79944]_  = \new_[79943]_  & \new_[79940]_ ;
  assign \new_[79945]_  = \new_[79944]_  & \new_[79937]_ ;
  assign \new_[79948]_  = ~A203 & ~A202;
  assign \new_[79951]_  = A266 & ~A265;
  assign \new_[79952]_  = \new_[79951]_  & \new_[79948]_ ;
  assign \new_[79955]_  = A268 & A267;
  assign \new_[79958]_  = A301 & ~A300;
  assign \new_[79959]_  = \new_[79958]_  & \new_[79955]_ ;
  assign \new_[79960]_  = \new_[79959]_  & \new_[79952]_ ;
  assign \new_[79964]_  = A167 & A168;
  assign \new_[79965]_  = A169 & \new_[79964]_ ;
  assign \new_[79968]_  = ~A199 & ~A166;
  assign \new_[79971]_  = ~A201 & A200;
  assign \new_[79972]_  = \new_[79971]_  & \new_[79968]_ ;
  assign \new_[79973]_  = \new_[79972]_  & \new_[79965]_ ;
  assign \new_[79976]_  = ~A203 & ~A202;
  assign \new_[79979]_  = A266 & ~A265;
  assign \new_[79980]_  = \new_[79979]_  & \new_[79976]_ ;
  assign \new_[79983]_  = A268 & A267;
  assign \new_[79986]_  = A302 & ~A300;
  assign \new_[79987]_  = \new_[79986]_  & \new_[79983]_ ;
  assign \new_[79988]_  = \new_[79987]_  & \new_[79980]_ ;
  assign \new_[79992]_  = A167 & A168;
  assign \new_[79993]_  = A169 & \new_[79992]_ ;
  assign \new_[79996]_  = ~A199 & ~A166;
  assign \new_[79999]_  = ~A201 & A200;
  assign \new_[80000]_  = \new_[79999]_  & \new_[79996]_ ;
  assign \new_[80001]_  = \new_[80000]_  & \new_[79993]_ ;
  assign \new_[80004]_  = ~A203 & ~A202;
  assign \new_[80007]_  = A266 & ~A265;
  assign \new_[80008]_  = \new_[80007]_  & \new_[80004]_ ;
  assign \new_[80011]_  = A268 & A267;
  assign \new_[80014]_  = A299 & A298;
  assign \new_[80015]_  = \new_[80014]_  & \new_[80011]_ ;
  assign \new_[80016]_  = \new_[80015]_  & \new_[80008]_ ;
  assign \new_[80020]_  = A167 & A168;
  assign \new_[80021]_  = A169 & \new_[80020]_ ;
  assign \new_[80024]_  = ~A199 & ~A166;
  assign \new_[80027]_  = ~A201 & A200;
  assign \new_[80028]_  = \new_[80027]_  & \new_[80024]_ ;
  assign \new_[80029]_  = \new_[80028]_  & \new_[80021]_ ;
  assign \new_[80032]_  = ~A203 & ~A202;
  assign \new_[80035]_  = A266 & ~A265;
  assign \new_[80036]_  = \new_[80035]_  & \new_[80032]_ ;
  assign \new_[80039]_  = A268 & A267;
  assign \new_[80042]_  = ~A299 & ~A298;
  assign \new_[80043]_  = \new_[80042]_  & \new_[80039]_ ;
  assign \new_[80044]_  = \new_[80043]_  & \new_[80036]_ ;
  assign \new_[80048]_  = A167 & A168;
  assign \new_[80049]_  = A169 & \new_[80048]_ ;
  assign \new_[80052]_  = ~A199 & ~A166;
  assign \new_[80055]_  = ~A201 & A200;
  assign \new_[80056]_  = \new_[80055]_  & \new_[80052]_ ;
  assign \new_[80057]_  = \new_[80056]_  & \new_[80049]_ ;
  assign \new_[80060]_  = ~A203 & ~A202;
  assign \new_[80063]_  = A266 & ~A265;
  assign \new_[80064]_  = \new_[80063]_  & \new_[80060]_ ;
  assign \new_[80067]_  = A269 & A267;
  assign \new_[80070]_  = A301 & ~A300;
  assign \new_[80071]_  = \new_[80070]_  & \new_[80067]_ ;
  assign \new_[80072]_  = \new_[80071]_  & \new_[80064]_ ;
  assign \new_[80076]_  = A167 & A168;
  assign \new_[80077]_  = A169 & \new_[80076]_ ;
  assign \new_[80080]_  = ~A199 & ~A166;
  assign \new_[80083]_  = ~A201 & A200;
  assign \new_[80084]_  = \new_[80083]_  & \new_[80080]_ ;
  assign \new_[80085]_  = \new_[80084]_  & \new_[80077]_ ;
  assign \new_[80088]_  = ~A203 & ~A202;
  assign \new_[80091]_  = A266 & ~A265;
  assign \new_[80092]_  = \new_[80091]_  & \new_[80088]_ ;
  assign \new_[80095]_  = A269 & A267;
  assign \new_[80098]_  = A302 & ~A300;
  assign \new_[80099]_  = \new_[80098]_  & \new_[80095]_ ;
  assign \new_[80100]_  = \new_[80099]_  & \new_[80092]_ ;
  assign \new_[80104]_  = A167 & A168;
  assign \new_[80105]_  = A169 & \new_[80104]_ ;
  assign \new_[80108]_  = ~A199 & ~A166;
  assign \new_[80111]_  = ~A201 & A200;
  assign \new_[80112]_  = \new_[80111]_  & \new_[80108]_ ;
  assign \new_[80113]_  = \new_[80112]_  & \new_[80105]_ ;
  assign \new_[80116]_  = ~A203 & ~A202;
  assign \new_[80119]_  = A266 & ~A265;
  assign \new_[80120]_  = \new_[80119]_  & \new_[80116]_ ;
  assign \new_[80123]_  = A269 & A267;
  assign \new_[80126]_  = A299 & A298;
  assign \new_[80127]_  = \new_[80126]_  & \new_[80123]_ ;
  assign \new_[80128]_  = \new_[80127]_  & \new_[80120]_ ;
  assign \new_[80132]_  = A167 & A168;
  assign \new_[80133]_  = A169 & \new_[80132]_ ;
  assign \new_[80136]_  = ~A199 & ~A166;
  assign \new_[80139]_  = ~A201 & A200;
  assign \new_[80140]_  = \new_[80139]_  & \new_[80136]_ ;
  assign \new_[80141]_  = \new_[80140]_  & \new_[80133]_ ;
  assign \new_[80144]_  = ~A203 & ~A202;
  assign \new_[80147]_  = A266 & ~A265;
  assign \new_[80148]_  = \new_[80147]_  & \new_[80144]_ ;
  assign \new_[80151]_  = A269 & A267;
  assign \new_[80154]_  = ~A299 & ~A298;
  assign \new_[80155]_  = \new_[80154]_  & \new_[80151]_ ;
  assign \new_[80156]_  = \new_[80155]_  & \new_[80148]_ ;
  assign \new_[80160]_  = A167 & A168;
  assign \new_[80161]_  = A169 & \new_[80160]_ ;
  assign \new_[80164]_  = ~A199 & ~A166;
  assign \new_[80167]_  = ~A201 & A200;
  assign \new_[80168]_  = \new_[80167]_  & \new_[80164]_ ;
  assign \new_[80169]_  = \new_[80168]_  & \new_[80161]_ ;
  assign \new_[80172]_  = ~A203 & ~A202;
  assign \new_[80175]_  = ~A266 & A265;
  assign \new_[80176]_  = \new_[80175]_  & \new_[80172]_ ;
  assign \new_[80179]_  = A268 & A267;
  assign \new_[80182]_  = A301 & ~A300;
  assign \new_[80183]_  = \new_[80182]_  & \new_[80179]_ ;
  assign \new_[80184]_  = \new_[80183]_  & \new_[80176]_ ;
  assign \new_[80188]_  = A167 & A168;
  assign \new_[80189]_  = A169 & \new_[80188]_ ;
  assign \new_[80192]_  = ~A199 & ~A166;
  assign \new_[80195]_  = ~A201 & A200;
  assign \new_[80196]_  = \new_[80195]_  & \new_[80192]_ ;
  assign \new_[80197]_  = \new_[80196]_  & \new_[80189]_ ;
  assign \new_[80200]_  = ~A203 & ~A202;
  assign \new_[80203]_  = ~A266 & A265;
  assign \new_[80204]_  = \new_[80203]_  & \new_[80200]_ ;
  assign \new_[80207]_  = A268 & A267;
  assign \new_[80210]_  = A302 & ~A300;
  assign \new_[80211]_  = \new_[80210]_  & \new_[80207]_ ;
  assign \new_[80212]_  = \new_[80211]_  & \new_[80204]_ ;
  assign \new_[80216]_  = A167 & A168;
  assign \new_[80217]_  = A169 & \new_[80216]_ ;
  assign \new_[80220]_  = ~A199 & ~A166;
  assign \new_[80223]_  = ~A201 & A200;
  assign \new_[80224]_  = \new_[80223]_  & \new_[80220]_ ;
  assign \new_[80225]_  = \new_[80224]_  & \new_[80217]_ ;
  assign \new_[80228]_  = ~A203 & ~A202;
  assign \new_[80231]_  = ~A266 & A265;
  assign \new_[80232]_  = \new_[80231]_  & \new_[80228]_ ;
  assign \new_[80235]_  = A268 & A267;
  assign \new_[80238]_  = A299 & A298;
  assign \new_[80239]_  = \new_[80238]_  & \new_[80235]_ ;
  assign \new_[80240]_  = \new_[80239]_  & \new_[80232]_ ;
  assign \new_[80244]_  = A167 & A168;
  assign \new_[80245]_  = A169 & \new_[80244]_ ;
  assign \new_[80248]_  = ~A199 & ~A166;
  assign \new_[80251]_  = ~A201 & A200;
  assign \new_[80252]_  = \new_[80251]_  & \new_[80248]_ ;
  assign \new_[80253]_  = \new_[80252]_  & \new_[80245]_ ;
  assign \new_[80256]_  = ~A203 & ~A202;
  assign \new_[80259]_  = ~A266 & A265;
  assign \new_[80260]_  = \new_[80259]_  & \new_[80256]_ ;
  assign \new_[80263]_  = A268 & A267;
  assign \new_[80266]_  = ~A299 & ~A298;
  assign \new_[80267]_  = \new_[80266]_  & \new_[80263]_ ;
  assign \new_[80268]_  = \new_[80267]_  & \new_[80260]_ ;
  assign \new_[80272]_  = A167 & A168;
  assign \new_[80273]_  = A169 & \new_[80272]_ ;
  assign \new_[80276]_  = ~A199 & ~A166;
  assign \new_[80279]_  = ~A201 & A200;
  assign \new_[80280]_  = \new_[80279]_  & \new_[80276]_ ;
  assign \new_[80281]_  = \new_[80280]_  & \new_[80273]_ ;
  assign \new_[80284]_  = ~A203 & ~A202;
  assign \new_[80287]_  = ~A266 & A265;
  assign \new_[80288]_  = \new_[80287]_  & \new_[80284]_ ;
  assign \new_[80291]_  = A269 & A267;
  assign \new_[80294]_  = A301 & ~A300;
  assign \new_[80295]_  = \new_[80294]_  & \new_[80291]_ ;
  assign \new_[80296]_  = \new_[80295]_  & \new_[80288]_ ;
  assign \new_[80300]_  = A167 & A168;
  assign \new_[80301]_  = A169 & \new_[80300]_ ;
  assign \new_[80304]_  = ~A199 & ~A166;
  assign \new_[80307]_  = ~A201 & A200;
  assign \new_[80308]_  = \new_[80307]_  & \new_[80304]_ ;
  assign \new_[80309]_  = \new_[80308]_  & \new_[80301]_ ;
  assign \new_[80312]_  = ~A203 & ~A202;
  assign \new_[80315]_  = ~A266 & A265;
  assign \new_[80316]_  = \new_[80315]_  & \new_[80312]_ ;
  assign \new_[80319]_  = A269 & A267;
  assign \new_[80322]_  = A302 & ~A300;
  assign \new_[80323]_  = \new_[80322]_  & \new_[80319]_ ;
  assign \new_[80324]_  = \new_[80323]_  & \new_[80316]_ ;
  assign \new_[80328]_  = A167 & A168;
  assign \new_[80329]_  = A169 & \new_[80328]_ ;
  assign \new_[80332]_  = ~A199 & ~A166;
  assign \new_[80335]_  = ~A201 & A200;
  assign \new_[80336]_  = \new_[80335]_  & \new_[80332]_ ;
  assign \new_[80337]_  = \new_[80336]_  & \new_[80329]_ ;
  assign \new_[80340]_  = ~A203 & ~A202;
  assign \new_[80343]_  = ~A266 & A265;
  assign \new_[80344]_  = \new_[80343]_  & \new_[80340]_ ;
  assign \new_[80347]_  = A269 & A267;
  assign \new_[80350]_  = A299 & A298;
  assign \new_[80351]_  = \new_[80350]_  & \new_[80347]_ ;
  assign \new_[80352]_  = \new_[80351]_  & \new_[80344]_ ;
  assign \new_[80356]_  = A167 & A168;
  assign \new_[80357]_  = A169 & \new_[80356]_ ;
  assign \new_[80360]_  = ~A199 & ~A166;
  assign \new_[80363]_  = ~A201 & A200;
  assign \new_[80364]_  = \new_[80363]_  & \new_[80360]_ ;
  assign \new_[80365]_  = \new_[80364]_  & \new_[80357]_ ;
  assign \new_[80368]_  = ~A203 & ~A202;
  assign \new_[80371]_  = ~A266 & A265;
  assign \new_[80372]_  = \new_[80371]_  & \new_[80368]_ ;
  assign \new_[80375]_  = A269 & A267;
  assign \new_[80378]_  = ~A299 & ~A298;
  assign \new_[80379]_  = \new_[80378]_  & \new_[80375]_ ;
  assign \new_[80380]_  = \new_[80379]_  & \new_[80372]_ ;
  assign \new_[80384]_  = A167 & A168;
  assign \new_[80385]_  = A169 & \new_[80384]_ ;
  assign \new_[80388]_  = A199 & ~A166;
  assign \new_[80391]_  = A201 & ~A200;
  assign \new_[80392]_  = \new_[80391]_  & \new_[80388]_ ;
  assign \new_[80393]_  = \new_[80392]_  & \new_[80385]_ ;
  assign \new_[80396]_  = ~A265 & A202;
  assign \new_[80399]_  = A267 & A266;
  assign \new_[80400]_  = \new_[80399]_  & \new_[80396]_ ;
  assign \new_[80403]_  = A300 & A268;
  assign \new_[80406]_  = ~A302 & ~A301;
  assign \new_[80407]_  = \new_[80406]_  & \new_[80403]_ ;
  assign \new_[80408]_  = \new_[80407]_  & \new_[80400]_ ;
  assign \new_[80412]_  = A167 & A168;
  assign \new_[80413]_  = A169 & \new_[80412]_ ;
  assign \new_[80416]_  = A199 & ~A166;
  assign \new_[80419]_  = A201 & ~A200;
  assign \new_[80420]_  = \new_[80419]_  & \new_[80416]_ ;
  assign \new_[80421]_  = \new_[80420]_  & \new_[80413]_ ;
  assign \new_[80424]_  = ~A265 & A202;
  assign \new_[80427]_  = A267 & A266;
  assign \new_[80428]_  = \new_[80427]_  & \new_[80424]_ ;
  assign \new_[80431]_  = A300 & A269;
  assign \new_[80434]_  = ~A302 & ~A301;
  assign \new_[80435]_  = \new_[80434]_  & \new_[80431]_ ;
  assign \new_[80436]_  = \new_[80435]_  & \new_[80428]_ ;
  assign \new_[80440]_  = A167 & A168;
  assign \new_[80441]_  = A169 & \new_[80440]_ ;
  assign \new_[80444]_  = A199 & ~A166;
  assign \new_[80447]_  = A201 & ~A200;
  assign \new_[80448]_  = \new_[80447]_  & \new_[80444]_ ;
  assign \new_[80449]_  = \new_[80448]_  & \new_[80441]_ ;
  assign \new_[80452]_  = ~A265 & A202;
  assign \new_[80455]_  = ~A267 & A266;
  assign \new_[80456]_  = \new_[80455]_  & \new_[80452]_ ;
  assign \new_[80459]_  = ~A269 & ~A268;
  assign \new_[80462]_  = A301 & ~A300;
  assign \new_[80463]_  = \new_[80462]_  & \new_[80459]_ ;
  assign \new_[80464]_  = \new_[80463]_  & \new_[80456]_ ;
  assign \new_[80468]_  = A167 & A168;
  assign \new_[80469]_  = A169 & \new_[80468]_ ;
  assign \new_[80472]_  = A199 & ~A166;
  assign \new_[80475]_  = A201 & ~A200;
  assign \new_[80476]_  = \new_[80475]_  & \new_[80472]_ ;
  assign \new_[80477]_  = \new_[80476]_  & \new_[80469]_ ;
  assign \new_[80480]_  = ~A265 & A202;
  assign \new_[80483]_  = ~A267 & A266;
  assign \new_[80484]_  = \new_[80483]_  & \new_[80480]_ ;
  assign \new_[80487]_  = ~A269 & ~A268;
  assign \new_[80490]_  = A302 & ~A300;
  assign \new_[80491]_  = \new_[80490]_  & \new_[80487]_ ;
  assign \new_[80492]_  = \new_[80491]_  & \new_[80484]_ ;
  assign \new_[80496]_  = A167 & A168;
  assign \new_[80497]_  = A169 & \new_[80496]_ ;
  assign \new_[80500]_  = A199 & ~A166;
  assign \new_[80503]_  = A201 & ~A200;
  assign \new_[80504]_  = \new_[80503]_  & \new_[80500]_ ;
  assign \new_[80505]_  = \new_[80504]_  & \new_[80497]_ ;
  assign \new_[80508]_  = ~A265 & A202;
  assign \new_[80511]_  = ~A267 & A266;
  assign \new_[80512]_  = \new_[80511]_  & \new_[80508]_ ;
  assign \new_[80515]_  = ~A269 & ~A268;
  assign \new_[80518]_  = A299 & A298;
  assign \new_[80519]_  = \new_[80518]_  & \new_[80515]_ ;
  assign \new_[80520]_  = \new_[80519]_  & \new_[80512]_ ;
  assign \new_[80524]_  = A167 & A168;
  assign \new_[80525]_  = A169 & \new_[80524]_ ;
  assign \new_[80528]_  = A199 & ~A166;
  assign \new_[80531]_  = A201 & ~A200;
  assign \new_[80532]_  = \new_[80531]_  & \new_[80528]_ ;
  assign \new_[80533]_  = \new_[80532]_  & \new_[80525]_ ;
  assign \new_[80536]_  = ~A265 & A202;
  assign \new_[80539]_  = ~A267 & A266;
  assign \new_[80540]_  = \new_[80539]_  & \new_[80536]_ ;
  assign \new_[80543]_  = ~A269 & ~A268;
  assign \new_[80546]_  = ~A299 & ~A298;
  assign \new_[80547]_  = \new_[80546]_  & \new_[80543]_ ;
  assign \new_[80548]_  = \new_[80547]_  & \new_[80540]_ ;
  assign \new_[80552]_  = A167 & A168;
  assign \new_[80553]_  = A169 & \new_[80552]_ ;
  assign \new_[80556]_  = A199 & ~A166;
  assign \new_[80559]_  = A201 & ~A200;
  assign \new_[80560]_  = \new_[80559]_  & \new_[80556]_ ;
  assign \new_[80561]_  = \new_[80560]_  & \new_[80553]_ ;
  assign \new_[80564]_  = A265 & A202;
  assign \new_[80567]_  = A267 & ~A266;
  assign \new_[80568]_  = \new_[80567]_  & \new_[80564]_ ;
  assign \new_[80571]_  = A300 & A268;
  assign \new_[80574]_  = ~A302 & ~A301;
  assign \new_[80575]_  = \new_[80574]_  & \new_[80571]_ ;
  assign \new_[80576]_  = \new_[80575]_  & \new_[80568]_ ;
  assign \new_[80580]_  = A167 & A168;
  assign \new_[80581]_  = A169 & \new_[80580]_ ;
  assign \new_[80584]_  = A199 & ~A166;
  assign \new_[80587]_  = A201 & ~A200;
  assign \new_[80588]_  = \new_[80587]_  & \new_[80584]_ ;
  assign \new_[80589]_  = \new_[80588]_  & \new_[80581]_ ;
  assign \new_[80592]_  = A265 & A202;
  assign \new_[80595]_  = A267 & ~A266;
  assign \new_[80596]_  = \new_[80595]_  & \new_[80592]_ ;
  assign \new_[80599]_  = A300 & A269;
  assign \new_[80602]_  = ~A302 & ~A301;
  assign \new_[80603]_  = \new_[80602]_  & \new_[80599]_ ;
  assign \new_[80604]_  = \new_[80603]_  & \new_[80596]_ ;
  assign \new_[80608]_  = A167 & A168;
  assign \new_[80609]_  = A169 & \new_[80608]_ ;
  assign \new_[80612]_  = A199 & ~A166;
  assign \new_[80615]_  = A201 & ~A200;
  assign \new_[80616]_  = \new_[80615]_  & \new_[80612]_ ;
  assign \new_[80617]_  = \new_[80616]_  & \new_[80609]_ ;
  assign \new_[80620]_  = A265 & A202;
  assign \new_[80623]_  = ~A267 & ~A266;
  assign \new_[80624]_  = \new_[80623]_  & \new_[80620]_ ;
  assign \new_[80627]_  = ~A269 & ~A268;
  assign \new_[80630]_  = A301 & ~A300;
  assign \new_[80631]_  = \new_[80630]_  & \new_[80627]_ ;
  assign \new_[80632]_  = \new_[80631]_  & \new_[80624]_ ;
  assign \new_[80636]_  = A167 & A168;
  assign \new_[80637]_  = A169 & \new_[80636]_ ;
  assign \new_[80640]_  = A199 & ~A166;
  assign \new_[80643]_  = A201 & ~A200;
  assign \new_[80644]_  = \new_[80643]_  & \new_[80640]_ ;
  assign \new_[80645]_  = \new_[80644]_  & \new_[80637]_ ;
  assign \new_[80648]_  = A265 & A202;
  assign \new_[80651]_  = ~A267 & ~A266;
  assign \new_[80652]_  = \new_[80651]_  & \new_[80648]_ ;
  assign \new_[80655]_  = ~A269 & ~A268;
  assign \new_[80658]_  = A302 & ~A300;
  assign \new_[80659]_  = \new_[80658]_  & \new_[80655]_ ;
  assign \new_[80660]_  = \new_[80659]_  & \new_[80652]_ ;
  assign \new_[80664]_  = A167 & A168;
  assign \new_[80665]_  = A169 & \new_[80664]_ ;
  assign \new_[80668]_  = A199 & ~A166;
  assign \new_[80671]_  = A201 & ~A200;
  assign \new_[80672]_  = \new_[80671]_  & \new_[80668]_ ;
  assign \new_[80673]_  = \new_[80672]_  & \new_[80665]_ ;
  assign \new_[80676]_  = A265 & A202;
  assign \new_[80679]_  = ~A267 & ~A266;
  assign \new_[80680]_  = \new_[80679]_  & \new_[80676]_ ;
  assign \new_[80683]_  = ~A269 & ~A268;
  assign \new_[80686]_  = A299 & A298;
  assign \new_[80687]_  = \new_[80686]_  & \new_[80683]_ ;
  assign \new_[80688]_  = \new_[80687]_  & \new_[80680]_ ;
  assign \new_[80692]_  = A167 & A168;
  assign \new_[80693]_  = A169 & \new_[80692]_ ;
  assign \new_[80696]_  = A199 & ~A166;
  assign \new_[80699]_  = A201 & ~A200;
  assign \new_[80700]_  = \new_[80699]_  & \new_[80696]_ ;
  assign \new_[80701]_  = \new_[80700]_  & \new_[80693]_ ;
  assign \new_[80704]_  = A265 & A202;
  assign \new_[80707]_  = ~A267 & ~A266;
  assign \new_[80708]_  = \new_[80707]_  & \new_[80704]_ ;
  assign \new_[80711]_  = ~A269 & ~A268;
  assign \new_[80714]_  = ~A299 & ~A298;
  assign \new_[80715]_  = \new_[80714]_  & \new_[80711]_ ;
  assign \new_[80716]_  = \new_[80715]_  & \new_[80708]_ ;
  assign \new_[80720]_  = A167 & A168;
  assign \new_[80721]_  = A169 & \new_[80720]_ ;
  assign \new_[80724]_  = A199 & ~A166;
  assign \new_[80727]_  = A201 & ~A200;
  assign \new_[80728]_  = \new_[80727]_  & \new_[80724]_ ;
  assign \new_[80729]_  = \new_[80728]_  & \new_[80721]_ ;
  assign \new_[80732]_  = ~A265 & A203;
  assign \new_[80735]_  = A267 & A266;
  assign \new_[80736]_  = \new_[80735]_  & \new_[80732]_ ;
  assign \new_[80739]_  = A300 & A268;
  assign \new_[80742]_  = ~A302 & ~A301;
  assign \new_[80743]_  = \new_[80742]_  & \new_[80739]_ ;
  assign \new_[80744]_  = \new_[80743]_  & \new_[80736]_ ;
  assign \new_[80748]_  = A167 & A168;
  assign \new_[80749]_  = A169 & \new_[80748]_ ;
  assign \new_[80752]_  = A199 & ~A166;
  assign \new_[80755]_  = A201 & ~A200;
  assign \new_[80756]_  = \new_[80755]_  & \new_[80752]_ ;
  assign \new_[80757]_  = \new_[80756]_  & \new_[80749]_ ;
  assign \new_[80760]_  = ~A265 & A203;
  assign \new_[80763]_  = A267 & A266;
  assign \new_[80764]_  = \new_[80763]_  & \new_[80760]_ ;
  assign \new_[80767]_  = A300 & A269;
  assign \new_[80770]_  = ~A302 & ~A301;
  assign \new_[80771]_  = \new_[80770]_  & \new_[80767]_ ;
  assign \new_[80772]_  = \new_[80771]_  & \new_[80764]_ ;
  assign \new_[80776]_  = A167 & A168;
  assign \new_[80777]_  = A169 & \new_[80776]_ ;
  assign \new_[80780]_  = A199 & ~A166;
  assign \new_[80783]_  = A201 & ~A200;
  assign \new_[80784]_  = \new_[80783]_  & \new_[80780]_ ;
  assign \new_[80785]_  = \new_[80784]_  & \new_[80777]_ ;
  assign \new_[80788]_  = ~A265 & A203;
  assign \new_[80791]_  = ~A267 & A266;
  assign \new_[80792]_  = \new_[80791]_  & \new_[80788]_ ;
  assign \new_[80795]_  = ~A269 & ~A268;
  assign \new_[80798]_  = A301 & ~A300;
  assign \new_[80799]_  = \new_[80798]_  & \new_[80795]_ ;
  assign \new_[80800]_  = \new_[80799]_  & \new_[80792]_ ;
  assign \new_[80804]_  = A167 & A168;
  assign \new_[80805]_  = A169 & \new_[80804]_ ;
  assign \new_[80808]_  = A199 & ~A166;
  assign \new_[80811]_  = A201 & ~A200;
  assign \new_[80812]_  = \new_[80811]_  & \new_[80808]_ ;
  assign \new_[80813]_  = \new_[80812]_  & \new_[80805]_ ;
  assign \new_[80816]_  = ~A265 & A203;
  assign \new_[80819]_  = ~A267 & A266;
  assign \new_[80820]_  = \new_[80819]_  & \new_[80816]_ ;
  assign \new_[80823]_  = ~A269 & ~A268;
  assign \new_[80826]_  = A302 & ~A300;
  assign \new_[80827]_  = \new_[80826]_  & \new_[80823]_ ;
  assign \new_[80828]_  = \new_[80827]_  & \new_[80820]_ ;
  assign \new_[80832]_  = A167 & A168;
  assign \new_[80833]_  = A169 & \new_[80832]_ ;
  assign \new_[80836]_  = A199 & ~A166;
  assign \new_[80839]_  = A201 & ~A200;
  assign \new_[80840]_  = \new_[80839]_  & \new_[80836]_ ;
  assign \new_[80841]_  = \new_[80840]_  & \new_[80833]_ ;
  assign \new_[80844]_  = ~A265 & A203;
  assign \new_[80847]_  = ~A267 & A266;
  assign \new_[80848]_  = \new_[80847]_  & \new_[80844]_ ;
  assign \new_[80851]_  = ~A269 & ~A268;
  assign \new_[80854]_  = A299 & A298;
  assign \new_[80855]_  = \new_[80854]_  & \new_[80851]_ ;
  assign \new_[80856]_  = \new_[80855]_  & \new_[80848]_ ;
  assign \new_[80860]_  = A167 & A168;
  assign \new_[80861]_  = A169 & \new_[80860]_ ;
  assign \new_[80864]_  = A199 & ~A166;
  assign \new_[80867]_  = A201 & ~A200;
  assign \new_[80868]_  = \new_[80867]_  & \new_[80864]_ ;
  assign \new_[80869]_  = \new_[80868]_  & \new_[80861]_ ;
  assign \new_[80872]_  = ~A265 & A203;
  assign \new_[80875]_  = ~A267 & A266;
  assign \new_[80876]_  = \new_[80875]_  & \new_[80872]_ ;
  assign \new_[80879]_  = ~A269 & ~A268;
  assign \new_[80882]_  = ~A299 & ~A298;
  assign \new_[80883]_  = \new_[80882]_  & \new_[80879]_ ;
  assign \new_[80884]_  = \new_[80883]_  & \new_[80876]_ ;
  assign \new_[80888]_  = A167 & A168;
  assign \new_[80889]_  = A169 & \new_[80888]_ ;
  assign \new_[80892]_  = A199 & ~A166;
  assign \new_[80895]_  = A201 & ~A200;
  assign \new_[80896]_  = \new_[80895]_  & \new_[80892]_ ;
  assign \new_[80897]_  = \new_[80896]_  & \new_[80889]_ ;
  assign \new_[80900]_  = A265 & A203;
  assign \new_[80903]_  = A267 & ~A266;
  assign \new_[80904]_  = \new_[80903]_  & \new_[80900]_ ;
  assign \new_[80907]_  = A300 & A268;
  assign \new_[80910]_  = ~A302 & ~A301;
  assign \new_[80911]_  = \new_[80910]_  & \new_[80907]_ ;
  assign \new_[80912]_  = \new_[80911]_  & \new_[80904]_ ;
  assign \new_[80916]_  = A167 & A168;
  assign \new_[80917]_  = A169 & \new_[80916]_ ;
  assign \new_[80920]_  = A199 & ~A166;
  assign \new_[80923]_  = A201 & ~A200;
  assign \new_[80924]_  = \new_[80923]_  & \new_[80920]_ ;
  assign \new_[80925]_  = \new_[80924]_  & \new_[80917]_ ;
  assign \new_[80928]_  = A265 & A203;
  assign \new_[80931]_  = A267 & ~A266;
  assign \new_[80932]_  = \new_[80931]_  & \new_[80928]_ ;
  assign \new_[80935]_  = A300 & A269;
  assign \new_[80938]_  = ~A302 & ~A301;
  assign \new_[80939]_  = \new_[80938]_  & \new_[80935]_ ;
  assign \new_[80940]_  = \new_[80939]_  & \new_[80932]_ ;
  assign \new_[80944]_  = A167 & A168;
  assign \new_[80945]_  = A169 & \new_[80944]_ ;
  assign \new_[80948]_  = A199 & ~A166;
  assign \new_[80951]_  = A201 & ~A200;
  assign \new_[80952]_  = \new_[80951]_  & \new_[80948]_ ;
  assign \new_[80953]_  = \new_[80952]_  & \new_[80945]_ ;
  assign \new_[80956]_  = A265 & A203;
  assign \new_[80959]_  = ~A267 & ~A266;
  assign \new_[80960]_  = \new_[80959]_  & \new_[80956]_ ;
  assign \new_[80963]_  = ~A269 & ~A268;
  assign \new_[80966]_  = A301 & ~A300;
  assign \new_[80967]_  = \new_[80966]_  & \new_[80963]_ ;
  assign \new_[80968]_  = \new_[80967]_  & \new_[80960]_ ;
  assign \new_[80972]_  = A167 & A168;
  assign \new_[80973]_  = A169 & \new_[80972]_ ;
  assign \new_[80976]_  = A199 & ~A166;
  assign \new_[80979]_  = A201 & ~A200;
  assign \new_[80980]_  = \new_[80979]_  & \new_[80976]_ ;
  assign \new_[80981]_  = \new_[80980]_  & \new_[80973]_ ;
  assign \new_[80984]_  = A265 & A203;
  assign \new_[80987]_  = ~A267 & ~A266;
  assign \new_[80988]_  = \new_[80987]_  & \new_[80984]_ ;
  assign \new_[80991]_  = ~A269 & ~A268;
  assign \new_[80994]_  = A302 & ~A300;
  assign \new_[80995]_  = \new_[80994]_  & \new_[80991]_ ;
  assign \new_[80996]_  = \new_[80995]_  & \new_[80988]_ ;
  assign \new_[81000]_  = A167 & A168;
  assign \new_[81001]_  = A169 & \new_[81000]_ ;
  assign \new_[81004]_  = A199 & ~A166;
  assign \new_[81007]_  = A201 & ~A200;
  assign \new_[81008]_  = \new_[81007]_  & \new_[81004]_ ;
  assign \new_[81009]_  = \new_[81008]_  & \new_[81001]_ ;
  assign \new_[81012]_  = A265 & A203;
  assign \new_[81015]_  = ~A267 & ~A266;
  assign \new_[81016]_  = \new_[81015]_  & \new_[81012]_ ;
  assign \new_[81019]_  = ~A269 & ~A268;
  assign \new_[81022]_  = A299 & A298;
  assign \new_[81023]_  = \new_[81022]_  & \new_[81019]_ ;
  assign \new_[81024]_  = \new_[81023]_  & \new_[81016]_ ;
  assign \new_[81028]_  = A167 & A168;
  assign \new_[81029]_  = A169 & \new_[81028]_ ;
  assign \new_[81032]_  = A199 & ~A166;
  assign \new_[81035]_  = A201 & ~A200;
  assign \new_[81036]_  = \new_[81035]_  & \new_[81032]_ ;
  assign \new_[81037]_  = \new_[81036]_  & \new_[81029]_ ;
  assign \new_[81040]_  = A265 & A203;
  assign \new_[81043]_  = ~A267 & ~A266;
  assign \new_[81044]_  = \new_[81043]_  & \new_[81040]_ ;
  assign \new_[81047]_  = ~A269 & ~A268;
  assign \new_[81050]_  = ~A299 & ~A298;
  assign \new_[81051]_  = \new_[81050]_  & \new_[81047]_ ;
  assign \new_[81052]_  = \new_[81051]_  & \new_[81044]_ ;
  assign \new_[81056]_  = A167 & A168;
  assign \new_[81057]_  = A169 & \new_[81056]_ ;
  assign \new_[81060]_  = A199 & ~A166;
  assign \new_[81063]_  = ~A201 & ~A200;
  assign \new_[81064]_  = \new_[81063]_  & \new_[81060]_ ;
  assign \new_[81065]_  = \new_[81064]_  & \new_[81057]_ ;
  assign \new_[81068]_  = ~A203 & ~A202;
  assign \new_[81071]_  = A266 & ~A265;
  assign \new_[81072]_  = \new_[81071]_  & \new_[81068]_ ;
  assign \new_[81075]_  = A268 & A267;
  assign \new_[81078]_  = A301 & ~A300;
  assign \new_[81079]_  = \new_[81078]_  & \new_[81075]_ ;
  assign \new_[81080]_  = \new_[81079]_  & \new_[81072]_ ;
  assign \new_[81084]_  = A167 & A168;
  assign \new_[81085]_  = A169 & \new_[81084]_ ;
  assign \new_[81088]_  = A199 & ~A166;
  assign \new_[81091]_  = ~A201 & ~A200;
  assign \new_[81092]_  = \new_[81091]_  & \new_[81088]_ ;
  assign \new_[81093]_  = \new_[81092]_  & \new_[81085]_ ;
  assign \new_[81096]_  = ~A203 & ~A202;
  assign \new_[81099]_  = A266 & ~A265;
  assign \new_[81100]_  = \new_[81099]_  & \new_[81096]_ ;
  assign \new_[81103]_  = A268 & A267;
  assign \new_[81106]_  = A302 & ~A300;
  assign \new_[81107]_  = \new_[81106]_  & \new_[81103]_ ;
  assign \new_[81108]_  = \new_[81107]_  & \new_[81100]_ ;
  assign \new_[81112]_  = A167 & A168;
  assign \new_[81113]_  = A169 & \new_[81112]_ ;
  assign \new_[81116]_  = A199 & ~A166;
  assign \new_[81119]_  = ~A201 & ~A200;
  assign \new_[81120]_  = \new_[81119]_  & \new_[81116]_ ;
  assign \new_[81121]_  = \new_[81120]_  & \new_[81113]_ ;
  assign \new_[81124]_  = ~A203 & ~A202;
  assign \new_[81127]_  = A266 & ~A265;
  assign \new_[81128]_  = \new_[81127]_  & \new_[81124]_ ;
  assign \new_[81131]_  = A268 & A267;
  assign \new_[81134]_  = A299 & A298;
  assign \new_[81135]_  = \new_[81134]_  & \new_[81131]_ ;
  assign \new_[81136]_  = \new_[81135]_  & \new_[81128]_ ;
  assign \new_[81140]_  = A167 & A168;
  assign \new_[81141]_  = A169 & \new_[81140]_ ;
  assign \new_[81144]_  = A199 & ~A166;
  assign \new_[81147]_  = ~A201 & ~A200;
  assign \new_[81148]_  = \new_[81147]_  & \new_[81144]_ ;
  assign \new_[81149]_  = \new_[81148]_  & \new_[81141]_ ;
  assign \new_[81152]_  = ~A203 & ~A202;
  assign \new_[81155]_  = A266 & ~A265;
  assign \new_[81156]_  = \new_[81155]_  & \new_[81152]_ ;
  assign \new_[81159]_  = A268 & A267;
  assign \new_[81162]_  = ~A299 & ~A298;
  assign \new_[81163]_  = \new_[81162]_  & \new_[81159]_ ;
  assign \new_[81164]_  = \new_[81163]_  & \new_[81156]_ ;
  assign \new_[81168]_  = A167 & A168;
  assign \new_[81169]_  = A169 & \new_[81168]_ ;
  assign \new_[81172]_  = A199 & ~A166;
  assign \new_[81175]_  = ~A201 & ~A200;
  assign \new_[81176]_  = \new_[81175]_  & \new_[81172]_ ;
  assign \new_[81177]_  = \new_[81176]_  & \new_[81169]_ ;
  assign \new_[81180]_  = ~A203 & ~A202;
  assign \new_[81183]_  = A266 & ~A265;
  assign \new_[81184]_  = \new_[81183]_  & \new_[81180]_ ;
  assign \new_[81187]_  = A269 & A267;
  assign \new_[81190]_  = A301 & ~A300;
  assign \new_[81191]_  = \new_[81190]_  & \new_[81187]_ ;
  assign \new_[81192]_  = \new_[81191]_  & \new_[81184]_ ;
  assign \new_[81196]_  = A167 & A168;
  assign \new_[81197]_  = A169 & \new_[81196]_ ;
  assign \new_[81200]_  = A199 & ~A166;
  assign \new_[81203]_  = ~A201 & ~A200;
  assign \new_[81204]_  = \new_[81203]_  & \new_[81200]_ ;
  assign \new_[81205]_  = \new_[81204]_  & \new_[81197]_ ;
  assign \new_[81208]_  = ~A203 & ~A202;
  assign \new_[81211]_  = A266 & ~A265;
  assign \new_[81212]_  = \new_[81211]_  & \new_[81208]_ ;
  assign \new_[81215]_  = A269 & A267;
  assign \new_[81218]_  = A302 & ~A300;
  assign \new_[81219]_  = \new_[81218]_  & \new_[81215]_ ;
  assign \new_[81220]_  = \new_[81219]_  & \new_[81212]_ ;
  assign \new_[81224]_  = A167 & A168;
  assign \new_[81225]_  = A169 & \new_[81224]_ ;
  assign \new_[81228]_  = A199 & ~A166;
  assign \new_[81231]_  = ~A201 & ~A200;
  assign \new_[81232]_  = \new_[81231]_  & \new_[81228]_ ;
  assign \new_[81233]_  = \new_[81232]_  & \new_[81225]_ ;
  assign \new_[81236]_  = ~A203 & ~A202;
  assign \new_[81239]_  = A266 & ~A265;
  assign \new_[81240]_  = \new_[81239]_  & \new_[81236]_ ;
  assign \new_[81243]_  = A269 & A267;
  assign \new_[81246]_  = A299 & A298;
  assign \new_[81247]_  = \new_[81246]_  & \new_[81243]_ ;
  assign \new_[81248]_  = \new_[81247]_  & \new_[81240]_ ;
  assign \new_[81252]_  = A167 & A168;
  assign \new_[81253]_  = A169 & \new_[81252]_ ;
  assign \new_[81256]_  = A199 & ~A166;
  assign \new_[81259]_  = ~A201 & ~A200;
  assign \new_[81260]_  = \new_[81259]_  & \new_[81256]_ ;
  assign \new_[81261]_  = \new_[81260]_  & \new_[81253]_ ;
  assign \new_[81264]_  = ~A203 & ~A202;
  assign \new_[81267]_  = A266 & ~A265;
  assign \new_[81268]_  = \new_[81267]_  & \new_[81264]_ ;
  assign \new_[81271]_  = A269 & A267;
  assign \new_[81274]_  = ~A299 & ~A298;
  assign \new_[81275]_  = \new_[81274]_  & \new_[81271]_ ;
  assign \new_[81276]_  = \new_[81275]_  & \new_[81268]_ ;
  assign \new_[81280]_  = A167 & A168;
  assign \new_[81281]_  = A169 & \new_[81280]_ ;
  assign \new_[81284]_  = A199 & ~A166;
  assign \new_[81287]_  = ~A201 & ~A200;
  assign \new_[81288]_  = \new_[81287]_  & \new_[81284]_ ;
  assign \new_[81289]_  = \new_[81288]_  & \new_[81281]_ ;
  assign \new_[81292]_  = ~A203 & ~A202;
  assign \new_[81295]_  = ~A266 & A265;
  assign \new_[81296]_  = \new_[81295]_  & \new_[81292]_ ;
  assign \new_[81299]_  = A268 & A267;
  assign \new_[81302]_  = A301 & ~A300;
  assign \new_[81303]_  = \new_[81302]_  & \new_[81299]_ ;
  assign \new_[81304]_  = \new_[81303]_  & \new_[81296]_ ;
  assign \new_[81308]_  = A167 & A168;
  assign \new_[81309]_  = A169 & \new_[81308]_ ;
  assign \new_[81312]_  = A199 & ~A166;
  assign \new_[81315]_  = ~A201 & ~A200;
  assign \new_[81316]_  = \new_[81315]_  & \new_[81312]_ ;
  assign \new_[81317]_  = \new_[81316]_  & \new_[81309]_ ;
  assign \new_[81320]_  = ~A203 & ~A202;
  assign \new_[81323]_  = ~A266 & A265;
  assign \new_[81324]_  = \new_[81323]_  & \new_[81320]_ ;
  assign \new_[81327]_  = A268 & A267;
  assign \new_[81330]_  = A302 & ~A300;
  assign \new_[81331]_  = \new_[81330]_  & \new_[81327]_ ;
  assign \new_[81332]_  = \new_[81331]_  & \new_[81324]_ ;
  assign \new_[81336]_  = A167 & A168;
  assign \new_[81337]_  = A169 & \new_[81336]_ ;
  assign \new_[81340]_  = A199 & ~A166;
  assign \new_[81343]_  = ~A201 & ~A200;
  assign \new_[81344]_  = \new_[81343]_  & \new_[81340]_ ;
  assign \new_[81345]_  = \new_[81344]_  & \new_[81337]_ ;
  assign \new_[81348]_  = ~A203 & ~A202;
  assign \new_[81351]_  = ~A266 & A265;
  assign \new_[81352]_  = \new_[81351]_  & \new_[81348]_ ;
  assign \new_[81355]_  = A268 & A267;
  assign \new_[81358]_  = A299 & A298;
  assign \new_[81359]_  = \new_[81358]_  & \new_[81355]_ ;
  assign \new_[81360]_  = \new_[81359]_  & \new_[81352]_ ;
  assign \new_[81364]_  = A167 & A168;
  assign \new_[81365]_  = A169 & \new_[81364]_ ;
  assign \new_[81368]_  = A199 & ~A166;
  assign \new_[81371]_  = ~A201 & ~A200;
  assign \new_[81372]_  = \new_[81371]_  & \new_[81368]_ ;
  assign \new_[81373]_  = \new_[81372]_  & \new_[81365]_ ;
  assign \new_[81376]_  = ~A203 & ~A202;
  assign \new_[81379]_  = ~A266 & A265;
  assign \new_[81380]_  = \new_[81379]_  & \new_[81376]_ ;
  assign \new_[81383]_  = A268 & A267;
  assign \new_[81386]_  = ~A299 & ~A298;
  assign \new_[81387]_  = \new_[81386]_  & \new_[81383]_ ;
  assign \new_[81388]_  = \new_[81387]_  & \new_[81380]_ ;
  assign \new_[81392]_  = A167 & A168;
  assign \new_[81393]_  = A169 & \new_[81392]_ ;
  assign \new_[81396]_  = A199 & ~A166;
  assign \new_[81399]_  = ~A201 & ~A200;
  assign \new_[81400]_  = \new_[81399]_  & \new_[81396]_ ;
  assign \new_[81401]_  = \new_[81400]_  & \new_[81393]_ ;
  assign \new_[81404]_  = ~A203 & ~A202;
  assign \new_[81407]_  = ~A266 & A265;
  assign \new_[81408]_  = \new_[81407]_  & \new_[81404]_ ;
  assign \new_[81411]_  = A269 & A267;
  assign \new_[81414]_  = A301 & ~A300;
  assign \new_[81415]_  = \new_[81414]_  & \new_[81411]_ ;
  assign \new_[81416]_  = \new_[81415]_  & \new_[81408]_ ;
  assign \new_[81420]_  = A167 & A168;
  assign \new_[81421]_  = A169 & \new_[81420]_ ;
  assign \new_[81424]_  = A199 & ~A166;
  assign \new_[81427]_  = ~A201 & ~A200;
  assign \new_[81428]_  = \new_[81427]_  & \new_[81424]_ ;
  assign \new_[81429]_  = \new_[81428]_  & \new_[81421]_ ;
  assign \new_[81432]_  = ~A203 & ~A202;
  assign \new_[81435]_  = ~A266 & A265;
  assign \new_[81436]_  = \new_[81435]_  & \new_[81432]_ ;
  assign \new_[81439]_  = A269 & A267;
  assign \new_[81442]_  = A302 & ~A300;
  assign \new_[81443]_  = \new_[81442]_  & \new_[81439]_ ;
  assign \new_[81444]_  = \new_[81443]_  & \new_[81436]_ ;
  assign \new_[81448]_  = A167 & A168;
  assign \new_[81449]_  = A169 & \new_[81448]_ ;
  assign \new_[81452]_  = A199 & ~A166;
  assign \new_[81455]_  = ~A201 & ~A200;
  assign \new_[81456]_  = \new_[81455]_  & \new_[81452]_ ;
  assign \new_[81457]_  = \new_[81456]_  & \new_[81449]_ ;
  assign \new_[81460]_  = ~A203 & ~A202;
  assign \new_[81463]_  = ~A266 & A265;
  assign \new_[81464]_  = \new_[81463]_  & \new_[81460]_ ;
  assign \new_[81467]_  = A269 & A267;
  assign \new_[81470]_  = A299 & A298;
  assign \new_[81471]_  = \new_[81470]_  & \new_[81467]_ ;
  assign \new_[81472]_  = \new_[81471]_  & \new_[81464]_ ;
  assign \new_[81476]_  = A167 & A168;
  assign \new_[81477]_  = A169 & \new_[81476]_ ;
  assign \new_[81480]_  = A199 & ~A166;
  assign \new_[81483]_  = ~A201 & ~A200;
  assign \new_[81484]_  = \new_[81483]_  & \new_[81480]_ ;
  assign \new_[81485]_  = \new_[81484]_  & \new_[81477]_ ;
  assign \new_[81488]_  = ~A203 & ~A202;
  assign \new_[81491]_  = ~A266 & A265;
  assign \new_[81492]_  = \new_[81491]_  & \new_[81488]_ ;
  assign \new_[81495]_  = A269 & A267;
  assign \new_[81498]_  = ~A299 & ~A298;
  assign \new_[81499]_  = \new_[81498]_  & \new_[81495]_ ;
  assign \new_[81500]_  = \new_[81499]_  & \new_[81492]_ ;
  assign \new_[81504]_  = ~A167 & A168;
  assign \new_[81505]_  = A169 & \new_[81504]_ ;
  assign \new_[81508]_  = A201 & A166;
  assign \new_[81511]_  = ~A203 & ~A202;
  assign \new_[81512]_  = \new_[81511]_  & \new_[81508]_ ;
  assign \new_[81513]_  = \new_[81512]_  & \new_[81505]_ ;
  assign \new_[81516]_  = ~A268 & A267;
  assign \new_[81519]_  = A298 & ~A269;
  assign \new_[81520]_  = \new_[81519]_  & \new_[81516]_ ;
  assign \new_[81523]_  = ~A300 & ~A299;
  assign \new_[81526]_  = ~A302 & ~A301;
  assign \new_[81527]_  = \new_[81526]_  & \new_[81523]_ ;
  assign \new_[81528]_  = \new_[81527]_  & \new_[81520]_ ;
  assign \new_[81532]_  = ~A167 & A168;
  assign \new_[81533]_  = A169 & \new_[81532]_ ;
  assign \new_[81536]_  = A201 & A166;
  assign \new_[81539]_  = ~A203 & ~A202;
  assign \new_[81540]_  = \new_[81539]_  & \new_[81536]_ ;
  assign \new_[81541]_  = \new_[81540]_  & \new_[81533]_ ;
  assign \new_[81544]_  = ~A268 & A267;
  assign \new_[81547]_  = ~A298 & ~A269;
  assign \new_[81548]_  = \new_[81547]_  & \new_[81544]_ ;
  assign \new_[81551]_  = ~A300 & A299;
  assign \new_[81554]_  = ~A302 & ~A301;
  assign \new_[81555]_  = \new_[81554]_  & \new_[81551]_ ;
  assign \new_[81556]_  = \new_[81555]_  & \new_[81548]_ ;
  assign \new_[81560]_  = ~A167 & A168;
  assign \new_[81561]_  = A169 & \new_[81560]_ ;
  assign \new_[81564]_  = ~A199 & A166;
  assign \new_[81567]_  = A201 & A200;
  assign \new_[81568]_  = \new_[81567]_  & \new_[81564]_ ;
  assign \new_[81569]_  = \new_[81568]_  & \new_[81561]_ ;
  assign \new_[81572]_  = ~A265 & A202;
  assign \new_[81575]_  = A267 & A266;
  assign \new_[81576]_  = \new_[81575]_  & \new_[81572]_ ;
  assign \new_[81579]_  = A300 & A268;
  assign \new_[81582]_  = ~A302 & ~A301;
  assign \new_[81583]_  = \new_[81582]_  & \new_[81579]_ ;
  assign \new_[81584]_  = \new_[81583]_  & \new_[81576]_ ;
  assign \new_[81588]_  = ~A167 & A168;
  assign \new_[81589]_  = A169 & \new_[81588]_ ;
  assign \new_[81592]_  = ~A199 & A166;
  assign \new_[81595]_  = A201 & A200;
  assign \new_[81596]_  = \new_[81595]_  & \new_[81592]_ ;
  assign \new_[81597]_  = \new_[81596]_  & \new_[81589]_ ;
  assign \new_[81600]_  = ~A265 & A202;
  assign \new_[81603]_  = A267 & A266;
  assign \new_[81604]_  = \new_[81603]_  & \new_[81600]_ ;
  assign \new_[81607]_  = A300 & A269;
  assign \new_[81610]_  = ~A302 & ~A301;
  assign \new_[81611]_  = \new_[81610]_  & \new_[81607]_ ;
  assign \new_[81612]_  = \new_[81611]_  & \new_[81604]_ ;
  assign \new_[81616]_  = ~A167 & A168;
  assign \new_[81617]_  = A169 & \new_[81616]_ ;
  assign \new_[81620]_  = ~A199 & A166;
  assign \new_[81623]_  = A201 & A200;
  assign \new_[81624]_  = \new_[81623]_  & \new_[81620]_ ;
  assign \new_[81625]_  = \new_[81624]_  & \new_[81617]_ ;
  assign \new_[81628]_  = ~A265 & A202;
  assign \new_[81631]_  = ~A267 & A266;
  assign \new_[81632]_  = \new_[81631]_  & \new_[81628]_ ;
  assign \new_[81635]_  = ~A269 & ~A268;
  assign \new_[81638]_  = A301 & ~A300;
  assign \new_[81639]_  = \new_[81638]_  & \new_[81635]_ ;
  assign \new_[81640]_  = \new_[81639]_  & \new_[81632]_ ;
  assign \new_[81644]_  = ~A167 & A168;
  assign \new_[81645]_  = A169 & \new_[81644]_ ;
  assign \new_[81648]_  = ~A199 & A166;
  assign \new_[81651]_  = A201 & A200;
  assign \new_[81652]_  = \new_[81651]_  & \new_[81648]_ ;
  assign \new_[81653]_  = \new_[81652]_  & \new_[81645]_ ;
  assign \new_[81656]_  = ~A265 & A202;
  assign \new_[81659]_  = ~A267 & A266;
  assign \new_[81660]_  = \new_[81659]_  & \new_[81656]_ ;
  assign \new_[81663]_  = ~A269 & ~A268;
  assign \new_[81666]_  = A302 & ~A300;
  assign \new_[81667]_  = \new_[81666]_  & \new_[81663]_ ;
  assign \new_[81668]_  = \new_[81667]_  & \new_[81660]_ ;
  assign \new_[81672]_  = ~A167 & A168;
  assign \new_[81673]_  = A169 & \new_[81672]_ ;
  assign \new_[81676]_  = ~A199 & A166;
  assign \new_[81679]_  = A201 & A200;
  assign \new_[81680]_  = \new_[81679]_  & \new_[81676]_ ;
  assign \new_[81681]_  = \new_[81680]_  & \new_[81673]_ ;
  assign \new_[81684]_  = ~A265 & A202;
  assign \new_[81687]_  = ~A267 & A266;
  assign \new_[81688]_  = \new_[81687]_  & \new_[81684]_ ;
  assign \new_[81691]_  = ~A269 & ~A268;
  assign \new_[81694]_  = A299 & A298;
  assign \new_[81695]_  = \new_[81694]_  & \new_[81691]_ ;
  assign \new_[81696]_  = \new_[81695]_  & \new_[81688]_ ;
  assign \new_[81700]_  = ~A167 & A168;
  assign \new_[81701]_  = A169 & \new_[81700]_ ;
  assign \new_[81704]_  = ~A199 & A166;
  assign \new_[81707]_  = A201 & A200;
  assign \new_[81708]_  = \new_[81707]_  & \new_[81704]_ ;
  assign \new_[81709]_  = \new_[81708]_  & \new_[81701]_ ;
  assign \new_[81712]_  = ~A265 & A202;
  assign \new_[81715]_  = ~A267 & A266;
  assign \new_[81716]_  = \new_[81715]_  & \new_[81712]_ ;
  assign \new_[81719]_  = ~A269 & ~A268;
  assign \new_[81722]_  = ~A299 & ~A298;
  assign \new_[81723]_  = \new_[81722]_  & \new_[81719]_ ;
  assign \new_[81724]_  = \new_[81723]_  & \new_[81716]_ ;
  assign \new_[81728]_  = ~A167 & A168;
  assign \new_[81729]_  = A169 & \new_[81728]_ ;
  assign \new_[81732]_  = ~A199 & A166;
  assign \new_[81735]_  = A201 & A200;
  assign \new_[81736]_  = \new_[81735]_  & \new_[81732]_ ;
  assign \new_[81737]_  = \new_[81736]_  & \new_[81729]_ ;
  assign \new_[81740]_  = A265 & A202;
  assign \new_[81743]_  = A267 & ~A266;
  assign \new_[81744]_  = \new_[81743]_  & \new_[81740]_ ;
  assign \new_[81747]_  = A300 & A268;
  assign \new_[81750]_  = ~A302 & ~A301;
  assign \new_[81751]_  = \new_[81750]_  & \new_[81747]_ ;
  assign \new_[81752]_  = \new_[81751]_  & \new_[81744]_ ;
  assign \new_[81756]_  = ~A167 & A168;
  assign \new_[81757]_  = A169 & \new_[81756]_ ;
  assign \new_[81760]_  = ~A199 & A166;
  assign \new_[81763]_  = A201 & A200;
  assign \new_[81764]_  = \new_[81763]_  & \new_[81760]_ ;
  assign \new_[81765]_  = \new_[81764]_  & \new_[81757]_ ;
  assign \new_[81768]_  = A265 & A202;
  assign \new_[81771]_  = A267 & ~A266;
  assign \new_[81772]_  = \new_[81771]_  & \new_[81768]_ ;
  assign \new_[81775]_  = A300 & A269;
  assign \new_[81778]_  = ~A302 & ~A301;
  assign \new_[81779]_  = \new_[81778]_  & \new_[81775]_ ;
  assign \new_[81780]_  = \new_[81779]_  & \new_[81772]_ ;
  assign \new_[81784]_  = ~A167 & A168;
  assign \new_[81785]_  = A169 & \new_[81784]_ ;
  assign \new_[81788]_  = ~A199 & A166;
  assign \new_[81791]_  = A201 & A200;
  assign \new_[81792]_  = \new_[81791]_  & \new_[81788]_ ;
  assign \new_[81793]_  = \new_[81792]_  & \new_[81785]_ ;
  assign \new_[81796]_  = A265 & A202;
  assign \new_[81799]_  = ~A267 & ~A266;
  assign \new_[81800]_  = \new_[81799]_  & \new_[81796]_ ;
  assign \new_[81803]_  = ~A269 & ~A268;
  assign \new_[81806]_  = A301 & ~A300;
  assign \new_[81807]_  = \new_[81806]_  & \new_[81803]_ ;
  assign \new_[81808]_  = \new_[81807]_  & \new_[81800]_ ;
  assign \new_[81812]_  = ~A167 & A168;
  assign \new_[81813]_  = A169 & \new_[81812]_ ;
  assign \new_[81816]_  = ~A199 & A166;
  assign \new_[81819]_  = A201 & A200;
  assign \new_[81820]_  = \new_[81819]_  & \new_[81816]_ ;
  assign \new_[81821]_  = \new_[81820]_  & \new_[81813]_ ;
  assign \new_[81824]_  = A265 & A202;
  assign \new_[81827]_  = ~A267 & ~A266;
  assign \new_[81828]_  = \new_[81827]_  & \new_[81824]_ ;
  assign \new_[81831]_  = ~A269 & ~A268;
  assign \new_[81834]_  = A302 & ~A300;
  assign \new_[81835]_  = \new_[81834]_  & \new_[81831]_ ;
  assign \new_[81836]_  = \new_[81835]_  & \new_[81828]_ ;
  assign \new_[81840]_  = ~A167 & A168;
  assign \new_[81841]_  = A169 & \new_[81840]_ ;
  assign \new_[81844]_  = ~A199 & A166;
  assign \new_[81847]_  = A201 & A200;
  assign \new_[81848]_  = \new_[81847]_  & \new_[81844]_ ;
  assign \new_[81849]_  = \new_[81848]_  & \new_[81841]_ ;
  assign \new_[81852]_  = A265 & A202;
  assign \new_[81855]_  = ~A267 & ~A266;
  assign \new_[81856]_  = \new_[81855]_  & \new_[81852]_ ;
  assign \new_[81859]_  = ~A269 & ~A268;
  assign \new_[81862]_  = A299 & A298;
  assign \new_[81863]_  = \new_[81862]_  & \new_[81859]_ ;
  assign \new_[81864]_  = \new_[81863]_  & \new_[81856]_ ;
  assign \new_[81868]_  = ~A167 & A168;
  assign \new_[81869]_  = A169 & \new_[81868]_ ;
  assign \new_[81872]_  = ~A199 & A166;
  assign \new_[81875]_  = A201 & A200;
  assign \new_[81876]_  = \new_[81875]_  & \new_[81872]_ ;
  assign \new_[81877]_  = \new_[81876]_  & \new_[81869]_ ;
  assign \new_[81880]_  = A265 & A202;
  assign \new_[81883]_  = ~A267 & ~A266;
  assign \new_[81884]_  = \new_[81883]_  & \new_[81880]_ ;
  assign \new_[81887]_  = ~A269 & ~A268;
  assign \new_[81890]_  = ~A299 & ~A298;
  assign \new_[81891]_  = \new_[81890]_  & \new_[81887]_ ;
  assign \new_[81892]_  = \new_[81891]_  & \new_[81884]_ ;
  assign \new_[81896]_  = ~A167 & A168;
  assign \new_[81897]_  = A169 & \new_[81896]_ ;
  assign \new_[81900]_  = ~A199 & A166;
  assign \new_[81903]_  = A201 & A200;
  assign \new_[81904]_  = \new_[81903]_  & \new_[81900]_ ;
  assign \new_[81905]_  = \new_[81904]_  & \new_[81897]_ ;
  assign \new_[81908]_  = ~A265 & A203;
  assign \new_[81911]_  = A267 & A266;
  assign \new_[81912]_  = \new_[81911]_  & \new_[81908]_ ;
  assign \new_[81915]_  = A300 & A268;
  assign \new_[81918]_  = ~A302 & ~A301;
  assign \new_[81919]_  = \new_[81918]_  & \new_[81915]_ ;
  assign \new_[81920]_  = \new_[81919]_  & \new_[81912]_ ;
  assign \new_[81924]_  = ~A167 & A168;
  assign \new_[81925]_  = A169 & \new_[81924]_ ;
  assign \new_[81928]_  = ~A199 & A166;
  assign \new_[81931]_  = A201 & A200;
  assign \new_[81932]_  = \new_[81931]_  & \new_[81928]_ ;
  assign \new_[81933]_  = \new_[81932]_  & \new_[81925]_ ;
  assign \new_[81936]_  = ~A265 & A203;
  assign \new_[81939]_  = A267 & A266;
  assign \new_[81940]_  = \new_[81939]_  & \new_[81936]_ ;
  assign \new_[81943]_  = A300 & A269;
  assign \new_[81946]_  = ~A302 & ~A301;
  assign \new_[81947]_  = \new_[81946]_  & \new_[81943]_ ;
  assign \new_[81948]_  = \new_[81947]_  & \new_[81940]_ ;
  assign \new_[81952]_  = ~A167 & A168;
  assign \new_[81953]_  = A169 & \new_[81952]_ ;
  assign \new_[81956]_  = ~A199 & A166;
  assign \new_[81959]_  = A201 & A200;
  assign \new_[81960]_  = \new_[81959]_  & \new_[81956]_ ;
  assign \new_[81961]_  = \new_[81960]_  & \new_[81953]_ ;
  assign \new_[81964]_  = ~A265 & A203;
  assign \new_[81967]_  = ~A267 & A266;
  assign \new_[81968]_  = \new_[81967]_  & \new_[81964]_ ;
  assign \new_[81971]_  = ~A269 & ~A268;
  assign \new_[81974]_  = A301 & ~A300;
  assign \new_[81975]_  = \new_[81974]_  & \new_[81971]_ ;
  assign \new_[81976]_  = \new_[81975]_  & \new_[81968]_ ;
  assign \new_[81980]_  = ~A167 & A168;
  assign \new_[81981]_  = A169 & \new_[81980]_ ;
  assign \new_[81984]_  = ~A199 & A166;
  assign \new_[81987]_  = A201 & A200;
  assign \new_[81988]_  = \new_[81987]_  & \new_[81984]_ ;
  assign \new_[81989]_  = \new_[81988]_  & \new_[81981]_ ;
  assign \new_[81992]_  = ~A265 & A203;
  assign \new_[81995]_  = ~A267 & A266;
  assign \new_[81996]_  = \new_[81995]_  & \new_[81992]_ ;
  assign \new_[81999]_  = ~A269 & ~A268;
  assign \new_[82002]_  = A302 & ~A300;
  assign \new_[82003]_  = \new_[82002]_  & \new_[81999]_ ;
  assign \new_[82004]_  = \new_[82003]_  & \new_[81996]_ ;
  assign \new_[82008]_  = ~A167 & A168;
  assign \new_[82009]_  = A169 & \new_[82008]_ ;
  assign \new_[82012]_  = ~A199 & A166;
  assign \new_[82015]_  = A201 & A200;
  assign \new_[82016]_  = \new_[82015]_  & \new_[82012]_ ;
  assign \new_[82017]_  = \new_[82016]_  & \new_[82009]_ ;
  assign \new_[82020]_  = ~A265 & A203;
  assign \new_[82023]_  = ~A267 & A266;
  assign \new_[82024]_  = \new_[82023]_  & \new_[82020]_ ;
  assign \new_[82027]_  = ~A269 & ~A268;
  assign \new_[82030]_  = A299 & A298;
  assign \new_[82031]_  = \new_[82030]_  & \new_[82027]_ ;
  assign \new_[82032]_  = \new_[82031]_  & \new_[82024]_ ;
  assign \new_[82036]_  = ~A167 & A168;
  assign \new_[82037]_  = A169 & \new_[82036]_ ;
  assign \new_[82040]_  = ~A199 & A166;
  assign \new_[82043]_  = A201 & A200;
  assign \new_[82044]_  = \new_[82043]_  & \new_[82040]_ ;
  assign \new_[82045]_  = \new_[82044]_  & \new_[82037]_ ;
  assign \new_[82048]_  = ~A265 & A203;
  assign \new_[82051]_  = ~A267 & A266;
  assign \new_[82052]_  = \new_[82051]_  & \new_[82048]_ ;
  assign \new_[82055]_  = ~A269 & ~A268;
  assign \new_[82058]_  = ~A299 & ~A298;
  assign \new_[82059]_  = \new_[82058]_  & \new_[82055]_ ;
  assign \new_[82060]_  = \new_[82059]_  & \new_[82052]_ ;
  assign \new_[82064]_  = ~A167 & A168;
  assign \new_[82065]_  = A169 & \new_[82064]_ ;
  assign \new_[82068]_  = ~A199 & A166;
  assign \new_[82071]_  = A201 & A200;
  assign \new_[82072]_  = \new_[82071]_  & \new_[82068]_ ;
  assign \new_[82073]_  = \new_[82072]_  & \new_[82065]_ ;
  assign \new_[82076]_  = A265 & A203;
  assign \new_[82079]_  = A267 & ~A266;
  assign \new_[82080]_  = \new_[82079]_  & \new_[82076]_ ;
  assign \new_[82083]_  = A300 & A268;
  assign \new_[82086]_  = ~A302 & ~A301;
  assign \new_[82087]_  = \new_[82086]_  & \new_[82083]_ ;
  assign \new_[82088]_  = \new_[82087]_  & \new_[82080]_ ;
  assign \new_[82092]_  = ~A167 & A168;
  assign \new_[82093]_  = A169 & \new_[82092]_ ;
  assign \new_[82096]_  = ~A199 & A166;
  assign \new_[82099]_  = A201 & A200;
  assign \new_[82100]_  = \new_[82099]_  & \new_[82096]_ ;
  assign \new_[82101]_  = \new_[82100]_  & \new_[82093]_ ;
  assign \new_[82104]_  = A265 & A203;
  assign \new_[82107]_  = A267 & ~A266;
  assign \new_[82108]_  = \new_[82107]_  & \new_[82104]_ ;
  assign \new_[82111]_  = A300 & A269;
  assign \new_[82114]_  = ~A302 & ~A301;
  assign \new_[82115]_  = \new_[82114]_  & \new_[82111]_ ;
  assign \new_[82116]_  = \new_[82115]_  & \new_[82108]_ ;
  assign \new_[82120]_  = ~A167 & A168;
  assign \new_[82121]_  = A169 & \new_[82120]_ ;
  assign \new_[82124]_  = ~A199 & A166;
  assign \new_[82127]_  = A201 & A200;
  assign \new_[82128]_  = \new_[82127]_  & \new_[82124]_ ;
  assign \new_[82129]_  = \new_[82128]_  & \new_[82121]_ ;
  assign \new_[82132]_  = A265 & A203;
  assign \new_[82135]_  = ~A267 & ~A266;
  assign \new_[82136]_  = \new_[82135]_  & \new_[82132]_ ;
  assign \new_[82139]_  = ~A269 & ~A268;
  assign \new_[82142]_  = A301 & ~A300;
  assign \new_[82143]_  = \new_[82142]_  & \new_[82139]_ ;
  assign \new_[82144]_  = \new_[82143]_  & \new_[82136]_ ;
  assign \new_[82148]_  = ~A167 & A168;
  assign \new_[82149]_  = A169 & \new_[82148]_ ;
  assign \new_[82152]_  = ~A199 & A166;
  assign \new_[82155]_  = A201 & A200;
  assign \new_[82156]_  = \new_[82155]_  & \new_[82152]_ ;
  assign \new_[82157]_  = \new_[82156]_  & \new_[82149]_ ;
  assign \new_[82160]_  = A265 & A203;
  assign \new_[82163]_  = ~A267 & ~A266;
  assign \new_[82164]_  = \new_[82163]_  & \new_[82160]_ ;
  assign \new_[82167]_  = ~A269 & ~A268;
  assign \new_[82170]_  = A302 & ~A300;
  assign \new_[82171]_  = \new_[82170]_  & \new_[82167]_ ;
  assign \new_[82172]_  = \new_[82171]_  & \new_[82164]_ ;
  assign \new_[82176]_  = ~A167 & A168;
  assign \new_[82177]_  = A169 & \new_[82176]_ ;
  assign \new_[82180]_  = ~A199 & A166;
  assign \new_[82183]_  = A201 & A200;
  assign \new_[82184]_  = \new_[82183]_  & \new_[82180]_ ;
  assign \new_[82185]_  = \new_[82184]_  & \new_[82177]_ ;
  assign \new_[82188]_  = A265 & A203;
  assign \new_[82191]_  = ~A267 & ~A266;
  assign \new_[82192]_  = \new_[82191]_  & \new_[82188]_ ;
  assign \new_[82195]_  = ~A269 & ~A268;
  assign \new_[82198]_  = A299 & A298;
  assign \new_[82199]_  = \new_[82198]_  & \new_[82195]_ ;
  assign \new_[82200]_  = \new_[82199]_  & \new_[82192]_ ;
  assign \new_[82204]_  = ~A167 & A168;
  assign \new_[82205]_  = A169 & \new_[82204]_ ;
  assign \new_[82208]_  = ~A199 & A166;
  assign \new_[82211]_  = A201 & A200;
  assign \new_[82212]_  = \new_[82211]_  & \new_[82208]_ ;
  assign \new_[82213]_  = \new_[82212]_  & \new_[82205]_ ;
  assign \new_[82216]_  = A265 & A203;
  assign \new_[82219]_  = ~A267 & ~A266;
  assign \new_[82220]_  = \new_[82219]_  & \new_[82216]_ ;
  assign \new_[82223]_  = ~A269 & ~A268;
  assign \new_[82226]_  = ~A299 & ~A298;
  assign \new_[82227]_  = \new_[82226]_  & \new_[82223]_ ;
  assign \new_[82228]_  = \new_[82227]_  & \new_[82220]_ ;
  assign \new_[82232]_  = ~A167 & A168;
  assign \new_[82233]_  = A169 & \new_[82232]_ ;
  assign \new_[82236]_  = ~A199 & A166;
  assign \new_[82239]_  = ~A201 & A200;
  assign \new_[82240]_  = \new_[82239]_  & \new_[82236]_ ;
  assign \new_[82241]_  = \new_[82240]_  & \new_[82233]_ ;
  assign \new_[82244]_  = ~A203 & ~A202;
  assign \new_[82247]_  = A266 & ~A265;
  assign \new_[82248]_  = \new_[82247]_  & \new_[82244]_ ;
  assign \new_[82251]_  = A268 & A267;
  assign \new_[82254]_  = A301 & ~A300;
  assign \new_[82255]_  = \new_[82254]_  & \new_[82251]_ ;
  assign \new_[82256]_  = \new_[82255]_  & \new_[82248]_ ;
  assign \new_[82260]_  = ~A167 & A168;
  assign \new_[82261]_  = A169 & \new_[82260]_ ;
  assign \new_[82264]_  = ~A199 & A166;
  assign \new_[82267]_  = ~A201 & A200;
  assign \new_[82268]_  = \new_[82267]_  & \new_[82264]_ ;
  assign \new_[82269]_  = \new_[82268]_  & \new_[82261]_ ;
  assign \new_[82272]_  = ~A203 & ~A202;
  assign \new_[82275]_  = A266 & ~A265;
  assign \new_[82276]_  = \new_[82275]_  & \new_[82272]_ ;
  assign \new_[82279]_  = A268 & A267;
  assign \new_[82282]_  = A302 & ~A300;
  assign \new_[82283]_  = \new_[82282]_  & \new_[82279]_ ;
  assign \new_[82284]_  = \new_[82283]_  & \new_[82276]_ ;
  assign \new_[82288]_  = ~A167 & A168;
  assign \new_[82289]_  = A169 & \new_[82288]_ ;
  assign \new_[82292]_  = ~A199 & A166;
  assign \new_[82295]_  = ~A201 & A200;
  assign \new_[82296]_  = \new_[82295]_  & \new_[82292]_ ;
  assign \new_[82297]_  = \new_[82296]_  & \new_[82289]_ ;
  assign \new_[82300]_  = ~A203 & ~A202;
  assign \new_[82303]_  = A266 & ~A265;
  assign \new_[82304]_  = \new_[82303]_  & \new_[82300]_ ;
  assign \new_[82307]_  = A268 & A267;
  assign \new_[82310]_  = A299 & A298;
  assign \new_[82311]_  = \new_[82310]_  & \new_[82307]_ ;
  assign \new_[82312]_  = \new_[82311]_  & \new_[82304]_ ;
  assign \new_[82316]_  = ~A167 & A168;
  assign \new_[82317]_  = A169 & \new_[82316]_ ;
  assign \new_[82320]_  = ~A199 & A166;
  assign \new_[82323]_  = ~A201 & A200;
  assign \new_[82324]_  = \new_[82323]_  & \new_[82320]_ ;
  assign \new_[82325]_  = \new_[82324]_  & \new_[82317]_ ;
  assign \new_[82328]_  = ~A203 & ~A202;
  assign \new_[82331]_  = A266 & ~A265;
  assign \new_[82332]_  = \new_[82331]_  & \new_[82328]_ ;
  assign \new_[82335]_  = A268 & A267;
  assign \new_[82338]_  = ~A299 & ~A298;
  assign \new_[82339]_  = \new_[82338]_  & \new_[82335]_ ;
  assign \new_[82340]_  = \new_[82339]_  & \new_[82332]_ ;
  assign \new_[82344]_  = ~A167 & A168;
  assign \new_[82345]_  = A169 & \new_[82344]_ ;
  assign \new_[82348]_  = ~A199 & A166;
  assign \new_[82351]_  = ~A201 & A200;
  assign \new_[82352]_  = \new_[82351]_  & \new_[82348]_ ;
  assign \new_[82353]_  = \new_[82352]_  & \new_[82345]_ ;
  assign \new_[82356]_  = ~A203 & ~A202;
  assign \new_[82359]_  = A266 & ~A265;
  assign \new_[82360]_  = \new_[82359]_  & \new_[82356]_ ;
  assign \new_[82363]_  = A269 & A267;
  assign \new_[82366]_  = A301 & ~A300;
  assign \new_[82367]_  = \new_[82366]_  & \new_[82363]_ ;
  assign \new_[82368]_  = \new_[82367]_  & \new_[82360]_ ;
  assign \new_[82372]_  = ~A167 & A168;
  assign \new_[82373]_  = A169 & \new_[82372]_ ;
  assign \new_[82376]_  = ~A199 & A166;
  assign \new_[82379]_  = ~A201 & A200;
  assign \new_[82380]_  = \new_[82379]_  & \new_[82376]_ ;
  assign \new_[82381]_  = \new_[82380]_  & \new_[82373]_ ;
  assign \new_[82384]_  = ~A203 & ~A202;
  assign \new_[82387]_  = A266 & ~A265;
  assign \new_[82388]_  = \new_[82387]_  & \new_[82384]_ ;
  assign \new_[82391]_  = A269 & A267;
  assign \new_[82394]_  = A302 & ~A300;
  assign \new_[82395]_  = \new_[82394]_  & \new_[82391]_ ;
  assign \new_[82396]_  = \new_[82395]_  & \new_[82388]_ ;
  assign \new_[82400]_  = ~A167 & A168;
  assign \new_[82401]_  = A169 & \new_[82400]_ ;
  assign \new_[82404]_  = ~A199 & A166;
  assign \new_[82407]_  = ~A201 & A200;
  assign \new_[82408]_  = \new_[82407]_  & \new_[82404]_ ;
  assign \new_[82409]_  = \new_[82408]_  & \new_[82401]_ ;
  assign \new_[82412]_  = ~A203 & ~A202;
  assign \new_[82415]_  = A266 & ~A265;
  assign \new_[82416]_  = \new_[82415]_  & \new_[82412]_ ;
  assign \new_[82419]_  = A269 & A267;
  assign \new_[82422]_  = A299 & A298;
  assign \new_[82423]_  = \new_[82422]_  & \new_[82419]_ ;
  assign \new_[82424]_  = \new_[82423]_  & \new_[82416]_ ;
  assign \new_[82428]_  = ~A167 & A168;
  assign \new_[82429]_  = A169 & \new_[82428]_ ;
  assign \new_[82432]_  = ~A199 & A166;
  assign \new_[82435]_  = ~A201 & A200;
  assign \new_[82436]_  = \new_[82435]_  & \new_[82432]_ ;
  assign \new_[82437]_  = \new_[82436]_  & \new_[82429]_ ;
  assign \new_[82440]_  = ~A203 & ~A202;
  assign \new_[82443]_  = A266 & ~A265;
  assign \new_[82444]_  = \new_[82443]_  & \new_[82440]_ ;
  assign \new_[82447]_  = A269 & A267;
  assign \new_[82450]_  = ~A299 & ~A298;
  assign \new_[82451]_  = \new_[82450]_  & \new_[82447]_ ;
  assign \new_[82452]_  = \new_[82451]_  & \new_[82444]_ ;
  assign \new_[82456]_  = ~A167 & A168;
  assign \new_[82457]_  = A169 & \new_[82456]_ ;
  assign \new_[82460]_  = ~A199 & A166;
  assign \new_[82463]_  = ~A201 & A200;
  assign \new_[82464]_  = \new_[82463]_  & \new_[82460]_ ;
  assign \new_[82465]_  = \new_[82464]_  & \new_[82457]_ ;
  assign \new_[82468]_  = ~A203 & ~A202;
  assign \new_[82471]_  = ~A266 & A265;
  assign \new_[82472]_  = \new_[82471]_  & \new_[82468]_ ;
  assign \new_[82475]_  = A268 & A267;
  assign \new_[82478]_  = A301 & ~A300;
  assign \new_[82479]_  = \new_[82478]_  & \new_[82475]_ ;
  assign \new_[82480]_  = \new_[82479]_  & \new_[82472]_ ;
  assign \new_[82484]_  = ~A167 & A168;
  assign \new_[82485]_  = A169 & \new_[82484]_ ;
  assign \new_[82488]_  = ~A199 & A166;
  assign \new_[82491]_  = ~A201 & A200;
  assign \new_[82492]_  = \new_[82491]_  & \new_[82488]_ ;
  assign \new_[82493]_  = \new_[82492]_  & \new_[82485]_ ;
  assign \new_[82496]_  = ~A203 & ~A202;
  assign \new_[82499]_  = ~A266 & A265;
  assign \new_[82500]_  = \new_[82499]_  & \new_[82496]_ ;
  assign \new_[82503]_  = A268 & A267;
  assign \new_[82506]_  = A302 & ~A300;
  assign \new_[82507]_  = \new_[82506]_  & \new_[82503]_ ;
  assign \new_[82508]_  = \new_[82507]_  & \new_[82500]_ ;
  assign \new_[82512]_  = ~A167 & A168;
  assign \new_[82513]_  = A169 & \new_[82512]_ ;
  assign \new_[82516]_  = ~A199 & A166;
  assign \new_[82519]_  = ~A201 & A200;
  assign \new_[82520]_  = \new_[82519]_  & \new_[82516]_ ;
  assign \new_[82521]_  = \new_[82520]_  & \new_[82513]_ ;
  assign \new_[82524]_  = ~A203 & ~A202;
  assign \new_[82527]_  = ~A266 & A265;
  assign \new_[82528]_  = \new_[82527]_  & \new_[82524]_ ;
  assign \new_[82531]_  = A268 & A267;
  assign \new_[82534]_  = A299 & A298;
  assign \new_[82535]_  = \new_[82534]_  & \new_[82531]_ ;
  assign \new_[82536]_  = \new_[82535]_  & \new_[82528]_ ;
  assign \new_[82540]_  = ~A167 & A168;
  assign \new_[82541]_  = A169 & \new_[82540]_ ;
  assign \new_[82544]_  = ~A199 & A166;
  assign \new_[82547]_  = ~A201 & A200;
  assign \new_[82548]_  = \new_[82547]_  & \new_[82544]_ ;
  assign \new_[82549]_  = \new_[82548]_  & \new_[82541]_ ;
  assign \new_[82552]_  = ~A203 & ~A202;
  assign \new_[82555]_  = ~A266 & A265;
  assign \new_[82556]_  = \new_[82555]_  & \new_[82552]_ ;
  assign \new_[82559]_  = A268 & A267;
  assign \new_[82562]_  = ~A299 & ~A298;
  assign \new_[82563]_  = \new_[82562]_  & \new_[82559]_ ;
  assign \new_[82564]_  = \new_[82563]_  & \new_[82556]_ ;
  assign \new_[82568]_  = ~A167 & A168;
  assign \new_[82569]_  = A169 & \new_[82568]_ ;
  assign \new_[82572]_  = ~A199 & A166;
  assign \new_[82575]_  = ~A201 & A200;
  assign \new_[82576]_  = \new_[82575]_  & \new_[82572]_ ;
  assign \new_[82577]_  = \new_[82576]_  & \new_[82569]_ ;
  assign \new_[82580]_  = ~A203 & ~A202;
  assign \new_[82583]_  = ~A266 & A265;
  assign \new_[82584]_  = \new_[82583]_  & \new_[82580]_ ;
  assign \new_[82587]_  = A269 & A267;
  assign \new_[82590]_  = A301 & ~A300;
  assign \new_[82591]_  = \new_[82590]_  & \new_[82587]_ ;
  assign \new_[82592]_  = \new_[82591]_  & \new_[82584]_ ;
  assign \new_[82596]_  = ~A167 & A168;
  assign \new_[82597]_  = A169 & \new_[82596]_ ;
  assign \new_[82600]_  = ~A199 & A166;
  assign \new_[82603]_  = ~A201 & A200;
  assign \new_[82604]_  = \new_[82603]_  & \new_[82600]_ ;
  assign \new_[82605]_  = \new_[82604]_  & \new_[82597]_ ;
  assign \new_[82608]_  = ~A203 & ~A202;
  assign \new_[82611]_  = ~A266 & A265;
  assign \new_[82612]_  = \new_[82611]_  & \new_[82608]_ ;
  assign \new_[82615]_  = A269 & A267;
  assign \new_[82618]_  = A302 & ~A300;
  assign \new_[82619]_  = \new_[82618]_  & \new_[82615]_ ;
  assign \new_[82620]_  = \new_[82619]_  & \new_[82612]_ ;
  assign \new_[82624]_  = ~A167 & A168;
  assign \new_[82625]_  = A169 & \new_[82624]_ ;
  assign \new_[82628]_  = ~A199 & A166;
  assign \new_[82631]_  = ~A201 & A200;
  assign \new_[82632]_  = \new_[82631]_  & \new_[82628]_ ;
  assign \new_[82633]_  = \new_[82632]_  & \new_[82625]_ ;
  assign \new_[82636]_  = ~A203 & ~A202;
  assign \new_[82639]_  = ~A266 & A265;
  assign \new_[82640]_  = \new_[82639]_  & \new_[82636]_ ;
  assign \new_[82643]_  = A269 & A267;
  assign \new_[82646]_  = A299 & A298;
  assign \new_[82647]_  = \new_[82646]_  & \new_[82643]_ ;
  assign \new_[82648]_  = \new_[82647]_  & \new_[82640]_ ;
  assign \new_[82652]_  = ~A167 & A168;
  assign \new_[82653]_  = A169 & \new_[82652]_ ;
  assign \new_[82656]_  = ~A199 & A166;
  assign \new_[82659]_  = ~A201 & A200;
  assign \new_[82660]_  = \new_[82659]_  & \new_[82656]_ ;
  assign \new_[82661]_  = \new_[82660]_  & \new_[82653]_ ;
  assign \new_[82664]_  = ~A203 & ~A202;
  assign \new_[82667]_  = ~A266 & A265;
  assign \new_[82668]_  = \new_[82667]_  & \new_[82664]_ ;
  assign \new_[82671]_  = A269 & A267;
  assign \new_[82674]_  = ~A299 & ~A298;
  assign \new_[82675]_  = \new_[82674]_  & \new_[82671]_ ;
  assign \new_[82676]_  = \new_[82675]_  & \new_[82668]_ ;
  assign \new_[82680]_  = ~A167 & A168;
  assign \new_[82681]_  = A169 & \new_[82680]_ ;
  assign \new_[82684]_  = A199 & A166;
  assign \new_[82687]_  = A201 & ~A200;
  assign \new_[82688]_  = \new_[82687]_  & \new_[82684]_ ;
  assign \new_[82689]_  = \new_[82688]_  & \new_[82681]_ ;
  assign \new_[82692]_  = ~A265 & A202;
  assign \new_[82695]_  = A267 & A266;
  assign \new_[82696]_  = \new_[82695]_  & \new_[82692]_ ;
  assign \new_[82699]_  = A300 & A268;
  assign \new_[82702]_  = ~A302 & ~A301;
  assign \new_[82703]_  = \new_[82702]_  & \new_[82699]_ ;
  assign \new_[82704]_  = \new_[82703]_  & \new_[82696]_ ;
  assign \new_[82708]_  = ~A167 & A168;
  assign \new_[82709]_  = A169 & \new_[82708]_ ;
  assign \new_[82712]_  = A199 & A166;
  assign \new_[82715]_  = A201 & ~A200;
  assign \new_[82716]_  = \new_[82715]_  & \new_[82712]_ ;
  assign \new_[82717]_  = \new_[82716]_  & \new_[82709]_ ;
  assign \new_[82720]_  = ~A265 & A202;
  assign \new_[82723]_  = A267 & A266;
  assign \new_[82724]_  = \new_[82723]_  & \new_[82720]_ ;
  assign \new_[82727]_  = A300 & A269;
  assign \new_[82730]_  = ~A302 & ~A301;
  assign \new_[82731]_  = \new_[82730]_  & \new_[82727]_ ;
  assign \new_[82732]_  = \new_[82731]_  & \new_[82724]_ ;
  assign \new_[82736]_  = ~A167 & A168;
  assign \new_[82737]_  = A169 & \new_[82736]_ ;
  assign \new_[82740]_  = A199 & A166;
  assign \new_[82743]_  = A201 & ~A200;
  assign \new_[82744]_  = \new_[82743]_  & \new_[82740]_ ;
  assign \new_[82745]_  = \new_[82744]_  & \new_[82737]_ ;
  assign \new_[82748]_  = ~A265 & A202;
  assign \new_[82751]_  = ~A267 & A266;
  assign \new_[82752]_  = \new_[82751]_  & \new_[82748]_ ;
  assign \new_[82755]_  = ~A269 & ~A268;
  assign \new_[82758]_  = A301 & ~A300;
  assign \new_[82759]_  = \new_[82758]_  & \new_[82755]_ ;
  assign \new_[82760]_  = \new_[82759]_  & \new_[82752]_ ;
  assign \new_[82764]_  = ~A167 & A168;
  assign \new_[82765]_  = A169 & \new_[82764]_ ;
  assign \new_[82768]_  = A199 & A166;
  assign \new_[82771]_  = A201 & ~A200;
  assign \new_[82772]_  = \new_[82771]_  & \new_[82768]_ ;
  assign \new_[82773]_  = \new_[82772]_  & \new_[82765]_ ;
  assign \new_[82776]_  = ~A265 & A202;
  assign \new_[82779]_  = ~A267 & A266;
  assign \new_[82780]_  = \new_[82779]_  & \new_[82776]_ ;
  assign \new_[82783]_  = ~A269 & ~A268;
  assign \new_[82786]_  = A302 & ~A300;
  assign \new_[82787]_  = \new_[82786]_  & \new_[82783]_ ;
  assign \new_[82788]_  = \new_[82787]_  & \new_[82780]_ ;
  assign \new_[82792]_  = ~A167 & A168;
  assign \new_[82793]_  = A169 & \new_[82792]_ ;
  assign \new_[82796]_  = A199 & A166;
  assign \new_[82799]_  = A201 & ~A200;
  assign \new_[82800]_  = \new_[82799]_  & \new_[82796]_ ;
  assign \new_[82801]_  = \new_[82800]_  & \new_[82793]_ ;
  assign \new_[82804]_  = ~A265 & A202;
  assign \new_[82807]_  = ~A267 & A266;
  assign \new_[82808]_  = \new_[82807]_  & \new_[82804]_ ;
  assign \new_[82811]_  = ~A269 & ~A268;
  assign \new_[82814]_  = A299 & A298;
  assign \new_[82815]_  = \new_[82814]_  & \new_[82811]_ ;
  assign \new_[82816]_  = \new_[82815]_  & \new_[82808]_ ;
  assign \new_[82820]_  = ~A167 & A168;
  assign \new_[82821]_  = A169 & \new_[82820]_ ;
  assign \new_[82824]_  = A199 & A166;
  assign \new_[82827]_  = A201 & ~A200;
  assign \new_[82828]_  = \new_[82827]_  & \new_[82824]_ ;
  assign \new_[82829]_  = \new_[82828]_  & \new_[82821]_ ;
  assign \new_[82832]_  = ~A265 & A202;
  assign \new_[82835]_  = ~A267 & A266;
  assign \new_[82836]_  = \new_[82835]_  & \new_[82832]_ ;
  assign \new_[82839]_  = ~A269 & ~A268;
  assign \new_[82842]_  = ~A299 & ~A298;
  assign \new_[82843]_  = \new_[82842]_  & \new_[82839]_ ;
  assign \new_[82844]_  = \new_[82843]_  & \new_[82836]_ ;
  assign \new_[82848]_  = ~A167 & A168;
  assign \new_[82849]_  = A169 & \new_[82848]_ ;
  assign \new_[82852]_  = A199 & A166;
  assign \new_[82855]_  = A201 & ~A200;
  assign \new_[82856]_  = \new_[82855]_  & \new_[82852]_ ;
  assign \new_[82857]_  = \new_[82856]_  & \new_[82849]_ ;
  assign \new_[82860]_  = A265 & A202;
  assign \new_[82863]_  = A267 & ~A266;
  assign \new_[82864]_  = \new_[82863]_  & \new_[82860]_ ;
  assign \new_[82867]_  = A300 & A268;
  assign \new_[82870]_  = ~A302 & ~A301;
  assign \new_[82871]_  = \new_[82870]_  & \new_[82867]_ ;
  assign \new_[82872]_  = \new_[82871]_  & \new_[82864]_ ;
  assign \new_[82876]_  = ~A167 & A168;
  assign \new_[82877]_  = A169 & \new_[82876]_ ;
  assign \new_[82880]_  = A199 & A166;
  assign \new_[82883]_  = A201 & ~A200;
  assign \new_[82884]_  = \new_[82883]_  & \new_[82880]_ ;
  assign \new_[82885]_  = \new_[82884]_  & \new_[82877]_ ;
  assign \new_[82888]_  = A265 & A202;
  assign \new_[82891]_  = A267 & ~A266;
  assign \new_[82892]_  = \new_[82891]_  & \new_[82888]_ ;
  assign \new_[82895]_  = A300 & A269;
  assign \new_[82898]_  = ~A302 & ~A301;
  assign \new_[82899]_  = \new_[82898]_  & \new_[82895]_ ;
  assign \new_[82900]_  = \new_[82899]_  & \new_[82892]_ ;
  assign \new_[82904]_  = ~A167 & A168;
  assign \new_[82905]_  = A169 & \new_[82904]_ ;
  assign \new_[82908]_  = A199 & A166;
  assign \new_[82911]_  = A201 & ~A200;
  assign \new_[82912]_  = \new_[82911]_  & \new_[82908]_ ;
  assign \new_[82913]_  = \new_[82912]_  & \new_[82905]_ ;
  assign \new_[82916]_  = A265 & A202;
  assign \new_[82919]_  = ~A267 & ~A266;
  assign \new_[82920]_  = \new_[82919]_  & \new_[82916]_ ;
  assign \new_[82923]_  = ~A269 & ~A268;
  assign \new_[82926]_  = A301 & ~A300;
  assign \new_[82927]_  = \new_[82926]_  & \new_[82923]_ ;
  assign \new_[82928]_  = \new_[82927]_  & \new_[82920]_ ;
  assign \new_[82932]_  = ~A167 & A168;
  assign \new_[82933]_  = A169 & \new_[82932]_ ;
  assign \new_[82936]_  = A199 & A166;
  assign \new_[82939]_  = A201 & ~A200;
  assign \new_[82940]_  = \new_[82939]_  & \new_[82936]_ ;
  assign \new_[82941]_  = \new_[82940]_  & \new_[82933]_ ;
  assign \new_[82944]_  = A265 & A202;
  assign \new_[82947]_  = ~A267 & ~A266;
  assign \new_[82948]_  = \new_[82947]_  & \new_[82944]_ ;
  assign \new_[82951]_  = ~A269 & ~A268;
  assign \new_[82954]_  = A302 & ~A300;
  assign \new_[82955]_  = \new_[82954]_  & \new_[82951]_ ;
  assign \new_[82956]_  = \new_[82955]_  & \new_[82948]_ ;
  assign \new_[82960]_  = ~A167 & A168;
  assign \new_[82961]_  = A169 & \new_[82960]_ ;
  assign \new_[82964]_  = A199 & A166;
  assign \new_[82967]_  = A201 & ~A200;
  assign \new_[82968]_  = \new_[82967]_  & \new_[82964]_ ;
  assign \new_[82969]_  = \new_[82968]_  & \new_[82961]_ ;
  assign \new_[82972]_  = A265 & A202;
  assign \new_[82975]_  = ~A267 & ~A266;
  assign \new_[82976]_  = \new_[82975]_  & \new_[82972]_ ;
  assign \new_[82979]_  = ~A269 & ~A268;
  assign \new_[82982]_  = A299 & A298;
  assign \new_[82983]_  = \new_[82982]_  & \new_[82979]_ ;
  assign \new_[82984]_  = \new_[82983]_  & \new_[82976]_ ;
  assign \new_[82988]_  = ~A167 & A168;
  assign \new_[82989]_  = A169 & \new_[82988]_ ;
  assign \new_[82992]_  = A199 & A166;
  assign \new_[82995]_  = A201 & ~A200;
  assign \new_[82996]_  = \new_[82995]_  & \new_[82992]_ ;
  assign \new_[82997]_  = \new_[82996]_  & \new_[82989]_ ;
  assign \new_[83000]_  = A265 & A202;
  assign \new_[83003]_  = ~A267 & ~A266;
  assign \new_[83004]_  = \new_[83003]_  & \new_[83000]_ ;
  assign \new_[83007]_  = ~A269 & ~A268;
  assign \new_[83010]_  = ~A299 & ~A298;
  assign \new_[83011]_  = \new_[83010]_  & \new_[83007]_ ;
  assign \new_[83012]_  = \new_[83011]_  & \new_[83004]_ ;
  assign \new_[83016]_  = ~A167 & A168;
  assign \new_[83017]_  = A169 & \new_[83016]_ ;
  assign \new_[83020]_  = A199 & A166;
  assign \new_[83023]_  = A201 & ~A200;
  assign \new_[83024]_  = \new_[83023]_  & \new_[83020]_ ;
  assign \new_[83025]_  = \new_[83024]_  & \new_[83017]_ ;
  assign \new_[83028]_  = ~A265 & A203;
  assign \new_[83031]_  = A267 & A266;
  assign \new_[83032]_  = \new_[83031]_  & \new_[83028]_ ;
  assign \new_[83035]_  = A300 & A268;
  assign \new_[83038]_  = ~A302 & ~A301;
  assign \new_[83039]_  = \new_[83038]_  & \new_[83035]_ ;
  assign \new_[83040]_  = \new_[83039]_  & \new_[83032]_ ;
  assign \new_[83044]_  = ~A167 & A168;
  assign \new_[83045]_  = A169 & \new_[83044]_ ;
  assign \new_[83048]_  = A199 & A166;
  assign \new_[83051]_  = A201 & ~A200;
  assign \new_[83052]_  = \new_[83051]_  & \new_[83048]_ ;
  assign \new_[83053]_  = \new_[83052]_  & \new_[83045]_ ;
  assign \new_[83056]_  = ~A265 & A203;
  assign \new_[83059]_  = A267 & A266;
  assign \new_[83060]_  = \new_[83059]_  & \new_[83056]_ ;
  assign \new_[83063]_  = A300 & A269;
  assign \new_[83066]_  = ~A302 & ~A301;
  assign \new_[83067]_  = \new_[83066]_  & \new_[83063]_ ;
  assign \new_[83068]_  = \new_[83067]_  & \new_[83060]_ ;
  assign \new_[83072]_  = ~A167 & A168;
  assign \new_[83073]_  = A169 & \new_[83072]_ ;
  assign \new_[83076]_  = A199 & A166;
  assign \new_[83079]_  = A201 & ~A200;
  assign \new_[83080]_  = \new_[83079]_  & \new_[83076]_ ;
  assign \new_[83081]_  = \new_[83080]_  & \new_[83073]_ ;
  assign \new_[83084]_  = ~A265 & A203;
  assign \new_[83087]_  = ~A267 & A266;
  assign \new_[83088]_  = \new_[83087]_  & \new_[83084]_ ;
  assign \new_[83091]_  = ~A269 & ~A268;
  assign \new_[83094]_  = A301 & ~A300;
  assign \new_[83095]_  = \new_[83094]_  & \new_[83091]_ ;
  assign \new_[83096]_  = \new_[83095]_  & \new_[83088]_ ;
  assign \new_[83100]_  = ~A167 & A168;
  assign \new_[83101]_  = A169 & \new_[83100]_ ;
  assign \new_[83104]_  = A199 & A166;
  assign \new_[83107]_  = A201 & ~A200;
  assign \new_[83108]_  = \new_[83107]_  & \new_[83104]_ ;
  assign \new_[83109]_  = \new_[83108]_  & \new_[83101]_ ;
  assign \new_[83112]_  = ~A265 & A203;
  assign \new_[83115]_  = ~A267 & A266;
  assign \new_[83116]_  = \new_[83115]_  & \new_[83112]_ ;
  assign \new_[83119]_  = ~A269 & ~A268;
  assign \new_[83122]_  = A302 & ~A300;
  assign \new_[83123]_  = \new_[83122]_  & \new_[83119]_ ;
  assign \new_[83124]_  = \new_[83123]_  & \new_[83116]_ ;
  assign \new_[83128]_  = ~A167 & A168;
  assign \new_[83129]_  = A169 & \new_[83128]_ ;
  assign \new_[83132]_  = A199 & A166;
  assign \new_[83135]_  = A201 & ~A200;
  assign \new_[83136]_  = \new_[83135]_  & \new_[83132]_ ;
  assign \new_[83137]_  = \new_[83136]_  & \new_[83129]_ ;
  assign \new_[83140]_  = ~A265 & A203;
  assign \new_[83143]_  = ~A267 & A266;
  assign \new_[83144]_  = \new_[83143]_  & \new_[83140]_ ;
  assign \new_[83147]_  = ~A269 & ~A268;
  assign \new_[83150]_  = A299 & A298;
  assign \new_[83151]_  = \new_[83150]_  & \new_[83147]_ ;
  assign \new_[83152]_  = \new_[83151]_  & \new_[83144]_ ;
  assign \new_[83156]_  = ~A167 & A168;
  assign \new_[83157]_  = A169 & \new_[83156]_ ;
  assign \new_[83160]_  = A199 & A166;
  assign \new_[83163]_  = A201 & ~A200;
  assign \new_[83164]_  = \new_[83163]_  & \new_[83160]_ ;
  assign \new_[83165]_  = \new_[83164]_  & \new_[83157]_ ;
  assign \new_[83168]_  = ~A265 & A203;
  assign \new_[83171]_  = ~A267 & A266;
  assign \new_[83172]_  = \new_[83171]_  & \new_[83168]_ ;
  assign \new_[83175]_  = ~A269 & ~A268;
  assign \new_[83178]_  = ~A299 & ~A298;
  assign \new_[83179]_  = \new_[83178]_  & \new_[83175]_ ;
  assign \new_[83180]_  = \new_[83179]_  & \new_[83172]_ ;
  assign \new_[83184]_  = ~A167 & A168;
  assign \new_[83185]_  = A169 & \new_[83184]_ ;
  assign \new_[83188]_  = A199 & A166;
  assign \new_[83191]_  = A201 & ~A200;
  assign \new_[83192]_  = \new_[83191]_  & \new_[83188]_ ;
  assign \new_[83193]_  = \new_[83192]_  & \new_[83185]_ ;
  assign \new_[83196]_  = A265 & A203;
  assign \new_[83199]_  = A267 & ~A266;
  assign \new_[83200]_  = \new_[83199]_  & \new_[83196]_ ;
  assign \new_[83203]_  = A300 & A268;
  assign \new_[83206]_  = ~A302 & ~A301;
  assign \new_[83207]_  = \new_[83206]_  & \new_[83203]_ ;
  assign \new_[83208]_  = \new_[83207]_  & \new_[83200]_ ;
  assign \new_[83212]_  = ~A167 & A168;
  assign \new_[83213]_  = A169 & \new_[83212]_ ;
  assign \new_[83216]_  = A199 & A166;
  assign \new_[83219]_  = A201 & ~A200;
  assign \new_[83220]_  = \new_[83219]_  & \new_[83216]_ ;
  assign \new_[83221]_  = \new_[83220]_  & \new_[83213]_ ;
  assign \new_[83224]_  = A265 & A203;
  assign \new_[83227]_  = A267 & ~A266;
  assign \new_[83228]_  = \new_[83227]_  & \new_[83224]_ ;
  assign \new_[83231]_  = A300 & A269;
  assign \new_[83234]_  = ~A302 & ~A301;
  assign \new_[83235]_  = \new_[83234]_  & \new_[83231]_ ;
  assign \new_[83236]_  = \new_[83235]_  & \new_[83228]_ ;
  assign \new_[83240]_  = ~A167 & A168;
  assign \new_[83241]_  = A169 & \new_[83240]_ ;
  assign \new_[83244]_  = A199 & A166;
  assign \new_[83247]_  = A201 & ~A200;
  assign \new_[83248]_  = \new_[83247]_  & \new_[83244]_ ;
  assign \new_[83249]_  = \new_[83248]_  & \new_[83241]_ ;
  assign \new_[83252]_  = A265 & A203;
  assign \new_[83255]_  = ~A267 & ~A266;
  assign \new_[83256]_  = \new_[83255]_  & \new_[83252]_ ;
  assign \new_[83259]_  = ~A269 & ~A268;
  assign \new_[83262]_  = A301 & ~A300;
  assign \new_[83263]_  = \new_[83262]_  & \new_[83259]_ ;
  assign \new_[83264]_  = \new_[83263]_  & \new_[83256]_ ;
  assign \new_[83268]_  = ~A167 & A168;
  assign \new_[83269]_  = A169 & \new_[83268]_ ;
  assign \new_[83272]_  = A199 & A166;
  assign \new_[83275]_  = A201 & ~A200;
  assign \new_[83276]_  = \new_[83275]_  & \new_[83272]_ ;
  assign \new_[83277]_  = \new_[83276]_  & \new_[83269]_ ;
  assign \new_[83280]_  = A265 & A203;
  assign \new_[83283]_  = ~A267 & ~A266;
  assign \new_[83284]_  = \new_[83283]_  & \new_[83280]_ ;
  assign \new_[83287]_  = ~A269 & ~A268;
  assign \new_[83290]_  = A302 & ~A300;
  assign \new_[83291]_  = \new_[83290]_  & \new_[83287]_ ;
  assign \new_[83292]_  = \new_[83291]_  & \new_[83284]_ ;
  assign \new_[83296]_  = ~A167 & A168;
  assign \new_[83297]_  = A169 & \new_[83296]_ ;
  assign \new_[83300]_  = A199 & A166;
  assign \new_[83303]_  = A201 & ~A200;
  assign \new_[83304]_  = \new_[83303]_  & \new_[83300]_ ;
  assign \new_[83305]_  = \new_[83304]_  & \new_[83297]_ ;
  assign \new_[83308]_  = A265 & A203;
  assign \new_[83311]_  = ~A267 & ~A266;
  assign \new_[83312]_  = \new_[83311]_  & \new_[83308]_ ;
  assign \new_[83315]_  = ~A269 & ~A268;
  assign \new_[83318]_  = A299 & A298;
  assign \new_[83319]_  = \new_[83318]_  & \new_[83315]_ ;
  assign \new_[83320]_  = \new_[83319]_  & \new_[83312]_ ;
  assign \new_[83324]_  = ~A167 & A168;
  assign \new_[83325]_  = A169 & \new_[83324]_ ;
  assign \new_[83328]_  = A199 & A166;
  assign \new_[83331]_  = A201 & ~A200;
  assign \new_[83332]_  = \new_[83331]_  & \new_[83328]_ ;
  assign \new_[83333]_  = \new_[83332]_  & \new_[83325]_ ;
  assign \new_[83336]_  = A265 & A203;
  assign \new_[83339]_  = ~A267 & ~A266;
  assign \new_[83340]_  = \new_[83339]_  & \new_[83336]_ ;
  assign \new_[83343]_  = ~A269 & ~A268;
  assign \new_[83346]_  = ~A299 & ~A298;
  assign \new_[83347]_  = \new_[83346]_  & \new_[83343]_ ;
  assign \new_[83348]_  = \new_[83347]_  & \new_[83340]_ ;
  assign \new_[83352]_  = ~A167 & A168;
  assign \new_[83353]_  = A169 & \new_[83352]_ ;
  assign \new_[83356]_  = A199 & A166;
  assign \new_[83359]_  = ~A201 & ~A200;
  assign \new_[83360]_  = \new_[83359]_  & \new_[83356]_ ;
  assign \new_[83361]_  = \new_[83360]_  & \new_[83353]_ ;
  assign \new_[83364]_  = ~A203 & ~A202;
  assign \new_[83367]_  = A266 & ~A265;
  assign \new_[83368]_  = \new_[83367]_  & \new_[83364]_ ;
  assign \new_[83371]_  = A268 & A267;
  assign \new_[83374]_  = A301 & ~A300;
  assign \new_[83375]_  = \new_[83374]_  & \new_[83371]_ ;
  assign \new_[83376]_  = \new_[83375]_  & \new_[83368]_ ;
  assign \new_[83380]_  = ~A167 & A168;
  assign \new_[83381]_  = A169 & \new_[83380]_ ;
  assign \new_[83384]_  = A199 & A166;
  assign \new_[83387]_  = ~A201 & ~A200;
  assign \new_[83388]_  = \new_[83387]_  & \new_[83384]_ ;
  assign \new_[83389]_  = \new_[83388]_  & \new_[83381]_ ;
  assign \new_[83392]_  = ~A203 & ~A202;
  assign \new_[83395]_  = A266 & ~A265;
  assign \new_[83396]_  = \new_[83395]_  & \new_[83392]_ ;
  assign \new_[83399]_  = A268 & A267;
  assign \new_[83402]_  = A302 & ~A300;
  assign \new_[83403]_  = \new_[83402]_  & \new_[83399]_ ;
  assign \new_[83404]_  = \new_[83403]_  & \new_[83396]_ ;
  assign \new_[83408]_  = ~A167 & A168;
  assign \new_[83409]_  = A169 & \new_[83408]_ ;
  assign \new_[83412]_  = A199 & A166;
  assign \new_[83415]_  = ~A201 & ~A200;
  assign \new_[83416]_  = \new_[83415]_  & \new_[83412]_ ;
  assign \new_[83417]_  = \new_[83416]_  & \new_[83409]_ ;
  assign \new_[83420]_  = ~A203 & ~A202;
  assign \new_[83423]_  = A266 & ~A265;
  assign \new_[83424]_  = \new_[83423]_  & \new_[83420]_ ;
  assign \new_[83427]_  = A268 & A267;
  assign \new_[83430]_  = A299 & A298;
  assign \new_[83431]_  = \new_[83430]_  & \new_[83427]_ ;
  assign \new_[83432]_  = \new_[83431]_  & \new_[83424]_ ;
  assign \new_[83436]_  = ~A167 & A168;
  assign \new_[83437]_  = A169 & \new_[83436]_ ;
  assign \new_[83440]_  = A199 & A166;
  assign \new_[83443]_  = ~A201 & ~A200;
  assign \new_[83444]_  = \new_[83443]_  & \new_[83440]_ ;
  assign \new_[83445]_  = \new_[83444]_  & \new_[83437]_ ;
  assign \new_[83448]_  = ~A203 & ~A202;
  assign \new_[83451]_  = A266 & ~A265;
  assign \new_[83452]_  = \new_[83451]_  & \new_[83448]_ ;
  assign \new_[83455]_  = A268 & A267;
  assign \new_[83458]_  = ~A299 & ~A298;
  assign \new_[83459]_  = \new_[83458]_  & \new_[83455]_ ;
  assign \new_[83460]_  = \new_[83459]_  & \new_[83452]_ ;
  assign \new_[83464]_  = ~A167 & A168;
  assign \new_[83465]_  = A169 & \new_[83464]_ ;
  assign \new_[83468]_  = A199 & A166;
  assign \new_[83471]_  = ~A201 & ~A200;
  assign \new_[83472]_  = \new_[83471]_  & \new_[83468]_ ;
  assign \new_[83473]_  = \new_[83472]_  & \new_[83465]_ ;
  assign \new_[83476]_  = ~A203 & ~A202;
  assign \new_[83479]_  = A266 & ~A265;
  assign \new_[83480]_  = \new_[83479]_  & \new_[83476]_ ;
  assign \new_[83483]_  = A269 & A267;
  assign \new_[83486]_  = A301 & ~A300;
  assign \new_[83487]_  = \new_[83486]_  & \new_[83483]_ ;
  assign \new_[83488]_  = \new_[83487]_  & \new_[83480]_ ;
  assign \new_[83492]_  = ~A167 & A168;
  assign \new_[83493]_  = A169 & \new_[83492]_ ;
  assign \new_[83496]_  = A199 & A166;
  assign \new_[83499]_  = ~A201 & ~A200;
  assign \new_[83500]_  = \new_[83499]_  & \new_[83496]_ ;
  assign \new_[83501]_  = \new_[83500]_  & \new_[83493]_ ;
  assign \new_[83504]_  = ~A203 & ~A202;
  assign \new_[83507]_  = A266 & ~A265;
  assign \new_[83508]_  = \new_[83507]_  & \new_[83504]_ ;
  assign \new_[83511]_  = A269 & A267;
  assign \new_[83514]_  = A302 & ~A300;
  assign \new_[83515]_  = \new_[83514]_  & \new_[83511]_ ;
  assign \new_[83516]_  = \new_[83515]_  & \new_[83508]_ ;
  assign \new_[83520]_  = ~A167 & A168;
  assign \new_[83521]_  = A169 & \new_[83520]_ ;
  assign \new_[83524]_  = A199 & A166;
  assign \new_[83527]_  = ~A201 & ~A200;
  assign \new_[83528]_  = \new_[83527]_  & \new_[83524]_ ;
  assign \new_[83529]_  = \new_[83528]_  & \new_[83521]_ ;
  assign \new_[83532]_  = ~A203 & ~A202;
  assign \new_[83535]_  = A266 & ~A265;
  assign \new_[83536]_  = \new_[83535]_  & \new_[83532]_ ;
  assign \new_[83539]_  = A269 & A267;
  assign \new_[83542]_  = A299 & A298;
  assign \new_[83543]_  = \new_[83542]_  & \new_[83539]_ ;
  assign \new_[83544]_  = \new_[83543]_  & \new_[83536]_ ;
  assign \new_[83548]_  = ~A167 & A168;
  assign \new_[83549]_  = A169 & \new_[83548]_ ;
  assign \new_[83552]_  = A199 & A166;
  assign \new_[83555]_  = ~A201 & ~A200;
  assign \new_[83556]_  = \new_[83555]_  & \new_[83552]_ ;
  assign \new_[83557]_  = \new_[83556]_  & \new_[83549]_ ;
  assign \new_[83560]_  = ~A203 & ~A202;
  assign \new_[83563]_  = A266 & ~A265;
  assign \new_[83564]_  = \new_[83563]_  & \new_[83560]_ ;
  assign \new_[83567]_  = A269 & A267;
  assign \new_[83570]_  = ~A299 & ~A298;
  assign \new_[83571]_  = \new_[83570]_  & \new_[83567]_ ;
  assign \new_[83572]_  = \new_[83571]_  & \new_[83564]_ ;
  assign \new_[83576]_  = ~A167 & A168;
  assign \new_[83577]_  = A169 & \new_[83576]_ ;
  assign \new_[83580]_  = A199 & A166;
  assign \new_[83583]_  = ~A201 & ~A200;
  assign \new_[83584]_  = \new_[83583]_  & \new_[83580]_ ;
  assign \new_[83585]_  = \new_[83584]_  & \new_[83577]_ ;
  assign \new_[83588]_  = ~A203 & ~A202;
  assign \new_[83591]_  = ~A266 & A265;
  assign \new_[83592]_  = \new_[83591]_  & \new_[83588]_ ;
  assign \new_[83595]_  = A268 & A267;
  assign \new_[83598]_  = A301 & ~A300;
  assign \new_[83599]_  = \new_[83598]_  & \new_[83595]_ ;
  assign \new_[83600]_  = \new_[83599]_  & \new_[83592]_ ;
  assign \new_[83604]_  = ~A167 & A168;
  assign \new_[83605]_  = A169 & \new_[83604]_ ;
  assign \new_[83608]_  = A199 & A166;
  assign \new_[83611]_  = ~A201 & ~A200;
  assign \new_[83612]_  = \new_[83611]_  & \new_[83608]_ ;
  assign \new_[83613]_  = \new_[83612]_  & \new_[83605]_ ;
  assign \new_[83616]_  = ~A203 & ~A202;
  assign \new_[83619]_  = ~A266 & A265;
  assign \new_[83620]_  = \new_[83619]_  & \new_[83616]_ ;
  assign \new_[83623]_  = A268 & A267;
  assign \new_[83626]_  = A302 & ~A300;
  assign \new_[83627]_  = \new_[83626]_  & \new_[83623]_ ;
  assign \new_[83628]_  = \new_[83627]_  & \new_[83620]_ ;
  assign \new_[83632]_  = ~A167 & A168;
  assign \new_[83633]_  = A169 & \new_[83632]_ ;
  assign \new_[83636]_  = A199 & A166;
  assign \new_[83639]_  = ~A201 & ~A200;
  assign \new_[83640]_  = \new_[83639]_  & \new_[83636]_ ;
  assign \new_[83641]_  = \new_[83640]_  & \new_[83633]_ ;
  assign \new_[83644]_  = ~A203 & ~A202;
  assign \new_[83647]_  = ~A266 & A265;
  assign \new_[83648]_  = \new_[83647]_  & \new_[83644]_ ;
  assign \new_[83651]_  = A268 & A267;
  assign \new_[83654]_  = A299 & A298;
  assign \new_[83655]_  = \new_[83654]_  & \new_[83651]_ ;
  assign \new_[83656]_  = \new_[83655]_  & \new_[83648]_ ;
  assign \new_[83660]_  = ~A167 & A168;
  assign \new_[83661]_  = A169 & \new_[83660]_ ;
  assign \new_[83664]_  = A199 & A166;
  assign \new_[83667]_  = ~A201 & ~A200;
  assign \new_[83668]_  = \new_[83667]_  & \new_[83664]_ ;
  assign \new_[83669]_  = \new_[83668]_  & \new_[83661]_ ;
  assign \new_[83672]_  = ~A203 & ~A202;
  assign \new_[83675]_  = ~A266 & A265;
  assign \new_[83676]_  = \new_[83675]_  & \new_[83672]_ ;
  assign \new_[83679]_  = A268 & A267;
  assign \new_[83682]_  = ~A299 & ~A298;
  assign \new_[83683]_  = \new_[83682]_  & \new_[83679]_ ;
  assign \new_[83684]_  = \new_[83683]_  & \new_[83676]_ ;
  assign \new_[83688]_  = ~A167 & A168;
  assign \new_[83689]_  = A169 & \new_[83688]_ ;
  assign \new_[83692]_  = A199 & A166;
  assign \new_[83695]_  = ~A201 & ~A200;
  assign \new_[83696]_  = \new_[83695]_  & \new_[83692]_ ;
  assign \new_[83697]_  = \new_[83696]_  & \new_[83689]_ ;
  assign \new_[83700]_  = ~A203 & ~A202;
  assign \new_[83703]_  = ~A266 & A265;
  assign \new_[83704]_  = \new_[83703]_  & \new_[83700]_ ;
  assign \new_[83707]_  = A269 & A267;
  assign \new_[83710]_  = A301 & ~A300;
  assign \new_[83711]_  = \new_[83710]_  & \new_[83707]_ ;
  assign \new_[83712]_  = \new_[83711]_  & \new_[83704]_ ;
  assign \new_[83716]_  = ~A167 & A168;
  assign \new_[83717]_  = A169 & \new_[83716]_ ;
  assign \new_[83720]_  = A199 & A166;
  assign \new_[83723]_  = ~A201 & ~A200;
  assign \new_[83724]_  = \new_[83723]_  & \new_[83720]_ ;
  assign \new_[83725]_  = \new_[83724]_  & \new_[83717]_ ;
  assign \new_[83728]_  = ~A203 & ~A202;
  assign \new_[83731]_  = ~A266 & A265;
  assign \new_[83732]_  = \new_[83731]_  & \new_[83728]_ ;
  assign \new_[83735]_  = A269 & A267;
  assign \new_[83738]_  = A302 & ~A300;
  assign \new_[83739]_  = \new_[83738]_  & \new_[83735]_ ;
  assign \new_[83740]_  = \new_[83739]_  & \new_[83732]_ ;
  assign \new_[83744]_  = ~A167 & A168;
  assign \new_[83745]_  = A169 & \new_[83744]_ ;
  assign \new_[83748]_  = A199 & A166;
  assign \new_[83751]_  = ~A201 & ~A200;
  assign \new_[83752]_  = \new_[83751]_  & \new_[83748]_ ;
  assign \new_[83753]_  = \new_[83752]_  & \new_[83745]_ ;
  assign \new_[83756]_  = ~A203 & ~A202;
  assign \new_[83759]_  = ~A266 & A265;
  assign \new_[83760]_  = \new_[83759]_  & \new_[83756]_ ;
  assign \new_[83763]_  = A269 & A267;
  assign \new_[83766]_  = A299 & A298;
  assign \new_[83767]_  = \new_[83766]_  & \new_[83763]_ ;
  assign \new_[83768]_  = \new_[83767]_  & \new_[83760]_ ;
  assign \new_[83772]_  = ~A167 & A168;
  assign \new_[83773]_  = A169 & \new_[83772]_ ;
  assign \new_[83776]_  = A199 & A166;
  assign \new_[83779]_  = ~A201 & ~A200;
  assign \new_[83780]_  = \new_[83779]_  & \new_[83776]_ ;
  assign \new_[83781]_  = \new_[83780]_  & \new_[83773]_ ;
  assign \new_[83784]_  = ~A203 & ~A202;
  assign \new_[83787]_  = ~A266 & A265;
  assign \new_[83788]_  = \new_[83787]_  & \new_[83784]_ ;
  assign \new_[83791]_  = A269 & A267;
  assign \new_[83794]_  = ~A299 & ~A298;
  assign \new_[83795]_  = \new_[83794]_  & \new_[83791]_ ;
  assign \new_[83796]_  = \new_[83795]_  & \new_[83788]_ ;
  assign \new_[83800]_  = ~A199 & ~A168;
  assign \new_[83801]_  = A169 & \new_[83800]_ ;
  assign \new_[83804]_  = ~A201 & A200;
  assign \new_[83807]_  = ~A203 & ~A202;
  assign \new_[83808]_  = \new_[83807]_  & \new_[83804]_ ;
  assign \new_[83809]_  = \new_[83808]_  & \new_[83801]_ ;
  assign \new_[83812]_  = ~A268 & A267;
  assign \new_[83815]_  = A298 & ~A269;
  assign \new_[83816]_  = \new_[83815]_  & \new_[83812]_ ;
  assign \new_[83819]_  = ~A300 & ~A299;
  assign \new_[83822]_  = ~A302 & ~A301;
  assign \new_[83823]_  = \new_[83822]_  & \new_[83819]_ ;
  assign \new_[83824]_  = \new_[83823]_  & \new_[83816]_ ;
  assign \new_[83828]_  = ~A199 & ~A168;
  assign \new_[83829]_  = A169 & \new_[83828]_ ;
  assign \new_[83832]_  = ~A201 & A200;
  assign \new_[83835]_  = ~A203 & ~A202;
  assign \new_[83836]_  = \new_[83835]_  & \new_[83832]_ ;
  assign \new_[83837]_  = \new_[83836]_  & \new_[83829]_ ;
  assign \new_[83840]_  = ~A268 & A267;
  assign \new_[83843]_  = ~A298 & ~A269;
  assign \new_[83844]_  = \new_[83843]_  & \new_[83840]_ ;
  assign \new_[83847]_  = ~A300 & A299;
  assign \new_[83850]_  = ~A302 & ~A301;
  assign \new_[83851]_  = \new_[83850]_  & \new_[83847]_ ;
  assign \new_[83852]_  = \new_[83851]_  & \new_[83844]_ ;
  assign \new_[83856]_  = A199 & ~A168;
  assign \new_[83857]_  = A169 & \new_[83856]_ ;
  assign \new_[83860]_  = ~A201 & ~A200;
  assign \new_[83863]_  = ~A203 & ~A202;
  assign \new_[83864]_  = \new_[83863]_  & \new_[83860]_ ;
  assign \new_[83865]_  = \new_[83864]_  & \new_[83857]_ ;
  assign \new_[83868]_  = ~A268 & A267;
  assign \new_[83871]_  = A298 & ~A269;
  assign \new_[83872]_  = \new_[83871]_  & \new_[83868]_ ;
  assign \new_[83875]_  = ~A300 & ~A299;
  assign \new_[83878]_  = ~A302 & ~A301;
  assign \new_[83879]_  = \new_[83878]_  & \new_[83875]_ ;
  assign \new_[83880]_  = \new_[83879]_  & \new_[83872]_ ;
  assign \new_[83884]_  = A199 & ~A168;
  assign \new_[83885]_  = A169 & \new_[83884]_ ;
  assign \new_[83888]_  = ~A201 & ~A200;
  assign \new_[83891]_  = ~A203 & ~A202;
  assign \new_[83892]_  = \new_[83891]_  & \new_[83888]_ ;
  assign \new_[83893]_  = \new_[83892]_  & \new_[83885]_ ;
  assign \new_[83896]_  = ~A268 & A267;
  assign \new_[83899]_  = ~A298 & ~A269;
  assign \new_[83900]_  = \new_[83899]_  & \new_[83896]_ ;
  assign \new_[83903]_  = ~A300 & A299;
  assign \new_[83906]_  = ~A302 & ~A301;
  assign \new_[83907]_  = \new_[83906]_  & \new_[83903]_ ;
  assign \new_[83908]_  = \new_[83907]_  & \new_[83900]_ ;
  assign \new_[83912]_  = A168 & ~A169;
  assign \new_[83913]_  = A170 & \new_[83912]_ ;
  assign \new_[83916]_  = A200 & ~A199;
  assign \new_[83919]_  = A202 & A201;
  assign \new_[83920]_  = \new_[83919]_  & \new_[83916]_ ;
  assign \new_[83921]_  = \new_[83920]_  & \new_[83913]_ ;
  assign \new_[83924]_  = ~A268 & A267;
  assign \new_[83927]_  = A298 & ~A269;
  assign \new_[83928]_  = \new_[83927]_  & \new_[83924]_ ;
  assign \new_[83931]_  = ~A300 & ~A299;
  assign \new_[83934]_  = ~A302 & ~A301;
  assign \new_[83935]_  = \new_[83934]_  & \new_[83931]_ ;
  assign \new_[83936]_  = \new_[83935]_  & \new_[83928]_ ;
  assign \new_[83940]_  = A168 & ~A169;
  assign \new_[83941]_  = A170 & \new_[83940]_ ;
  assign \new_[83944]_  = A200 & ~A199;
  assign \new_[83947]_  = A202 & A201;
  assign \new_[83948]_  = \new_[83947]_  & \new_[83944]_ ;
  assign \new_[83949]_  = \new_[83948]_  & \new_[83941]_ ;
  assign \new_[83952]_  = ~A268 & A267;
  assign \new_[83955]_  = ~A298 & ~A269;
  assign \new_[83956]_  = \new_[83955]_  & \new_[83952]_ ;
  assign \new_[83959]_  = ~A300 & A299;
  assign \new_[83962]_  = ~A302 & ~A301;
  assign \new_[83963]_  = \new_[83962]_  & \new_[83959]_ ;
  assign \new_[83964]_  = \new_[83963]_  & \new_[83956]_ ;
  assign \new_[83968]_  = A168 & ~A169;
  assign \new_[83969]_  = A170 & \new_[83968]_ ;
  assign \new_[83972]_  = A200 & ~A199;
  assign \new_[83975]_  = A203 & A201;
  assign \new_[83976]_  = \new_[83975]_  & \new_[83972]_ ;
  assign \new_[83977]_  = \new_[83976]_  & \new_[83969]_ ;
  assign \new_[83980]_  = ~A268 & A267;
  assign \new_[83983]_  = A298 & ~A269;
  assign \new_[83984]_  = \new_[83983]_  & \new_[83980]_ ;
  assign \new_[83987]_  = ~A300 & ~A299;
  assign \new_[83990]_  = ~A302 & ~A301;
  assign \new_[83991]_  = \new_[83990]_  & \new_[83987]_ ;
  assign \new_[83992]_  = \new_[83991]_  & \new_[83984]_ ;
  assign \new_[83996]_  = A168 & ~A169;
  assign \new_[83997]_  = A170 & \new_[83996]_ ;
  assign \new_[84000]_  = A200 & ~A199;
  assign \new_[84003]_  = A203 & A201;
  assign \new_[84004]_  = \new_[84003]_  & \new_[84000]_ ;
  assign \new_[84005]_  = \new_[84004]_  & \new_[83997]_ ;
  assign \new_[84008]_  = ~A268 & A267;
  assign \new_[84011]_  = ~A298 & ~A269;
  assign \new_[84012]_  = \new_[84011]_  & \new_[84008]_ ;
  assign \new_[84015]_  = ~A300 & A299;
  assign \new_[84018]_  = ~A302 & ~A301;
  assign \new_[84019]_  = \new_[84018]_  & \new_[84015]_ ;
  assign \new_[84020]_  = \new_[84019]_  & \new_[84012]_ ;
  assign \new_[84024]_  = A168 & ~A169;
  assign \new_[84025]_  = A170 & \new_[84024]_ ;
  assign \new_[84028]_  = A200 & ~A199;
  assign \new_[84031]_  = ~A202 & ~A201;
  assign \new_[84032]_  = \new_[84031]_  & \new_[84028]_ ;
  assign \new_[84033]_  = \new_[84032]_  & \new_[84025]_ ;
  assign \new_[84036]_  = A267 & ~A203;
  assign \new_[84039]_  = ~A269 & ~A268;
  assign \new_[84040]_  = \new_[84039]_  & \new_[84036]_ ;
  assign \new_[84043]_  = ~A299 & A298;
  assign \new_[84046]_  = A301 & A300;
  assign \new_[84047]_  = \new_[84046]_  & \new_[84043]_ ;
  assign \new_[84048]_  = \new_[84047]_  & \new_[84040]_ ;
  assign \new_[84052]_  = A168 & ~A169;
  assign \new_[84053]_  = A170 & \new_[84052]_ ;
  assign \new_[84056]_  = A200 & ~A199;
  assign \new_[84059]_  = ~A202 & ~A201;
  assign \new_[84060]_  = \new_[84059]_  & \new_[84056]_ ;
  assign \new_[84061]_  = \new_[84060]_  & \new_[84053]_ ;
  assign \new_[84064]_  = A267 & ~A203;
  assign \new_[84067]_  = ~A269 & ~A268;
  assign \new_[84068]_  = \new_[84067]_  & \new_[84064]_ ;
  assign \new_[84071]_  = ~A299 & A298;
  assign \new_[84074]_  = A302 & A300;
  assign \new_[84075]_  = \new_[84074]_  & \new_[84071]_ ;
  assign \new_[84076]_  = \new_[84075]_  & \new_[84068]_ ;
  assign \new_[84080]_  = A168 & ~A169;
  assign \new_[84081]_  = A170 & \new_[84080]_ ;
  assign \new_[84084]_  = A200 & ~A199;
  assign \new_[84087]_  = ~A202 & ~A201;
  assign \new_[84088]_  = \new_[84087]_  & \new_[84084]_ ;
  assign \new_[84089]_  = \new_[84088]_  & \new_[84081]_ ;
  assign \new_[84092]_  = A267 & ~A203;
  assign \new_[84095]_  = ~A269 & ~A268;
  assign \new_[84096]_  = \new_[84095]_  & \new_[84092]_ ;
  assign \new_[84099]_  = A299 & ~A298;
  assign \new_[84102]_  = A301 & A300;
  assign \new_[84103]_  = \new_[84102]_  & \new_[84099]_ ;
  assign \new_[84104]_  = \new_[84103]_  & \new_[84096]_ ;
  assign \new_[84108]_  = A168 & ~A169;
  assign \new_[84109]_  = A170 & \new_[84108]_ ;
  assign \new_[84112]_  = A200 & ~A199;
  assign \new_[84115]_  = ~A202 & ~A201;
  assign \new_[84116]_  = \new_[84115]_  & \new_[84112]_ ;
  assign \new_[84117]_  = \new_[84116]_  & \new_[84109]_ ;
  assign \new_[84120]_  = A267 & ~A203;
  assign \new_[84123]_  = ~A269 & ~A268;
  assign \new_[84124]_  = \new_[84123]_  & \new_[84120]_ ;
  assign \new_[84127]_  = A299 & ~A298;
  assign \new_[84130]_  = A302 & A300;
  assign \new_[84131]_  = \new_[84130]_  & \new_[84127]_ ;
  assign \new_[84132]_  = \new_[84131]_  & \new_[84124]_ ;
  assign \new_[84136]_  = A168 & ~A169;
  assign \new_[84137]_  = A170 & \new_[84136]_ ;
  assign \new_[84140]_  = A200 & ~A199;
  assign \new_[84143]_  = ~A202 & ~A201;
  assign \new_[84144]_  = \new_[84143]_  & \new_[84140]_ ;
  assign \new_[84145]_  = \new_[84144]_  & \new_[84137]_ ;
  assign \new_[84148]_  = ~A267 & ~A203;
  assign \new_[84151]_  = A298 & A268;
  assign \new_[84152]_  = \new_[84151]_  & \new_[84148]_ ;
  assign \new_[84155]_  = ~A300 & ~A299;
  assign \new_[84158]_  = ~A302 & ~A301;
  assign \new_[84159]_  = \new_[84158]_  & \new_[84155]_ ;
  assign \new_[84160]_  = \new_[84159]_  & \new_[84152]_ ;
  assign \new_[84164]_  = A168 & ~A169;
  assign \new_[84165]_  = A170 & \new_[84164]_ ;
  assign \new_[84168]_  = A200 & ~A199;
  assign \new_[84171]_  = ~A202 & ~A201;
  assign \new_[84172]_  = \new_[84171]_  & \new_[84168]_ ;
  assign \new_[84173]_  = \new_[84172]_  & \new_[84165]_ ;
  assign \new_[84176]_  = ~A267 & ~A203;
  assign \new_[84179]_  = ~A298 & A268;
  assign \new_[84180]_  = \new_[84179]_  & \new_[84176]_ ;
  assign \new_[84183]_  = ~A300 & A299;
  assign \new_[84186]_  = ~A302 & ~A301;
  assign \new_[84187]_  = \new_[84186]_  & \new_[84183]_ ;
  assign \new_[84188]_  = \new_[84187]_  & \new_[84180]_ ;
  assign \new_[84192]_  = A168 & ~A169;
  assign \new_[84193]_  = A170 & \new_[84192]_ ;
  assign \new_[84196]_  = A200 & ~A199;
  assign \new_[84199]_  = ~A202 & ~A201;
  assign \new_[84200]_  = \new_[84199]_  & \new_[84196]_ ;
  assign \new_[84201]_  = \new_[84200]_  & \new_[84193]_ ;
  assign \new_[84204]_  = ~A267 & ~A203;
  assign \new_[84207]_  = A298 & A269;
  assign \new_[84208]_  = \new_[84207]_  & \new_[84204]_ ;
  assign \new_[84211]_  = ~A300 & ~A299;
  assign \new_[84214]_  = ~A302 & ~A301;
  assign \new_[84215]_  = \new_[84214]_  & \new_[84211]_ ;
  assign \new_[84216]_  = \new_[84215]_  & \new_[84208]_ ;
  assign \new_[84220]_  = A168 & ~A169;
  assign \new_[84221]_  = A170 & \new_[84220]_ ;
  assign \new_[84224]_  = A200 & ~A199;
  assign \new_[84227]_  = ~A202 & ~A201;
  assign \new_[84228]_  = \new_[84227]_  & \new_[84224]_ ;
  assign \new_[84229]_  = \new_[84228]_  & \new_[84221]_ ;
  assign \new_[84232]_  = ~A267 & ~A203;
  assign \new_[84235]_  = ~A298 & A269;
  assign \new_[84236]_  = \new_[84235]_  & \new_[84232]_ ;
  assign \new_[84239]_  = ~A300 & A299;
  assign \new_[84242]_  = ~A302 & ~A301;
  assign \new_[84243]_  = \new_[84242]_  & \new_[84239]_ ;
  assign \new_[84244]_  = \new_[84243]_  & \new_[84236]_ ;
  assign \new_[84248]_  = A168 & ~A169;
  assign \new_[84249]_  = A170 & \new_[84248]_ ;
  assign \new_[84252]_  = A200 & ~A199;
  assign \new_[84255]_  = ~A202 & ~A201;
  assign \new_[84256]_  = \new_[84255]_  & \new_[84252]_ ;
  assign \new_[84257]_  = \new_[84256]_  & \new_[84249]_ ;
  assign \new_[84260]_  = A265 & ~A203;
  assign \new_[84263]_  = A298 & A266;
  assign \new_[84264]_  = \new_[84263]_  & \new_[84260]_ ;
  assign \new_[84267]_  = ~A300 & ~A299;
  assign \new_[84270]_  = ~A302 & ~A301;
  assign \new_[84271]_  = \new_[84270]_  & \new_[84267]_ ;
  assign \new_[84272]_  = \new_[84271]_  & \new_[84264]_ ;
  assign \new_[84276]_  = A168 & ~A169;
  assign \new_[84277]_  = A170 & \new_[84276]_ ;
  assign \new_[84280]_  = A200 & ~A199;
  assign \new_[84283]_  = ~A202 & ~A201;
  assign \new_[84284]_  = \new_[84283]_  & \new_[84280]_ ;
  assign \new_[84285]_  = \new_[84284]_  & \new_[84277]_ ;
  assign \new_[84288]_  = A265 & ~A203;
  assign \new_[84291]_  = ~A298 & A266;
  assign \new_[84292]_  = \new_[84291]_  & \new_[84288]_ ;
  assign \new_[84295]_  = ~A300 & A299;
  assign \new_[84298]_  = ~A302 & ~A301;
  assign \new_[84299]_  = \new_[84298]_  & \new_[84295]_ ;
  assign \new_[84300]_  = \new_[84299]_  & \new_[84292]_ ;
  assign \new_[84304]_  = A168 & ~A169;
  assign \new_[84305]_  = A170 & \new_[84304]_ ;
  assign \new_[84308]_  = A200 & ~A199;
  assign \new_[84311]_  = ~A202 & ~A201;
  assign \new_[84312]_  = \new_[84311]_  & \new_[84308]_ ;
  assign \new_[84313]_  = \new_[84312]_  & \new_[84305]_ ;
  assign \new_[84316]_  = ~A265 & ~A203;
  assign \new_[84319]_  = A298 & ~A266;
  assign \new_[84320]_  = \new_[84319]_  & \new_[84316]_ ;
  assign \new_[84323]_  = ~A300 & ~A299;
  assign \new_[84326]_  = ~A302 & ~A301;
  assign \new_[84327]_  = \new_[84326]_  & \new_[84323]_ ;
  assign \new_[84328]_  = \new_[84327]_  & \new_[84320]_ ;
  assign \new_[84332]_  = A168 & ~A169;
  assign \new_[84333]_  = A170 & \new_[84332]_ ;
  assign \new_[84336]_  = A200 & ~A199;
  assign \new_[84339]_  = ~A202 & ~A201;
  assign \new_[84340]_  = \new_[84339]_  & \new_[84336]_ ;
  assign \new_[84341]_  = \new_[84340]_  & \new_[84333]_ ;
  assign \new_[84344]_  = ~A265 & ~A203;
  assign \new_[84347]_  = ~A298 & ~A266;
  assign \new_[84348]_  = \new_[84347]_  & \new_[84344]_ ;
  assign \new_[84351]_  = ~A300 & A299;
  assign \new_[84354]_  = ~A302 & ~A301;
  assign \new_[84355]_  = \new_[84354]_  & \new_[84351]_ ;
  assign \new_[84356]_  = \new_[84355]_  & \new_[84348]_ ;
  assign \new_[84360]_  = A168 & ~A169;
  assign \new_[84361]_  = A170 & \new_[84360]_ ;
  assign \new_[84364]_  = ~A200 & A199;
  assign \new_[84367]_  = A202 & A201;
  assign \new_[84368]_  = \new_[84367]_  & \new_[84364]_ ;
  assign \new_[84369]_  = \new_[84368]_  & \new_[84361]_ ;
  assign \new_[84372]_  = ~A268 & A267;
  assign \new_[84375]_  = A298 & ~A269;
  assign \new_[84376]_  = \new_[84375]_  & \new_[84372]_ ;
  assign \new_[84379]_  = ~A300 & ~A299;
  assign \new_[84382]_  = ~A302 & ~A301;
  assign \new_[84383]_  = \new_[84382]_  & \new_[84379]_ ;
  assign \new_[84384]_  = \new_[84383]_  & \new_[84376]_ ;
  assign \new_[84388]_  = A168 & ~A169;
  assign \new_[84389]_  = A170 & \new_[84388]_ ;
  assign \new_[84392]_  = ~A200 & A199;
  assign \new_[84395]_  = A202 & A201;
  assign \new_[84396]_  = \new_[84395]_  & \new_[84392]_ ;
  assign \new_[84397]_  = \new_[84396]_  & \new_[84389]_ ;
  assign \new_[84400]_  = ~A268 & A267;
  assign \new_[84403]_  = ~A298 & ~A269;
  assign \new_[84404]_  = \new_[84403]_  & \new_[84400]_ ;
  assign \new_[84407]_  = ~A300 & A299;
  assign \new_[84410]_  = ~A302 & ~A301;
  assign \new_[84411]_  = \new_[84410]_  & \new_[84407]_ ;
  assign \new_[84412]_  = \new_[84411]_  & \new_[84404]_ ;
  assign \new_[84416]_  = A168 & ~A169;
  assign \new_[84417]_  = A170 & \new_[84416]_ ;
  assign \new_[84420]_  = ~A200 & A199;
  assign \new_[84423]_  = A203 & A201;
  assign \new_[84424]_  = \new_[84423]_  & \new_[84420]_ ;
  assign \new_[84425]_  = \new_[84424]_  & \new_[84417]_ ;
  assign \new_[84428]_  = ~A268 & A267;
  assign \new_[84431]_  = A298 & ~A269;
  assign \new_[84432]_  = \new_[84431]_  & \new_[84428]_ ;
  assign \new_[84435]_  = ~A300 & ~A299;
  assign \new_[84438]_  = ~A302 & ~A301;
  assign \new_[84439]_  = \new_[84438]_  & \new_[84435]_ ;
  assign \new_[84440]_  = \new_[84439]_  & \new_[84432]_ ;
  assign \new_[84444]_  = A168 & ~A169;
  assign \new_[84445]_  = A170 & \new_[84444]_ ;
  assign \new_[84448]_  = ~A200 & A199;
  assign \new_[84451]_  = A203 & A201;
  assign \new_[84452]_  = \new_[84451]_  & \new_[84448]_ ;
  assign \new_[84453]_  = \new_[84452]_  & \new_[84445]_ ;
  assign \new_[84456]_  = ~A268 & A267;
  assign \new_[84459]_  = ~A298 & ~A269;
  assign \new_[84460]_  = \new_[84459]_  & \new_[84456]_ ;
  assign \new_[84463]_  = ~A300 & A299;
  assign \new_[84466]_  = ~A302 & ~A301;
  assign \new_[84467]_  = \new_[84466]_  & \new_[84463]_ ;
  assign \new_[84468]_  = \new_[84467]_  & \new_[84460]_ ;
  assign \new_[84472]_  = A168 & ~A169;
  assign \new_[84473]_  = A170 & \new_[84472]_ ;
  assign \new_[84476]_  = ~A200 & A199;
  assign \new_[84479]_  = ~A202 & ~A201;
  assign \new_[84480]_  = \new_[84479]_  & \new_[84476]_ ;
  assign \new_[84481]_  = \new_[84480]_  & \new_[84473]_ ;
  assign \new_[84484]_  = A267 & ~A203;
  assign \new_[84487]_  = ~A269 & ~A268;
  assign \new_[84488]_  = \new_[84487]_  & \new_[84484]_ ;
  assign \new_[84491]_  = ~A299 & A298;
  assign \new_[84494]_  = A301 & A300;
  assign \new_[84495]_  = \new_[84494]_  & \new_[84491]_ ;
  assign \new_[84496]_  = \new_[84495]_  & \new_[84488]_ ;
  assign \new_[84500]_  = A168 & ~A169;
  assign \new_[84501]_  = A170 & \new_[84500]_ ;
  assign \new_[84504]_  = ~A200 & A199;
  assign \new_[84507]_  = ~A202 & ~A201;
  assign \new_[84508]_  = \new_[84507]_  & \new_[84504]_ ;
  assign \new_[84509]_  = \new_[84508]_  & \new_[84501]_ ;
  assign \new_[84512]_  = A267 & ~A203;
  assign \new_[84515]_  = ~A269 & ~A268;
  assign \new_[84516]_  = \new_[84515]_  & \new_[84512]_ ;
  assign \new_[84519]_  = ~A299 & A298;
  assign \new_[84522]_  = A302 & A300;
  assign \new_[84523]_  = \new_[84522]_  & \new_[84519]_ ;
  assign \new_[84524]_  = \new_[84523]_  & \new_[84516]_ ;
  assign \new_[84528]_  = A168 & ~A169;
  assign \new_[84529]_  = A170 & \new_[84528]_ ;
  assign \new_[84532]_  = ~A200 & A199;
  assign \new_[84535]_  = ~A202 & ~A201;
  assign \new_[84536]_  = \new_[84535]_  & \new_[84532]_ ;
  assign \new_[84537]_  = \new_[84536]_  & \new_[84529]_ ;
  assign \new_[84540]_  = A267 & ~A203;
  assign \new_[84543]_  = ~A269 & ~A268;
  assign \new_[84544]_  = \new_[84543]_  & \new_[84540]_ ;
  assign \new_[84547]_  = A299 & ~A298;
  assign \new_[84550]_  = A301 & A300;
  assign \new_[84551]_  = \new_[84550]_  & \new_[84547]_ ;
  assign \new_[84552]_  = \new_[84551]_  & \new_[84544]_ ;
  assign \new_[84556]_  = A168 & ~A169;
  assign \new_[84557]_  = A170 & \new_[84556]_ ;
  assign \new_[84560]_  = ~A200 & A199;
  assign \new_[84563]_  = ~A202 & ~A201;
  assign \new_[84564]_  = \new_[84563]_  & \new_[84560]_ ;
  assign \new_[84565]_  = \new_[84564]_  & \new_[84557]_ ;
  assign \new_[84568]_  = A267 & ~A203;
  assign \new_[84571]_  = ~A269 & ~A268;
  assign \new_[84572]_  = \new_[84571]_  & \new_[84568]_ ;
  assign \new_[84575]_  = A299 & ~A298;
  assign \new_[84578]_  = A302 & A300;
  assign \new_[84579]_  = \new_[84578]_  & \new_[84575]_ ;
  assign \new_[84580]_  = \new_[84579]_  & \new_[84572]_ ;
  assign \new_[84584]_  = A168 & ~A169;
  assign \new_[84585]_  = A170 & \new_[84584]_ ;
  assign \new_[84588]_  = ~A200 & A199;
  assign \new_[84591]_  = ~A202 & ~A201;
  assign \new_[84592]_  = \new_[84591]_  & \new_[84588]_ ;
  assign \new_[84593]_  = \new_[84592]_  & \new_[84585]_ ;
  assign \new_[84596]_  = ~A267 & ~A203;
  assign \new_[84599]_  = A298 & A268;
  assign \new_[84600]_  = \new_[84599]_  & \new_[84596]_ ;
  assign \new_[84603]_  = ~A300 & ~A299;
  assign \new_[84606]_  = ~A302 & ~A301;
  assign \new_[84607]_  = \new_[84606]_  & \new_[84603]_ ;
  assign \new_[84608]_  = \new_[84607]_  & \new_[84600]_ ;
  assign \new_[84612]_  = A168 & ~A169;
  assign \new_[84613]_  = A170 & \new_[84612]_ ;
  assign \new_[84616]_  = ~A200 & A199;
  assign \new_[84619]_  = ~A202 & ~A201;
  assign \new_[84620]_  = \new_[84619]_  & \new_[84616]_ ;
  assign \new_[84621]_  = \new_[84620]_  & \new_[84613]_ ;
  assign \new_[84624]_  = ~A267 & ~A203;
  assign \new_[84627]_  = ~A298 & A268;
  assign \new_[84628]_  = \new_[84627]_  & \new_[84624]_ ;
  assign \new_[84631]_  = ~A300 & A299;
  assign \new_[84634]_  = ~A302 & ~A301;
  assign \new_[84635]_  = \new_[84634]_  & \new_[84631]_ ;
  assign \new_[84636]_  = \new_[84635]_  & \new_[84628]_ ;
  assign \new_[84640]_  = A168 & ~A169;
  assign \new_[84641]_  = A170 & \new_[84640]_ ;
  assign \new_[84644]_  = ~A200 & A199;
  assign \new_[84647]_  = ~A202 & ~A201;
  assign \new_[84648]_  = \new_[84647]_  & \new_[84644]_ ;
  assign \new_[84649]_  = \new_[84648]_  & \new_[84641]_ ;
  assign \new_[84652]_  = ~A267 & ~A203;
  assign \new_[84655]_  = A298 & A269;
  assign \new_[84656]_  = \new_[84655]_  & \new_[84652]_ ;
  assign \new_[84659]_  = ~A300 & ~A299;
  assign \new_[84662]_  = ~A302 & ~A301;
  assign \new_[84663]_  = \new_[84662]_  & \new_[84659]_ ;
  assign \new_[84664]_  = \new_[84663]_  & \new_[84656]_ ;
  assign \new_[84668]_  = A168 & ~A169;
  assign \new_[84669]_  = A170 & \new_[84668]_ ;
  assign \new_[84672]_  = ~A200 & A199;
  assign \new_[84675]_  = ~A202 & ~A201;
  assign \new_[84676]_  = \new_[84675]_  & \new_[84672]_ ;
  assign \new_[84677]_  = \new_[84676]_  & \new_[84669]_ ;
  assign \new_[84680]_  = ~A267 & ~A203;
  assign \new_[84683]_  = ~A298 & A269;
  assign \new_[84684]_  = \new_[84683]_  & \new_[84680]_ ;
  assign \new_[84687]_  = ~A300 & A299;
  assign \new_[84690]_  = ~A302 & ~A301;
  assign \new_[84691]_  = \new_[84690]_  & \new_[84687]_ ;
  assign \new_[84692]_  = \new_[84691]_  & \new_[84684]_ ;
  assign \new_[84696]_  = A168 & ~A169;
  assign \new_[84697]_  = A170 & \new_[84696]_ ;
  assign \new_[84700]_  = ~A200 & A199;
  assign \new_[84703]_  = ~A202 & ~A201;
  assign \new_[84704]_  = \new_[84703]_  & \new_[84700]_ ;
  assign \new_[84705]_  = \new_[84704]_  & \new_[84697]_ ;
  assign \new_[84708]_  = A265 & ~A203;
  assign \new_[84711]_  = A298 & A266;
  assign \new_[84712]_  = \new_[84711]_  & \new_[84708]_ ;
  assign \new_[84715]_  = ~A300 & ~A299;
  assign \new_[84718]_  = ~A302 & ~A301;
  assign \new_[84719]_  = \new_[84718]_  & \new_[84715]_ ;
  assign \new_[84720]_  = \new_[84719]_  & \new_[84712]_ ;
  assign \new_[84724]_  = A168 & ~A169;
  assign \new_[84725]_  = A170 & \new_[84724]_ ;
  assign \new_[84728]_  = ~A200 & A199;
  assign \new_[84731]_  = ~A202 & ~A201;
  assign \new_[84732]_  = \new_[84731]_  & \new_[84728]_ ;
  assign \new_[84733]_  = \new_[84732]_  & \new_[84725]_ ;
  assign \new_[84736]_  = A265 & ~A203;
  assign \new_[84739]_  = ~A298 & A266;
  assign \new_[84740]_  = \new_[84739]_  & \new_[84736]_ ;
  assign \new_[84743]_  = ~A300 & A299;
  assign \new_[84746]_  = ~A302 & ~A301;
  assign \new_[84747]_  = \new_[84746]_  & \new_[84743]_ ;
  assign \new_[84748]_  = \new_[84747]_  & \new_[84740]_ ;
  assign \new_[84752]_  = A168 & ~A169;
  assign \new_[84753]_  = A170 & \new_[84752]_ ;
  assign \new_[84756]_  = ~A200 & A199;
  assign \new_[84759]_  = ~A202 & ~A201;
  assign \new_[84760]_  = \new_[84759]_  & \new_[84756]_ ;
  assign \new_[84761]_  = \new_[84760]_  & \new_[84753]_ ;
  assign \new_[84764]_  = ~A265 & ~A203;
  assign \new_[84767]_  = A298 & ~A266;
  assign \new_[84768]_  = \new_[84767]_  & \new_[84764]_ ;
  assign \new_[84771]_  = ~A300 & ~A299;
  assign \new_[84774]_  = ~A302 & ~A301;
  assign \new_[84775]_  = \new_[84774]_  & \new_[84771]_ ;
  assign \new_[84776]_  = \new_[84775]_  & \new_[84768]_ ;
  assign \new_[84780]_  = A168 & ~A169;
  assign \new_[84781]_  = A170 & \new_[84780]_ ;
  assign \new_[84784]_  = ~A200 & A199;
  assign \new_[84787]_  = ~A202 & ~A201;
  assign \new_[84788]_  = \new_[84787]_  & \new_[84784]_ ;
  assign \new_[84789]_  = \new_[84788]_  & \new_[84781]_ ;
  assign \new_[84792]_  = ~A265 & ~A203;
  assign \new_[84795]_  = ~A298 & ~A266;
  assign \new_[84796]_  = \new_[84795]_  & \new_[84792]_ ;
  assign \new_[84799]_  = ~A300 & A299;
  assign \new_[84802]_  = ~A302 & ~A301;
  assign \new_[84803]_  = \new_[84802]_  & \new_[84799]_ ;
  assign \new_[84804]_  = \new_[84803]_  & \new_[84796]_ ;
  assign \new_[84808]_  = ~A168 & ~A169;
  assign \new_[84809]_  = A170 & \new_[84808]_ ;
  assign \new_[84812]_  = ~A166 & A167;
  assign \new_[84815]_  = ~A202 & A201;
  assign \new_[84816]_  = \new_[84815]_  & \new_[84812]_ ;
  assign \new_[84817]_  = \new_[84816]_  & \new_[84809]_ ;
  assign \new_[84820]_  = A267 & ~A203;
  assign \new_[84823]_  = ~A269 & ~A268;
  assign \new_[84824]_  = \new_[84823]_  & \new_[84820]_ ;
  assign \new_[84827]_  = ~A299 & A298;
  assign \new_[84830]_  = A301 & A300;
  assign \new_[84831]_  = \new_[84830]_  & \new_[84827]_ ;
  assign \new_[84832]_  = \new_[84831]_  & \new_[84824]_ ;
  assign \new_[84836]_  = ~A168 & ~A169;
  assign \new_[84837]_  = A170 & \new_[84836]_ ;
  assign \new_[84840]_  = ~A166 & A167;
  assign \new_[84843]_  = ~A202 & A201;
  assign \new_[84844]_  = \new_[84843]_  & \new_[84840]_ ;
  assign \new_[84845]_  = \new_[84844]_  & \new_[84837]_ ;
  assign \new_[84848]_  = A267 & ~A203;
  assign \new_[84851]_  = ~A269 & ~A268;
  assign \new_[84852]_  = \new_[84851]_  & \new_[84848]_ ;
  assign \new_[84855]_  = ~A299 & A298;
  assign \new_[84858]_  = A302 & A300;
  assign \new_[84859]_  = \new_[84858]_  & \new_[84855]_ ;
  assign \new_[84860]_  = \new_[84859]_  & \new_[84852]_ ;
  assign \new_[84864]_  = ~A168 & ~A169;
  assign \new_[84865]_  = A170 & \new_[84864]_ ;
  assign \new_[84868]_  = ~A166 & A167;
  assign \new_[84871]_  = ~A202 & A201;
  assign \new_[84872]_  = \new_[84871]_  & \new_[84868]_ ;
  assign \new_[84873]_  = \new_[84872]_  & \new_[84865]_ ;
  assign \new_[84876]_  = A267 & ~A203;
  assign \new_[84879]_  = ~A269 & ~A268;
  assign \new_[84880]_  = \new_[84879]_  & \new_[84876]_ ;
  assign \new_[84883]_  = A299 & ~A298;
  assign \new_[84886]_  = A301 & A300;
  assign \new_[84887]_  = \new_[84886]_  & \new_[84883]_ ;
  assign \new_[84888]_  = \new_[84887]_  & \new_[84880]_ ;
  assign \new_[84892]_  = ~A168 & ~A169;
  assign \new_[84893]_  = A170 & \new_[84892]_ ;
  assign \new_[84896]_  = ~A166 & A167;
  assign \new_[84899]_  = ~A202 & A201;
  assign \new_[84900]_  = \new_[84899]_  & \new_[84896]_ ;
  assign \new_[84901]_  = \new_[84900]_  & \new_[84893]_ ;
  assign \new_[84904]_  = A267 & ~A203;
  assign \new_[84907]_  = ~A269 & ~A268;
  assign \new_[84908]_  = \new_[84907]_  & \new_[84904]_ ;
  assign \new_[84911]_  = A299 & ~A298;
  assign \new_[84914]_  = A302 & A300;
  assign \new_[84915]_  = \new_[84914]_  & \new_[84911]_ ;
  assign \new_[84916]_  = \new_[84915]_  & \new_[84908]_ ;
  assign \new_[84920]_  = ~A168 & ~A169;
  assign \new_[84921]_  = A170 & \new_[84920]_ ;
  assign \new_[84924]_  = ~A166 & A167;
  assign \new_[84927]_  = ~A202 & A201;
  assign \new_[84928]_  = \new_[84927]_  & \new_[84924]_ ;
  assign \new_[84929]_  = \new_[84928]_  & \new_[84921]_ ;
  assign \new_[84932]_  = ~A267 & ~A203;
  assign \new_[84935]_  = A298 & A268;
  assign \new_[84936]_  = \new_[84935]_  & \new_[84932]_ ;
  assign \new_[84939]_  = ~A300 & ~A299;
  assign \new_[84942]_  = ~A302 & ~A301;
  assign \new_[84943]_  = \new_[84942]_  & \new_[84939]_ ;
  assign \new_[84944]_  = \new_[84943]_  & \new_[84936]_ ;
  assign \new_[84948]_  = ~A168 & ~A169;
  assign \new_[84949]_  = A170 & \new_[84948]_ ;
  assign \new_[84952]_  = ~A166 & A167;
  assign \new_[84955]_  = ~A202 & A201;
  assign \new_[84956]_  = \new_[84955]_  & \new_[84952]_ ;
  assign \new_[84957]_  = \new_[84956]_  & \new_[84949]_ ;
  assign \new_[84960]_  = ~A267 & ~A203;
  assign \new_[84963]_  = ~A298 & A268;
  assign \new_[84964]_  = \new_[84963]_  & \new_[84960]_ ;
  assign \new_[84967]_  = ~A300 & A299;
  assign \new_[84970]_  = ~A302 & ~A301;
  assign \new_[84971]_  = \new_[84970]_  & \new_[84967]_ ;
  assign \new_[84972]_  = \new_[84971]_  & \new_[84964]_ ;
  assign \new_[84976]_  = ~A168 & ~A169;
  assign \new_[84977]_  = A170 & \new_[84976]_ ;
  assign \new_[84980]_  = ~A166 & A167;
  assign \new_[84983]_  = ~A202 & A201;
  assign \new_[84984]_  = \new_[84983]_  & \new_[84980]_ ;
  assign \new_[84985]_  = \new_[84984]_  & \new_[84977]_ ;
  assign \new_[84988]_  = ~A267 & ~A203;
  assign \new_[84991]_  = A298 & A269;
  assign \new_[84992]_  = \new_[84991]_  & \new_[84988]_ ;
  assign \new_[84995]_  = ~A300 & ~A299;
  assign \new_[84998]_  = ~A302 & ~A301;
  assign \new_[84999]_  = \new_[84998]_  & \new_[84995]_ ;
  assign \new_[85000]_  = \new_[84999]_  & \new_[84992]_ ;
  assign \new_[85004]_  = ~A168 & ~A169;
  assign \new_[85005]_  = A170 & \new_[85004]_ ;
  assign \new_[85008]_  = ~A166 & A167;
  assign \new_[85011]_  = ~A202 & A201;
  assign \new_[85012]_  = \new_[85011]_  & \new_[85008]_ ;
  assign \new_[85013]_  = \new_[85012]_  & \new_[85005]_ ;
  assign \new_[85016]_  = ~A267 & ~A203;
  assign \new_[85019]_  = ~A298 & A269;
  assign \new_[85020]_  = \new_[85019]_  & \new_[85016]_ ;
  assign \new_[85023]_  = ~A300 & A299;
  assign \new_[85026]_  = ~A302 & ~A301;
  assign \new_[85027]_  = \new_[85026]_  & \new_[85023]_ ;
  assign \new_[85028]_  = \new_[85027]_  & \new_[85020]_ ;
  assign \new_[85032]_  = ~A168 & ~A169;
  assign \new_[85033]_  = A170 & \new_[85032]_ ;
  assign \new_[85036]_  = ~A166 & A167;
  assign \new_[85039]_  = ~A202 & A201;
  assign \new_[85040]_  = \new_[85039]_  & \new_[85036]_ ;
  assign \new_[85041]_  = \new_[85040]_  & \new_[85033]_ ;
  assign \new_[85044]_  = A265 & ~A203;
  assign \new_[85047]_  = A298 & A266;
  assign \new_[85048]_  = \new_[85047]_  & \new_[85044]_ ;
  assign \new_[85051]_  = ~A300 & ~A299;
  assign \new_[85054]_  = ~A302 & ~A301;
  assign \new_[85055]_  = \new_[85054]_  & \new_[85051]_ ;
  assign \new_[85056]_  = \new_[85055]_  & \new_[85048]_ ;
  assign \new_[85060]_  = ~A168 & ~A169;
  assign \new_[85061]_  = A170 & \new_[85060]_ ;
  assign \new_[85064]_  = ~A166 & A167;
  assign \new_[85067]_  = ~A202 & A201;
  assign \new_[85068]_  = \new_[85067]_  & \new_[85064]_ ;
  assign \new_[85069]_  = \new_[85068]_  & \new_[85061]_ ;
  assign \new_[85072]_  = A265 & ~A203;
  assign \new_[85075]_  = ~A298 & A266;
  assign \new_[85076]_  = \new_[85075]_  & \new_[85072]_ ;
  assign \new_[85079]_  = ~A300 & A299;
  assign \new_[85082]_  = ~A302 & ~A301;
  assign \new_[85083]_  = \new_[85082]_  & \new_[85079]_ ;
  assign \new_[85084]_  = \new_[85083]_  & \new_[85076]_ ;
  assign \new_[85088]_  = ~A168 & ~A169;
  assign \new_[85089]_  = A170 & \new_[85088]_ ;
  assign \new_[85092]_  = ~A166 & A167;
  assign \new_[85095]_  = ~A202 & A201;
  assign \new_[85096]_  = \new_[85095]_  & \new_[85092]_ ;
  assign \new_[85097]_  = \new_[85096]_  & \new_[85089]_ ;
  assign \new_[85100]_  = ~A265 & ~A203;
  assign \new_[85103]_  = A298 & ~A266;
  assign \new_[85104]_  = \new_[85103]_  & \new_[85100]_ ;
  assign \new_[85107]_  = ~A300 & ~A299;
  assign \new_[85110]_  = ~A302 & ~A301;
  assign \new_[85111]_  = \new_[85110]_  & \new_[85107]_ ;
  assign \new_[85112]_  = \new_[85111]_  & \new_[85104]_ ;
  assign \new_[85116]_  = ~A168 & ~A169;
  assign \new_[85117]_  = A170 & \new_[85116]_ ;
  assign \new_[85120]_  = ~A166 & A167;
  assign \new_[85123]_  = ~A202 & A201;
  assign \new_[85124]_  = \new_[85123]_  & \new_[85120]_ ;
  assign \new_[85125]_  = \new_[85124]_  & \new_[85117]_ ;
  assign \new_[85128]_  = ~A265 & ~A203;
  assign \new_[85131]_  = ~A298 & ~A266;
  assign \new_[85132]_  = \new_[85131]_  & \new_[85128]_ ;
  assign \new_[85135]_  = ~A300 & A299;
  assign \new_[85138]_  = ~A302 & ~A301;
  assign \new_[85139]_  = \new_[85138]_  & \new_[85135]_ ;
  assign \new_[85140]_  = \new_[85139]_  & \new_[85132]_ ;
  assign \new_[85144]_  = ~A168 & ~A169;
  assign \new_[85145]_  = A170 & \new_[85144]_ ;
  assign \new_[85148]_  = ~A166 & A167;
  assign \new_[85151]_  = A202 & ~A201;
  assign \new_[85152]_  = \new_[85151]_  & \new_[85148]_ ;
  assign \new_[85153]_  = \new_[85152]_  & \new_[85145]_ ;
  assign \new_[85156]_  = ~A268 & A267;
  assign \new_[85159]_  = A298 & ~A269;
  assign \new_[85160]_  = \new_[85159]_  & \new_[85156]_ ;
  assign \new_[85163]_  = ~A300 & ~A299;
  assign \new_[85166]_  = ~A302 & ~A301;
  assign \new_[85167]_  = \new_[85166]_  & \new_[85163]_ ;
  assign \new_[85168]_  = \new_[85167]_  & \new_[85160]_ ;
  assign \new_[85172]_  = ~A168 & ~A169;
  assign \new_[85173]_  = A170 & \new_[85172]_ ;
  assign \new_[85176]_  = ~A166 & A167;
  assign \new_[85179]_  = A202 & ~A201;
  assign \new_[85180]_  = \new_[85179]_  & \new_[85176]_ ;
  assign \new_[85181]_  = \new_[85180]_  & \new_[85173]_ ;
  assign \new_[85184]_  = ~A268 & A267;
  assign \new_[85187]_  = ~A298 & ~A269;
  assign \new_[85188]_  = \new_[85187]_  & \new_[85184]_ ;
  assign \new_[85191]_  = ~A300 & A299;
  assign \new_[85194]_  = ~A302 & ~A301;
  assign \new_[85195]_  = \new_[85194]_  & \new_[85191]_ ;
  assign \new_[85196]_  = \new_[85195]_  & \new_[85188]_ ;
  assign \new_[85200]_  = ~A168 & ~A169;
  assign \new_[85201]_  = A170 & \new_[85200]_ ;
  assign \new_[85204]_  = ~A166 & A167;
  assign \new_[85207]_  = A203 & ~A201;
  assign \new_[85208]_  = \new_[85207]_  & \new_[85204]_ ;
  assign \new_[85209]_  = \new_[85208]_  & \new_[85201]_ ;
  assign \new_[85212]_  = ~A268 & A267;
  assign \new_[85215]_  = A298 & ~A269;
  assign \new_[85216]_  = \new_[85215]_  & \new_[85212]_ ;
  assign \new_[85219]_  = ~A300 & ~A299;
  assign \new_[85222]_  = ~A302 & ~A301;
  assign \new_[85223]_  = \new_[85222]_  & \new_[85219]_ ;
  assign \new_[85224]_  = \new_[85223]_  & \new_[85216]_ ;
  assign \new_[85228]_  = ~A168 & ~A169;
  assign \new_[85229]_  = A170 & \new_[85228]_ ;
  assign \new_[85232]_  = ~A166 & A167;
  assign \new_[85235]_  = A203 & ~A201;
  assign \new_[85236]_  = \new_[85235]_  & \new_[85232]_ ;
  assign \new_[85237]_  = \new_[85236]_  & \new_[85229]_ ;
  assign \new_[85240]_  = ~A268 & A267;
  assign \new_[85243]_  = ~A298 & ~A269;
  assign \new_[85244]_  = \new_[85243]_  & \new_[85240]_ ;
  assign \new_[85247]_  = ~A300 & A299;
  assign \new_[85250]_  = ~A302 & ~A301;
  assign \new_[85251]_  = \new_[85250]_  & \new_[85247]_ ;
  assign \new_[85252]_  = \new_[85251]_  & \new_[85244]_ ;
  assign \new_[85256]_  = ~A168 & ~A169;
  assign \new_[85257]_  = A170 & \new_[85256]_ ;
  assign \new_[85260]_  = ~A166 & A167;
  assign \new_[85263]_  = A200 & A199;
  assign \new_[85264]_  = \new_[85263]_  & \new_[85260]_ ;
  assign \new_[85265]_  = \new_[85264]_  & \new_[85257]_ ;
  assign \new_[85268]_  = ~A268 & A267;
  assign \new_[85271]_  = A298 & ~A269;
  assign \new_[85272]_  = \new_[85271]_  & \new_[85268]_ ;
  assign \new_[85275]_  = ~A300 & ~A299;
  assign \new_[85278]_  = ~A302 & ~A301;
  assign \new_[85279]_  = \new_[85278]_  & \new_[85275]_ ;
  assign \new_[85280]_  = \new_[85279]_  & \new_[85272]_ ;
  assign \new_[85284]_  = ~A168 & ~A169;
  assign \new_[85285]_  = A170 & \new_[85284]_ ;
  assign \new_[85288]_  = ~A166 & A167;
  assign \new_[85291]_  = A200 & A199;
  assign \new_[85292]_  = \new_[85291]_  & \new_[85288]_ ;
  assign \new_[85293]_  = \new_[85292]_  & \new_[85285]_ ;
  assign \new_[85296]_  = ~A268 & A267;
  assign \new_[85299]_  = ~A298 & ~A269;
  assign \new_[85300]_  = \new_[85299]_  & \new_[85296]_ ;
  assign \new_[85303]_  = ~A300 & A299;
  assign \new_[85306]_  = ~A302 & ~A301;
  assign \new_[85307]_  = \new_[85306]_  & \new_[85303]_ ;
  assign \new_[85308]_  = \new_[85307]_  & \new_[85300]_ ;
  assign \new_[85312]_  = ~A168 & ~A169;
  assign \new_[85313]_  = A170 & \new_[85312]_ ;
  assign \new_[85316]_  = ~A166 & A167;
  assign \new_[85319]_  = A200 & ~A199;
  assign \new_[85320]_  = \new_[85319]_  & \new_[85316]_ ;
  assign \new_[85321]_  = \new_[85320]_  & \new_[85313]_ ;
  assign \new_[85324]_  = A202 & A201;
  assign \new_[85327]_  = A266 & ~A265;
  assign \new_[85328]_  = \new_[85327]_  & \new_[85324]_ ;
  assign \new_[85331]_  = A268 & A267;
  assign \new_[85334]_  = A301 & ~A300;
  assign \new_[85335]_  = \new_[85334]_  & \new_[85331]_ ;
  assign \new_[85336]_  = \new_[85335]_  & \new_[85328]_ ;
  assign \new_[85340]_  = ~A168 & ~A169;
  assign \new_[85341]_  = A170 & \new_[85340]_ ;
  assign \new_[85344]_  = ~A166 & A167;
  assign \new_[85347]_  = A200 & ~A199;
  assign \new_[85348]_  = \new_[85347]_  & \new_[85344]_ ;
  assign \new_[85349]_  = \new_[85348]_  & \new_[85341]_ ;
  assign \new_[85352]_  = A202 & A201;
  assign \new_[85355]_  = A266 & ~A265;
  assign \new_[85356]_  = \new_[85355]_  & \new_[85352]_ ;
  assign \new_[85359]_  = A268 & A267;
  assign \new_[85362]_  = A302 & ~A300;
  assign \new_[85363]_  = \new_[85362]_  & \new_[85359]_ ;
  assign \new_[85364]_  = \new_[85363]_  & \new_[85356]_ ;
  assign \new_[85368]_  = ~A168 & ~A169;
  assign \new_[85369]_  = A170 & \new_[85368]_ ;
  assign \new_[85372]_  = ~A166 & A167;
  assign \new_[85375]_  = A200 & ~A199;
  assign \new_[85376]_  = \new_[85375]_  & \new_[85372]_ ;
  assign \new_[85377]_  = \new_[85376]_  & \new_[85369]_ ;
  assign \new_[85380]_  = A202 & A201;
  assign \new_[85383]_  = A266 & ~A265;
  assign \new_[85384]_  = \new_[85383]_  & \new_[85380]_ ;
  assign \new_[85387]_  = A268 & A267;
  assign \new_[85390]_  = A299 & A298;
  assign \new_[85391]_  = \new_[85390]_  & \new_[85387]_ ;
  assign \new_[85392]_  = \new_[85391]_  & \new_[85384]_ ;
  assign \new_[85396]_  = ~A168 & ~A169;
  assign \new_[85397]_  = A170 & \new_[85396]_ ;
  assign \new_[85400]_  = ~A166 & A167;
  assign \new_[85403]_  = A200 & ~A199;
  assign \new_[85404]_  = \new_[85403]_  & \new_[85400]_ ;
  assign \new_[85405]_  = \new_[85404]_  & \new_[85397]_ ;
  assign \new_[85408]_  = A202 & A201;
  assign \new_[85411]_  = A266 & ~A265;
  assign \new_[85412]_  = \new_[85411]_  & \new_[85408]_ ;
  assign \new_[85415]_  = A268 & A267;
  assign \new_[85418]_  = ~A299 & ~A298;
  assign \new_[85419]_  = \new_[85418]_  & \new_[85415]_ ;
  assign \new_[85420]_  = \new_[85419]_  & \new_[85412]_ ;
  assign \new_[85424]_  = ~A168 & ~A169;
  assign \new_[85425]_  = A170 & \new_[85424]_ ;
  assign \new_[85428]_  = ~A166 & A167;
  assign \new_[85431]_  = A200 & ~A199;
  assign \new_[85432]_  = \new_[85431]_  & \new_[85428]_ ;
  assign \new_[85433]_  = \new_[85432]_  & \new_[85425]_ ;
  assign \new_[85436]_  = A202 & A201;
  assign \new_[85439]_  = A266 & ~A265;
  assign \new_[85440]_  = \new_[85439]_  & \new_[85436]_ ;
  assign \new_[85443]_  = A269 & A267;
  assign \new_[85446]_  = A301 & ~A300;
  assign \new_[85447]_  = \new_[85446]_  & \new_[85443]_ ;
  assign \new_[85448]_  = \new_[85447]_  & \new_[85440]_ ;
  assign \new_[85452]_  = ~A168 & ~A169;
  assign \new_[85453]_  = A170 & \new_[85452]_ ;
  assign \new_[85456]_  = ~A166 & A167;
  assign \new_[85459]_  = A200 & ~A199;
  assign \new_[85460]_  = \new_[85459]_  & \new_[85456]_ ;
  assign \new_[85461]_  = \new_[85460]_  & \new_[85453]_ ;
  assign \new_[85464]_  = A202 & A201;
  assign \new_[85467]_  = A266 & ~A265;
  assign \new_[85468]_  = \new_[85467]_  & \new_[85464]_ ;
  assign \new_[85471]_  = A269 & A267;
  assign \new_[85474]_  = A302 & ~A300;
  assign \new_[85475]_  = \new_[85474]_  & \new_[85471]_ ;
  assign \new_[85476]_  = \new_[85475]_  & \new_[85468]_ ;
  assign \new_[85480]_  = ~A168 & ~A169;
  assign \new_[85481]_  = A170 & \new_[85480]_ ;
  assign \new_[85484]_  = ~A166 & A167;
  assign \new_[85487]_  = A200 & ~A199;
  assign \new_[85488]_  = \new_[85487]_  & \new_[85484]_ ;
  assign \new_[85489]_  = \new_[85488]_  & \new_[85481]_ ;
  assign \new_[85492]_  = A202 & A201;
  assign \new_[85495]_  = A266 & ~A265;
  assign \new_[85496]_  = \new_[85495]_  & \new_[85492]_ ;
  assign \new_[85499]_  = A269 & A267;
  assign \new_[85502]_  = A299 & A298;
  assign \new_[85503]_  = \new_[85502]_  & \new_[85499]_ ;
  assign \new_[85504]_  = \new_[85503]_  & \new_[85496]_ ;
  assign \new_[85508]_  = ~A168 & ~A169;
  assign \new_[85509]_  = A170 & \new_[85508]_ ;
  assign \new_[85512]_  = ~A166 & A167;
  assign \new_[85515]_  = A200 & ~A199;
  assign \new_[85516]_  = \new_[85515]_  & \new_[85512]_ ;
  assign \new_[85517]_  = \new_[85516]_  & \new_[85509]_ ;
  assign \new_[85520]_  = A202 & A201;
  assign \new_[85523]_  = A266 & ~A265;
  assign \new_[85524]_  = \new_[85523]_  & \new_[85520]_ ;
  assign \new_[85527]_  = A269 & A267;
  assign \new_[85530]_  = ~A299 & ~A298;
  assign \new_[85531]_  = \new_[85530]_  & \new_[85527]_ ;
  assign \new_[85532]_  = \new_[85531]_  & \new_[85524]_ ;
  assign \new_[85536]_  = ~A168 & ~A169;
  assign \new_[85537]_  = A170 & \new_[85536]_ ;
  assign \new_[85540]_  = ~A166 & A167;
  assign \new_[85543]_  = A200 & ~A199;
  assign \new_[85544]_  = \new_[85543]_  & \new_[85540]_ ;
  assign \new_[85545]_  = \new_[85544]_  & \new_[85537]_ ;
  assign \new_[85548]_  = A202 & A201;
  assign \new_[85551]_  = ~A266 & A265;
  assign \new_[85552]_  = \new_[85551]_  & \new_[85548]_ ;
  assign \new_[85555]_  = A268 & A267;
  assign \new_[85558]_  = A301 & ~A300;
  assign \new_[85559]_  = \new_[85558]_  & \new_[85555]_ ;
  assign \new_[85560]_  = \new_[85559]_  & \new_[85552]_ ;
  assign \new_[85564]_  = ~A168 & ~A169;
  assign \new_[85565]_  = A170 & \new_[85564]_ ;
  assign \new_[85568]_  = ~A166 & A167;
  assign \new_[85571]_  = A200 & ~A199;
  assign \new_[85572]_  = \new_[85571]_  & \new_[85568]_ ;
  assign \new_[85573]_  = \new_[85572]_  & \new_[85565]_ ;
  assign \new_[85576]_  = A202 & A201;
  assign \new_[85579]_  = ~A266 & A265;
  assign \new_[85580]_  = \new_[85579]_  & \new_[85576]_ ;
  assign \new_[85583]_  = A268 & A267;
  assign \new_[85586]_  = A302 & ~A300;
  assign \new_[85587]_  = \new_[85586]_  & \new_[85583]_ ;
  assign \new_[85588]_  = \new_[85587]_  & \new_[85580]_ ;
  assign \new_[85592]_  = ~A168 & ~A169;
  assign \new_[85593]_  = A170 & \new_[85592]_ ;
  assign \new_[85596]_  = ~A166 & A167;
  assign \new_[85599]_  = A200 & ~A199;
  assign \new_[85600]_  = \new_[85599]_  & \new_[85596]_ ;
  assign \new_[85601]_  = \new_[85600]_  & \new_[85593]_ ;
  assign \new_[85604]_  = A202 & A201;
  assign \new_[85607]_  = ~A266 & A265;
  assign \new_[85608]_  = \new_[85607]_  & \new_[85604]_ ;
  assign \new_[85611]_  = A268 & A267;
  assign \new_[85614]_  = A299 & A298;
  assign \new_[85615]_  = \new_[85614]_  & \new_[85611]_ ;
  assign \new_[85616]_  = \new_[85615]_  & \new_[85608]_ ;
  assign \new_[85620]_  = ~A168 & ~A169;
  assign \new_[85621]_  = A170 & \new_[85620]_ ;
  assign \new_[85624]_  = ~A166 & A167;
  assign \new_[85627]_  = A200 & ~A199;
  assign \new_[85628]_  = \new_[85627]_  & \new_[85624]_ ;
  assign \new_[85629]_  = \new_[85628]_  & \new_[85621]_ ;
  assign \new_[85632]_  = A202 & A201;
  assign \new_[85635]_  = ~A266 & A265;
  assign \new_[85636]_  = \new_[85635]_  & \new_[85632]_ ;
  assign \new_[85639]_  = A268 & A267;
  assign \new_[85642]_  = ~A299 & ~A298;
  assign \new_[85643]_  = \new_[85642]_  & \new_[85639]_ ;
  assign \new_[85644]_  = \new_[85643]_  & \new_[85636]_ ;
  assign \new_[85648]_  = ~A168 & ~A169;
  assign \new_[85649]_  = A170 & \new_[85648]_ ;
  assign \new_[85652]_  = ~A166 & A167;
  assign \new_[85655]_  = A200 & ~A199;
  assign \new_[85656]_  = \new_[85655]_  & \new_[85652]_ ;
  assign \new_[85657]_  = \new_[85656]_  & \new_[85649]_ ;
  assign \new_[85660]_  = A202 & A201;
  assign \new_[85663]_  = ~A266 & A265;
  assign \new_[85664]_  = \new_[85663]_  & \new_[85660]_ ;
  assign \new_[85667]_  = A269 & A267;
  assign \new_[85670]_  = A301 & ~A300;
  assign \new_[85671]_  = \new_[85670]_  & \new_[85667]_ ;
  assign \new_[85672]_  = \new_[85671]_  & \new_[85664]_ ;
  assign \new_[85676]_  = ~A168 & ~A169;
  assign \new_[85677]_  = A170 & \new_[85676]_ ;
  assign \new_[85680]_  = ~A166 & A167;
  assign \new_[85683]_  = A200 & ~A199;
  assign \new_[85684]_  = \new_[85683]_  & \new_[85680]_ ;
  assign \new_[85685]_  = \new_[85684]_  & \new_[85677]_ ;
  assign \new_[85688]_  = A202 & A201;
  assign \new_[85691]_  = ~A266 & A265;
  assign \new_[85692]_  = \new_[85691]_  & \new_[85688]_ ;
  assign \new_[85695]_  = A269 & A267;
  assign \new_[85698]_  = A302 & ~A300;
  assign \new_[85699]_  = \new_[85698]_  & \new_[85695]_ ;
  assign \new_[85700]_  = \new_[85699]_  & \new_[85692]_ ;
  assign \new_[85704]_  = ~A168 & ~A169;
  assign \new_[85705]_  = A170 & \new_[85704]_ ;
  assign \new_[85708]_  = ~A166 & A167;
  assign \new_[85711]_  = A200 & ~A199;
  assign \new_[85712]_  = \new_[85711]_  & \new_[85708]_ ;
  assign \new_[85713]_  = \new_[85712]_  & \new_[85705]_ ;
  assign \new_[85716]_  = A202 & A201;
  assign \new_[85719]_  = ~A266 & A265;
  assign \new_[85720]_  = \new_[85719]_  & \new_[85716]_ ;
  assign \new_[85723]_  = A269 & A267;
  assign \new_[85726]_  = A299 & A298;
  assign \new_[85727]_  = \new_[85726]_  & \new_[85723]_ ;
  assign \new_[85728]_  = \new_[85727]_  & \new_[85720]_ ;
  assign \new_[85732]_  = ~A168 & ~A169;
  assign \new_[85733]_  = A170 & \new_[85732]_ ;
  assign \new_[85736]_  = ~A166 & A167;
  assign \new_[85739]_  = A200 & ~A199;
  assign \new_[85740]_  = \new_[85739]_  & \new_[85736]_ ;
  assign \new_[85741]_  = \new_[85740]_  & \new_[85733]_ ;
  assign \new_[85744]_  = A202 & A201;
  assign \new_[85747]_  = ~A266 & A265;
  assign \new_[85748]_  = \new_[85747]_  & \new_[85744]_ ;
  assign \new_[85751]_  = A269 & A267;
  assign \new_[85754]_  = ~A299 & ~A298;
  assign \new_[85755]_  = \new_[85754]_  & \new_[85751]_ ;
  assign \new_[85756]_  = \new_[85755]_  & \new_[85748]_ ;
  assign \new_[85760]_  = ~A168 & ~A169;
  assign \new_[85761]_  = A170 & \new_[85760]_ ;
  assign \new_[85764]_  = ~A166 & A167;
  assign \new_[85767]_  = A200 & ~A199;
  assign \new_[85768]_  = \new_[85767]_  & \new_[85764]_ ;
  assign \new_[85769]_  = \new_[85768]_  & \new_[85761]_ ;
  assign \new_[85772]_  = A203 & A201;
  assign \new_[85775]_  = A266 & ~A265;
  assign \new_[85776]_  = \new_[85775]_  & \new_[85772]_ ;
  assign \new_[85779]_  = A268 & A267;
  assign \new_[85782]_  = A301 & ~A300;
  assign \new_[85783]_  = \new_[85782]_  & \new_[85779]_ ;
  assign \new_[85784]_  = \new_[85783]_  & \new_[85776]_ ;
  assign \new_[85788]_  = ~A168 & ~A169;
  assign \new_[85789]_  = A170 & \new_[85788]_ ;
  assign \new_[85792]_  = ~A166 & A167;
  assign \new_[85795]_  = A200 & ~A199;
  assign \new_[85796]_  = \new_[85795]_  & \new_[85792]_ ;
  assign \new_[85797]_  = \new_[85796]_  & \new_[85789]_ ;
  assign \new_[85800]_  = A203 & A201;
  assign \new_[85803]_  = A266 & ~A265;
  assign \new_[85804]_  = \new_[85803]_  & \new_[85800]_ ;
  assign \new_[85807]_  = A268 & A267;
  assign \new_[85810]_  = A302 & ~A300;
  assign \new_[85811]_  = \new_[85810]_  & \new_[85807]_ ;
  assign \new_[85812]_  = \new_[85811]_  & \new_[85804]_ ;
  assign \new_[85816]_  = ~A168 & ~A169;
  assign \new_[85817]_  = A170 & \new_[85816]_ ;
  assign \new_[85820]_  = ~A166 & A167;
  assign \new_[85823]_  = A200 & ~A199;
  assign \new_[85824]_  = \new_[85823]_  & \new_[85820]_ ;
  assign \new_[85825]_  = \new_[85824]_  & \new_[85817]_ ;
  assign \new_[85828]_  = A203 & A201;
  assign \new_[85831]_  = A266 & ~A265;
  assign \new_[85832]_  = \new_[85831]_  & \new_[85828]_ ;
  assign \new_[85835]_  = A268 & A267;
  assign \new_[85838]_  = A299 & A298;
  assign \new_[85839]_  = \new_[85838]_  & \new_[85835]_ ;
  assign \new_[85840]_  = \new_[85839]_  & \new_[85832]_ ;
  assign \new_[85844]_  = ~A168 & ~A169;
  assign \new_[85845]_  = A170 & \new_[85844]_ ;
  assign \new_[85848]_  = ~A166 & A167;
  assign \new_[85851]_  = A200 & ~A199;
  assign \new_[85852]_  = \new_[85851]_  & \new_[85848]_ ;
  assign \new_[85853]_  = \new_[85852]_  & \new_[85845]_ ;
  assign \new_[85856]_  = A203 & A201;
  assign \new_[85859]_  = A266 & ~A265;
  assign \new_[85860]_  = \new_[85859]_  & \new_[85856]_ ;
  assign \new_[85863]_  = A268 & A267;
  assign \new_[85866]_  = ~A299 & ~A298;
  assign \new_[85867]_  = \new_[85866]_  & \new_[85863]_ ;
  assign \new_[85868]_  = \new_[85867]_  & \new_[85860]_ ;
  assign \new_[85872]_  = ~A168 & ~A169;
  assign \new_[85873]_  = A170 & \new_[85872]_ ;
  assign \new_[85876]_  = ~A166 & A167;
  assign \new_[85879]_  = A200 & ~A199;
  assign \new_[85880]_  = \new_[85879]_  & \new_[85876]_ ;
  assign \new_[85881]_  = \new_[85880]_  & \new_[85873]_ ;
  assign \new_[85884]_  = A203 & A201;
  assign \new_[85887]_  = A266 & ~A265;
  assign \new_[85888]_  = \new_[85887]_  & \new_[85884]_ ;
  assign \new_[85891]_  = A269 & A267;
  assign \new_[85894]_  = A301 & ~A300;
  assign \new_[85895]_  = \new_[85894]_  & \new_[85891]_ ;
  assign \new_[85896]_  = \new_[85895]_  & \new_[85888]_ ;
  assign \new_[85900]_  = ~A168 & ~A169;
  assign \new_[85901]_  = A170 & \new_[85900]_ ;
  assign \new_[85904]_  = ~A166 & A167;
  assign \new_[85907]_  = A200 & ~A199;
  assign \new_[85908]_  = \new_[85907]_  & \new_[85904]_ ;
  assign \new_[85909]_  = \new_[85908]_  & \new_[85901]_ ;
  assign \new_[85912]_  = A203 & A201;
  assign \new_[85915]_  = A266 & ~A265;
  assign \new_[85916]_  = \new_[85915]_  & \new_[85912]_ ;
  assign \new_[85919]_  = A269 & A267;
  assign \new_[85922]_  = A302 & ~A300;
  assign \new_[85923]_  = \new_[85922]_  & \new_[85919]_ ;
  assign \new_[85924]_  = \new_[85923]_  & \new_[85916]_ ;
  assign \new_[85928]_  = ~A168 & ~A169;
  assign \new_[85929]_  = A170 & \new_[85928]_ ;
  assign \new_[85932]_  = ~A166 & A167;
  assign \new_[85935]_  = A200 & ~A199;
  assign \new_[85936]_  = \new_[85935]_  & \new_[85932]_ ;
  assign \new_[85937]_  = \new_[85936]_  & \new_[85929]_ ;
  assign \new_[85940]_  = A203 & A201;
  assign \new_[85943]_  = A266 & ~A265;
  assign \new_[85944]_  = \new_[85943]_  & \new_[85940]_ ;
  assign \new_[85947]_  = A269 & A267;
  assign \new_[85950]_  = A299 & A298;
  assign \new_[85951]_  = \new_[85950]_  & \new_[85947]_ ;
  assign \new_[85952]_  = \new_[85951]_  & \new_[85944]_ ;
  assign \new_[85956]_  = ~A168 & ~A169;
  assign \new_[85957]_  = A170 & \new_[85956]_ ;
  assign \new_[85960]_  = ~A166 & A167;
  assign \new_[85963]_  = A200 & ~A199;
  assign \new_[85964]_  = \new_[85963]_  & \new_[85960]_ ;
  assign \new_[85965]_  = \new_[85964]_  & \new_[85957]_ ;
  assign \new_[85968]_  = A203 & A201;
  assign \new_[85971]_  = A266 & ~A265;
  assign \new_[85972]_  = \new_[85971]_  & \new_[85968]_ ;
  assign \new_[85975]_  = A269 & A267;
  assign \new_[85978]_  = ~A299 & ~A298;
  assign \new_[85979]_  = \new_[85978]_  & \new_[85975]_ ;
  assign \new_[85980]_  = \new_[85979]_  & \new_[85972]_ ;
  assign \new_[85984]_  = ~A168 & ~A169;
  assign \new_[85985]_  = A170 & \new_[85984]_ ;
  assign \new_[85988]_  = ~A166 & A167;
  assign \new_[85991]_  = A200 & ~A199;
  assign \new_[85992]_  = \new_[85991]_  & \new_[85988]_ ;
  assign \new_[85993]_  = \new_[85992]_  & \new_[85985]_ ;
  assign \new_[85996]_  = A203 & A201;
  assign \new_[85999]_  = ~A266 & A265;
  assign \new_[86000]_  = \new_[85999]_  & \new_[85996]_ ;
  assign \new_[86003]_  = A268 & A267;
  assign \new_[86006]_  = A301 & ~A300;
  assign \new_[86007]_  = \new_[86006]_  & \new_[86003]_ ;
  assign \new_[86008]_  = \new_[86007]_  & \new_[86000]_ ;
  assign \new_[86012]_  = ~A168 & ~A169;
  assign \new_[86013]_  = A170 & \new_[86012]_ ;
  assign \new_[86016]_  = ~A166 & A167;
  assign \new_[86019]_  = A200 & ~A199;
  assign \new_[86020]_  = \new_[86019]_  & \new_[86016]_ ;
  assign \new_[86021]_  = \new_[86020]_  & \new_[86013]_ ;
  assign \new_[86024]_  = A203 & A201;
  assign \new_[86027]_  = ~A266 & A265;
  assign \new_[86028]_  = \new_[86027]_  & \new_[86024]_ ;
  assign \new_[86031]_  = A268 & A267;
  assign \new_[86034]_  = A302 & ~A300;
  assign \new_[86035]_  = \new_[86034]_  & \new_[86031]_ ;
  assign \new_[86036]_  = \new_[86035]_  & \new_[86028]_ ;
  assign \new_[86040]_  = ~A168 & ~A169;
  assign \new_[86041]_  = A170 & \new_[86040]_ ;
  assign \new_[86044]_  = ~A166 & A167;
  assign \new_[86047]_  = A200 & ~A199;
  assign \new_[86048]_  = \new_[86047]_  & \new_[86044]_ ;
  assign \new_[86049]_  = \new_[86048]_  & \new_[86041]_ ;
  assign \new_[86052]_  = A203 & A201;
  assign \new_[86055]_  = ~A266 & A265;
  assign \new_[86056]_  = \new_[86055]_  & \new_[86052]_ ;
  assign \new_[86059]_  = A268 & A267;
  assign \new_[86062]_  = A299 & A298;
  assign \new_[86063]_  = \new_[86062]_  & \new_[86059]_ ;
  assign \new_[86064]_  = \new_[86063]_  & \new_[86056]_ ;
  assign \new_[86068]_  = ~A168 & ~A169;
  assign \new_[86069]_  = A170 & \new_[86068]_ ;
  assign \new_[86072]_  = ~A166 & A167;
  assign \new_[86075]_  = A200 & ~A199;
  assign \new_[86076]_  = \new_[86075]_  & \new_[86072]_ ;
  assign \new_[86077]_  = \new_[86076]_  & \new_[86069]_ ;
  assign \new_[86080]_  = A203 & A201;
  assign \new_[86083]_  = ~A266 & A265;
  assign \new_[86084]_  = \new_[86083]_  & \new_[86080]_ ;
  assign \new_[86087]_  = A268 & A267;
  assign \new_[86090]_  = ~A299 & ~A298;
  assign \new_[86091]_  = \new_[86090]_  & \new_[86087]_ ;
  assign \new_[86092]_  = \new_[86091]_  & \new_[86084]_ ;
  assign \new_[86096]_  = ~A168 & ~A169;
  assign \new_[86097]_  = A170 & \new_[86096]_ ;
  assign \new_[86100]_  = ~A166 & A167;
  assign \new_[86103]_  = A200 & ~A199;
  assign \new_[86104]_  = \new_[86103]_  & \new_[86100]_ ;
  assign \new_[86105]_  = \new_[86104]_  & \new_[86097]_ ;
  assign \new_[86108]_  = A203 & A201;
  assign \new_[86111]_  = ~A266 & A265;
  assign \new_[86112]_  = \new_[86111]_  & \new_[86108]_ ;
  assign \new_[86115]_  = A269 & A267;
  assign \new_[86118]_  = A301 & ~A300;
  assign \new_[86119]_  = \new_[86118]_  & \new_[86115]_ ;
  assign \new_[86120]_  = \new_[86119]_  & \new_[86112]_ ;
  assign \new_[86124]_  = ~A168 & ~A169;
  assign \new_[86125]_  = A170 & \new_[86124]_ ;
  assign \new_[86128]_  = ~A166 & A167;
  assign \new_[86131]_  = A200 & ~A199;
  assign \new_[86132]_  = \new_[86131]_  & \new_[86128]_ ;
  assign \new_[86133]_  = \new_[86132]_  & \new_[86125]_ ;
  assign \new_[86136]_  = A203 & A201;
  assign \new_[86139]_  = ~A266 & A265;
  assign \new_[86140]_  = \new_[86139]_  & \new_[86136]_ ;
  assign \new_[86143]_  = A269 & A267;
  assign \new_[86146]_  = A302 & ~A300;
  assign \new_[86147]_  = \new_[86146]_  & \new_[86143]_ ;
  assign \new_[86148]_  = \new_[86147]_  & \new_[86140]_ ;
  assign \new_[86152]_  = ~A168 & ~A169;
  assign \new_[86153]_  = A170 & \new_[86152]_ ;
  assign \new_[86156]_  = ~A166 & A167;
  assign \new_[86159]_  = A200 & ~A199;
  assign \new_[86160]_  = \new_[86159]_  & \new_[86156]_ ;
  assign \new_[86161]_  = \new_[86160]_  & \new_[86153]_ ;
  assign \new_[86164]_  = A203 & A201;
  assign \new_[86167]_  = ~A266 & A265;
  assign \new_[86168]_  = \new_[86167]_  & \new_[86164]_ ;
  assign \new_[86171]_  = A269 & A267;
  assign \new_[86174]_  = A299 & A298;
  assign \new_[86175]_  = \new_[86174]_  & \new_[86171]_ ;
  assign \new_[86176]_  = \new_[86175]_  & \new_[86168]_ ;
  assign \new_[86180]_  = ~A168 & ~A169;
  assign \new_[86181]_  = A170 & \new_[86180]_ ;
  assign \new_[86184]_  = ~A166 & A167;
  assign \new_[86187]_  = A200 & ~A199;
  assign \new_[86188]_  = \new_[86187]_  & \new_[86184]_ ;
  assign \new_[86189]_  = \new_[86188]_  & \new_[86181]_ ;
  assign \new_[86192]_  = A203 & A201;
  assign \new_[86195]_  = ~A266 & A265;
  assign \new_[86196]_  = \new_[86195]_  & \new_[86192]_ ;
  assign \new_[86199]_  = A269 & A267;
  assign \new_[86202]_  = ~A299 & ~A298;
  assign \new_[86203]_  = \new_[86202]_  & \new_[86199]_ ;
  assign \new_[86204]_  = \new_[86203]_  & \new_[86196]_ ;
  assign \new_[86208]_  = ~A168 & ~A169;
  assign \new_[86209]_  = A170 & \new_[86208]_ ;
  assign \new_[86212]_  = ~A166 & A167;
  assign \new_[86215]_  = ~A200 & A199;
  assign \new_[86216]_  = \new_[86215]_  & \new_[86212]_ ;
  assign \new_[86217]_  = \new_[86216]_  & \new_[86209]_ ;
  assign \new_[86220]_  = A202 & A201;
  assign \new_[86223]_  = A266 & ~A265;
  assign \new_[86224]_  = \new_[86223]_  & \new_[86220]_ ;
  assign \new_[86227]_  = A268 & A267;
  assign \new_[86230]_  = A301 & ~A300;
  assign \new_[86231]_  = \new_[86230]_  & \new_[86227]_ ;
  assign \new_[86232]_  = \new_[86231]_  & \new_[86224]_ ;
  assign \new_[86236]_  = ~A168 & ~A169;
  assign \new_[86237]_  = A170 & \new_[86236]_ ;
  assign \new_[86240]_  = ~A166 & A167;
  assign \new_[86243]_  = ~A200 & A199;
  assign \new_[86244]_  = \new_[86243]_  & \new_[86240]_ ;
  assign \new_[86245]_  = \new_[86244]_  & \new_[86237]_ ;
  assign \new_[86248]_  = A202 & A201;
  assign \new_[86251]_  = A266 & ~A265;
  assign \new_[86252]_  = \new_[86251]_  & \new_[86248]_ ;
  assign \new_[86255]_  = A268 & A267;
  assign \new_[86258]_  = A302 & ~A300;
  assign \new_[86259]_  = \new_[86258]_  & \new_[86255]_ ;
  assign \new_[86260]_  = \new_[86259]_  & \new_[86252]_ ;
  assign \new_[86264]_  = ~A168 & ~A169;
  assign \new_[86265]_  = A170 & \new_[86264]_ ;
  assign \new_[86268]_  = ~A166 & A167;
  assign \new_[86271]_  = ~A200 & A199;
  assign \new_[86272]_  = \new_[86271]_  & \new_[86268]_ ;
  assign \new_[86273]_  = \new_[86272]_  & \new_[86265]_ ;
  assign \new_[86276]_  = A202 & A201;
  assign \new_[86279]_  = A266 & ~A265;
  assign \new_[86280]_  = \new_[86279]_  & \new_[86276]_ ;
  assign \new_[86283]_  = A268 & A267;
  assign \new_[86286]_  = A299 & A298;
  assign \new_[86287]_  = \new_[86286]_  & \new_[86283]_ ;
  assign \new_[86288]_  = \new_[86287]_  & \new_[86280]_ ;
  assign \new_[86292]_  = ~A168 & ~A169;
  assign \new_[86293]_  = A170 & \new_[86292]_ ;
  assign \new_[86296]_  = ~A166 & A167;
  assign \new_[86299]_  = ~A200 & A199;
  assign \new_[86300]_  = \new_[86299]_  & \new_[86296]_ ;
  assign \new_[86301]_  = \new_[86300]_  & \new_[86293]_ ;
  assign \new_[86304]_  = A202 & A201;
  assign \new_[86307]_  = A266 & ~A265;
  assign \new_[86308]_  = \new_[86307]_  & \new_[86304]_ ;
  assign \new_[86311]_  = A268 & A267;
  assign \new_[86314]_  = ~A299 & ~A298;
  assign \new_[86315]_  = \new_[86314]_  & \new_[86311]_ ;
  assign \new_[86316]_  = \new_[86315]_  & \new_[86308]_ ;
  assign \new_[86320]_  = ~A168 & ~A169;
  assign \new_[86321]_  = A170 & \new_[86320]_ ;
  assign \new_[86324]_  = ~A166 & A167;
  assign \new_[86327]_  = ~A200 & A199;
  assign \new_[86328]_  = \new_[86327]_  & \new_[86324]_ ;
  assign \new_[86329]_  = \new_[86328]_  & \new_[86321]_ ;
  assign \new_[86332]_  = A202 & A201;
  assign \new_[86335]_  = A266 & ~A265;
  assign \new_[86336]_  = \new_[86335]_  & \new_[86332]_ ;
  assign \new_[86339]_  = A269 & A267;
  assign \new_[86342]_  = A301 & ~A300;
  assign \new_[86343]_  = \new_[86342]_  & \new_[86339]_ ;
  assign \new_[86344]_  = \new_[86343]_  & \new_[86336]_ ;
  assign \new_[86348]_  = ~A168 & ~A169;
  assign \new_[86349]_  = A170 & \new_[86348]_ ;
  assign \new_[86352]_  = ~A166 & A167;
  assign \new_[86355]_  = ~A200 & A199;
  assign \new_[86356]_  = \new_[86355]_  & \new_[86352]_ ;
  assign \new_[86357]_  = \new_[86356]_  & \new_[86349]_ ;
  assign \new_[86360]_  = A202 & A201;
  assign \new_[86363]_  = A266 & ~A265;
  assign \new_[86364]_  = \new_[86363]_  & \new_[86360]_ ;
  assign \new_[86367]_  = A269 & A267;
  assign \new_[86370]_  = A302 & ~A300;
  assign \new_[86371]_  = \new_[86370]_  & \new_[86367]_ ;
  assign \new_[86372]_  = \new_[86371]_  & \new_[86364]_ ;
  assign \new_[86376]_  = ~A168 & ~A169;
  assign \new_[86377]_  = A170 & \new_[86376]_ ;
  assign \new_[86380]_  = ~A166 & A167;
  assign \new_[86383]_  = ~A200 & A199;
  assign \new_[86384]_  = \new_[86383]_  & \new_[86380]_ ;
  assign \new_[86385]_  = \new_[86384]_  & \new_[86377]_ ;
  assign \new_[86388]_  = A202 & A201;
  assign \new_[86391]_  = A266 & ~A265;
  assign \new_[86392]_  = \new_[86391]_  & \new_[86388]_ ;
  assign \new_[86395]_  = A269 & A267;
  assign \new_[86398]_  = A299 & A298;
  assign \new_[86399]_  = \new_[86398]_  & \new_[86395]_ ;
  assign \new_[86400]_  = \new_[86399]_  & \new_[86392]_ ;
  assign \new_[86404]_  = ~A168 & ~A169;
  assign \new_[86405]_  = A170 & \new_[86404]_ ;
  assign \new_[86408]_  = ~A166 & A167;
  assign \new_[86411]_  = ~A200 & A199;
  assign \new_[86412]_  = \new_[86411]_  & \new_[86408]_ ;
  assign \new_[86413]_  = \new_[86412]_  & \new_[86405]_ ;
  assign \new_[86416]_  = A202 & A201;
  assign \new_[86419]_  = A266 & ~A265;
  assign \new_[86420]_  = \new_[86419]_  & \new_[86416]_ ;
  assign \new_[86423]_  = A269 & A267;
  assign \new_[86426]_  = ~A299 & ~A298;
  assign \new_[86427]_  = \new_[86426]_  & \new_[86423]_ ;
  assign \new_[86428]_  = \new_[86427]_  & \new_[86420]_ ;
  assign \new_[86432]_  = ~A168 & ~A169;
  assign \new_[86433]_  = A170 & \new_[86432]_ ;
  assign \new_[86436]_  = ~A166 & A167;
  assign \new_[86439]_  = ~A200 & A199;
  assign \new_[86440]_  = \new_[86439]_  & \new_[86436]_ ;
  assign \new_[86441]_  = \new_[86440]_  & \new_[86433]_ ;
  assign \new_[86444]_  = A202 & A201;
  assign \new_[86447]_  = ~A266 & A265;
  assign \new_[86448]_  = \new_[86447]_  & \new_[86444]_ ;
  assign \new_[86451]_  = A268 & A267;
  assign \new_[86454]_  = A301 & ~A300;
  assign \new_[86455]_  = \new_[86454]_  & \new_[86451]_ ;
  assign \new_[86456]_  = \new_[86455]_  & \new_[86448]_ ;
  assign \new_[86460]_  = ~A168 & ~A169;
  assign \new_[86461]_  = A170 & \new_[86460]_ ;
  assign \new_[86464]_  = ~A166 & A167;
  assign \new_[86467]_  = ~A200 & A199;
  assign \new_[86468]_  = \new_[86467]_  & \new_[86464]_ ;
  assign \new_[86469]_  = \new_[86468]_  & \new_[86461]_ ;
  assign \new_[86472]_  = A202 & A201;
  assign \new_[86475]_  = ~A266 & A265;
  assign \new_[86476]_  = \new_[86475]_  & \new_[86472]_ ;
  assign \new_[86479]_  = A268 & A267;
  assign \new_[86482]_  = A302 & ~A300;
  assign \new_[86483]_  = \new_[86482]_  & \new_[86479]_ ;
  assign \new_[86484]_  = \new_[86483]_  & \new_[86476]_ ;
  assign \new_[86488]_  = ~A168 & ~A169;
  assign \new_[86489]_  = A170 & \new_[86488]_ ;
  assign \new_[86492]_  = ~A166 & A167;
  assign \new_[86495]_  = ~A200 & A199;
  assign \new_[86496]_  = \new_[86495]_  & \new_[86492]_ ;
  assign \new_[86497]_  = \new_[86496]_  & \new_[86489]_ ;
  assign \new_[86500]_  = A202 & A201;
  assign \new_[86503]_  = ~A266 & A265;
  assign \new_[86504]_  = \new_[86503]_  & \new_[86500]_ ;
  assign \new_[86507]_  = A268 & A267;
  assign \new_[86510]_  = A299 & A298;
  assign \new_[86511]_  = \new_[86510]_  & \new_[86507]_ ;
  assign \new_[86512]_  = \new_[86511]_  & \new_[86504]_ ;
  assign \new_[86516]_  = ~A168 & ~A169;
  assign \new_[86517]_  = A170 & \new_[86516]_ ;
  assign \new_[86520]_  = ~A166 & A167;
  assign \new_[86523]_  = ~A200 & A199;
  assign \new_[86524]_  = \new_[86523]_  & \new_[86520]_ ;
  assign \new_[86525]_  = \new_[86524]_  & \new_[86517]_ ;
  assign \new_[86528]_  = A202 & A201;
  assign \new_[86531]_  = ~A266 & A265;
  assign \new_[86532]_  = \new_[86531]_  & \new_[86528]_ ;
  assign \new_[86535]_  = A268 & A267;
  assign \new_[86538]_  = ~A299 & ~A298;
  assign \new_[86539]_  = \new_[86538]_  & \new_[86535]_ ;
  assign \new_[86540]_  = \new_[86539]_  & \new_[86532]_ ;
  assign \new_[86544]_  = ~A168 & ~A169;
  assign \new_[86545]_  = A170 & \new_[86544]_ ;
  assign \new_[86548]_  = ~A166 & A167;
  assign \new_[86551]_  = ~A200 & A199;
  assign \new_[86552]_  = \new_[86551]_  & \new_[86548]_ ;
  assign \new_[86553]_  = \new_[86552]_  & \new_[86545]_ ;
  assign \new_[86556]_  = A202 & A201;
  assign \new_[86559]_  = ~A266 & A265;
  assign \new_[86560]_  = \new_[86559]_  & \new_[86556]_ ;
  assign \new_[86563]_  = A269 & A267;
  assign \new_[86566]_  = A301 & ~A300;
  assign \new_[86567]_  = \new_[86566]_  & \new_[86563]_ ;
  assign \new_[86568]_  = \new_[86567]_  & \new_[86560]_ ;
  assign \new_[86572]_  = ~A168 & ~A169;
  assign \new_[86573]_  = A170 & \new_[86572]_ ;
  assign \new_[86576]_  = ~A166 & A167;
  assign \new_[86579]_  = ~A200 & A199;
  assign \new_[86580]_  = \new_[86579]_  & \new_[86576]_ ;
  assign \new_[86581]_  = \new_[86580]_  & \new_[86573]_ ;
  assign \new_[86584]_  = A202 & A201;
  assign \new_[86587]_  = ~A266 & A265;
  assign \new_[86588]_  = \new_[86587]_  & \new_[86584]_ ;
  assign \new_[86591]_  = A269 & A267;
  assign \new_[86594]_  = A302 & ~A300;
  assign \new_[86595]_  = \new_[86594]_  & \new_[86591]_ ;
  assign \new_[86596]_  = \new_[86595]_  & \new_[86588]_ ;
  assign \new_[86600]_  = ~A168 & ~A169;
  assign \new_[86601]_  = A170 & \new_[86600]_ ;
  assign \new_[86604]_  = ~A166 & A167;
  assign \new_[86607]_  = ~A200 & A199;
  assign \new_[86608]_  = \new_[86607]_  & \new_[86604]_ ;
  assign \new_[86609]_  = \new_[86608]_  & \new_[86601]_ ;
  assign \new_[86612]_  = A202 & A201;
  assign \new_[86615]_  = ~A266 & A265;
  assign \new_[86616]_  = \new_[86615]_  & \new_[86612]_ ;
  assign \new_[86619]_  = A269 & A267;
  assign \new_[86622]_  = A299 & A298;
  assign \new_[86623]_  = \new_[86622]_  & \new_[86619]_ ;
  assign \new_[86624]_  = \new_[86623]_  & \new_[86616]_ ;
  assign \new_[86628]_  = ~A168 & ~A169;
  assign \new_[86629]_  = A170 & \new_[86628]_ ;
  assign \new_[86632]_  = ~A166 & A167;
  assign \new_[86635]_  = ~A200 & A199;
  assign \new_[86636]_  = \new_[86635]_  & \new_[86632]_ ;
  assign \new_[86637]_  = \new_[86636]_  & \new_[86629]_ ;
  assign \new_[86640]_  = A202 & A201;
  assign \new_[86643]_  = ~A266 & A265;
  assign \new_[86644]_  = \new_[86643]_  & \new_[86640]_ ;
  assign \new_[86647]_  = A269 & A267;
  assign \new_[86650]_  = ~A299 & ~A298;
  assign \new_[86651]_  = \new_[86650]_  & \new_[86647]_ ;
  assign \new_[86652]_  = \new_[86651]_  & \new_[86644]_ ;
  assign \new_[86656]_  = ~A168 & ~A169;
  assign \new_[86657]_  = A170 & \new_[86656]_ ;
  assign \new_[86660]_  = ~A166 & A167;
  assign \new_[86663]_  = ~A200 & A199;
  assign \new_[86664]_  = \new_[86663]_  & \new_[86660]_ ;
  assign \new_[86665]_  = \new_[86664]_  & \new_[86657]_ ;
  assign \new_[86668]_  = A203 & A201;
  assign \new_[86671]_  = A266 & ~A265;
  assign \new_[86672]_  = \new_[86671]_  & \new_[86668]_ ;
  assign \new_[86675]_  = A268 & A267;
  assign \new_[86678]_  = A301 & ~A300;
  assign \new_[86679]_  = \new_[86678]_  & \new_[86675]_ ;
  assign \new_[86680]_  = \new_[86679]_  & \new_[86672]_ ;
  assign \new_[86684]_  = ~A168 & ~A169;
  assign \new_[86685]_  = A170 & \new_[86684]_ ;
  assign \new_[86688]_  = ~A166 & A167;
  assign \new_[86691]_  = ~A200 & A199;
  assign \new_[86692]_  = \new_[86691]_  & \new_[86688]_ ;
  assign \new_[86693]_  = \new_[86692]_  & \new_[86685]_ ;
  assign \new_[86696]_  = A203 & A201;
  assign \new_[86699]_  = A266 & ~A265;
  assign \new_[86700]_  = \new_[86699]_  & \new_[86696]_ ;
  assign \new_[86703]_  = A268 & A267;
  assign \new_[86706]_  = A302 & ~A300;
  assign \new_[86707]_  = \new_[86706]_  & \new_[86703]_ ;
  assign \new_[86708]_  = \new_[86707]_  & \new_[86700]_ ;
  assign \new_[86712]_  = ~A168 & ~A169;
  assign \new_[86713]_  = A170 & \new_[86712]_ ;
  assign \new_[86716]_  = ~A166 & A167;
  assign \new_[86719]_  = ~A200 & A199;
  assign \new_[86720]_  = \new_[86719]_  & \new_[86716]_ ;
  assign \new_[86721]_  = \new_[86720]_  & \new_[86713]_ ;
  assign \new_[86724]_  = A203 & A201;
  assign \new_[86727]_  = A266 & ~A265;
  assign \new_[86728]_  = \new_[86727]_  & \new_[86724]_ ;
  assign \new_[86731]_  = A268 & A267;
  assign \new_[86734]_  = A299 & A298;
  assign \new_[86735]_  = \new_[86734]_  & \new_[86731]_ ;
  assign \new_[86736]_  = \new_[86735]_  & \new_[86728]_ ;
  assign \new_[86740]_  = ~A168 & ~A169;
  assign \new_[86741]_  = A170 & \new_[86740]_ ;
  assign \new_[86744]_  = ~A166 & A167;
  assign \new_[86747]_  = ~A200 & A199;
  assign \new_[86748]_  = \new_[86747]_  & \new_[86744]_ ;
  assign \new_[86749]_  = \new_[86748]_  & \new_[86741]_ ;
  assign \new_[86752]_  = A203 & A201;
  assign \new_[86755]_  = A266 & ~A265;
  assign \new_[86756]_  = \new_[86755]_  & \new_[86752]_ ;
  assign \new_[86759]_  = A268 & A267;
  assign \new_[86762]_  = ~A299 & ~A298;
  assign \new_[86763]_  = \new_[86762]_  & \new_[86759]_ ;
  assign \new_[86764]_  = \new_[86763]_  & \new_[86756]_ ;
  assign \new_[86768]_  = ~A168 & ~A169;
  assign \new_[86769]_  = A170 & \new_[86768]_ ;
  assign \new_[86772]_  = ~A166 & A167;
  assign \new_[86775]_  = ~A200 & A199;
  assign \new_[86776]_  = \new_[86775]_  & \new_[86772]_ ;
  assign \new_[86777]_  = \new_[86776]_  & \new_[86769]_ ;
  assign \new_[86780]_  = A203 & A201;
  assign \new_[86783]_  = A266 & ~A265;
  assign \new_[86784]_  = \new_[86783]_  & \new_[86780]_ ;
  assign \new_[86787]_  = A269 & A267;
  assign \new_[86790]_  = A301 & ~A300;
  assign \new_[86791]_  = \new_[86790]_  & \new_[86787]_ ;
  assign \new_[86792]_  = \new_[86791]_  & \new_[86784]_ ;
  assign \new_[86796]_  = ~A168 & ~A169;
  assign \new_[86797]_  = A170 & \new_[86796]_ ;
  assign \new_[86800]_  = ~A166 & A167;
  assign \new_[86803]_  = ~A200 & A199;
  assign \new_[86804]_  = \new_[86803]_  & \new_[86800]_ ;
  assign \new_[86805]_  = \new_[86804]_  & \new_[86797]_ ;
  assign \new_[86808]_  = A203 & A201;
  assign \new_[86811]_  = A266 & ~A265;
  assign \new_[86812]_  = \new_[86811]_  & \new_[86808]_ ;
  assign \new_[86815]_  = A269 & A267;
  assign \new_[86818]_  = A302 & ~A300;
  assign \new_[86819]_  = \new_[86818]_  & \new_[86815]_ ;
  assign \new_[86820]_  = \new_[86819]_  & \new_[86812]_ ;
  assign \new_[86824]_  = ~A168 & ~A169;
  assign \new_[86825]_  = A170 & \new_[86824]_ ;
  assign \new_[86828]_  = ~A166 & A167;
  assign \new_[86831]_  = ~A200 & A199;
  assign \new_[86832]_  = \new_[86831]_  & \new_[86828]_ ;
  assign \new_[86833]_  = \new_[86832]_  & \new_[86825]_ ;
  assign \new_[86836]_  = A203 & A201;
  assign \new_[86839]_  = A266 & ~A265;
  assign \new_[86840]_  = \new_[86839]_  & \new_[86836]_ ;
  assign \new_[86843]_  = A269 & A267;
  assign \new_[86846]_  = A299 & A298;
  assign \new_[86847]_  = \new_[86846]_  & \new_[86843]_ ;
  assign \new_[86848]_  = \new_[86847]_  & \new_[86840]_ ;
  assign \new_[86852]_  = ~A168 & ~A169;
  assign \new_[86853]_  = A170 & \new_[86852]_ ;
  assign \new_[86856]_  = ~A166 & A167;
  assign \new_[86859]_  = ~A200 & A199;
  assign \new_[86860]_  = \new_[86859]_  & \new_[86856]_ ;
  assign \new_[86861]_  = \new_[86860]_  & \new_[86853]_ ;
  assign \new_[86864]_  = A203 & A201;
  assign \new_[86867]_  = A266 & ~A265;
  assign \new_[86868]_  = \new_[86867]_  & \new_[86864]_ ;
  assign \new_[86871]_  = A269 & A267;
  assign \new_[86874]_  = ~A299 & ~A298;
  assign \new_[86875]_  = \new_[86874]_  & \new_[86871]_ ;
  assign \new_[86876]_  = \new_[86875]_  & \new_[86868]_ ;
  assign \new_[86880]_  = ~A168 & ~A169;
  assign \new_[86881]_  = A170 & \new_[86880]_ ;
  assign \new_[86884]_  = ~A166 & A167;
  assign \new_[86887]_  = ~A200 & A199;
  assign \new_[86888]_  = \new_[86887]_  & \new_[86884]_ ;
  assign \new_[86889]_  = \new_[86888]_  & \new_[86881]_ ;
  assign \new_[86892]_  = A203 & A201;
  assign \new_[86895]_  = ~A266 & A265;
  assign \new_[86896]_  = \new_[86895]_  & \new_[86892]_ ;
  assign \new_[86899]_  = A268 & A267;
  assign \new_[86902]_  = A301 & ~A300;
  assign \new_[86903]_  = \new_[86902]_  & \new_[86899]_ ;
  assign \new_[86904]_  = \new_[86903]_  & \new_[86896]_ ;
  assign \new_[86908]_  = ~A168 & ~A169;
  assign \new_[86909]_  = A170 & \new_[86908]_ ;
  assign \new_[86912]_  = ~A166 & A167;
  assign \new_[86915]_  = ~A200 & A199;
  assign \new_[86916]_  = \new_[86915]_  & \new_[86912]_ ;
  assign \new_[86917]_  = \new_[86916]_  & \new_[86909]_ ;
  assign \new_[86920]_  = A203 & A201;
  assign \new_[86923]_  = ~A266 & A265;
  assign \new_[86924]_  = \new_[86923]_  & \new_[86920]_ ;
  assign \new_[86927]_  = A268 & A267;
  assign \new_[86930]_  = A302 & ~A300;
  assign \new_[86931]_  = \new_[86930]_  & \new_[86927]_ ;
  assign \new_[86932]_  = \new_[86931]_  & \new_[86924]_ ;
  assign \new_[86936]_  = ~A168 & ~A169;
  assign \new_[86937]_  = A170 & \new_[86936]_ ;
  assign \new_[86940]_  = ~A166 & A167;
  assign \new_[86943]_  = ~A200 & A199;
  assign \new_[86944]_  = \new_[86943]_  & \new_[86940]_ ;
  assign \new_[86945]_  = \new_[86944]_  & \new_[86937]_ ;
  assign \new_[86948]_  = A203 & A201;
  assign \new_[86951]_  = ~A266 & A265;
  assign \new_[86952]_  = \new_[86951]_  & \new_[86948]_ ;
  assign \new_[86955]_  = A268 & A267;
  assign \new_[86958]_  = A299 & A298;
  assign \new_[86959]_  = \new_[86958]_  & \new_[86955]_ ;
  assign \new_[86960]_  = \new_[86959]_  & \new_[86952]_ ;
  assign \new_[86964]_  = ~A168 & ~A169;
  assign \new_[86965]_  = A170 & \new_[86964]_ ;
  assign \new_[86968]_  = ~A166 & A167;
  assign \new_[86971]_  = ~A200 & A199;
  assign \new_[86972]_  = \new_[86971]_  & \new_[86968]_ ;
  assign \new_[86973]_  = \new_[86972]_  & \new_[86965]_ ;
  assign \new_[86976]_  = A203 & A201;
  assign \new_[86979]_  = ~A266 & A265;
  assign \new_[86980]_  = \new_[86979]_  & \new_[86976]_ ;
  assign \new_[86983]_  = A268 & A267;
  assign \new_[86986]_  = ~A299 & ~A298;
  assign \new_[86987]_  = \new_[86986]_  & \new_[86983]_ ;
  assign \new_[86988]_  = \new_[86987]_  & \new_[86980]_ ;
  assign \new_[86992]_  = ~A168 & ~A169;
  assign \new_[86993]_  = A170 & \new_[86992]_ ;
  assign \new_[86996]_  = ~A166 & A167;
  assign \new_[86999]_  = ~A200 & A199;
  assign \new_[87000]_  = \new_[86999]_  & \new_[86996]_ ;
  assign \new_[87001]_  = \new_[87000]_  & \new_[86993]_ ;
  assign \new_[87004]_  = A203 & A201;
  assign \new_[87007]_  = ~A266 & A265;
  assign \new_[87008]_  = \new_[87007]_  & \new_[87004]_ ;
  assign \new_[87011]_  = A269 & A267;
  assign \new_[87014]_  = A301 & ~A300;
  assign \new_[87015]_  = \new_[87014]_  & \new_[87011]_ ;
  assign \new_[87016]_  = \new_[87015]_  & \new_[87008]_ ;
  assign \new_[87020]_  = ~A168 & ~A169;
  assign \new_[87021]_  = A170 & \new_[87020]_ ;
  assign \new_[87024]_  = ~A166 & A167;
  assign \new_[87027]_  = ~A200 & A199;
  assign \new_[87028]_  = \new_[87027]_  & \new_[87024]_ ;
  assign \new_[87029]_  = \new_[87028]_  & \new_[87021]_ ;
  assign \new_[87032]_  = A203 & A201;
  assign \new_[87035]_  = ~A266 & A265;
  assign \new_[87036]_  = \new_[87035]_  & \new_[87032]_ ;
  assign \new_[87039]_  = A269 & A267;
  assign \new_[87042]_  = A302 & ~A300;
  assign \new_[87043]_  = \new_[87042]_  & \new_[87039]_ ;
  assign \new_[87044]_  = \new_[87043]_  & \new_[87036]_ ;
  assign \new_[87048]_  = ~A168 & ~A169;
  assign \new_[87049]_  = A170 & \new_[87048]_ ;
  assign \new_[87052]_  = ~A166 & A167;
  assign \new_[87055]_  = ~A200 & A199;
  assign \new_[87056]_  = \new_[87055]_  & \new_[87052]_ ;
  assign \new_[87057]_  = \new_[87056]_  & \new_[87049]_ ;
  assign \new_[87060]_  = A203 & A201;
  assign \new_[87063]_  = ~A266 & A265;
  assign \new_[87064]_  = \new_[87063]_  & \new_[87060]_ ;
  assign \new_[87067]_  = A269 & A267;
  assign \new_[87070]_  = A299 & A298;
  assign \new_[87071]_  = \new_[87070]_  & \new_[87067]_ ;
  assign \new_[87072]_  = \new_[87071]_  & \new_[87064]_ ;
  assign \new_[87076]_  = ~A168 & ~A169;
  assign \new_[87077]_  = A170 & \new_[87076]_ ;
  assign \new_[87080]_  = ~A166 & A167;
  assign \new_[87083]_  = ~A200 & A199;
  assign \new_[87084]_  = \new_[87083]_  & \new_[87080]_ ;
  assign \new_[87085]_  = \new_[87084]_  & \new_[87077]_ ;
  assign \new_[87088]_  = A203 & A201;
  assign \new_[87091]_  = ~A266 & A265;
  assign \new_[87092]_  = \new_[87091]_  & \new_[87088]_ ;
  assign \new_[87095]_  = A269 & A267;
  assign \new_[87098]_  = ~A299 & ~A298;
  assign \new_[87099]_  = \new_[87098]_  & \new_[87095]_ ;
  assign \new_[87100]_  = \new_[87099]_  & \new_[87092]_ ;
  assign \new_[87104]_  = ~A168 & ~A169;
  assign \new_[87105]_  = A170 & \new_[87104]_ ;
  assign \new_[87108]_  = ~A166 & A167;
  assign \new_[87111]_  = ~A200 & ~A199;
  assign \new_[87112]_  = \new_[87111]_  & \new_[87108]_ ;
  assign \new_[87113]_  = \new_[87112]_  & \new_[87105]_ ;
  assign \new_[87116]_  = ~A268 & A267;
  assign \new_[87119]_  = A298 & ~A269;
  assign \new_[87120]_  = \new_[87119]_  & \new_[87116]_ ;
  assign \new_[87123]_  = ~A300 & ~A299;
  assign \new_[87126]_  = ~A302 & ~A301;
  assign \new_[87127]_  = \new_[87126]_  & \new_[87123]_ ;
  assign \new_[87128]_  = \new_[87127]_  & \new_[87120]_ ;
  assign \new_[87132]_  = ~A168 & ~A169;
  assign \new_[87133]_  = A170 & \new_[87132]_ ;
  assign \new_[87136]_  = ~A166 & A167;
  assign \new_[87139]_  = ~A200 & ~A199;
  assign \new_[87140]_  = \new_[87139]_  & \new_[87136]_ ;
  assign \new_[87141]_  = \new_[87140]_  & \new_[87133]_ ;
  assign \new_[87144]_  = ~A268 & A267;
  assign \new_[87147]_  = ~A298 & ~A269;
  assign \new_[87148]_  = \new_[87147]_  & \new_[87144]_ ;
  assign \new_[87151]_  = ~A300 & A299;
  assign \new_[87154]_  = ~A302 & ~A301;
  assign \new_[87155]_  = \new_[87154]_  & \new_[87151]_ ;
  assign \new_[87156]_  = \new_[87155]_  & \new_[87148]_ ;
  assign \new_[87160]_  = ~A168 & ~A169;
  assign \new_[87161]_  = A170 & \new_[87160]_ ;
  assign \new_[87164]_  = A166 & ~A167;
  assign \new_[87167]_  = ~A202 & A201;
  assign \new_[87168]_  = \new_[87167]_  & \new_[87164]_ ;
  assign \new_[87169]_  = \new_[87168]_  & \new_[87161]_ ;
  assign \new_[87172]_  = A267 & ~A203;
  assign \new_[87175]_  = ~A269 & ~A268;
  assign \new_[87176]_  = \new_[87175]_  & \new_[87172]_ ;
  assign \new_[87179]_  = ~A299 & A298;
  assign \new_[87182]_  = A301 & A300;
  assign \new_[87183]_  = \new_[87182]_  & \new_[87179]_ ;
  assign \new_[87184]_  = \new_[87183]_  & \new_[87176]_ ;
  assign \new_[87188]_  = ~A168 & ~A169;
  assign \new_[87189]_  = A170 & \new_[87188]_ ;
  assign \new_[87192]_  = A166 & ~A167;
  assign \new_[87195]_  = ~A202 & A201;
  assign \new_[87196]_  = \new_[87195]_  & \new_[87192]_ ;
  assign \new_[87197]_  = \new_[87196]_  & \new_[87189]_ ;
  assign \new_[87200]_  = A267 & ~A203;
  assign \new_[87203]_  = ~A269 & ~A268;
  assign \new_[87204]_  = \new_[87203]_  & \new_[87200]_ ;
  assign \new_[87207]_  = ~A299 & A298;
  assign \new_[87210]_  = A302 & A300;
  assign \new_[87211]_  = \new_[87210]_  & \new_[87207]_ ;
  assign \new_[87212]_  = \new_[87211]_  & \new_[87204]_ ;
  assign \new_[87216]_  = ~A168 & ~A169;
  assign \new_[87217]_  = A170 & \new_[87216]_ ;
  assign \new_[87220]_  = A166 & ~A167;
  assign \new_[87223]_  = ~A202 & A201;
  assign \new_[87224]_  = \new_[87223]_  & \new_[87220]_ ;
  assign \new_[87225]_  = \new_[87224]_  & \new_[87217]_ ;
  assign \new_[87228]_  = A267 & ~A203;
  assign \new_[87231]_  = ~A269 & ~A268;
  assign \new_[87232]_  = \new_[87231]_  & \new_[87228]_ ;
  assign \new_[87235]_  = A299 & ~A298;
  assign \new_[87238]_  = A301 & A300;
  assign \new_[87239]_  = \new_[87238]_  & \new_[87235]_ ;
  assign \new_[87240]_  = \new_[87239]_  & \new_[87232]_ ;
  assign \new_[87244]_  = ~A168 & ~A169;
  assign \new_[87245]_  = A170 & \new_[87244]_ ;
  assign \new_[87248]_  = A166 & ~A167;
  assign \new_[87251]_  = ~A202 & A201;
  assign \new_[87252]_  = \new_[87251]_  & \new_[87248]_ ;
  assign \new_[87253]_  = \new_[87252]_  & \new_[87245]_ ;
  assign \new_[87256]_  = A267 & ~A203;
  assign \new_[87259]_  = ~A269 & ~A268;
  assign \new_[87260]_  = \new_[87259]_  & \new_[87256]_ ;
  assign \new_[87263]_  = A299 & ~A298;
  assign \new_[87266]_  = A302 & A300;
  assign \new_[87267]_  = \new_[87266]_  & \new_[87263]_ ;
  assign \new_[87268]_  = \new_[87267]_  & \new_[87260]_ ;
  assign \new_[87272]_  = ~A168 & ~A169;
  assign \new_[87273]_  = A170 & \new_[87272]_ ;
  assign \new_[87276]_  = A166 & ~A167;
  assign \new_[87279]_  = ~A202 & A201;
  assign \new_[87280]_  = \new_[87279]_  & \new_[87276]_ ;
  assign \new_[87281]_  = \new_[87280]_  & \new_[87273]_ ;
  assign \new_[87284]_  = ~A267 & ~A203;
  assign \new_[87287]_  = A298 & A268;
  assign \new_[87288]_  = \new_[87287]_  & \new_[87284]_ ;
  assign \new_[87291]_  = ~A300 & ~A299;
  assign \new_[87294]_  = ~A302 & ~A301;
  assign \new_[87295]_  = \new_[87294]_  & \new_[87291]_ ;
  assign \new_[87296]_  = \new_[87295]_  & \new_[87288]_ ;
  assign \new_[87300]_  = ~A168 & ~A169;
  assign \new_[87301]_  = A170 & \new_[87300]_ ;
  assign \new_[87304]_  = A166 & ~A167;
  assign \new_[87307]_  = ~A202 & A201;
  assign \new_[87308]_  = \new_[87307]_  & \new_[87304]_ ;
  assign \new_[87309]_  = \new_[87308]_  & \new_[87301]_ ;
  assign \new_[87312]_  = ~A267 & ~A203;
  assign \new_[87315]_  = ~A298 & A268;
  assign \new_[87316]_  = \new_[87315]_  & \new_[87312]_ ;
  assign \new_[87319]_  = ~A300 & A299;
  assign \new_[87322]_  = ~A302 & ~A301;
  assign \new_[87323]_  = \new_[87322]_  & \new_[87319]_ ;
  assign \new_[87324]_  = \new_[87323]_  & \new_[87316]_ ;
  assign \new_[87328]_  = ~A168 & ~A169;
  assign \new_[87329]_  = A170 & \new_[87328]_ ;
  assign \new_[87332]_  = A166 & ~A167;
  assign \new_[87335]_  = ~A202 & A201;
  assign \new_[87336]_  = \new_[87335]_  & \new_[87332]_ ;
  assign \new_[87337]_  = \new_[87336]_  & \new_[87329]_ ;
  assign \new_[87340]_  = ~A267 & ~A203;
  assign \new_[87343]_  = A298 & A269;
  assign \new_[87344]_  = \new_[87343]_  & \new_[87340]_ ;
  assign \new_[87347]_  = ~A300 & ~A299;
  assign \new_[87350]_  = ~A302 & ~A301;
  assign \new_[87351]_  = \new_[87350]_  & \new_[87347]_ ;
  assign \new_[87352]_  = \new_[87351]_  & \new_[87344]_ ;
  assign \new_[87356]_  = ~A168 & ~A169;
  assign \new_[87357]_  = A170 & \new_[87356]_ ;
  assign \new_[87360]_  = A166 & ~A167;
  assign \new_[87363]_  = ~A202 & A201;
  assign \new_[87364]_  = \new_[87363]_  & \new_[87360]_ ;
  assign \new_[87365]_  = \new_[87364]_  & \new_[87357]_ ;
  assign \new_[87368]_  = ~A267 & ~A203;
  assign \new_[87371]_  = ~A298 & A269;
  assign \new_[87372]_  = \new_[87371]_  & \new_[87368]_ ;
  assign \new_[87375]_  = ~A300 & A299;
  assign \new_[87378]_  = ~A302 & ~A301;
  assign \new_[87379]_  = \new_[87378]_  & \new_[87375]_ ;
  assign \new_[87380]_  = \new_[87379]_  & \new_[87372]_ ;
  assign \new_[87384]_  = ~A168 & ~A169;
  assign \new_[87385]_  = A170 & \new_[87384]_ ;
  assign \new_[87388]_  = A166 & ~A167;
  assign \new_[87391]_  = ~A202 & A201;
  assign \new_[87392]_  = \new_[87391]_  & \new_[87388]_ ;
  assign \new_[87393]_  = \new_[87392]_  & \new_[87385]_ ;
  assign \new_[87396]_  = A265 & ~A203;
  assign \new_[87399]_  = A298 & A266;
  assign \new_[87400]_  = \new_[87399]_  & \new_[87396]_ ;
  assign \new_[87403]_  = ~A300 & ~A299;
  assign \new_[87406]_  = ~A302 & ~A301;
  assign \new_[87407]_  = \new_[87406]_  & \new_[87403]_ ;
  assign \new_[87408]_  = \new_[87407]_  & \new_[87400]_ ;
  assign \new_[87412]_  = ~A168 & ~A169;
  assign \new_[87413]_  = A170 & \new_[87412]_ ;
  assign \new_[87416]_  = A166 & ~A167;
  assign \new_[87419]_  = ~A202 & A201;
  assign \new_[87420]_  = \new_[87419]_  & \new_[87416]_ ;
  assign \new_[87421]_  = \new_[87420]_  & \new_[87413]_ ;
  assign \new_[87424]_  = A265 & ~A203;
  assign \new_[87427]_  = ~A298 & A266;
  assign \new_[87428]_  = \new_[87427]_  & \new_[87424]_ ;
  assign \new_[87431]_  = ~A300 & A299;
  assign \new_[87434]_  = ~A302 & ~A301;
  assign \new_[87435]_  = \new_[87434]_  & \new_[87431]_ ;
  assign \new_[87436]_  = \new_[87435]_  & \new_[87428]_ ;
  assign \new_[87440]_  = ~A168 & ~A169;
  assign \new_[87441]_  = A170 & \new_[87440]_ ;
  assign \new_[87444]_  = A166 & ~A167;
  assign \new_[87447]_  = ~A202 & A201;
  assign \new_[87448]_  = \new_[87447]_  & \new_[87444]_ ;
  assign \new_[87449]_  = \new_[87448]_  & \new_[87441]_ ;
  assign \new_[87452]_  = ~A265 & ~A203;
  assign \new_[87455]_  = A298 & ~A266;
  assign \new_[87456]_  = \new_[87455]_  & \new_[87452]_ ;
  assign \new_[87459]_  = ~A300 & ~A299;
  assign \new_[87462]_  = ~A302 & ~A301;
  assign \new_[87463]_  = \new_[87462]_  & \new_[87459]_ ;
  assign \new_[87464]_  = \new_[87463]_  & \new_[87456]_ ;
  assign \new_[87468]_  = ~A168 & ~A169;
  assign \new_[87469]_  = A170 & \new_[87468]_ ;
  assign \new_[87472]_  = A166 & ~A167;
  assign \new_[87475]_  = ~A202 & A201;
  assign \new_[87476]_  = \new_[87475]_  & \new_[87472]_ ;
  assign \new_[87477]_  = \new_[87476]_  & \new_[87469]_ ;
  assign \new_[87480]_  = ~A265 & ~A203;
  assign \new_[87483]_  = ~A298 & ~A266;
  assign \new_[87484]_  = \new_[87483]_  & \new_[87480]_ ;
  assign \new_[87487]_  = ~A300 & A299;
  assign \new_[87490]_  = ~A302 & ~A301;
  assign \new_[87491]_  = \new_[87490]_  & \new_[87487]_ ;
  assign \new_[87492]_  = \new_[87491]_  & \new_[87484]_ ;
  assign \new_[87496]_  = ~A168 & ~A169;
  assign \new_[87497]_  = A170 & \new_[87496]_ ;
  assign \new_[87500]_  = A166 & ~A167;
  assign \new_[87503]_  = A202 & ~A201;
  assign \new_[87504]_  = \new_[87503]_  & \new_[87500]_ ;
  assign \new_[87505]_  = \new_[87504]_  & \new_[87497]_ ;
  assign \new_[87508]_  = ~A268 & A267;
  assign \new_[87511]_  = A298 & ~A269;
  assign \new_[87512]_  = \new_[87511]_  & \new_[87508]_ ;
  assign \new_[87515]_  = ~A300 & ~A299;
  assign \new_[87518]_  = ~A302 & ~A301;
  assign \new_[87519]_  = \new_[87518]_  & \new_[87515]_ ;
  assign \new_[87520]_  = \new_[87519]_  & \new_[87512]_ ;
  assign \new_[87524]_  = ~A168 & ~A169;
  assign \new_[87525]_  = A170 & \new_[87524]_ ;
  assign \new_[87528]_  = A166 & ~A167;
  assign \new_[87531]_  = A202 & ~A201;
  assign \new_[87532]_  = \new_[87531]_  & \new_[87528]_ ;
  assign \new_[87533]_  = \new_[87532]_  & \new_[87525]_ ;
  assign \new_[87536]_  = ~A268 & A267;
  assign \new_[87539]_  = ~A298 & ~A269;
  assign \new_[87540]_  = \new_[87539]_  & \new_[87536]_ ;
  assign \new_[87543]_  = ~A300 & A299;
  assign \new_[87546]_  = ~A302 & ~A301;
  assign \new_[87547]_  = \new_[87546]_  & \new_[87543]_ ;
  assign \new_[87548]_  = \new_[87547]_  & \new_[87540]_ ;
  assign \new_[87552]_  = ~A168 & ~A169;
  assign \new_[87553]_  = A170 & \new_[87552]_ ;
  assign \new_[87556]_  = A166 & ~A167;
  assign \new_[87559]_  = A203 & ~A201;
  assign \new_[87560]_  = \new_[87559]_  & \new_[87556]_ ;
  assign \new_[87561]_  = \new_[87560]_  & \new_[87553]_ ;
  assign \new_[87564]_  = ~A268 & A267;
  assign \new_[87567]_  = A298 & ~A269;
  assign \new_[87568]_  = \new_[87567]_  & \new_[87564]_ ;
  assign \new_[87571]_  = ~A300 & ~A299;
  assign \new_[87574]_  = ~A302 & ~A301;
  assign \new_[87575]_  = \new_[87574]_  & \new_[87571]_ ;
  assign \new_[87576]_  = \new_[87575]_  & \new_[87568]_ ;
  assign \new_[87580]_  = ~A168 & ~A169;
  assign \new_[87581]_  = A170 & \new_[87580]_ ;
  assign \new_[87584]_  = A166 & ~A167;
  assign \new_[87587]_  = A203 & ~A201;
  assign \new_[87588]_  = \new_[87587]_  & \new_[87584]_ ;
  assign \new_[87589]_  = \new_[87588]_  & \new_[87581]_ ;
  assign \new_[87592]_  = ~A268 & A267;
  assign \new_[87595]_  = ~A298 & ~A269;
  assign \new_[87596]_  = \new_[87595]_  & \new_[87592]_ ;
  assign \new_[87599]_  = ~A300 & A299;
  assign \new_[87602]_  = ~A302 & ~A301;
  assign \new_[87603]_  = \new_[87602]_  & \new_[87599]_ ;
  assign \new_[87604]_  = \new_[87603]_  & \new_[87596]_ ;
  assign \new_[87608]_  = ~A168 & ~A169;
  assign \new_[87609]_  = A170 & \new_[87608]_ ;
  assign \new_[87612]_  = A166 & ~A167;
  assign \new_[87615]_  = A200 & A199;
  assign \new_[87616]_  = \new_[87615]_  & \new_[87612]_ ;
  assign \new_[87617]_  = \new_[87616]_  & \new_[87609]_ ;
  assign \new_[87620]_  = ~A268 & A267;
  assign \new_[87623]_  = A298 & ~A269;
  assign \new_[87624]_  = \new_[87623]_  & \new_[87620]_ ;
  assign \new_[87627]_  = ~A300 & ~A299;
  assign \new_[87630]_  = ~A302 & ~A301;
  assign \new_[87631]_  = \new_[87630]_  & \new_[87627]_ ;
  assign \new_[87632]_  = \new_[87631]_  & \new_[87624]_ ;
  assign \new_[87636]_  = ~A168 & ~A169;
  assign \new_[87637]_  = A170 & \new_[87636]_ ;
  assign \new_[87640]_  = A166 & ~A167;
  assign \new_[87643]_  = A200 & A199;
  assign \new_[87644]_  = \new_[87643]_  & \new_[87640]_ ;
  assign \new_[87645]_  = \new_[87644]_  & \new_[87637]_ ;
  assign \new_[87648]_  = ~A268 & A267;
  assign \new_[87651]_  = ~A298 & ~A269;
  assign \new_[87652]_  = \new_[87651]_  & \new_[87648]_ ;
  assign \new_[87655]_  = ~A300 & A299;
  assign \new_[87658]_  = ~A302 & ~A301;
  assign \new_[87659]_  = \new_[87658]_  & \new_[87655]_ ;
  assign \new_[87660]_  = \new_[87659]_  & \new_[87652]_ ;
  assign \new_[87664]_  = ~A168 & ~A169;
  assign \new_[87665]_  = A170 & \new_[87664]_ ;
  assign \new_[87668]_  = A166 & ~A167;
  assign \new_[87671]_  = A200 & ~A199;
  assign \new_[87672]_  = \new_[87671]_  & \new_[87668]_ ;
  assign \new_[87673]_  = \new_[87672]_  & \new_[87665]_ ;
  assign \new_[87676]_  = A202 & A201;
  assign \new_[87679]_  = A266 & ~A265;
  assign \new_[87680]_  = \new_[87679]_  & \new_[87676]_ ;
  assign \new_[87683]_  = A268 & A267;
  assign \new_[87686]_  = A301 & ~A300;
  assign \new_[87687]_  = \new_[87686]_  & \new_[87683]_ ;
  assign \new_[87688]_  = \new_[87687]_  & \new_[87680]_ ;
  assign \new_[87692]_  = ~A168 & ~A169;
  assign \new_[87693]_  = A170 & \new_[87692]_ ;
  assign \new_[87696]_  = A166 & ~A167;
  assign \new_[87699]_  = A200 & ~A199;
  assign \new_[87700]_  = \new_[87699]_  & \new_[87696]_ ;
  assign \new_[87701]_  = \new_[87700]_  & \new_[87693]_ ;
  assign \new_[87704]_  = A202 & A201;
  assign \new_[87707]_  = A266 & ~A265;
  assign \new_[87708]_  = \new_[87707]_  & \new_[87704]_ ;
  assign \new_[87711]_  = A268 & A267;
  assign \new_[87714]_  = A302 & ~A300;
  assign \new_[87715]_  = \new_[87714]_  & \new_[87711]_ ;
  assign \new_[87716]_  = \new_[87715]_  & \new_[87708]_ ;
  assign \new_[87720]_  = ~A168 & ~A169;
  assign \new_[87721]_  = A170 & \new_[87720]_ ;
  assign \new_[87724]_  = A166 & ~A167;
  assign \new_[87727]_  = A200 & ~A199;
  assign \new_[87728]_  = \new_[87727]_  & \new_[87724]_ ;
  assign \new_[87729]_  = \new_[87728]_  & \new_[87721]_ ;
  assign \new_[87732]_  = A202 & A201;
  assign \new_[87735]_  = A266 & ~A265;
  assign \new_[87736]_  = \new_[87735]_  & \new_[87732]_ ;
  assign \new_[87739]_  = A268 & A267;
  assign \new_[87742]_  = A299 & A298;
  assign \new_[87743]_  = \new_[87742]_  & \new_[87739]_ ;
  assign \new_[87744]_  = \new_[87743]_  & \new_[87736]_ ;
  assign \new_[87748]_  = ~A168 & ~A169;
  assign \new_[87749]_  = A170 & \new_[87748]_ ;
  assign \new_[87752]_  = A166 & ~A167;
  assign \new_[87755]_  = A200 & ~A199;
  assign \new_[87756]_  = \new_[87755]_  & \new_[87752]_ ;
  assign \new_[87757]_  = \new_[87756]_  & \new_[87749]_ ;
  assign \new_[87760]_  = A202 & A201;
  assign \new_[87763]_  = A266 & ~A265;
  assign \new_[87764]_  = \new_[87763]_  & \new_[87760]_ ;
  assign \new_[87767]_  = A268 & A267;
  assign \new_[87770]_  = ~A299 & ~A298;
  assign \new_[87771]_  = \new_[87770]_  & \new_[87767]_ ;
  assign \new_[87772]_  = \new_[87771]_  & \new_[87764]_ ;
  assign \new_[87776]_  = ~A168 & ~A169;
  assign \new_[87777]_  = A170 & \new_[87776]_ ;
  assign \new_[87780]_  = A166 & ~A167;
  assign \new_[87783]_  = A200 & ~A199;
  assign \new_[87784]_  = \new_[87783]_  & \new_[87780]_ ;
  assign \new_[87785]_  = \new_[87784]_  & \new_[87777]_ ;
  assign \new_[87788]_  = A202 & A201;
  assign \new_[87791]_  = A266 & ~A265;
  assign \new_[87792]_  = \new_[87791]_  & \new_[87788]_ ;
  assign \new_[87795]_  = A269 & A267;
  assign \new_[87798]_  = A301 & ~A300;
  assign \new_[87799]_  = \new_[87798]_  & \new_[87795]_ ;
  assign \new_[87800]_  = \new_[87799]_  & \new_[87792]_ ;
  assign \new_[87804]_  = ~A168 & ~A169;
  assign \new_[87805]_  = A170 & \new_[87804]_ ;
  assign \new_[87808]_  = A166 & ~A167;
  assign \new_[87811]_  = A200 & ~A199;
  assign \new_[87812]_  = \new_[87811]_  & \new_[87808]_ ;
  assign \new_[87813]_  = \new_[87812]_  & \new_[87805]_ ;
  assign \new_[87816]_  = A202 & A201;
  assign \new_[87819]_  = A266 & ~A265;
  assign \new_[87820]_  = \new_[87819]_  & \new_[87816]_ ;
  assign \new_[87823]_  = A269 & A267;
  assign \new_[87826]_  = A302 & ~A300;
  assign \new_[87827]_  = \new_[87826]_  & \new_[87823]_ ;
  assign \new_[87828]_  = \new_[87827]_  & \new_[87820]_ ;
  assign \new_[87832]_  = ~A168 & ~A169;
  assign \new_[87833]_  = A170 & \new_[87832]_ ;
  assign \new_[87836]_  = A166 & ~A167;
  assign \new_[87839]_  = A200 & ~A199;
  assign \new_[87840]_  = \new_[87839]_  & \new_[87836]_ ;
  assign \new_[87841]_  = \new_[87840]_  & \new_[87833]_ ;
  assign \new_[87844]_  = A202 & A201;
  assign \new_[87847]_  = A266 & ~A265;
  assign \new_[87848]_  = \new_[87847]_  & \new_[87844]_ ;
  assign \new_[87851]_  = A269 & A267;
  assign \new_[87854]_  = A299 & A298;
  assign \new_[87855]_  = \new_[87854]_  & \new_[87851]_ ;
  assign \new_[87856]_  = \new_[87855]_  & \new_[87848]_ ;
  assign \new_[87860]_  = ~A168 & ~A169;
  assign \new_[87861]_  = A170 & \new_[87860]_ ;
  assign \new_[87864]_  = A166 & ~A167;
  assign \new_[87867]_  = A200 & ~A199;
  assign \new_[87868]_  = \new_[87867]_  & \new_[87864]_ ;
  assign \new_[87869]_  = \new_[87868]_  & \new_[87861]_ ;
  assign \new_[87872]_  = A202 & A201;
  assign \new_[87875]_  = A266 & ~A265;
  assign \new_[87876]_  = \new_[87875]_  & \new_[87872]_ ;
  assign \new_[87879]_  = A269 & A267;
  assign \new_[87882]_  = ~A299 & ~A298;
  assign \new_[87883]_  = \new_[87882]_  & \new_[87879]_ ;
  assign \new_[87884]_  = \new_[87883]_  & \new_[87876]_ ;
  assign \new_[87888]_  = ~A168 & ~A169;
  assign \new_[87889]_  = A170 & \new_[87888]_ ;
  assign \new_[87892]_  = A166 & ~A167;
  assign \new_[87895]_  = A200 & ~A199;
  assign \new_[87896]_  = \new_[87895]_  & \new_[87892]_ ;
  assign \new_[87897]_  = \new_[87896]_  & \new_[87889]_ ;
  assign \new_[87900]_  = A202 & A201;
  assign \new_[87903]_  = ~A266 & A265;
  assign \new_[87904]_  = \new_[87903]_  & \new_[87900]_ ;
  assign \new_[87907]_  = A268 & A267;
  assign \new_[87910]_  = A301 & ~A300;
  assign \new_[87911]_  = \new_[87910]_  & \new_[87907]_ ;
  assign \new_[87912]_  = \new_[87911]_  & \new_[87904]_ ;
  assign \new_[87916]_  = ~A168 & ~A169;
  assign \new_[87917]_  = A170 & \new_[87916]_ ;
  assign \new_[87920]_  = A166 & ~A167;
  assign \new_[87923]_  = A200 & ~A199;
  assign \new_[87924]_  = \new_[87923]_  & \new_[87920]_ ;
  assign \new_[87925]_  = \new_[87924]_  & \new_[87917]_ ;
  assign \new_[87928]_  = A202 & A201;
  assign \new_[87931]_  = ~A266 & A265;
  assign \new_[87932]_  = \new_[87931]_  & \new_[87928]_ ;
  assign \new_[87935]_  = A268 & A267;
  assign \new_[87938]_  = A302 & ~A300;
  assign \new_[87939]_  = \new_[87938]_  & \new_[87935]_ ;
  assign \new_[87940]_  = \new_[87939]_  & \new_[87932]_ ;
  assign \new_[87944]_  = ~A168 & ~A169;
  assign \new_[87945]_  = A170 & \new_[87944]_ ;
  assign \new_[87948]_  = A166 & ~A167;
  assign \new_[87951]_  = A200 & ~A199;
  assign \new_[87952]_  = \new_[87951]_  & \new_[87948]_ ;
  assign \new_[87953]_  = \new_[87952]_  & \new_[87945]_ ;
  assign \new_[87956]_  = A202 & A201;
  assign \new_[87959]_  = ~A266 & A265;
  assign \new_[87960]_  = \new_[87959]_  & \new_[87956]_ ;
  assign \new_[87963]_  = A268 & A267;
  assign \new_[87966]_  = A299 & A298;
  assign \new_[87967]_  = \new_[87966]_  & \new_[87963]_ ;
  assign \new_[87968]_  = \new_[87967]_  & \new_[87960]_ ;
  assign \new_[87972]_  = ~A168 & ~A169;
  assign \new_[87973]_  = A170 & \new_[87972]_ ;
  assign \new_[87976]_  = A166 & ~A167;
  assign \new_[87979]_  = A200 & ~A199;
  assign \new_[87980]_  = \new_[87979]_  & \new_[87976]_ ;
  assign \new_[87981]_  = \new_[87980]_  & \new_[87973]_ ;
  assign \new_[87984]_  = A202 & A201;
  assign \new_[87987]_  = ~A266 & A265;
  assign \new_[87988]_  = \new_[87987]_  & \new_[87984]_ ;
  assign \new_[87991]_  = A268 & A267;
  assign \new_[87994]_  = ~A299 & ~A298;
  assign \new_[87995]_  = \new_[87994]_  & \new_[87991]_ ;
  assign \new_[87996]_  = \new_[87995]_  & \new_[87988]_ ;
  assign \new_[88000]_  = ~A168 & ~A169;
  assign \new_[88001]_  = A170 & \new_[88000]_ ;
  assign \new_[88004]_  = A166 & ~A167;
  assign \new_[88007]_  = A200 & ~A199;
  assign \new_[88008]_  = \new_[88007]_  & \new_[88004]_ ;
  assign \new_[88009]_  = \new_[88008]_  & \new_[88001]_ ;
  assign \new_[88012]_  = A202 & A201;
  assign \new_[88015]_  = ~A266 & A265;
  assign \new_[88016]_  = \new_[88015]_  & \new_[88012]_ ;
  assign \new_[88019]_  = A269 & A267;
  assign \new_[88022]_  = A301 & ~A300;
  assign \new_[88023]_  = \new_[88022]_  & \new_[88019]_ ;
  assign \new_[88024]_  = \new_[88023]_  & \new_[88016]_ ;
  assign \new_[88028]_  = ~A168 & ~A169;
  assign \new_[88029]_  = A170 & \new_[88028]_ ;
  assign \new_[88032]_  = A166 & ~A167;
  assign \new_[88035]_  = A200 & ~A199;
  assign \new_[88036]_  = \new_[88035]_  & \new_[88032]_ ;
  assign \new_[88037]_  = \new_[88036]_  & \new_[88029]_ ;
  assign \new_[88040]_  = A202 & A201;
  assign \new_[88043]_  = ~A266 & A265;
  assign \new_[88044]_  = \new_[88043]_  & \new_[88040]_ ;
  assign \new_[88047]_  = A269 & A267;
  assign \new_[88050]_  = A302 & ~A300;
  assign \new_[88051]_  = \new_[88050]_  & \new_[88047]_ ;
  assign \new_[88052]_  = \new_[88051]_  & \new_[88044]_ ;
  assign \new_[88056]_  = ~A168 & ~A169;
  assign \new_[88057]_  = A170 & \new_[88056]_ ;
  assign \new_[88060]_  = A166 & ~A167;
  assign \new_[88063]_  = A200 & ~A199;
  assign \new_[88064]_  = \new_[88063]_  & \new_[88060]_ ;
  assign \new_[88065]_  = \new_[88064]_  & \new_[88057]_ ;
  assign \new_[88068]_  = A202 & A201;
  assign \new_[88071]_  = ~A266 & A265;
  assign \new_[88072]_  = \new_[88071]_  & \new_[88068]_ ;
  assign \new_[88075]_  = A269 & A267;
  assign \new_[88078]_  = A299 & A298;
  assign \new_[88079]_  = \new_[88078]_  & \new_[88075]_ ;
  assign \new_[88080]_  = \new_[88079]_  & \new_[88072]_ ;
  assign \new_[88084]_  = ~A168 & ~A169;
  assign \new_[88085]_  = A170 & \new_[88084]_ ;
  assign \new_[88088]_  = A166 & ~A167;
  assign \new_[88091]_  = A200 & ~A199;
  assign \new_[88092]_  = \new_[88091]_  & \new_[88088]_ ;
  assign \new_[88093]_  = \new_[88092]_  & \new_[88085]_ ;
  assign \new_[88096]_  = A202 & A201;
  assign \new_[88099]_  = ~A266 & A265;
  assign \new_[88100]_  = \new_[88099]_  & \new_[88096]_ ;
  assign \new_[88103]_  = A269 & A267;
  assign \new_[88106]_  = ~A299 & ~A298;
  assign \new_[88107]_  = \new_[88106]_  & \new_[88103]_ ;
  assign \new_[88108]_  = \new_[88107]_  & \new_[88100]_ ;
  assign \new_[88112]_  = ~A168 & ~A169;
  assign \new_[88113]_  = A170 & \new_[88112]_ ;
  assign \new_[88116]_  = A166 & ~A167;
  assign \new_[88119]_  = A200 & ~A199;
  assign \new_[88120]_  = \new_[88119]_  & \new_[88116]_ ;
  assign \new_[88121]_  = \new_[88120]_  & \new_[88113]_ ;
  assign \new_[88124]_  = A203 & A201;
  assign \new_[88127]_  = A266 & ~A265;
  assign \new_[88128]_  = \new_[88127]_  & \new_[88124]_ ;
  assign \new_[88131]_  = A268 & A267;
  assign \new_[88134]_  = A301 & ~A300;
  assign \new_[88135]_  = \new_[88134]_  & \new_[88131]_ ;
  assign \new_[88136]_  = \new_[88135]_  & \new_[88128]_ ;
  assign \new_[88140]_  = ~A168 & ~A169;
  assign \new_[88141]_  = A170 & \new_[88140]_ ;
  assign \new_[88144]_  = A166 & ~A167;
  assign \new_[88147]_  = A200 & ~A199;
  assign \new_[88148]_  = \new_[88147]_  & \new_[88144]_ ;
  assign \new_[88149]_  = \new_[88148]_  & \new_[88141]_ ;
  assign \new_[88152]_  = A203 & A201;
  assign \new_[88155]_  = A266 & ~A265;
  assign \new_[88156]_  = \new_[88155]_  & \new_[88152]_ ;
  assign \new_[88159]_  = A268 & A267;
  assign \new_[88162]_  = A302 & ~A300;
  assign \new_[88163]_  = \new_[88162]_  & \new_[88159]_ ;
  assign \new_[88164]_  = \new_[88163]_  & \new_[88156]_ ;
  assign \new_[88168]_  = ~A168 & ~A169;
  assign \new_[88169]_  = A170 & \new_[88168]_ ;
  assign \new_[88172]_  = A166 & ~A167;
  assign \new_[88175]_  = A200 & ~A199;
  assign \new_[88176]_  = \new_[88175]_  & \new_[88172]_ ;
  assign \new_[88177]_  = \new_[88176]_  & \new_[88169]_ ;
  assign \new_[88180]_  = A203 & A201;
  assign \new_[88183]_  = A266 & ~A265;
  assign \new_[88184]_  = \new_[88183]_  & \new_[88180]_ ;
  assign \new_[88187]_  = A268 & A267;
  assign \new_[88190]_  = A299 & A298;
  assign \new_[88191]_  = \new_[88190]_  & \new_[88187]_ ;
  assign \new_[88192]_  = \new_[88191]_  & \new_[88184]_ ;
  assign \new_[88196]_  = ~A168 & ~A169;
  assign \new_[88197]_  = A170 & \new_[88196]_ ;
  assign \new_[88200]_  = A166 & ~A167;
  assign \new_[88203]_  = A200 & ~A199;
  assign \new_[88204]_  = \new_[88203]_  & \new_[88200]_ ;
  assign \new_[88205]_  = \new_[88204]_  & \new_[88197]_ ;
  assign \new_[88208]_  = A203 & A201;
  assign \new_[88211]_  = A266 & ~A265;
  assign \new_[88212]_  = \new_[88211]_  & \new_[88208]_ ;
  assign \new_[88215]_  = A268 & A267;
  assign \new_[88218]_  = ~A299 & ~A298;
  assign \new_[88219]_  = \new_[88218]_  & \new_[88215]_ ;
  assign \new_[88220]_  = \new_[88219]_  & \new_[88212]_ ;
  assign \new_[88224]_  = ~A168 & ~A169;
  assign \new_[88225]_  = A170 & \new_[88224]_ ;
  assign \new_[88228]_  = A166 & ~A167;
  assign \new_[88231]_  = A200 & ~A199;
  assign \new_[88232]_  = \new_[88231]_  & \new_[88228]_ ;
  assign \new_[88233]_  = \new_[88232]_  & \new_[88225]_ ;
  assign \new_[88236]_  = A203 & A201;
  assign \new_[88239]_  = A266 & ~A265;
  assign \new_[88240]_  = \new_[88239]_  & \new_[88236]_ ;
  assign \new_[88243]_  = A269 & A267;
  assign \new_[88246]_  = A301 & ~A300;
  assign \new_[88247]_  = \new_[88246]_  & \new_[88243]_ ;
  assign \new_[88248]_  = \new_[88247]_  & \new_[88240]_ ;
  assign \new_[88252]_  = ~A168 & ~A169;
  assign \new_[88253]_  = A170 & \new_[88252]_ ;
  assign \new_[88256]_  = A166 & ~A167;
  assign \new_[88259]_  = A200 & ~A199;
  assign \new_[88260]_  = \new_[88259]_  & \new_[88256]_ ;
  assign \new_[88261]_  = \new_[88260]_  & \new_[88253]_ ;
  assign \new_[88264]_  = A203 & A201;
  assign \new_[88267]_  = A266 & ~A265;
  assign \new_[88268]_  = \new_[88267]_  & \new_[88264]_ ;
  assign \new_[88271]_  = A269 & A267;
  assign \new_[88274]_  = A302 & ~A300;
  assign \new_[88275]_  = \new_[88274]_  & \new_[88271]_ ;
  assign \new_[88276]_  = \new_[88275]_  & \new_[88268]_ ;
  assign \new_[88280]_  = ~A168 & ~A169;
  assign \new_[88281]_  = A170 & \new_[88280]_ ;
  assign \new_[88284]_  = A166 & ~A167;
  assign \new_[88287]_  = A200 & ~A199;
  assign \new_[88288]_  = \new_[88287]_  & \new_[88284]_ ;
  assign \new_[88289]_  = \new_[88288]_  & \new_[88281]_ ;
  assign \new_[88292]_  = A203 & A201;
  assign \new_[88295]_  = A266 & ~A265;
  assign \new_[88296]_  = \new_[88295]_  & \new_[88292]_ ;
  assign \new_[88299]_  = A269 & A267;
  assign \new_[88302]_  = A299 & A298;
  assign \new_[88303]_  = \new_[88302]_  & \new_[88299]_ ;
  assign \new_[88304]_  = \new_[88303]_  & \new_[88296]_ ;
  assign \new_[88308]_  = ~A168 & ~A169;
  assign \new_[88309]_  = A170 & \new_[88308]_ ;
  assign \new_[88312]_  = A166 & ~A167;
  assign \new_[88315]_  = A200 & ~A199;
  assign \new_[88316]_  = \new_[88315]_  & \new_[88312]_ ;
  assign \new_[88317]_  = \new_[88316]_  & \new_[88309]_ ;
  assign \new_[88320]_  = A203 & A201;
  assign \new_[88323]_  = A266 & ~A265;
  assign \new_[88324]_  = \new_[88323]_  & \new_[88320]_ ;
  assign \new_[88327]_  = A269 & A267;
  assign \new_[88330]_  = ~A299 & ~A298;
  assign \new_[88331]_  = \new_[88330]_  & \new_[88327]_ ;
  assign \new_[88332]_  = \new_[88331]_  & \new_[88324]_ ;
  assign \new_[88336]_  = ~A168 & ~A169;
  assign \new_[88337]_  = A170 & \new_[88336]_ ;
  assign \new_[88340]_  = A166 & ~A167;
  assign \new_[88343]_  = A200 & ~A199;
  assign \new_[88344]_  = \new_[88343]_  & \new_[88340]_ ;
  assign \new_[88345]_  = \new_[88344]_  & \new_[88337]_ ;
  assign \new_[88348]_  = A203 & A201;
  assign \new_[88351]_  = ~A266 & A265;
  assign \new_[88352]_  = \new_[88351]_  & \new_[88348]_ ;
  assign \new_[88355]_  = A268 & A267;
  assign \new_[88358]_  = A301 & ~A300;
  assign \new_[88359]_  = \new_[88358]_  & \new_[88355]_ ;
  assign \new_[88360]_  = \new_[88359]_  & \new_[88352]_ ;
  assign \new_[88364]_  = ~A168 & ~A169;
  assign \new_[88365]_  = A170 & \new_[88364]_ ;
  assign \new_[88368]_  = A166 & ~A167;
  assign \new_[88371]_  = A200 & ~A199;
  assign \new_[88372]_  = \new_[88371]_  & \new_[88368]_ ;
  assign \new_[88373]_  = \new_[88372]_  & \new_[88365]_ ;
  assign \new_[88376]_  = A203 & A201;
  assign \new_[88379]_  = ~A266 & A265;
  assign \new_[88380]_  = \new_[88379]_  & \new_[88376]_ ;
  assign \new_[88383]_  = A268 & A267;
  assign \new_[88386]_  = A302 & ~A300;
  assign \new_[88387]_  = \new_[88386]_  & \new_[88383]_ ;
  assign \new_[88388]_  = \new_[88387]_  & \new_[88380]_ ;
  assign \new_[88392]_  = ~A168 & ~A169;
  assign \new_[88393]_  = A170 & \new_[88392]_ ;
  assign \new_[88396]_  = A166 & ~A167;
  assign \new_[88399]_  = A200 & ~A199;
  assign \new_[88400]_  = \new_[88399]_  & \new_[88396]_ ;
  assign \new_[88401]_  = \new_[88400]_  & \new_[88393]_ ;
  assign \new_[88404]_  = A203 & A201;
  assign \new_[88407]_  = ~A266 & A265;
  assign \new_[88408]_  = \new_[88407]_  & \new_[88404]_ ;
  assign \new_[88411]_  = A268 & A267;
  assign \new_[88414]_  = A299 & A298;
  assign \new_[88415]_  = \new_[88414]_  & \new_[88411]_ ;
  assign \new_[88416]_  = \new_[88415]_  & \new_[88408]_ ;
  assign \new_[88420]_  = ~A168 & ~A169;
  assign \new_[88421]_  = A170 & \new_[88420]_ ;
  assign \new_[88424]_  = A166 & ~A167;
  assign \new_[88427]_  = A200 & ~A199;
  assign \new_[88428]_  = \new_[88427]_  & \new_[88424]_ ;
  assign \new_[88429]_  = \new_[88428]_  & \new_[88421]_ ;
  assign \new_[88432]_  = A203 & A201;
  assign \new_[88435]_  = ~A266 & A265;
  assign \new_[88436]_  = \new_[88435]_  & \new_[88432]_ ;
  assign \new_[88439]_  = A268 & A267;
  assign \new_[88442]_  = ~A299 & ~A298;
  assign \new_[88443]_  = \new_[88442]_  & \new_[88439]_ ;
  assign \new_[88444]_  = \new_[88443]_  & \new_[88436]_ ;
  assign \new_[88448]_  = ~A168 & ~A169;
  assign \new_[88449]_  = A170 & \new_[88448]_ ;
  assign \new_[88452]_  = A166 & ~A167;
  assign \new_[88455]_  = A200 & ~A199;
  assign \new_[88456]_  = \new_[88455]_  & \new_[88452]_ ;
  assign \new_[88457]_  = \new_[88456]_  & \new_[88449]_ ;
  assign \new_[88460]_  = A203 & A201;
  assign \new_[88463]_  = ~A266 & A265;
  assign \new_[88464]_  = \new_[88463]_  & \new_[88460]_ ;
  assign \new_[88467]_  = A269 & A267;
  assign \new_[88470]_  = A301 & ~A300;
  assign \new_[88471]_  = \new_[88470]_  & \new_[88467]_ ;
  assign \new_[88472]_  = \new_[88471]_  & \new_[88464]_ ;
  assign \new_[88476]_  = ~A168 & ~A169;
  assign \new_[88477]_  = A170 & \new_[88476]_ ;
  assign \new_[88480]_  = A166 & ~A167;
  assign \new_[88483]_  = A200 & ~A199;
  assign \new_[88484]_  = \new_[88483]_  & \new_[88480]_ ;
  assign \new_[88485]_  = \new_[88484]_  & \new_[88477]_ ;
  assign \new_[88488]_  = A203 & A201;
  assign \new_[88491]_  = ~A266 & A265;
  assign \new_[88492]_  = \new_[88491]_  & \new_[88488]_ ;
  assign \new_[88495]_  = A269 & A267;
  assign \new_[88498]_  = A302 & ~A300;
  assign \new_[88499]_  = \new_[88498]_  & \new_[88495]_ ;
  assign \new_[88500]_  = \new_[88499]_  & \new_[88492]_ ;
  assign \new_[88504]_  = ~A168 & ~A169;
  assign \new_[88505]_  = A170 & \new_[88504]_ ;
  assign \new_[88508]_  = A166 & ~A167;
  assign \new_[88511]_  = A200 & ~A199;
  assign \new_[88512]_  = \new_[88511]_  & \new_[88508]_ ;
  assign \new_[88513]_  = \new_[88512]_  & \new_[88505]_ ;
  assign \new_[88516]_  = A203 & A201;
  assign \new_[88519]_  = ~A266 & A265;
  assign \new_[88520]_  = \new_[88519]_  & \new_[88516]_ ;
  assign \new_[88523]_  = A269 & A267;
  assign \new_[88526]_  = A299 & A298;
  assign \new_[88527]_  = \new_[88526]_  & \new_[88523]_ ;
  assign \new_[88528]_  = \new_[88527]_  & \new_[88520]_ ;
  assign \new_[88532]_  = ~A168 & ~A169;
  assign \new_[88533]_  = A170 & \new_[88532]_ ;
  assign \new_[88536]_  = A166 & ~A167;
  assign \new_[88539]_  = A200 & ~A199;
  assign \new_[88540]_  = \new_[88539]_  & \new_[88536]_ ;
  assign \new_[88541]_  = \new_[88540]_  & \new_[88533]_ ;
  assign \new_[88544]_  = A203 & A201;
  assign \new_[88547]_  = ~A266 & A265;
  assign \new_[88548]_  = \new_[88547]_  & \new_[88544]_ ;
  assign \new_[88551]_  = A269 & A267;
  assign \new_[88554]_  = ~A299 & ~A298;
  assign \new_[88555]_  = \new_[88554]_  & \new_[88551]_ ;
  assign \new_[88556]_  = \new_[88555]_  & \new_[88548]_ ;
  assign \new_[88560]_  = ~A168 & ~A169;
  assign \new_[88561]_  = A170 & \new_[88560]_ ;
  assign \new_[88564]_  = A166 & ~A167;
  assign \new_[88567]_  = ~A200 & A199;
  assign \new_[88568]_  = \new_[88567]_  & \new_[88564]_ ;
  assign \new_[88569]_  = \new_[88568]_  & \new_[88561]_ ;
  assign \new_[88572]_  = A202 & A201;
  assign \new_[88575]_  = A266 & ~A265;
  assign \new_[88576]_  = \new_[88575]_  & \new_[88572]_ ;
  assign \new_[88579]_  = A268 & A267;
  assign \new_[88582]_  = A301 & ~A300;
  assign \new_[88583]_  = \new_[88582]_  & \new_[88579]_ ;
  assign \new_[88584]_  = \new_[88583]_  & \new_[88576]_ ;
  assign \new_[88588]_  = ~A168 & ~A169;
  assign \new_[88589]_  = A170 & \new_[88588]_ ;
  assign \new_[88592]_  = A166 & ~A167;
  assign \new_[88595]_  = ~A200 & A199;
  assign \new_[88596]_  = \new_[88595]_  & \new_[88592]_ ;
  assign \new_[88597]_  = \new_[88596]_  & \new_[88589]_ ;
  assign \new_[88600]_  = A202 & A201;
  assign \new_[88603]_  = A266 & ~A265;
  assign \new_[88604]_  = \new_[88603]_  & \new_[88600]_ ;
  assign \new_[88607]_  = A268 & A267;
  assign \new_[88610]_  = A302 & ~A300;
  assign \new_[88611]_  = \new_[88610]_  & \new_[88607]_ ;
  assign \new_[88612]_  = \new_[88611]_  & \new_[88604]_ ;
  assign \new_[88616]_  = ~A168 & ~A169;
  assign \new_[88617]_  = A170 & \new_[88616]_ ;
  assign \new_[88620]_  = A166 & ~A167;
  assign \new_[88623]_  = ~A200 & A199;
  assign \new_[88624]_  = \new_[88623]_  & \new_[88620]_ ;
  assign \new_[88625]_  = \new_[88624]_  & \new_[88617]_ ;
  assign \new_[88628]_  = A202 & A201;
  assign \new_[88631]_  = A266 & ~A265;
  assign \new_[88632]_  = \new_[88631]_  & \new_[88628]_ ;
  assign \new_[88635]_  = A268 & A267;
  assign \new_[88638]_  = A299 & A298;
  assign \new_[88639]_  = \new_[88638]_  & \new_[88635]_ ;
  assign \new_[88640]_  = \new_[88639]_  & \new_[88632]_ ;
  assign \new_[88644]_  = ~A168 & ~A169;
  assign \new_[88645]_  = A170 & \new_[88644]_ ;
  assign \new_[88648]_  = A166 & ~A167;
  assign \new_[88651]_  = ~A200 & A199;
  assign \new_[88652]_  = \new_[88651]_  & \new_[88648]_ ;
  assign \new_[88653]_  = \new_[88652]_  & \new_[88645]_ ;
  assign \new_[88656]_  = A202 & A201;
  assign \new_[88659]_  = A266 & ~A265;
  assign \new_[88660]_  = \new_[88659]_  & \new_[88656]_ ;
  assign \new_[88663]_  = A268 & A267;
  assign \new_[88666]_  = ~A299 & ~A298;
  assign \new_[88667]_  = \new_[88666]_  & \new_[88663]_ ;
  assign \new_[88668]_  = \new_[88667]_  & \new_[88660]_ ;
  assign \new_[88672]_  = ~A168 & ~A169;
  assign \new_[88673]_  = A170 & \new_[88672]_ ;
  assign \new_[88676]_  = A166 & ~A167;
  assign \new_[88679]_  = ~A200 & A199;
  assign \new_[88680]_  = \new_[88679]_  & \new_[88676]_ ;
  assign \new_[88681]_  = \new_[88680]_  & \new_[88673]_ ;
  assign \new_[88684]_  = A202 & A201;
  assign \new_[88687]_  = A266 & ~A265;
  assign \new_[88688]_  = \new_[88687]_  & \new_[88684]_ ;
  assign \new_[88691]_  = A269 & A267;
  assign \new_[88694]_  = A301 & ~A300;
  assign \new_[88695]_  = \new_[88694]_  & \new_[88691]_ ;
  assign \new_[88696]_  = \new_[88695]_  & \new_[88688]_ ;
  assign \new_[88700]_  = ~A168 & ~A169;
  assign \new_[88701]_  = A170 & \new_[88700]_ ;
  assign \new_[88704]_  = A166 & ~A167;
  assign \new_[88707]_  = ~A200 & A199;
  assign \new_[88708]_  = \new_[88707]_  & \new_[88704]_ ;
  assign \new_[88709]_  = \new_[88708]_  & \new_[88701]_ ;
  assign \new_[88712]_  = A202 & A201;
  assign \new_[88715]_  = A266 & ~A265;
  assign \new_[88716]_  = \new_[88715]_  & \new_[88712]_ ;
  assign \new_[88719]_  = A269 & A267;
  assign \new_[88722]_  = A302 & ~A300;
  assign \new_[88723]_  = \new_[88722]_  & \new_[88719]_ ;
  assign \new_[88724]_  = \new_[88723]_  & \new_[88716]_ ;
  assign \new_[88728]_  = ~A168 & ~A169;
  assign \new_[88729]_  = A170 & \new_[88728]_ ;
  assign \new_[88732]_  = A166 & ~A167;
  assign \new_[88735]_  = ~A200 & A199;
  assign \new_[88736]_  = \new_[88735]_  & \new_[88732]_ ;
  assign \new_[88737]_  = \new_[88736]_  & \new_[88729]_ ;
  assign \new_[88740]_  = A202 & A201;
  assign \new_[88743]_  = A266 & ~A265;
  assign \new_[88744]_  = \new_[88743]_  & \new_[88740]_ ;
  assign \new_[88747]_  = A269 & A267;
  assign \new_[88750]_  = A299 & A298;
  assign \new_[88751]_  = \new_[88750]_  & \new_[88747]_ ;
  assign \new_[88752]_  = \new_[88751]_  & \new_[88744]_ ;
  assign \new_[88756]_  = ~A168 & ~A169;
  assign \new_[88757]_  = A170 & \new_[88756]_ ;
  assign \new_[88760]_  = A166 & ~A167;
  assign \new_[88763]_  = ~A200 & A199;
  assign \new_[88764]_  = \new_[88763]_  & \new_[88760]_ ;
  assign \new_[88765]_  = \new_[88764]_  & \new_[88757]_ ;
  assign \new_[88768]_  = A202 & A201;
  assign \new_[88771]_  = A266 & ~A265;
  assign \new_[88772]_  = \new_[88771]_  & \new_[88768]_ ;
  assign \new_[88775]_  = A269 & A267;
  assign \new_[88778]_  = ~A299 & ~A298;
  assign \new_[88779]_  = \new_[88778]_  & \new_[88775]_ ;
  assign \new_[88780]_  = \new_[88779]_  & \new_[88772]_ ;
  assign \new_[88784]_  = ~A168 & ~A169;
  assign \new_[88785]_  = A170 & \new_[88784]_ ;
  assign \new_[88788]_  = A166 & ~A167;
  assign \new_[88791]_  = ~A200 & A199;
  assign \new_[88792]_  = \new_[88791]_  & \new_[88788]_ ;
  assign \new_[88793]_  = \new_[88792]_  & \new_[88785]_ ;
  assign \new_[88796]_  = A202 & A201;
  assign \new_[88799]_  = ~A266 & A265;
  assign \new_[88800]_  = \new_[88799]_  & \new_[88796]_ ;
  assign \new_[88803]_  = A268 & A267;
  assign \new_[88806]_  = A301 & ~A300;
  assign \new_[88807]_  = \new_[88806]_  & \new_[88803]_ ;
  assign \new_[88808]_  = \new_[88807]_  & \new_[88800]_ ;
  assign \new_[88812]_  = ~A168 & ~A169;
  assign \new_[88813]_  = A170 & \new_[88812]_ ;
  assign \new_[88816]_  = A166 & ~A167;
  assign \new_[88819]_  = ~A200 & A199;
  assign \new_[88820]_  = \new_[88819]_  & \new_[88816]_ ;
  assign \new_[88821]_  = \new_[88820]_  & \new_[88813]_ ;
  assign \new_[88824]_  = A202 & A201;
  assign \new_[88827]_  = ~A266 & A265;
  assign \new_[88828]_  = \new_[88827]_  & \new_[88824]_ ;
  assign \new_[88831]_  = A268 & A267;
  assign \new_[88834]_  = A302 & ~A300;
  assign \new_[88835]_  = \new_[88834]_  & \new_[88831]_ ;
  assign \new_[88836]_  = \new_[88835]_  & \new_[88828]_ ;
  assign \new_[88840]_  = ~A168 & ~A169;
  assign \new_[88841]_  = A170 & \new_[88840]_ ;
  assign \new_[88844]_  = A166 & ~A167;
  assign \new_[88847]_  = ~A200 & A199;
  assign \new_[88848]_  = \new_[88847]_  & \new_[88844]_ ;
  assign \new_[88849]_  = \new_[88848]_  & \new_[88841]_ ;
  assign \new_[88852]_  = A202 & A201;
  assign \new_[88855]_  = ~A266 & A265;
  assign \new_[88856]_  = \new_[88855]_  & \new_[88852]_ ;
  assign \new_[88859]_  = A268 & A267;
  assign \new_[88862]_  = A299 & A298;
  assign \new_[88863]_  = \new_[88862]_  & \new_[88859]_ ;
  assign \new_[88864]_  = \new_[88863]_  & \new_[88856]_ ;
  assign \new_[88868]_  = ~A168 & ~A169;
  assign \new_[88869]_  = A170 & \new_[88868]_ ;
  assign \new_[88872]_  = A166 & ~A167;
  assign \new_[88875]_  = ~A200 & A199;
  assign \new_[88876]_  = \new_[88875]_  & \new_[88872]_ ;
  assign \new_[88877]_  = \new_[88876]_  & \new_[88869]_ ;
  assign \new_[88880]_  = A202 & A201;
  assign \new_[88883]_  = ~A266 & A265;
  assign \new_[88884]_  = \new_[88883]_  & \new_[88880]_ ;
  assign \new_[88887]_  = A268 & A267;
  assign \new_[88890]_  = ~A299 & ~A298;
  assign \new_[88891]_  = \new_[88890]_  & \new_[88887]_ ;
  assign \new_[88892]_  = \new_[88891]_  & \new_[88884]_ ;
  assign \new_[88896]_  = ~A168 & ~A169;
  assign \new_[88897]_  = A170 & \new_[88896]_ ;
  assign \new_[88900]_  = A166 & ~A167;
  assign \new_[88903]_  = ~A200 & A199;
  assign \new_[88904]_  = \new_[88903]_  & \new_[88900]_ ;
  assign \new_[88905]_  = \new_[88904]_  & \new_[88897]_ ;
  assign \new_[88908]_  = A202 & A201;
  assign \new_[88911]_  = ~A266 & A265;
  assign \new_[88912]_  = \new_[88911]_  & \new_[88908]_ ;
  assign \new_[88915]_  = A269 & A267;
  assign \new_[88918]_  = A301 & ~A300;
  assign \new_[88919]_  = \new_[88918]_  & \new_[88915]_ ;
  assign \new_[88920]_  = \new_[88919]_  & \new_[88912]_ ;
  assign \new_[88924]_  = ~A168 & ~A169;
  assign \new_[88925]_  = A170 & \new_[88924]_ ;
  assign \new_[88928]_  = A166 & ~A167;
  assign \new_[88931]_  = ~A200 & A199;
  assign \new_[88932]_  = \new_[88931]_  & \new_[88928]_ ;
  assign \new_[88933]_  = \new_[88932]_  & \new_[88925]_ ;
  assign \new_[88936]_  = A202 & A201;
  assign \new_[88939]_  = ~A266 & A265;
  assign \new_[88940]_  = \new_[88939]_  & \new_[88936]_ ;
  assign \new_[88943]_  = A269 & A267;
  assign \new_[88946]_  = A302 & ~A300;
  assign \new_[88947]_  = \new_[88946]_  & \new_[88943]_ ;
  assign \new_[88948]_  = \new_[88947]_  & \new_[88940]_ ;
  assign \new_[88952]_  = ~A168 & ~A169;
  assign \new_[88953]_  = A170 & \new_[88952]_ ;
  assign \new_[88956]_  = A166 & ~A167;
  assign \new_[88959]_  = ~A200 & A199;
  assign \new_[88960]_  = \new_[88959]_  & \new_[88956]_ ;
  assign \new_[88961]_  = \new_[88960]_  & \new_[88953]_ ;
  assign \new_[88964]_  = A202 & A201;
  assign \new_[88967]_  = ~A266 & A265;
  assign \new_[88968]_  = \new_[88967]_  & \new_[88964]_ ;
  assign \new_[88971]_  = A269 & A267;
  assign \new_[88974]_  = A299 & A298;
  assign \new_[88975]_  = \new_[88974]_  & \new_[88971]_ ;
  assign \new_[88976]_  = \new_[88975]_  & \new_[88968]_ ;
  assign \new_[88980]_  = ~A168 & ~A169;
  assign \new_[88981]_  = A170 & \new_[88980]_ ;
  assign \new_[88984]_  = A166 & ~A167;
  assign \new_[88987]_  = ~A200 & A199;
  assign \new_[88988]_  = \new_[88987]_  & \new_[88984]_ ;
  assign \new_[88989]_  = \new_[88988]_  & \new_[88981]_ ;
  assign \new_[88992]_  = A202 & A201;
  assign \new_[88995]_  = ~A266 & A265;
  assign \new_[88996]_  = \new_[88995]_  & \new_[88992]_ ;
  assign \new_[88999]_  = A269 & A267;
  assign \new_[89002]_  = ~A299 & ~A298;
  assign \new_[89003]_  = \new_[89002]_  & \new_[88999]_ ;
  assign \new_[89004]_  = \new_[89003]_  & \new_[88996]_ ;
  assign \new_[89008]_  = ~A168 & ~A169;
  assign \new_[89009]_  = A170 & \new_[89008]_ ;
  assign \new_[89012]_  = A166 & ~A167;
  assign \new_[89015]_  = ~A200 & A199;
  assign \new_[89016]_  = \new_[89015]_  & \new_[89012]_ ;
  assign \new_[89017]_  = \new_[89016]_  & \new_[89009]_ ;
  assign \new_[89020]_  = A203 & A201;
  assign \new_[89023]_  = A266 & ~A265;
  assign \new_[89024]_  = \new_[89023]_  & \new_[89020]_ ;
  assign \new_[89027]_  = A268 & A267;
  assign \new_[89030]_  = A301 & ~A300;
  assign \new_[89031]_  = \new_[89030]_  & \new_[89027]_ ;
  assign \new_[89032]_  = \new_[89031]_  & \new_[89024]_ ;
  assign \new_[89036]_  = ~A168 & ~A169;
  assign \new_[89037]_  = A170 & \new_[89036]_ ;
  assign \new_[89040]_  = A166 & ~A167;
  assign \new_[89043]_  = ~A200 & A199;
  assign \new_[89044]_  = \new_[89043]_  & \new_[89040]_ ;
  assign \new_[89045]_  = \new_[89044]_  & \new_[89037]_ ;
  assign \new_[89048]_  = A203 & A201;
  assign \new_[89051]_  = A266 & ~A265;
  assign \new_[89052]_  = \new_[89051]_  & \new_[89048]_ ;
  assign \new_[89055]_  = A268 & A267;
  assign \new_[89058]_  = A302 & ~A300;
  assign \new_[89059]_  = \new_[89058]_  & \new_[89055]_ ;
  assign \new_[89060]_  = \new_[89059]_  & \new_[89052]_ ;
  assign \new_[89064]_  = ~A168 & ~A169;
  assign \new_[89065]_  = A170 & \new_[89064]_ ;
  assign \new_[89068]_  = A166 & ~A167;
  assign \new_[89071]_  = ~A200 & A199;
  assign \new_[89072]_  = \new_[89071]_  & \new_[89068]_ ;
  assign \new_[89073]_  = \new_[89072]_  & \new_[89065]_ ;
  assign \new_[89076]_  = A203 & A201;
  assign \new_[89079]_  = A266 & ~A265;
  assign \new_[89080]_  = \new_[89079]_  & \new_[89076]_ ;
  assign \new_[89083]_  = A268 & A267;
  assign \new_[89086]_  = A299 & A298;
  assign \new_[89087]_  = \new_[89086]_  & \new_[89083]_ ;
  assign \new_[89088]_  = \new_[89087]_  & \new_[89080]_ ;
  assign \new_[89092]_  = ~A168 & ~A169;
  assign \new_[89093]_  = A170 & \new_[89092]_ ;
  assign \new_[89096]_  = A166 & ~A167;
  assign \new_[89099]_  = ~A200 & A199;
  assign \new_[89100]_  = \new_[89099]_  & \new_[89096]_ ;
  assign \new_[89101]_  = \new_[89100]_  & \new_[89093]_ ;
  assign \new_[89104]_  = A203 & A201;
  assign \new_[89107]_  = A266 & ~A265;
  assign \new_[89108]_  = \new_[89107]_  & \new_[89104]_ ;
  assign \new_[89111]_  = A268 & A267;
  assign \new_[89114]_  = ~A299 & ~A298;
  assign \new_[89115]_  = \new_[89114]_  & \new_[89111]_ ;
  assign \new_[89116]_  = \new_[89115]_  & \new_[89108]_ ;
  assign \new_[89120]_  = ~A168 & ~A169;
  assign \new_[89121]_  = A170 & \new_[89120]_ ;
  assign \new_[89124]_  = A166 & ~A167;
  assign \new_[89127]_  = ~A200 & A199;
  assign \new_[89128]_  = \new_[89127]_  & \new_[89124]_ ;
  assign \new_[89129]_  = \new_[89128]_  & \new_[89121]_ ;
  assign \new_[89132]_  = A203 & A201;
  assign \new_[89135]_  = A266 & ~A265;
  assign \new_[89136]_  = \new_[89135]_  & \new_[89132]_ ;
  assign \new_[89139]_  = A269 & A267;
  assign \new_[89142]_  = A301 & ~A300;
  assign \new_[89143]_  = \new_[89142]_  & \new_[89139]_ ;
  assign \new_[89144]_  = \new_[89143]_  & \new_[89136]_ ;
  assign \new_[89148]_  = ~A168 & ~A169;
  assign \new_[89149]_  = A170 & \new_[89148]_ ;
  assign \new_[89152]_  = A166 & ~A167;
  assign \new_[89155]_  = ~A200 & A199;
  assign \new_[89156]_  = \new_[89155]_  & \new_[89152]_ ;
  assign \new_[89157]_  = \new_[89156]_  & \new_[89149]_ ;
  assign \new_[89160]_  = A203 & A201;
  assign \new_[89163]_  = A266 & ~A265;
  assign \new_[89164]_  = \new_[89163]_  & \new_[89160]_ ;
  assign \new_[89167]_  = A269 & A267;
  assign \new_[89170]_  = A302 & ~A300;
  assign \new_[89171]_  = \new_[89170]_  & \new_[89167]_ ;
  assign \new_[89172]_  = \new_[89171]_  & \new_[89164]_ ;
  assign \new_[89176]_  = ~A168 & ~A169;
  assign \new_[89177]_  = A170 & \new_[89176]_ ;
  assign \new_[89180]_  = A166 & ~A167;
  assign \new_[89183]_  = ~A200 & A199;
  assign \new_[89184]_  = \new_[89183]_  & \new_[89180]_ ;
  assign \new_[89185]_  = \new_[89184]_  & \new_[89177]_ ;
  assign \new_[89188]_  = A203 & A201;
  assign \new_[89191]_  = A266 & ~A265;
  assign \new_[89192]_  = \new_[89191]_  & \new_[89188]_ ;
  assign \new_[89195]_  = A269 & A267;
  assign \new_[89198]_  = A299 & A298;
  assign \new_[89199]_  = \new_[89198]_  & \new_[89195]_ ;
  assign \new_[89200]_  = \new_[89199]_  & \new_[89192]_ ;
  assign \new_[89204]_  = ~A168 & ~A169;
  assign \new_[89205]_  = A170 & \new_[89204]_ ;
  assign \new_[89208]_  = A166 & ~A167;
  assign \new_[89211]_  = ~A200 & A199;
  assign \new_[89212]_  = \new_[89211]_  & \new_[89208]_ ;
  assign \new_[89213]_  = \new_[89212]_  & \new_[89205]_ ;
  assign \new_[89216]_  = A203 & A201;
  assign \new_[89219]_  = A266 & ~A265;
  assign \new_[89220]_  = \new_[89219]_  & \new_[89216]_ ;
  assign \new_[89223]_  = A269 & A267;
  assign \new_[89226]_  = ~A299 & ~A298;
  assign \new_[89227]_  = \new_[89226]_  & \new_[89223]_ ;
  assign \new_[89228]_  = \new_[89227]_  & \new_[89220]_ ;
  assign \new_[89232]_  = ~A168 & ~A169;
  assign \new_[89233]_  = A170 & \new_[89232]_ ;
  assign \new_[89236]_  = A166 & ~A167;
  assign \new_[89239]_  = ~A200 & A199;
  assign \new_[89240]_  = \new_[89239]_  & \new_[89236]_ ;
  assign \new_[89241]_  = \new_[89240]_  & \new_[89233]_ ;
  assign \new_[89244]_  = A203 & A201;
  assign \new_[89247]_  = ~A266 & A265;
  assign \new_[89248]_  = \new_[89247]_  & \new_[89244]_ ;
  assign \new_[89251]_  = A268 & A267;
  assign \new_[89254]_  = A301 & ~A300;
  assign \new_[89255]_  = \new_[89254]_  & \new_[89251]_ ;
  assign \new_[89256]_  = \new_[89255]_  & \new_[89248]_ ;
  assign \new_[89260]_  = ~A168 & ~A169;
  assign \new_[89261]_  = A170 & \new_[89260]_ ;
  assign \new_[89264]_  = A166 & ~A167;
  assign \new_[89267]_  = ~A200 & A199;
  assign \new_[89268]_  = \new_[89267]_  & \new_[89264]_ ;
  assign \new_[89269]_  = \new_[89268]_  & \new_[89261]_ ;
  assign \new_[89272]_  = A203 & A201;
  assign \new_[89275]_  = ~A266 & A265;
  assign \new_[89276]_  = \new_[89275]_  & \new_[89272]_ ;
  assign \new_[89279]_  = A268 & A267;
  assign \new_[89282]_  = A302 & ~A300;
  assign \new_[89283]_  = \new_[89282]_  & \new_[89279]_ ;
  assign \new_[89284]_  = \new_[89283]_  & \new_[89276]_ ;
  assign \new_[89288]_  = ~A168 & ~A169;
  assign \new_[89289]_  = A170 & \new_[89288]_ ;
  assign \new_[89292]_  = A166 & ~A167;
  assign \new_[89295]_  = ~A200 & A199;
  assign \new_[89296]_  = \new_[89295]_  & \new_[89292]_ ;
  assign \new_[89297]_  = \new_[89296]_  & \new_[89289]_ ;
  assign \new_[89300]_  = A203 & A201;
  assign \new_[89303]_  = ~A266 & A265;
  assign \new_[89304]_  = \new_[89303]_  & \new_[89300]_ ;
  assign \new_[89307]_  = A268 & A267;
  assign \new_[89310]_  = A299 & A298;
  assign \new_[89311]_  = \new_[89310]_  & \new_[89307]_ ;
  assign \new_[89312]_  = \new_[89311]_  & \new_[89304]_ ;
  assign \new_[89316]_  = ~A168 & ~A169;
  assign \new_[89317]_  = A170 & \new_[89316]_ ;
  assign \new_[89320]_  = A166 & ~A167;
  assign \new_[89323]_  = ~A200 & A199;
  assign \new_[89324]_  = \new_[89323]_  & \new_[89320]_ ;
  assign \new_[89325]_  = \new_[89324]_  & \new_[89317]_ ;
  assign \new_[89328]_  = A203 & A201;
  assign \new_[89331]_  = ~A266 & A265;
  assign \new_[89332]_  = \new_[89331]_  & \new_[89328]_ ;
  assign \new_[89335]_  = A268 & A267;
  assign \new_[89338]_  = ~A299 & ~A298;
  assign \new_[89339]_  = \new_[89338]_  & \new_[89335]_ ;
  assign \new_[89340]_  = \new_[89339]_  & \new_[89332]_ ;
  assign \new_[89344]_  = ~A168 & ~A169;
  assign \new_[89345]_  = A170 & \new_[89344]_ ;
  assign \new_[89348]_  = A166 & ~A167;
  assign \new_[89351]_  = ~A200 & A199;
  assign \new_[89352]_  = \new_[89351]_  & \new_[89348]_ ;
  assign \new_[89353]_  = \new_[89352]_  & \new_[89345]_ ;
  assign \new_[89356]_  = A203 & A201;
  assign \new_[89359]_  = ~A266 & A265;
  assign \new_[89360]_  = \new_[89359]_  & \new_[89356]_ ;
  assign \new_[89363]_  = A269 & A267;
  assign \new_[89366]_  = A301 & ~A300;
  assign \new_[89367]_  = \new_[89366]_  & \new_[89363]_ ;
  assign \new_[89368]_  = \new_[89367]_  & \new_[89360]_ ;
  assign \new_[89372]_  = ~A168 & ~A169;
  assign \new_[89373]_  = A170 & \new_[89372]_ ;
  assign \new_[89376]_  = A166 & ~A167;
  assign \new_[89379]_  = ~A200 & A199;
  assign \new_[89380]_  = \new_[89379]_  & \new_[89376]_ ;
  assign \new_[89381]_  = \new_[89380]_  & \new_[89373]_ ;
  assign \new_[89384]_  = A203 & A201;
  assign \new_[89387]_  = ~A266 & A265;
  assign \new_[89388]_  = \new_[89387]_  & \new_[89384]_ ;
  assign \new_[89391]_  = A269 & A267;
  assign \new_[89394]_  = A302 & ~A300;
  assign \new_[89395]_  = \new_[89394]_  & \new_[89391]_ ;
  assign \new_[89396]_  = \new_[89395]_  & \new_[89388]_ ;
  assign \new_[89400]_  = ~A168 & ~A169;
  assign \new_[89401]_  = A170 & \new_[89400]_ ;
  assign \new_[89404]_  = A166 & ~A167;
  assign \new_[89407]_  = ~A200 & A199;
  assign \new_[89408]_  = \new_[89407]_  & \new_[89404]_ ;
  assign \new_[89409]_  = \new_[89408]_  & \new_[89401]_ ;
  assign \new_[89412]_  = A203 & A201;
  assign \new_[89415]_  = ~A266 & A265;
  assign \new_[89416]_  = \new_[89415]_  & \new_[89412]_ ;
  assign \new_[89419]_  = A269 & A267;
  assign \new_[89422]_  = A299 & A298;
  assign \new_[89423]_  = \new_[89422]_  & \new_[89419]_ ;
  assign \new_[89424]_  = \new_[89423]_  & \new_[89416]_ ;
  assign \new_[89428]_  = ~A168 & ~A169;
  assign \new_[89429]_  = A170 & \new_[89428]_ ;
  assign \new_[89432]_  = A166 & ~A167;
  assign \new_[89435]_  = ~A200 & A199;
  assign \new_[89436]_  = \new_[89435]_  & \new_[89432]_ ;
  assign \new_[89437]_  = \new_[89436]_  & \new_[89429]_ ;
  assign \new_[89440]_  = A203 & A201;
  assign \new_[89443]_  = ~A266 & A265;
  assign \new_[89444]_  = \new_[89443]_  & \new_[89440]_ ;
  assign \new_[89447]_  = A269 & A267;
  assign \new_[89450]_  = ~A299 & ~A298;
  assign \new_[89451]_  = \new_[89450]_  & \new_[89447]_ ;
  assign \new_[89452]_  = \new_[89451]_  & \new_[89444]_ ;
  assign \new_[89456]_  = ~A168 & ~A169;
  assign \new_[89457]_  = A170 & \new_[89456]_ ;
  assign \new_[89460]_  = A166 & ~A167;
  assign \new_[89463]_  = ~A200 & ~A199;
  assign \new_[89464]_  = \new_[89463]_  & \new_[89460]_ ;
  assign \new_[89465]_  = \new_[89464]_  & \new_[89457]_ ;
  assign \new_[89468]_  = ~A268 & A267;
  assign \new_[89471]_  = A298 & ~A269;
  assign \new_[89472]_  = \new_[89471]_  & \new_[89468]_ ;
  assign \new_[89475]_  = ~A300 & ~A299;
  assign \new_[89478]_  = ~A302 & ~A301;
  assign \new_[89479]_  = \new_[89478]_  & \new_[89475]_ ;
  assign \new_[89480]_  = \new_[89479]_  & \new_[89472]_ ;
  assign \new_[89484]_  = ~A168 & ~A169;
  assign \new_[89485]_  = A170 & \new_[89484]_ ;
  assign \new_[89488]_  = A166 & ~A167;
  assign \new_[89491]_  = ~A200 & ~A199;
  assign \new_[89492]_  = \new_[89491]_  & \new_[89488]_ ;
  assign \new_[89493]_  = \new_[89492]_  & \new_[89485]_ ;
  assign \new_[89496]_  = ~A268 & A267;
  assign \new_[89499]_  = ~A298 & ~A269;
  assign \new_[89500]_  = \new_[89499]_  & \new_[89496]_ ;
  assign \new_[89503]_  = ~A300 & A299;
  assign \new_[89506]_  = ~A302 & ~A301;
  assign \new_[89507]_  = \new_[89506]_  & \new_[89503]_ ;
  assign \new_[89508]_  = \new_[89507]_  & \new_[89500]_ ;
  assign \new_[89511]_  = A168 & ~A170;
  assign \new_[89514]_  = ~A166 & A167;
  assign \new_[89515]_  = \new_[89514]_  & \new_[89511]_ ;
  assign \new_[89518]_  = A200 & ~A199;
  assign \new_[89521]_  = A202 & A201;
  assign \new_[89522]_  = \new_[89521]_  & \new_[89518]_ ;
  assign \new_[89523]_  = \new_[89522]_  & \new_[89515]_ ;
  assign \new_[89526]_  = A266 & ~A265;
  assign \new_[89529]_  = ~A268 & ~A267;
  assign \new_[89530]_  = \new_[89529]_  & \new_[89526]_ ;
  assign \new_[89533]_  = A300 & ~A269;
  assign \new_[89536]_  = ~A302 & ~A301;
  assign \new_[89537]_  = \new_[89536]_  & \new_[89533]_ ;
  assign \new_[89538]_  = \new_[89537]_  & \new_[89530]_ ;
  assign \new_[89541]_  = A168 & ~A170;
  assign \new_[89544]_  = ~A166 & A167;
  assign \new_[89545]_  = \new_[89544]_  & \new_[89541]_ ;
  assign \new_[89548]_  = A200 & ~A199;
  assign \new_[89551]_  = A202 & A201;
  assign \new_[89552]_  = \new_[89551]_  & \new_[89548]_ ;
  assign \new_[89553]_  = \new_[89552]_  & \new_[89545]_ ;
  assign \new_[89556]_  = ~A266 & A265;
  assign \new_[89559]_  = ~A268 & ~A267;
  assign \new_[89560]_  = \new_[89559]_  & \new_[89556]_ ;
  assign \new_[89563]_  = A300 & ~A269;
  assign \new_[89566]_  = ~A302 & ~A301;
  assign \new_[89567]_  = \new_[89566]_  & \new_[89563]_ ;
  assign \new_[89568]_  = \new_[89567]_  & \new_[89560]_ ;
  assign \new_[89571]_  = A168 & ~A170;
  assign \new_[89574]_  = ~A166 & A167;
  assign \new_[89575]_  = \new_[89574]_  & \new_[89571]_ ;
  assign \new_[89578]_  = A200 & ~A199;
  assign \new_[89581]_  = A203 & A201;
  assign \new_[89582]_  = \new_[89581]_  & \new_[89578]_ ;
  assign \new_[89583]_  = \new_[89582]_  & \new_[89575]_ ;
  assign \new_[89586]_  = A266 & ~A265;
  assign \new_[89589]_  = ~A268 & ~A267;
  assign \new_[89590]_  = \new_[89589]_  & \new_[89586]_ ;
  assign \new_[89593]_  = A300 & ~A269;
  assign \new_[89596]_  = ~A302 & ~A301;
  assign \new_[89597]_  = \new_[89596]_  & \new_[89593]_ ;
  assign \new_[89598]_  = \new_[89597]_  & \new_[89590]_ ;
  assign \new_[89601]_  = A168 & ~A170;
  assign \new_[89604]_  = ~A166 & A167;
  assign \new_[89605]_  = \new_[89604]_  & \new_[89601]_ ;
  assign \new_[89608]_  = A200 & ~A199;
  assign \new_[89611]_  = A203 & A201;
  assign \new_[89612]_  = \new_[89611]_  & \new_[89608]_ ;
  assign \new_[89613]_  = \new_[89612]_  & \new_[89605]_ ;
  assign \new_[89616]_  = ~A266 & A265;
  assign \new_[89619]_  = ~A268 & ~A267;
  assign \new_[89620]_  = \new_[89619]_  & \new_[89616]_ ;
  assign \new_[89623]_  = A300 & ~A269;
  assign \new_[89626]_  = ~A302 & ~A301;
  assign \new_[89627]_  = \new_[89626]_  & \new_[89623]_ ;
  assign \new_[89628]_  = \new_[89627]_  & \new_[89620]_ ;
  assign \new_[89631]_  = A168 & ~A170;
  assign \new_[89634]_  = ~A166 & A167;
  assign \new_[89635]_  = \new_[89634]_  & \new_[89631]_ ;
  assign \new_[89638]_  = A200 & ~A199;
  assign \new_[89641]_  = ~A202 & ~A201;
  assign \new_[89642]_  = \new_[89641]_  & \new_[89638]_ ;
  assign \new_[89643]_  = \new_[89642]_  & \new_[89635]_ ;
  assign \new_[89646]_  = ~A265 & ~A203;
  assign \new_[89649]_  = A267 & A266;
  assign \new_[89650]_  = \new_[89649]_  & \new_[89646]_ ;
  assign \new_[89653]_  = A300 & A268;
  assign \new_[89656]_  = ~A302 & ~A301;
  assign \new_[89657]_  = \new_[89656]_  & \new_[89653]_ ;
  assign \new_[89658]_  = \new_[89657]_  & \new_[89650]_ ;
  assign \new_[89661]_  = A168 & ~A170;
  assign \new_[89664]_  = ~A166 & A167;
  assign \new_[89665]_  = \new_[89664]_  & \new_[89661]_ ;
  assign \new_[89668]_  = A200 & ~A199;
  assign \new_[89671]_  = ~A202 & ~A201;
  assign \new_[89672]_  = \new_[89671]_  & \new_[89668]_ ;
  assign \new_[89673]_  = \new_[89672]_  & \new_[89665]_ ;
  assign \new_[89676]_  = ~A265 & ~A203;
  assign \new_[89679]_  = A267 & A266;
  assign \new_[89680]_  = \new_[89679]_  & \new_[89676]_ ;
  assign \new_[89683]_  = A300 & A269;
  assign \new_[89686]_  = ~A302 & ~A301;
  assign \new_[89687]_  = \new_[89686]_  & \new_[89683]_ ;
  assign \new_[89688]_  = \new_[89687]_  & \new_[89680]_ ;
  assign \new_[89691]_  = A168 & ~A170;
  assign \new_[89694]_  = ~A166 & A167;
  assign \new_[89695]_  = \new_[89694]_  & \new_[89691]_ ;
  assign \new_[89698]_  = A200 & ~A199;
  assign \new_[89701]_  = ~A202 & ~A201;
  assign \new_[89702]_  = \new_[89701]_  & \new_[89698]_ ;
  assign \new_[89703]_  = \new_[89702]_  & \new_[89695]_ ;
  assign \new_[89706]_  = ~A265 & ~A203;
  assign \new_[89709]_  = ~A267 & A266;
  assign \new_[89710]_  = \new_[89709]_  & \new_[89706]_ ;
  assign \new_[89713]_  = ~A269 & ~A268;
  assign \new_[89716]_  = A301 & ~A300;
  assign \new_[89717]_  = \new_[89716]_  & \new_[89713]_ ;
  assign \new_[89718]_  = \new_[89717]_  & \new_[89710]_ ;
  assign \new_[89721]_  = A168 & ~A170;
  assign \new_[89724]_  = ~A166 & A167;
  assign \new_[89725]_  = \new_[89724]_  & \new_[89721]_ ;
  assign \new_[89728]_  = A200 & ~A199;
  assign \new_[89731]_  = ~A202 & ~A201;
  assign \new_[89732]_  = \new_[89731]_  & \new_[89728]_ ;
  assign \new_[89733]_  = \new_[89732]_  & \new_[89725]_ ;
  assign \new_[89736]_  = ~A265 & ~A203;
  assign \new_[89739]_  = ~A267 & A266;
  assign \new_[89740]_  = \new_[89739]_  & \new_[89736]_ ;
  assign \new_[89743]_  = ~A269 & ~A268;
  assign \new_[89746]_  = A302 & ~A300;
  assign \new_[89747]_  = \new_[89746]_  & \new_[89743]_ ;
  assign \new_[89748]_  = \new_[89747]_  & \new_[89740]_ ;
  assign \new_[89751]_  = A168 & ~A170;
  assign \new_[89754]_  = ~A166 & A167;
  assign \new_[89755]_  = \new_[89754]_  & \new_[89751]_ ;
  assign \new_[89758]_  = A200 & ~A199;
  assign \new_[89761]_  = ~A202 & ~A201;
  assign \new_[89762]_  = \new_[89761]_  & \new_[89758]_ ;
  assign \new_[89763]_  = \new_[89762]_  & \new_[89755]_ ;
  assign \new_[89766]_  = ~A265 & ~A203;
  assign \new_[89769]_  = ~A267 & A266;
  assign \new_[89770]_  = \new_[89769]_  & \new_[89766]_ ;
  assign \new_[89773]_  = ~A269 & ~A268;
  assign \new_[89776]_  = A299 & A298;
  assign \new_[89777]_  = \new_[89776]_  & \new_[89773]_ ;
  assign \new_[89778]_  = \new_[89777]_  & \new_[89770]_ ;
  assign \new_[89781]_  = A168 & ~A170;
  assign \new_[89784]_  = ~A166 & A167;
  assign \new_[89785]_  = \new_[89784]_  & \new_[89781]_ ;
  assign \new_[89788]_  = A200 & ~A199;
  assign \new_[89791]_  = ~A202 & ~A201;
  assign \new_[89792]_  = \new_[89791]_  & \new_[89788]_ ;
  assign \new_[89793]_  = \new_[89792]_  & \new_[89785]_ ;
  assign \new_[89796]_  = ~A265 & ~A203;
  assign \new_[89799]_  = ~A267 & A266;
  assign \new_[89800]_  = \new_[89799]_  & \new_[89796]_ ;
  assign \new_[89803]_  = ~A269 & ~A268;
  assign \new_[89806]_  = ~A299 & ~A298;
  assign \new_[89807]_  = \new_[89806]_  & \new_[89803]_ ;
  assign \new_[89808]_  = \new_[89807]_  & \new_[89800]_ ;
  assign \new_[89811]_  = A168 & ~A170;
  assign \new_[89814]_  = ~A166 & A167;
  assign \new_[89815]_  = \new_[89814]_  & \new_[89811]_ ;
  assign \new_[89818]_  = A200 & ~A199;
  assign \new_[89821]_  = ~A202 & ~A201;
  assign \new_[89822]_  = \new_[89821]_  & \new_[89818]_ ;
  assign \new_[89823]_  = \new_[89822]_  & \new_[89815]_ ;
  assign \new_[89826]_  = A265 & ~A203;
  assign \new_[89829]_  = A267 & ~A266;
  assign \new_[89830]_  = \new_[89829]_  & \new_[89826]_ ;
  assign \new_[89833]_  = A300 & A268;
  assign \new_[89836]_  = ~A302 & ~A301;
  assign \new_[89837]_  = \new_[89836]_  & \new_[89833]_ ;
  assign \new_[89838]_  = \new_[89837]_  & \new_[89830]_ ;
  assign \new_[89841]_  = A168 & ~A170;
  assign \new_[89844]_  = ~A166 & A167;
  assign \new_[89845]_  = \new_[89844]_  & \new_[89841]_ ;
  assign \new_[89848]_  = A200 & ~A199;
  assign \new_[89851]_  = ~A202 & ~A201;
  assign \new_[89852]_  = \new_[89851]_  & \new_[89848]_ ;
  assign \new_[89853]_  = \new_[89852]_  & \new_[89845]_ ;
  assign \new_[89856]_  = A265 & ~A203;
  assign \new_[89859]_  = A267 & ~A266;
  assign \new_[89860]_  = \new_[89859]_  & \new_[89856]_ ;
  assign \new_[89863]_  = A300 & A269;
  assign \new_[89866]_  = ~A302 & ~A301;
  assign \new_[89867]_  = \new_[89866]_  & \new_[89863]_ ;
  assign \new_[89868]_  = \new_[89867]_  & \new_[89860]_ ;
  assign \new_[89871]_  = A168 & ~A170;
  assign \new_[89874]_  = ~A166 & A167;
  assign \new_[89875]_  = \new_[89874]_  & \new_[89871]_ ;
  assign \new_[89878]_  = A200 & ~A199;
  assign \new_[89881]_  = ~A202 & ~A201;
  assign \new_[89882]_  = \new_[89881]_  & \new_[89878]_ ;
  assign \new_[89883]_  = \new_[89882]_  & \new_[89875]_ ;
  assign \new_[89886]_  = A265 & ~A203;
  assign \new_[89889]_  = ~A267 & ~A266;
  assign \new_[89890]_  = \new_[89889]_  & \new_[89886]_ ;
  assign \new_[89893]_  = ~A269 & ~A268;
  assign \new_[89896]_  = A301 & ~A300;
  assign \new_[89897]_  = \new_[89896]_  & \new_[89893]_ ;
  assign \new_[89898]_  = \new_[89897]_  & \new_[89890]_ ;
  assign \new_[89901]_  = A168 & ~A170;
  assign \new_[89904]_  = ~A166 & A167;
  assign \new_[89905]_  = \new_[89904]_  & \new_[89901]_ ;
  assign \new_[89908]_  = A200 & ~A199;
  assign \new_[89911]_  = ~A202 & ~A201;
  assign \new_[89912]_  = \new_[89911]_  & \new_[89908]_ ;
  assign \new_[89913]_  = \new_[89912]_  & \new_[89905]_ ;
  assign \new_[89916]_  = A265 & ~A203;
  assign \new_[89919]_  = ~A267 & ~A266;
  assign \new_[89920]_  = \new_[89919]_  & \new_[89916]_ ;
  assign \new_[89923]_  = ~A269 & ~A268;
  assign \new_[89926]_  = A302 & ~A300;
  assign \new_[89927]_  = \new_[89926]_  & \new_[89923]_ ;
  assign \new_[89928]_  = \new_[89927]_  & \new_[89920]_ ;
  assign \new_[89931]_  = A168 & ~A170;
  assign \new_[89934]_  = ~A166 & A167;
  assign \new_[89935]_  = \new_[89934]_  & \new_[89931]_ ;
  assign \new_[89938]_  = A200 & ~A199;
  assign \new_[89941]_  = ~A202 & ~A201;
  assign \new_[89942]_  = \new_[89941]_  & \new_[89938]_ ;
  assign \new_[89943]_  = \new_[89942]_  & \new_[89935]_ ;
  assign \new_[89946]_  = A265 & ~A203;
  assign \new_[89949]_  = ~A267 & ~A266;
  assign \new_[89950]_  = \new_[89949]_  & \new_[89946]_ ;
  assign \new_[89953]_  = ~A269 & ~A268;
  assign \new_[89956]_  = A299 & A298;
  assign \new_[89957]_  = \new_[89956]_  & \new_[89953]_ ;
  assign \new_[89958]_  = \new_[89957]_  & \new_[89950]_ ;
  assign \new_[89961]_  = A168 & ~A170;
  assign \new_[89964]_  = ~A166 & A167;
  assign \new_[89965]_  = \new_[89964]_  & \new_[89961]_ ;
  assign \new_[89968]_  = A200 & ~A199;
  assign \new_[89971]_  = ~A202 & ~A201;
  assign \new_[89972]_  = \new_[89971]_  & \new_[89968]_ ;
  assign \new_[89973]_  = \new_[89972]_  & \new_[89965]_ ;
  assign \new_[89976]_  = A265 & ~A203;
  assign \new_[89979]_  = ~A267 & ~A266;
  assign \new_[89980]_  = \new_[89979]_  & \new_[89976]_ ;
  assign \new_[89983]_  = ~A269 & ~A268;
  assign \new_[89986]_  = ~A299 & ~A298;
  assign \new_[89987]_  = \new_[89986]_  & \new_[89983]_ ;
  assign \new_[89988]_  = \new_[89987]_  & \new_[89980]_ ;
  assign \new_[89991]_  = A168 & ~A170;
  assign \new_[89994]_  = ~A166 & A167;
  assign \new_[89995]_  = \new_[89994]_  & \new_[89991]_ ;
  assign \new_[89998]_  = ~A200 & A199;
  assign \new_[90001]_  = A202 & A201;
  assign \new_[90002]_  = \new_[90001]_  & \new_[89998]_ ;
  assign \new_[90003]_  = \new_[90002]_  & \new_[89995]_ ;
  assign \new_[90006]_  = A266 & ~A265;
  assign \new_[90009]_  = ~A268 & ~A267;
  assign \new_[90010]_  = \new_[90009]_  & \new_[90006]_ ;
  assign \new_[90013]_  = A300 & ~A269;
  assign \new_[90016]_  = ~A302 & ~A301;
  assign \new_[90017]_  = \new_[90016]_  & \new_[90013]_ ;
  assign \new_[90018]_  = \new_[90017]_  & \new_[90010]_ ;
  assign \new_[90021]_  = A168 & ~A170;
  assign \new_[90024]_  = ~A166 & A167;
  assign \new_[90025]_  = \new_[90024]_  & \new_[90021]_ ;
  assign \new_[90028]_  = ~A200 & A199;
  assign \new_[90031]_  = A202 & A201;
  assign \new_[90032]_  = \new_[90031]_  & \new_[90028]_ ;
  assign \new_[90033]_  = \new_[90032]_  & \new_[90025]_ ;
  assign \new_[90036]_  = ~A266 & A265;
  assign \new_[90039]_  = ~A268 & ~A267;
  assign \new_[90040]_  = \new_[90039]_  & \new_[90036]_ ;
  assign \new_[90043]_  = A300 & ~A269;
  assign \new_[90046]_  = ~A302 & ~A301;
  assign \new_[90047]_  = \new_[90046]_  & \new_[90043]_ ;
  assign \new_[90048]_  = \new_[90047]_  & \new_[90040]_ ;
  assign \new_[90051]_  = A168 & ~A170;
  assign \new_[90054]_  = ~A166 & A167;
  assign \new_[90055]_  = \new_[90054]_  & \new_[90051]_ ;
  assign \new_[90058]_  = ~A200 & A199;
  assign \new_[90061]_  = A203 & A201;
  assign \new_[90062]_  = \new_[90061]_  & \new_[90058]_ ;
  assign \new_[90063]_  = \new_[90062]_  & \new_[90055]_ ;
  assign \new_[90066]_  = A266 & ~A265;
  assign \new_[90069]_  = ~A268 & ~A267;
  assign \new_[90070]_  = \new_[90069]_  & \new_[90066]_ ;
  assign \new_[90073]_  = A300 & ~A269;
  assign \new_[90076]_  = ~A302 & ~A301;
  assign \new_[90077]_  = \new_[90076]_  & \new_[90073]_ ;
  assign \new_[90078]_  = \new_[90077]_  & \new_[90070]_ ;
  assign \new_[90081]_  = A168 & ~A170;
  assign \new_[90084]_  = ~A166 & A167;
  assign \new_[90085]_  = \new_[90084]_  & \new_[90081]_ ;
  assign \new_[90088]_  = ~A200 & A199;
  assign \new_[90091]_  = A203 & A201;
  assign \new_[90092]_  = \new_[90091]_  & \new_[90088]_ ;
  assign \new_[90093]_  = \new_[90092]_  & \new_[90085]_ ;
  assign \new_[90096]_  = ~A266 & A265;
  assign \new_[90099]_  = ~A268 & ~A267;
  assign \new_[90100]_  = \new_[90099]_  & \new_[90096]_ ;
  assign \new_[90103]_  = A300 & ~A269;
  assign \new_[90106]_  = ~A302 & ~A301;
  assign \new_[90107]_  = \new_[90106]_  & \new_[90103]_ ;
  assign \new_[90108]_  = \new_[90107]_  & \new_[90100]_ ;
  assign \new_[90111]_  = A168 & ~A170;
  assign \new_[90114]_  = ~A166 & A167;
  assign \new_[90115]_  = \new_[90114]_  & \new_[90111]_ ;
  assign \new_[90118]_  = ~A200 & A199;
  assign \new_[90121]_  = ~A202 & ~A201;
  assign \new_[90122]_  = \new_[90121]_  & \new_[90118]_ ;
  assign \new_[90123]_  = \new_[90122]_  & \new_[90115]_ ;
  assign \new_[90126]_  = ~A265 & ~A203;
  assign \new_[90129]_  = A267 & A266;
  assign \new_[90130]_  = \new_[90129]_  & \new_[90126]_ ;
  assign \new_[90133]_  = A300 & A268;
  assign \new_[90136]_  = ~A302 & ~A301;
  assign \new_[90137]_  = \new_[90136]_  & \new_[90133]_ ;
  assign \new_[90138]_  = \new_[90137]_  & \new_[90130]_ ;
  assign \new_[90141]_  = A168 & ~A170;
  assign \new_[90144]_  = ~A166 & A167;
  assign \new_[90145]_  = \new_[90144]_  & \new_[90141]_ ;
  assign \new_[90148]_  = ~A200 & A199;
  assign \new_[90151]_  = ~A202 & ~A201;
  assign \new_[90152]_  = \new_[90151]_  & \new_[90148]_ ;
  assign \new_[90153]_  = \new_[90152]_  & \new_[90145]_ ;
  assign \new_[90156]_  = ~A265 & ~A203;
  assign \new_[90159]_  = A267 & A266;
  assign \new_[90160]_  = \new_[90159]_  & \new_[90156]_ ;
  assign \new_[90163]_  = A300 & A269;
  assign \new_[90166]_  = ~A302 & ~A301;
  assign \new_[90167]_  = \new_[90166]_  & \new_[90163]_ ;
  assign \new_[90168]_  = \new_[90167]_  & \new_[90160]_ ;
  assign \new_[90171]_  = A168 & ~A170;
  assign \new_[90174]_  = ~A166 & A167;
  assign \new_[90175]_  = \new_[90174]_  & \new_[90171]_ ;
  assign \new_[90178]_  = ~A200 & A199;
  assign \new_[90181]_  = ~A202 & ~A201;
  assign \new_[90182]_  = \new_[90181]_  & \new_[90178]_ ;
  assign \new_[90183]_  = \new_[90182]_  & \new_[90175]_ ;
  assign \new_[90186]_  = ~A265 & ~A203;
  assign \new_[90189]_  = ~A267 & A266;
  assign \new_[90190]_  = \new_[90189]_  & \new_[90186]_ ;
  assign \new_[90193]_  = ~A269 & ~A268;
  assign \new_[90196]_  = A301 & ~A300;
  assign \new_[90197]_  = \new_[90196]_  & \new_[90193]_ ;
  assign \new_[90198]_  = \new_[90197]_  & \new_[90190]_ ;
  assign \new_[90201]_  = A168 & ~A170;
  assign \new_[90204]_  = ~A166 & A167;
  assign \new_[90205]_  = \new_[90204]_  & \new_[90201]_ ;
  assign \new_[90208]_  = ~A200 & A199;
  assign \new_[90211]_  = ~A202 & ~A201;
  assign \new_[90212]_  = \new_[90211]_  & \new_[90208]_ ;
  assign \new_[90213]_  = \new_[90212]_  & \new_[90205]_ ;
  assign \new_[90216]_  = ~A265 & ~A203;
  assign \new_[90219]_  = ~A267 & A266;
  assign \new_[90220]_  = \new_[90219]_  & \new_[90216]_ ;
  assign \new_[90223]_  = ~A269 & ~A268;
  assign \new_[90226]_  = A302 & ~A300;
  assign \new_[90227]_  = \new_[90226]_  & \new_[90223]_ ;
  assign \new_[90228]_  = \new_[90227]_  & \new_[90220]_ ;
  assign \new_[90231]_  = A168 & ~A170;
  assign \new_[90234]_  = ~A166 & A167;
  assign \new_[90235]_  = \new_[90234]_  & \new_[90231]_ ;
  assign \new_[90238]_  = ~A200 & A199;
  assign \new_[90241]_  = ~A202 & ~A201;
  assign \new_[90242]_  = \new_[90241]_  & \new_[90238]_ ;
  assign \new_[90243]_  = \new_[90242]_  & \new_[90235]_ ;
  assign \new_[90246]_  = ~A265 & ~A203;
  assign \new_[90249]_  = ~A267 & A266;
  assign \new_[90250]_  = \new_[90249]_  & \new_[90246]_ ;
  assign \new_[90253]_  = ~A269 & ~A268;
  assign \new_[90256]_  = A299 & A298;
  assign \new_[90257]_  = \new_[90256]_  & \new_[90253]_ ;
  assign \new_[90258]_  = \new_[90257]_  & \new_[90250]_ ;
  assign \new_[90261]_  = A168 & ~A170;
  assign \new_[90264]_  = ~A166 & A167;
  assign \new_[90265]_  = \new_[90264]_  & \new_[90261]_ ;
  assign \new_[90268]_  = ~A200 & A199;
  assign \new_[90271]_  = ~A202 & ~A201;
  assign \new_[90272]_  = \new_[90271]_  & \new_[90268]_ ;
  assign \new_[90273]_  = \new_[90272]_  & \new_[90265]_ ;
  assign \new_[90276]_  = ~A265 & ~A203;
  assign \new_[90279]_  = ~A267 & A266;
  assign \new_[90280]_  = \new_[90279]_  & \new_[90276]_ ;
  assign \new_[90283]_  = ~A269 & ~A268;
  assign \new_[90286]_  = ~A299 & ~A298;
  assign \new_[90287]_  = \new_[90286]_  & \new_[90283]_ ;
  assign \new_[90288]_  = \new_[90287]_  & \new_[90280]_ ;
  assign \new_[90291]_  = A168 & ~A170;
  assign \new_[90294]_  = ~A166 & A167;
  assign \new_[90295]_  = \new_[90294]_  & \new_[90291]_ ;
  assign \new_[90298]_  = ~A200 & A199;
  assign \new_[90301]_  = ~A202 & ~A201;
  assign \new_[90302]_  = \new_[90301]_  & \new_[90298]_ ;
  assign \new_[90303]_  = \new_[90302]_  & \new_[90295]_ ;
  assign \new_[90306]_  = A265 & ~A203;
  assign \new_[90309]_  = A267 & ~A266;
  assign \new_[90310]_  = \new_[90309]_  & \new_[90306]_ ;
  assign \new_[90313]_  = A300 & A268;
  assign \new_[90316]_  = ~A302 & ~A301;
  assign \new_[90317]_  = \new_[90316]_  & \new_[90313]_ ;
  assign \new_[90318]_  = \new_[90317]_  & \new_[90310]_ ;
  assign \new_[90321]_  = A168 & ~A170;
  assign \new_[90324]_  = ~A166 & A167;
  assign \new_[90325]_  = \new_[90324]_  & \new_[90321]_ ;
  assign \new_[90328]_  = ~A200 & A199;
  assign \new_[90331]_  = ~A202 & ~A201;
  assign \new_[90332]_  = \new_[90331]_  & \new_[90328]_ ;
  assign \new_[90333]_  = \new_[90332]_  & \new_[90325]_ ;
  assign \new_[90336]_  = A265 & ~A203;
  assign \new_[90339]_  = A267 & ~A266;
  assign \new_[90340]_  = \new_[90339]_  & \new_[90336]_ ;
  assign \new_[90343]_  = A300 & A269;
  assign \new_[90346]_  = ~A302 & ~A301;
  assign \new_[90347]_  = \new_[90346]_  & \new_[90343]_ ;
  assign \new_[90348]_  = \new_[90347]_  & \new_[90340]_ ;
  assign \new_[90351]_  = A168 & ~A170;
  assign \new_[90354]_  = ~A166 & A167;
  assign \new_[90355]_  = \new_[90354]_  & \new_[90351]_ ;
  assign \new_[90358]_  = ~A200 & A199;
  assign \new_[90361]_  = ~A202 & ~A201;
  assign \new_[90362]_  = \new_[90361]_  & \new_[90358]_ ;
  assign \new_[90363]_  = \new_[90362]_  & \new_[90355]_ ;
  assign \new_[90366]_  = A265 & ~A203;
  assign \new_[90369]_  = ~A267 & ~A266;
  assign \new_[90370]_  = \new_[90369]_  & \new_[90366]_ ;
  assign \new_[90373]_  = ~A269 & ~A268;
  assign \new_[90376]_  = A301 & ~A300;
  assign \new_[90377]_  = \new_[90376]_  & \new_[90373]_ ;
  assign \new_[90378]_  = \new_[90377]_  & \new_[90370]_ ;
  assign \new_[90381]_  = A168 & ~A170;
  assign \new_[90384]_  = ~A166 & A167;
  assign \new_[90385]_  = \new_[90384]_  & \new_[90381]_ ;
  assign \new_[90388]_  = ~A200 & A199;
  assign \new_[90391]_  = ~A202 & ~A201;
  assign \new_[90392]_  = \new_[90391]_  & \new_[90388]_ ;
  assign \new_[90393]_  = \new_[90392]_  & \new_[90385]_ ;
  assign \new_[90396]_  = A265 & ~A203;
  assign \new_[90399]_  = ~A267 & ~A266;
  assign \new_[90400]_  = \new_[90399]_  & \new_[90396]_ ;
  assign \new_[90403]_  = ~A269 & ~A268;
  assign \new_[90406]_  = A302 & ~A300;
  assign \new_[90407]_  = \new_[90406]_  & \new_[90403]_ ;
  assign \new_[90408]_  = \new_[90407]_  & \new_[90400]_ ;
  assign \new_[90411]_  = A168 & ~A170;
  assign \new_[90414]_  = ~A166 & A167;
  assign \new_[90415]_  = \new_[90414]_  & \new_[90411]_ ;
  assign \new_[90418]_  = ~A200 & A199;
  assign \new_[90421]_  = ~A202 & ~A201;
  assign \new_[90422]_  = \new_[90421]_  & \new_[90418]_ ;
  assign \new_[90423]_  = \new_[90422]_  & \new_[90415]_ ;
  assign \new_[90426]_  = A265 & ~A203;
  assign \new_[90429]_  = ~A267 & ~A266;
  assign \new_[90430]_  = \new_[90429]_  & \new_[90426]_ ;
  assign \new_[90433]_  = ~A269 & ~A268;
  assign \new_[90436]_  = A299 & A298;
  assign \new_[90437]_  = \new_[90436]_  & \new_[90433]_ ;
  assign \new_[90438]_  = \new_[90437]_  & \new_[90430]_ ;
  assign \new_[90441]_  = A168 & ~A170;
  assign \new_[90444]_  = ~A166 & A167;
  assign \new_[90445]_  = \new_[90444]_  & \new_[90441]_ ;
  assign \new_[90448]_  = ~A200 & A199;
  assign \new_[90451]_  = ~A202 & ~A201;
  assign \new_[90452]_  = \new_[90451]_  & \new_[90448]_ ;
  assign \new_[90453]_  = \new_[90452]_  & \new_[90445]_ ;
  assign \new_[90456]_  = A265 & ~A203;
  assign \new_[90459]_  = ~A267 & ~A266;
  assign \new_[90460]_  = \new_[90459]_  & \new_[90456]_ ;
  assign \new_[90463]_  = ~A269 & ~A268;
  assign \new_[90466]_  = ~A299 & ~A298;
  assign \new_[90467]_  = \new_[90466]_  & \new_[90463]_ ;
  assign \new_[90468]_  = \new_[90467]_  & \new_[90460]_ ;
  assign \new_[90471]_  = A168 & ~A170;
  assign \new_[90474]_  = A166 & ~A167;
  assign \new_[90475]_  = \new_[90474]_  & \new_[90471]_ ;
  assign \new_[90478]_  = A200 & ~A199;
  assign \new_[90481]_  = A202 & A201;
  assign \new_[90482]_  = \new_[90481]_  & \new_[90478]_ ;
  assign \new_[90483]_  = \new_[90482]_  & \new_[90475]_ ;
  assign \new_[90486]_  = A266 & ~A265;
  assign \new_[90489]_  = ~A268 & ~A267;
  assign \new_[90490]_  = \new_[90489]_  & \new_[90486]_ ;
  assign \new_[90493]_  = A300 & ~A269;
  assign \new_[90496]_  = ~A302 & ~A301;
  assign \new_[90497]_  = \new_[90496]_  & \new_[90493]_ ;
  assign \new_[90498]_  = \new_[90497]_  & \new_[90490]_ ;
  assign \new_[90501]_  = A168 & ~A170;
  assign \new_[90504]_  = A166 & ~A167;
  assign \new_[90505]_  = \new_[90504]_  & \new_[90501]_ ;
  assign \new_[90508]_  = A200 & ~A199;
  assign \new_[90511]_  = A202 & A201;
  assign \new_[90512]_  = \new_[90511]_  & \new_[90508]_ ;
  assign \new_[90513]_  = \new_[90512]_  & \new_[90505]_ ;
  assign \new_[90516]_  = ~A266 & A265;
  assign \new_[90519]_  = ~A268 & ~A267;
  assign \new_[90520]_  = \new_[90519]_  & \new_[90516]_ ;
  assign \new_[90523]_  = A300 & ~A269;
  assign \new_[90526]_  = ~A302 & ~A301;
  assign \new_[90527]_  = \new_[90526]_  & \new_[90523]_ ;
  assign \new_[90528]_  = \new_[90527]_  & \new_[90520]_ ;
  assign \new_[90531]_  = A168 & ~A170;
  assign \new_[90534]_  = A166 & ~A167;
  assign \new_[90535]_  = \new_[90534]_  & \new_[90531]_ ;
  assign \new_[90538]_  = A200 & ~A199;
  assign \new_[90541]_  = A203 & A201;
  assign \new_[90542]_  = \new_[90541]_  & \new_[90538]_ ;
  assign \new_[90543]_  = \new_[90542]_  & \new_[90535]_ ;
  assign \new_[90546]_  = A266 & ~A265;
  assign \new_[90549]_  = ~A268 & ~A267;
  assign \new_[90550]_  = \new_[90549]_  & \new_[90546]_ ;
  assign \new_[90553]_  = A300 & ~A269;
  assign \new_[90556]_  = ~A302 & ~A301;
  assign \new_[90557]_  = \new_[90556]_  & \new_[90553]_ ;
  assign \new_[90558]_  = \new_[90557]_  & \new_[90550]_ ;
  assign \new_[90561]_  = A168 & ~A170;
  assign \new_[90564]_  = A166 & ~A167;
  assign \new_[90565]_  = \new_[90564]_  & \new_[90561]_ ;
  assign \new_[90568]_  = A200 & ~A199;
  assign \new_[90571]_  = A203 & A201;
  assign \new_[90572]_  = \new_[90571]_  & \new_[90568]_ ;
  assign \new_[90573]_  = \new_[90572]_  & \new_[90565]_ ;
  assign \new_[90576]_  = ~A266 & A265;
  assign \new_[90579]_  = ~A268 & ~A267;
  assign \new_[90580]_  = \new_[90579]_  & \new_[90576]_ ;
  assign \new_[90583]_  = A300 & ~A269;
  assign \new_[90586]_  = ~A302 & ~A301;
  assign \new_[90587]_  = \new_[90586]_  & \new_[90583]_ ;
  assign \new_[90588]_  = \new_[90587]_  & \new_[90580]_ ;
  assign \new_[90591]_  = A168 & ~A170;
  assign \new_[90594]_  = A166 & ~A167;
  assign \new_[90595]_  = \new_[90594]_  & \new_[90591]_ ;
  assign \new_[90598]_  = A200 & ~A199;
  assign \new_[90601]_  = ~A202 & ~A201;
  assign \new_[90602]_  = \new_[90601]_  & \new_[90598]_ ;
  assign \new_[90603]_  = \new_[90602]_  & \new_[90595]_ ;
  assign \new_[90606]_  = ~A265 & ~A203;
  assign \new_[90609]_  = A267 & A266;
  assign \new_[90610]_  = \new_[90609]_  & \new_[90606]_ ;
  assign \new_[90613]_  = A300 & A268;
  assign \new_[90616]_  = ~A302 & ~A301;
  assign \new_[90617]_  = \new_[90616]_  & \new_[90613]_ ;
  assign \new_[90618]_  = \new_[90617]_  & \new_[90610]_ ;
  assign \new_[90621]_  = A168 & ~A170;
  assign \new_[90624]_  = A166 & ~A167;
  assign \new_[90625]_  = \new_[90624]_  & \new_[90621]_ ;
  assign \new_[90628]_  = A200 & ~A199;
  assign \new_[90631]_  = ~A202 & ~A201;
  assign \new_[90632]_  = \new_[90631]_  & \new_[90628]_ ;
  assign \new_[90633]_  = \new_[90632]_  & \new_[90625]_ ;
  assign \new_[90636]_  = ~A265 & ~A203;
  assign \new_[90639]_  = A267 & A266;
  assign \new_[90640]_  = \new_[90639]_  & \new_[90636]_ ;
  assign \new_[90643]_  = A300 & A269;
  assign \new_[90646]_  = ~A302 & ~A301;
  assign \new_[90647]_  = \new_[90646]_  & \new_[90643]_ ;
  assign \new_[90648]_  = \new_[90647]_  & \new_[90640]_ ;
  assign \new_[90651]_  = A168 & ~A170;
  assign \new_[90654]_  = A166 & ~A167;
  assign \new_[90655]_  = \new_[90654]_  & \new_[90651]_ ;
  assign \new_[90658]_  = A200 & ~A199;
  assign \new_[90661]_  = ~A202 & ~A201;
  assign \new_[90662]_  = \new_[90661]_  & \new_[90658]_ ;
  assign \new_[90663]_  = \new_[90662]_  & \new_[90655]_ ;
  assign \new_[90666]_  = ~A265 & ~A203;
  assign \new_[90669]_  = ~A267 & A266;
  assign \new_[90670]_  = \new_[90669]_  & \new_[90666]_ ;
  assign \new_[90673]_  = ~A269 & ~A268;
  assign \new_[90676]_  = A301 & ~A300;
  assign \new_[90677]_  = \new_[90676]_  & \new_[90673]_ ;
  assign \new_[90678]_  = \new_[90677]_  & \new_[90670]_ ;
  assign \new_[90681]_  = A168 & ~A170;
  assign \new_[90684]_  = A166 & ~A167;
  assign \new_[90685]_  = \new_[90684]_  & \new_[90681]_ ;
  assign \new_[90688]_  = A200 & ~A199;
  assign \new_[90691]_  = ~A202 & ~A201;
  assign \new_[90692]_  = \new_[90691]_  & \new_[90688]_ ;
  assign \new_[90693]_  = \new_[90692]_  & \new_[90685]_ ;
  assign \new_[90696]_  = ~A265 & ~A203;
  assign \new_[90699]_  = ~A267 & A266;
  assign \new_[90700]_  = \new_[90699]_  & \new_[90696]_ ;
  assign \new_[90703]_  = ~A269 & ~A268;
  assign \new_[90706]_  = A302 & ~A300;
  assign \new_[90707]_  = \new_[90706]_  & \new_[90703]_ ;
  assign \new_[90708]_  = \new_[90707]_  & \new_[90700]_ ;
  assign \new_[90711]_  = A168 & ~A170;
  assign \new_[90714]_  = A166 & ~A167;
  assign \new_[90715]_  = \new_[90714]_  & \new_[90711]_ ;
  assign \new_[90718]_  = A200 & ~A199;
  assign \new_[90721]_  = ~A202 & ~A201;
  assign \new_[90722]_  = \new_[90721]_  & \new_[90718]_ ;
  assign \new_[90723]_  = \new_[90722]_  & \new_[90715]_ ;
  assign \new_[90726]_  = ~A265 & ~A203;
  assign \new_[90729]_  = ~A267 & A266;
  assign \new_[90730]_  = \new_[90729]_  & \new_[90726]_ ;
  assign \new_[90733]_  = ~A269 & ~A268;
  assign \new_[90736]_  = A299 & A298;
  assign \new_[90737]_  = \new_[90736]_  & \new_[90733]_ ;
  assign \new_[90738]_  = \new_[90737]_  & \new_[90730]_ ;
  assign \new_[90741]_  = A168 & ~A170;
  assign \new_[90744]_  = A166 & ~A167;
  assign \new_[90745]_  = \new_[90744]_  & \new_[90741]_ ;
  assign \new_[90748]_  = A200 & ~A199;
  assign \new_[90751]_  = ~A202 & ~A201;
  assign \new_[90752]_  = \new_[90751]_  & \new_[90748]_ ;
  assign \new_[90753]_  = \new_[90752]_  & \new_[90745]_ ;
  assign \new_[90756]_  = ~A265 & ~A203;
  assign \new_[90759]_  = ~A267 & A266;
  assign \new_[90760]_  = \new_[90759]_  & \new_[90756]_ ;
  assign \new_[90763]_  = ~A269 & ~A268;
  assign \new_[90766]_  = ~A299 & ~A298;
  assign \new_[90767]_  = \new_[90766]_  & \new_[90763]_ ;
  assign \new_[90768]_  = \new_[90767]_  & \new_[90760]_ ;
  assign \new_[90771]_  = A168 & ~A170;
  assign \new_[90774]_  = A166 & ~A167;
  assign \new_[90775]_  = \new_[90774]_  & \new_[90771]_ ;
  assign \new_[90778]_  = A200 & ~A199;
  assign \new_[90781]_  = ~A202 & ~A201;
  assign \new_[90782]_  = \new_[90781]_  & \new_[90778]_ ;
  assign \new_[90783]_  = \new_[90782]_  & \new_[90775]_ ;
  assign \new_[90786]_  = A265 & ~A203;
  assign \new_[90789]_  = A267 & ~A266;
  assign \new_[90790]_  = \new_[90789]_  & \new_[90786]_ ;
  assign \new_[90793]_  = A300 & A268;
  assign \new_[90796]_  = ~A302 & ~A301;
  assign \new_[90797]_  = \new_[90796]_  & \new_[90793]_ ;
  assign \new_[90798]_  = \new_[90797]_  & \new_[90790]_ ;
  assign \new_[90801]_  = A168 & ~A170;
  assign \new_[90804]_  = A166 & ~A167;
  assign \new_[90805]_  = \new_[90804]_  & \new_[90801]_ ;
  assign \new_[90808]_  = A200 & ~A199;
  assign \new_[90811]_  = ~A202 & ~A201;
  assign \new_[90812]_  = \new_[90811]_  & \new_[90808]_ ;
  assign \new_[90813]_  = \new_[90812]_  & \new_[90805]_ ;
  assign \new_[90816]_  = A265 & ~A203;
  assign \new_[90819]_  = A267 & ~A266;
  assign \new_[90820]_  = \new_[90819]_  & \new_[90816]_ ;
  assign \new_[90823]_  = A300 & A269;
  assign \new_[90826]_  = ~A302 & ~A301;
  assign \new_[90827]_  = \new_[90826]_  & \new_[90823]_ ;
  assign \new_[90828]_  = \new_[90827]_  & \new_[90820]_ ;
  assign \new_[90831]_  = A168 & ~A170;
  assign \new_[90834]_  = A166 & ~A167;
  assign \new_[90835]_  = \new_[90834]_  & \new_[90831]_ ;
  assign \new_[90838]_  = A200 & ~A199;
  assign \new_[90841]_  = ~A202 & ~A201;
  assign \new_[90842]_  = \new_[90841]_  & \new_[90838]_ ;
  assign \new_[90843]_  = \new_[90842]_  & \new_[90835]_ ;
  assign \new_[90846]_  = A265 & ~A203;
  assign \new_[90849]_  = ~A267 & ~A266;
  assign \new_[90850]_  = \new_[90849]_  & \new_[90846]_ ;
  assign \new_[90853]_  = ~A269 & ~A268;
  assign \new_[90856]_  = A301 & ~A300;
  assign \new_[90857]_  = \new_[90856]_  & \new_[90853]_ ;
  assign \new_[90858]_  = \new_[90857]_  & \new_[90850]_ ;
  assign \new_[90861]_  = A168 & ~A170;
  assign \new_[90864]_  = A166 & ~A167;
  assign \new_[90865]_  = \new_[90864]_  & \new_[90861]_ ;
  assign \new_[90868]_  = A200 & ~A199;
  assign \new_[90871]_  = ~A202 & ~A201;
  assign \new_[90872]_  = \new_[90871]_  & \new_[90868]_ ;
  assign \new_[90873]_  = \new_[90872]_  & \new_[90865]_ ;
  assign \new_[90876]_  = A265 & ~A203;
  assign \new_[90879]_  = ~A267 & ~A266;
  assign \new_[90880]_  = \new_[90879]_  & \new_[90876]_ ;
  assign \new_[90883]_  = ~A269 & ~A268;
  assign \new_[90886]_  = A302 & ~A300;
  assign \new_[90887]_  = \new_[90886]_  & \new_[90883]_ ;
  assign \new_[90888]_  = \new_[90887]_  & \new_[90880]_ ;
  assign \new_[90891]_  = A168 & ~A170;
  assign \new_[90894]_  = A166 & ~A167;
  assign \new_[90895]_  = \new_[90894]_  & \new_[90891]_ ;
  assign \new_[90898]_  = A200 & ~A199;
  assign \new_[90901]_  = ~A202 & ~A201;
  assign \new_[90902]_  = \new_[90901]_  & \new_[90898]_ ;
  assign \new_[90903]_  = \new_[90902]_  & \new_[90895]_ ;
  assign \new_[90906]_  = A265 & ~A203;
  assign \new_[90909]_  = ~A267 & ~A266;
  assign \new_[90910]_  = \new_[90909]_  & \new_[90906]_ ;
  assign \new_[90913]_  = ~A269 & ~A268;
  assign \new_[90916]_  = A299 & A298;
  assign \new_[90917]_  = \new_[90916]_  & \new_[90913]_ ;
  assign \new_[90918]_  = \new_[90917]_  & \new_[90910]_ ;
  assign \new_[90921]_  = A168 & ~A170;
  assign \new_[90924]_  = A166 & ~A167;
  assign \new_[90925]_  = \new_[90924]_  & \new_[90921]_ ;
  assign \new_[90928]_  = A200 & ~A199;
  assign \new_[90931]_  = ~A202 & ~A201;
  assign \new_[90932]_  = \new_[90931]_  & \new_[90928]_ ;
  assign \new_[90933]_  = \new_[90932]_  & \new_[90925]_ ;
  assign \new_[90936]_  = A265 & ~A203;
  assign \new_[90939]_  = ~A267 & ~A266;
  assign \new_[90940]_  = \new_[90939]_  & \new_[90936]_ ;
  assign \new_[90943]_  = ~A269 & ~A268;
  assign \new_[90946]_  = ~A299 & ~A298;
  assign \new_[90947]_  = \new_[90946]_  & \new_[90943]_ ;
  assign \new_[90948]_  = \new_[90947]_  & \new_[90940]_ ;
  assign \new_[90951]_  = A168 & ~A170;
  assign \new_[90954]_  = A166 & ~A167;
  assign \new_[90955]_  = \new_[90954]_  & \new_[90951]_ ;
  assign \new_[90958]_  = ~A200 & A199;
  assign \new_[90961]_  = A202 & A201;
  assign \new_[90962]_  = \new_[90961]_  & \new_[90958]_ ;
  assign \new_[90963]_  = \new_[90962]_  & \new_[90955]_ ;
  assign \new_[90966]_  = A266 & ~A265;
  assign \new_[90969]_  = ~A268 & ~A267;
  assign \new_[90970]_  = \new_[90969]_  & \new_[90966]_ ;
  assign \new_[90973]_  = A300 & ~A269;
  assign \new_[90976]_  = ~A302 & ~A301;
  assign \new_[90977]_  = \new_[90976]_  & \new_[90973]_ ;
  assign \new_[90978]_  = \new_[90977]_  & \new_[90970]_ ;
  assign \new_[90981]_  = A168 & ~A170;
  assign \new_[90984]_  = A166 & ~A167;
  assign \new_[90985]_  = \new_[90984]_  & \new_[90981]_ ;
  assign \new_[90988]_  = ~A200 & A199;
  assign \new_[90991]_  = A202 & A201;
  assign \new_[90992]_  = \new_[90991]_  & \new_[90988]_ ;
  assign \new_[90993]_  = \new_[90992]_  & \new_[90985]_ ;
  assign \new_[90996]_  = ~A266 & A265;
  assign \new_[90999]_  = ~A268 & ~A267;
  assign \new_[91000]_  = \new_[90999]_  & \new_[90996]_ ;
  assign \new_[91003]_  = A300 & ~A269;
  assign \new_[91006]_  = ~A302 & ~A301;
  assign \new_[91007]_  = \new_[91006]_  & \new_[91003]_ ;
  assign \new_[91008]_  = \new_[91007]_  & \new_[91000]_ ;
  assign \new_[91011]_  = A168 & ~A170;
  assign \new_[91014]_  = A166 & ~A167;
  assign \new_[91015]_  = \new_[91014]_  & \new_[91011]_ ;
  assign \new_[91018]_  = ~A200 & A199;
  assign \new_[91021]_  = A203 & A201;
  assign \new_[91022]_  = \new_[91021]_  & \new_[91018]_ ;
  assign \new_[91023]_  = \new_[91022]_  & \new_[91015]_ ;
  assign \new_[91026]_  = A266 & ~A265;
  assign \new_[91029]_  = ~A268 & ~A267;
  assign \new_[91030]_  = \new_[91029]_  & \new_[91026]_ ;
  assign \new_[91033]_  = A300 & ~A269;
  assign \new_[91036]_  = ~A302 & ~A301;
  assign \new_[91037]_  = \new_[91036]_  & \new_[91033]_ ;
  assign \new_[91038]_  = \new_[91037]_  & \new_[91030]_ ;
  assign \new_[91041]_  = A168 & ~A170;
  assign \new_[91044]_  = A166 & ~A167;
  assign \new_[91045]_  = \new_[91044]_  & \new_[91041]_ ;
  assign \new_[91048]_  = ~A200 & A199;
  assign \new_[91051]_  = A203 & A201;
  assign \new_[91052]_  = \new_[91051]_  & \new_[91048]_ ;
  assign \new_[91053]_  = \new_[91052]_  & \new_[91045]_ ;
  assign \new_[91056]_  = ~A266 & A265;
  assign \new_[91059]_  = ~A268 & ~A267;
  assign \new_[91060]_  = \new_[91059]_  & \new_[91056]_ ;
  assign \new_[91063]_  = A300 & ~A269;
  assign \new_[91066]_  = ~A302 & ~A301;
  assign \new_[91067]_  = \new_[91066]_  & \new_[91063]_ ;
  assign \new_[91068]_  = \new_[91067]_  & \new_[91060]_ ;
  assign \new_[91071]_  = A168 & ~A170;
  assign \new_[91074]_  = A166 & ~A167;
  assign \new_[91075]_  = \new_[91074]_  & \new_[91071]_ ;
  assign \new_[91078]_  = ~A200 & A199;
  assign \new_[91081]_  = ~A202 & ~A201;
  assign \new_[91082]_  = \new_[91081]_  & \new_[91078]_ ;
  assign \new_[91083]_  = \new_[91082]_  & \new_[91075]_ ;
  assign \new_[91086]_  = ~A265 & ~A203;
  assign \new_[91089]_  = A267 & A266;
  assign \new_[91090]_  = \new_[91089]_  & \new_[91086]_ ;
  assign \new_[91093]_  = A300 & A268;
  assign \new_[91096]_  = ~A302 & ~A301;
  assign \new_[91097]_  = \new_[91096]_  & \new_[91093]_ ;
  assign \new_[91098]_  = \new_[91097]_  & \new_[91090]_ ;
  assign \new_[91101]_  = A168 & ~A170;
  assign \new_[91104]_  = A166 & ~A167;
  assign \new_[91105]_  = \new_[91104]_  & \new_[91101]_ ;
  assign \new_[91108]_  = ~A200 & A199;
  assign \new_[91111]_  = ~A202 & ~A201;
  assign \new_[91112]_  = \new_[91111]_  & \new_[91108]_ ;
  assign \new_[91113]_  = \new_[91112]_  & \new_[91105]_ ;
  assign \new_[91116]_  = ~A265 & ~A203;
  assign \new_[91119]_  = A267 & A266;
  assign \new_[91120]_  = \new_[91119]_  & \new_[91116]_ ;
  assign \new_[91123]_  = A300 & A269;
  assign \new_[91126]_  = ~A302 & ~A301;
  assign \new_[91127]_  = \new_[91126]_  & \new_[91123]_ ;
  assign \new_[91128]_  = \new_[91127]_  & \new_[91120]_ ;
  assign \new_[91131]_  = A168 & ~A170;
  assign \new_[91134]_  = A166 & ~A167;
  assign \new_[91135]_  = \new_[91134]_  & \new_[91131]_ ;
  assign \new_[91138]_  = ~A200 & A199;
  assign \new_[91141]_  = ~A202 & ~A201;
  assign \new_[91142]_  = \new_[91141]_  & \new_[91138]_ ;
  assign \new_[91143]_  = \new_[91142]_  & \new_[91135]_ ;
  assign \new_[91146]_  = ~A265 & ~A203;
  assign \new_[91149]_  = ~A267 & A266;
  assign \new_[91150]_  = \new_[91149]_  & \new_[91146]_ ;
  assign \new_[91153]_  = ~A269 & ~A268;
  assign \new_[91156]_  = A301 & ~A300;
  assign \new_[91157]_  = \new_[91156]_  & \new_[91153]_ ;
  assign \new_[91158]_  = \new_[91157]_  & \new_[91150]_ ;
  assign \new_[91161]_  = A168 & ~A170;
  assign \new_[91164]_  = A166 & ~A167;
  assign \new_[91165]_  = \new_[91164]_  & \new_[91161]_ ;
  assign \new_[91168]_  = ~A200 & A199;
  assign \new_[91171]_  = ~A202 & ~A201;
  assign \new_[91172]_  = \new_[91171]_  & \new_[91168]_ ;
  assign \new_[91173]_  = \new_[91172]_  & \new_[91165]_ ;
  assign \new_[91176]_  = ~A265 & ~A203;
  assign \new_[91179]_  = ~A267 & A266;
  assign \new_[91180]_  = \new_[91179]_  & \new_[91176]_ ;
  assign \new_[91183]_  = ~A269 & ~A268;
  assign \new_[91186]_  = A302 & ~A300;
  assign \new_[91187]_  = \new_[91186]_  & \new_[91183]_ ;
  assign \new_[91188]_  = \new_[91187]_  & \new_[91180]_ ;
  assign \new_[91191]_  = A168 & ~A170;
  assign \new_[91194]_  = A166 & ~A167;
  assign \new_[91195]_  = \new_[91194]_  & \new_[91191]_ ;
  assign \new_[91198]_  = ~A200 & A199;
  assign \new_[91201]_  = ~A202 & ~A201;
  assign \new_[91202]_  = \new_[91201]_  & \new_[91198]_ ;
  assign \new_[91203]_  = \new_[91202]_  & \new_[91195]_ ;
  assign \new_[91206]_  = ~A265 & ~A203;
  assign \new_[91209]_  = ~A267 & A266;
  assign \new_[91210]_  = \new_[91209]_  & \new_[91206]_ ;
  assign \new_[91213]_  = ~A269 & ~A268;
  assign \new_[91216]_  = A299 & A298;
  assign \new_[91217]_  = \new_[91216]_  & \new_[91213]_ ;
  assign \new_[91218]_  = \new_[91217]_  & \new_[91210]_ ;
  assign \new_[91221]_  = A168 & ~A170;
  assign \new_[91224]_  = A166 & ~A167;
  assign \new_[91225]_  = \new_[91224]_  & \new_[91221]_ ;
  assign \new_[91228]_  = ~A200 & A199;
  assign \new_[91231]_  = ~A202 & ~A201;
  assign \new_[91232]_  = \new_[91231]_  & \new_[91228]_ ;
  assign \new_[91233]_  = \new_[91232]_  & \new_[91225]_ ;
  assign \new_[91236]_  = ~A265 & ~A203;
  assign \new_[91239]_  = ~A267 & A266;
  assign \new_[91240]_  = \new_[91239]_  & \new_[91236]_ ;
  assign \new_[91243]_  = ~A269 & ~A268;
  assign \new_[91246]_  = ~A299 & ~A298;
  assign \new_[91247]_  = \new_[91246]_  & \new_[91243]_ ;
  assign \new_[91248]_  = \new_[91247]_  & \new_[91240]_ ;
  assign \new_[91251]_  = A168 & ~A170;
  assign \new_[91254]_  = A166 & ~A167;
  assign \new_[91255]_  = \new_[91254]_  & \new_[91251]_ ;
  assign \new_[91258]_  = ~A200 & A199;
  assign \new_[91261]_  = ~A202 & ~A201;
  assign \new_[91262]_  = \new_[91261]_  & \new_[91258]_ ;
  assign \new_[91263]_  = \new_[91262]_  & \new_[91255]_ ;
  assign \new_[91266]_  = A265 & ~A203;
  assign \new_[91269]_  = A267 & ~A266;
  assign \new_[91270]_  = \new_[91269]_  & \new_[91266]_ ;
  assign \new_[91273]_  = A300 & A268;
  assign \new_[91276]_  = ~A302 & ~A301;
  assign \new_[91277]_  = \new_[91276]_  & \new_[91273]_ ;
  assign \new_[91278]_  = \new_[91277]_  & \new_[91270]_ ;
  assign \new_[91281]_  = A168 & ~A170;
  assign \new_[91284]_  = A166 & ~A167;
  assign \new_[91285]_  = \new_[91284]_  & \new_[91281]_ ;
  assign \new_[91288]_  = ~A200 & A199;
  assign \new_[91291]_  = ~A202 & ~A201;
  assign \new_[91292]_  = \new_[91291]_  & \new_[91288]_ ;
  assign \new_[91293]_  = \new_[91292]_  & \new_[91285]_ ;
  assign \new_[91296]_  = A265 & ~A203;
  assign \new_[91299]_  = A267 & ~A266;
  assign \new_[91300]_  = \new_[91299]_  & \new_[91296]_ ;
  assign \new_[91303]_  = A300 & A269;
  assign \new_[91306]_  = ~A302 & ~A301;
  assign \new_[91307]_  = \new_[91306]_  & \new_[91303]_ ;
  assign \new_[91308]_  = \new_[91307]_  & \new_[91300]_ ;
  assign \new_[91311]_  = A168 & ~A170;
  assign \new_[91314]_  = A166 & ~A167;
  assign \new_[91315]_  = \new_[91314]_  & \new_[91311]_ ;
  assign \new_[91318]_  = ~A200 & A199;
  assign \new_[91321]_  = ~A202 & ~A201;
  assign \new_[91322]_  = \new_[91321]_  & \new_[91318]_ ;
  assign \new_[91323]_  = \new_[91322]_  & \new_[91315]_ ;
  assign \new_[91326]_  = A265 & ~A203;
  assign \new_[91329]_  = ~A267 & ~A266;
  assign \new_[91330]_  = \new_[91329]_  & \new_[91326]_ ;
  assign \new_[91333]_  = ~A269 & ~A268;
  assign \new_[91336]_  = A301 & ~A300;
  assign \new_[91337]_  = \new_[91336]_  & \new_[91333]_ ;
  assign \new_[91338]_  = \new_[91337]_  & \new_[91330]_ ;
  assign \new_[91341]_  = A168 & ~A170;
  assign \new_[91344]_  = A166 & ~A167;
  assign \new_[91345]_  = \new_[91344]_  & \new_[91341]_ ;
  assign \new_[91348]_  = ~A200 & A199;
  assign \new_[91351]_  = ~A202 & ~A201;
  assign \new_[91352]_  = \new_[91351]_  & \new_[91348]_ ;
  assign \new_[91353]_  = \new_[91352]_  & \new_[91345]_ ;
  assign \new_[91356]_  = A265 & ~A203;
  assign \new_[91359]_  = ~A267 & ~A266;
  assign \new_[91360]_  = \new_[91359]_  & \new_[91356]_ ;
  assign \new_[91363]_  = ~A269 & ~A268;
  assign \new_[91366]_  = A302 & ~A300;
  assign \new_[91367]_  = \new_[91366]_  & \new_[91363]_ ;
  assign \new_[91368]_  = \new_[91367]_  & \new_[91360]_ ;
  assign \new_[91371]_  = A168 & ~A170;
  assign \new_[91374]_  = A166 & ~A167;
  assign \new_[91375]_  = \new_[91374]_  & \new_[91371]_ ;
  assign \new_[91378]_  = ~A200 & A199;
  assign \new_[91381]_  = ~A202 & ~A201;
  assign \new_[91382]_  = \new_[91381]_  & \new_[91378]_ ;
  assign \new_[91383]_  = \new_[91382]_  & \new_[91375]_ ;
  assign \new_[91386]_  = A265 & ~A203;
  assign \new_[91389]_  = ~A267 & ~A266;
  assign \new_[91390]_  = \new_[91389]_  & \new_[91386]_ ;
  assign \new_[91393]_  = ~A269 & ~A268;
  assign \new_[91396]_  = A299 & A298;
  assign \new_[91397]_  = \new_[91396]_  & \new_[91393]_ ;
  assign \new_[91398]_  = \new_[91397]_  & \new_[91390]_ ;
  assign \new_[91401]_  = A168 & ~A170;
  assign \new_[91404]_  = A166 & ~A167;
  assign \new_[91405]_  = \new_[91404]_  & \new_[91401]_ ;
  assign \new_[91408]_  = ~A200 & A199;
  assign \new_[91411]_  = ~A202 & ~A201;
  assign \new_[91412]_  = \new_[91411]_  & \new_[91408]_ ;
  assign \new_[91413]_  = \new_[91412]_  & \new_[91405]_ ;
  assign \new_[91416]_  = A265 & ~A203;
  assign \new_[91419]_  = ~A267 & ~A266;
  assign \new_[91420]_  = \new_[91419]_  & \new_[91416]_ ;
  assign \new_[91423]_  = ~A269 & ~A268;
  assign \new_[91426]_  = ~A299 & ~A298;
  assign \new_[91427]_  = \new_[91426]_  & \new_[91423]_ ;
  assign \new_[91428]_  = \new_[91427]_  & \new_[91420]_ ;
  assign \new_[91431]_  = A168 & A169;
  assign \new_[91434]_  = ~A166 & A167;
  assign \new_[91435]_  = \new_[91434]_  & \new_[91431]_ ;
  assign \new_[91438]_  = A200 & ~A199;
  assign \new_[91441]_  = A202 & A201;
  assign \new_[91442]_  = \new_[91441]_  & \new_[91438]_ ;
  assign \new_[91443]_  = \new_[91442]_  & \new_[91435]_ ;
  assign \new_[91446]_  = A266 & ~A265;
  assign \new_[91449]_  = ~A268 & ~A267;
  assign \new_[91450]_  = \new_[91449]_  & \new_[91446]_ ;
  assign \new_[91453]_  = A300 & ~A269;
  assign \new_[91456]_  = ~A302 & ~A301;
  assign \new_[91457]_  = \new_[91456]_  & \new_[91453]_ ;
  assign \new_[91458]_  = \new_[91457]_  & \new_[91450]_ ;
  assign \new_[91461]_  = A168 & A169;
  assign \new_[91464]_  = ~A166 & A167;
  assign \new_[91465]_  = \new_[91464]_  & \new_[91461]_ ;
  assign \new_[91468]_  = A200 & ~A199;
  assign \new_[91471]_  = A202 & A201;
  assign \new_[91472]_  = \new_[91471]_  & \new_[91468]_ ;
  assign \new_[91473]_  = \new_[91472]_  & \new_[91465]_ ;
  assign \new_[91476]_  = ~A266 & A265;
  assign \new_[91479]_  = ~A268 & ~A267;
  assign \new_[91480]_  = \new_[91479]_  & \new_[91476]_ ;
  assign \new_[91483]_  = A300 & ~A269;
  assign \new_[91486]_  = ~A302 & ~A301;
  assign \new_[91487]_  = \new_[91486]_  & \new_[91483]_ ;
  assign \new_[91488]_  = \new_[91487]_  & \new_[91480]_ ;
  assign \new_[91491]_  = A168 & A169;
  assign \new_[91494]_  = ~A166 & A167;
  assign \new_[91495]_  = \new_[91494]_  & \new_[91491]_ ;
  assign \new_[91498]_  = A200 & ~A199;
  assign \new_[91501]_  = A203 & A201;
  assign \new_[91502]_  = \new_[91501]_  & \new_[91498]_ ;
  assign \new_[91503]_  = \new_[91502]_  & \new_[91495]_ ;
  assign \new_[91506]_  = A266 & ~A265;
  assign \new_[91509]_  = ~A268 & ~A267;
  assign \new_[91510]_  = \new_[91509]_  & \new_[91506]_ ;
  assign \new_[91513]_  = A300 & ~A269;
  assign \new_[91516]_  = ~A302 & ~A301;
  assign \new_[91517]_  = \new_[91516]_  & \new_[91513]_ ;
  assign \new_[91518]_  = \new_[91517]_  & \new_[91510]_ ;
  assign \new_[91521]_  = A168 & A169;
  assign \new_[91524]_  = ~A166 & A167;
  assign \new_[91525]_  = \new_[91524]_  & \new_[91521]_ ;
  assign \new_[91528]_  = A200 & ~A199;
  assign \new_[91531]_  = A203 & A201;
  assign \new_[91532]_  = \new_[91531]_  & \new_[91528]_ ;
  assign \new_[91533]_  = \new_[91532]_  & \new_[91525]_ ;
  assign \new_[91536]_  = ~A266 & A265;
  assign \new_[91539]_  = ~A268 & ~A267;
  assign \new_[91540]_  = \new_[91539]_  & \new_[91536]_ ;
  assign \new_[91543]_  = A300 & ~A269;
  assign \new_[91546]_  = ~A302 & ~A301;
  assign \new_[91547]_  = \new_[91546]_  & \new_[91543]_ ;
  assign \new_[91548]_  = \new_[91547]_  & \new_[91540]_ ;
  assign \new_[91551]_  = A168 & A169;
  assign \new_[91554]_  = ~A166 & A167;
  assign \new_[91555]_  = \new_[91554]_  & \new_[91551]_ ;
  assign \new_[91558]_  = A200 & ~A199;
  assign \new_[91561]_  = ~A202 & ~A201;
  assign \new_[91562]_  = \new_[91561]_  & \new_[91558]_ ;
  assign \new_[91563]_  = \new_[91562]_  & \new_[91555]_ ;
  assign \new_[91566]_  = ~A265 & ~A203;
  assign \new_[91569]_  = A267 & A266;
  assign \new_[91570]_  = \new_[91569]_  & \new_[91566]_ ;
  assign \new_[91573]_  = A300 & A268;
  assign \new_[91576]_  = ~A302 & ~A301;
  assign \new_[91577]_  = \new_[91576]_  & \new_[91573]_ ;
  assign \new_[91578]_  = \new_[91577]_  & \new_[91570]_ ;
  assign \new_[91581]_  = A168 & A169;
  assign \new_[91584]_  = ~A166 & A167;
  assign \new_[91585]_  = \new_[91584]_  & \new_[91581]_ ;
  assign \new_[91588]_  = A200 & ~A199;
  assign \new_[91591]_  = ~A202 & ~A201;
  assign \new_[91592]_  = \new_[91591]_  & \new_[91588]_ ;
  assign \new_[91593]_  = \new_[91592]_  & \new_[91585]_ ;
  assign \new_[91596]_  = ~A265 & ~A203;
  assign \new_[91599]_  = A267 & A266;
  assign \new_[91600]_  = \new_[91599]_  & \new_[91596]_ ;
  assign \new_[91603]_  = A300 & A269;
  assign \new_[91606]_  = ~A302 & ~A301;
  assign \new_[91607]_  = \new_[91606]_  & \new_[91603]_ ;
  assign \new_[91608]_  = \new_[91607]_  & \new_[91600]_ ;
  assign \new_[91611]_  = A168 & A169;
  assign \new_[91614]_  = ~A166 & A167;
  assign \new_[91615]_  = \new_[91614]_  & \new_[91611]_ ;
  assign \new_[91618]_  = A200 & ~A199;
  assign \new_[91621]_  = ~A202 & ~A201;
  assign \new_[91622]_  = \new_[91621]_  & \new_[91618]_ ;
  assign \new_[91623]_  = \new_[91622]_  & \new_[91615]_ ;
  assign \new_[91626]_  = ~A265 & ~A203;
  assign \new_[91629]_  = ~A267 & A266;
  assign \new_[91630]_  = \new_[91629]_  & \new_[91626]_ ;
  assign \new_[91633]_  = ~A269 & ~A268;
  assign \new_[91636]_  = A301 & ~A300;
  assign \new_[91637]_  = \new_[91636]_  & \new_[91633]_ ;
  assign \new_[91638]_  = \new_[91637]_  & \new_[91630]_ ;
  assign \new_[91641]_  = A168 & A169;
  assign \new_[91644]_  = ~A166 & A167;
  assign \new_[91645]_  = \new_[91644]_  & \new_[91641]_ ;
  assign \new_[91648]_  = A200 & ~A199;
  assign \new_[91651]_  = ~A202 & ~A201;
  assign \new_[91652]_  = \new_[91651]_  & \new_[91648]_ ;
  assign \new_[91653]_  = \new_[91652]_  & \new_[91645]_ ;
  assign \new_[91656]_  = ~A265 & ~A203;
  assign \new_[91659]_  = ~A267 & A266;
  assign \new_[91660]_  = \new_[91659]_  & \new_[91656]_ ;
  assign \new_[91663]_  = ~A269 & ~A268;
  assign \new_[91666]_  = A302 & ~A300;
  assign \new_[91667]_  = \new_[91666]_  & \new_[91663]_ ;
  assign \new_[91668]_  = \new_[91667]_  & \new_[91660]_ ;
  assign \new_[91671]_  = A168 & A169;
  assign \new_[91674]_  = ~A166 & A167;
  assign \new_[91675]_  = \new_[91674]_  & \new_[91671]_ ;
  assign \new_[91678]_  = A200 & ~A199;
  assign \new_[91681]_  = ~A202 & ~A201;
  assign \new_[91682]_  = \new_[91681]_  & \new_[91678]_ ;
  assign \new_[91683]_  = \new_[91682]_  & \new_[91675]_ ;
  assign \new_[91686]_  = ~A265 & ~A203;
  assign \new_[91689]_  = ~A267 & A266;
  assign \new_[91690]_  = \new_[91689]_  & \new_[91686]_ ;
  assign \new_[91693]_  = ~A269 & ~A268;
  assign \new_[91696]_  = A299 & A298;
  assign \new_[91697]_  = \new_[91696]_  & \new_[91693]_ ;
  assign \new_[91698]_  = \new_[91697]_  & \new_[91690]_ ;
  assign \new_[91701]_  = A168 & A169;
  assign \new_[91704]_  = ~A166 & A167;
  assign \new_[91705]_  = \new_[91704]_  & \new_[91701]_ ;
  assign \new_[91708]_  = A200 & ~A199;
  assign \new_[91711]_  = ~A202 & ~A201;
  assign \new_[91712]_  = \new_[91711]_  & \new_[91708]_ ;
  assign \new_[91713]_  = \new_[91712]_  & \new_[91705]_ ;
  assign \new_[91716]_  = ~A265 & ~A203;
  assign \new_[91719]_  = ~A267 & A266;
  assign \new_[91720]_  = \new_[91719]_  & \new_[91716]_ ;
  assign \new_[91723]_  = ~A269 & ~A268;
  assign \new_[91726]_  = ~A299 & ~A298;
  assign \new_[91727]_  = \new_[91726]_  & \new_[91723]_ ;
  assign \new_[91728]_  = \new_[91727]_  & \new_[91720]_ ;
  assign \new_[91731]_  = A168 & A169;
  assign \new_[91734]_  = ~A166 & A167;
  assign \new_[91735]_  = \new_[91734]_  & \new_[91731]_ ;
  assign \new_[91738]_  = A200 & ~A199;
  assign \new_[91741]_  = ~A202 & ~A201;
  assign \new_[91742]_  = \new_[91741]_  & \new_[91738]_ ;
  assign \new_[91743]_  = \new_[91742]_  & \new_[91735]_ ;
  assign \new_[91746]_  = A265 & ~A203;
  assign \new_[91749]_  = A267 & ~A266;
  assign \new_[91750]_  = \new_[91749]_  & \new_[91746]_ ;
  assign \new_[91753]_  = A300 & A268;
  assign \new_[91756]_  = ~A302 & ~A301;
  assign \new_[91757]_  = \new_[91756]_  & \new_[91753]_ ;
  assign \new_[91758]_  = \new_[91757]_  & \new_[91750]_ ;
  assign \new_[91761]_  = A168 & A169;
  assign \new_[91764]_  = ~A166 & A167;
  assign \new_[91765]_  = \new_[91764]_  & \new_[91761]_ ;
  assign \new_[91768]_  = A200 & ~A199;
  assign \new_[91771]_  = ~A202 & ~A201;
  assign \new_[91772]_  = \new_[91771]_  & \new_[91768]_ ;
  assign \new_[91773]_  = \new_[91772]_  & \new_[91765]_ ;
  assign \new_[91776]_  = A265 & ~A203;
  assign \new_[91779]_  = A267 & ~A266;
  assign \new_[91780]_  = \new_[91779]_  & \new_[91776]_ ;
  assign \new_[91783]_  = A300 & A269;
  assign \new_[91786]_  = ~A302 & ~A301;
  assign \new_[91787]_  = \new_[91786]_  & \new_[91783]_ ;
  assign \new_[91788]_  = \new_[91787]_  & \new_[91780]_ ;
  assign \new_[91791]_  = A168 & A169;
  assign \new_[91794]_  = ~A166 & A167;
  assign \new_[91795]_  = \new_[91794]_  & \new_[91791]_ ;
  assign \new_[91798]_  = A200 & ~A199;
  assign \new_[91801]_  = ~A202 & ~A201;
  assign \new_[91802]_  = \new_[91801]_  & \new_[91798]_ ;
  assign \new_[91803]_  = \new_[91802]_  & \new_[91795]_ ;
  assign \new_[91806]_  = A265 & ~A203;
  assign \new_[91809]_  = ~A267 & ~A266;
  assign \new_[91810]_  = \new_[91809]_  & \new_[91806]_ ;
  assign \new_[91813]_  = ~A269 & ~A268;
  assign \new_[91816]_  = A301 & ~A300;
  assign \new_[91817]_  = \new_[91816]_  & \new_[91813]_ ;
  assign \new_[91818]_  = \new_[91817]_  & \new_[91810]_ ;
  assign \new_[91821]_  = A168 & A169;
  assign \new_[91824]_  = ~A166 & A167;
  assign \new_[91825]_  = \new_[91824]_  & \new_[91821]_ ;
  assign \new_[91828]_  = A200 & ~A199;
  assign \new_[91831]_  = ~A202 & ~A201;
  assign \new_[91832]_  = \new_[91831]_  & \new_[91828]_ ;
  assign \new_[91833]_  = \new_[91832]_  & \new_[91825]_ ;
  assign \new_[91836]_  = A265 & ~A203;
  assign \new_[91839]_  = ~A267 & ~A266;
  assign \new_[91840]_  = \new_[91839]_  & \new_[91836]_ ;
  assign \new_[91843]_  = ~A269 & ~A268;
  assign \new_[91846]_  = A302 & ~A300;
  assign \new_[91847]_  = \new_[91846]_  & \new_[91843]_ ;
  assign \new_[91848]_  = \new_[91847]_  & \new_[91840]_ ;
  assign \new_[91851]_  = A168 & A169;
  assign \new_[91854]_  = ~A166 & A167;
  assign \new_[91855]_  = \new_[91854]_  & \new_[91851]_ ;
  assign \new_[91858]_  = A200 & ~A199;
  assign \new_[91861]_  = ~A202 & ~A201;
  assign \new_[91862]_  = \new_[91861]_  & \new_[91858]_ ;
  assign \new_[91863]_  = \new_[91862]_  & \new_[91855]_ ;
  assign \new_[91866]_  = A265 & ~A203;
  assign \new_[91869]_  = ~A267 & ~A266;
  assign \new_[91870]_  = \new_[91869]_  & \new_[91866]_ ;
  assign \new_[91873]_  = ~A269 & ~A268;
  assign \new_[91876]_  = A299 & A298;
  assign \new_[91877]_  = \new_[91876]_  & \new_[91873]_ ;
  assign \new_[91878]_  = \new_[91877]_  & \new_[91870]_ ;
  assign \new_[91881]_  = A168 & A169;
  assign \new_[91884]_  = ~A166 & A167;
  assign \new_[91885]_  = \new_[91884]_  & \new_[91881]_ ;
  assign \new_[91888]_  = A200 & ~A199;
  assign \new_[91891]_  = ~A202 & ~A201;
  assign \new_[91892]_  = \new_[91891]_  & \new_[91888]_ ;
  assign \new_[91893]_  = \new_[91892]_  & \new_[91885]_ ;
  assign \new_[91896]_  = A265 & ~A203;
  assign \new_[91899]_  = ~A267 & ~A266;
  assign \new_[91900]_  = \new_[91899]_  & \new_[91896]_ ;
  assign \new_[91903]_  = ~A269 & ~A268;
  assign \new_[91906]_  = ~A299 & ~A298;
  assign \new_[91907]_  = \new_[91906]_  & \new_[91903]_ ;
  assign \new_[91908]_  = \new_[91907]_  & \new_[91900]_ ;
  assign \new_[91911]_  = A168 & A169;
  assign \new_[91914]_  = ~A166 & A167;
  assign \new_[91915]_  = \new_[91914]_  & \new_[91911]_ ;
  assign \new_[91918]_  = ~A200 & A199;
  assign \new_[91921]_  = A202 & A201;
  assign \new_[91922]_  = \new_[91921]_  & \new_[91918]_ ;
  assign \new_[91923]_  = \new_[91922]_  & \new_[91915]_ ;
  assign \new_[91926]_  = A266 & ~A265;
  assign \new_[91929]_  = ~A268 & ~A267;
  assign \new_[91930]_  = \new_[91929]_  & \new_[91926]_ ;
  assign \new_[91933]_  = A300 & ~A269;
  assign \new_[91936]_  = ~A302 & ~A301;
  assign \new_[91937]_  = \new_[91936]_  & \new_[91933]_ ;
  assign \new_[91938]_  = \new_[91937]_  & \new_[91930]_ ;
  assign \new_[91941]_  = A168 & A169;
  assign \new_[91944]_  = ~A166 & A167;
  assign \new_[91945]_  = \new_[91944]_  & \new_[91941]_ ;
  assign \new_[91948]_  = ~A200 & A199;
  assign \new_[91951]_  = A202 & A201;
  assign \new_[91952]_  = \new_[91951]_  & \new_[91948]_ ;
  assign \new_[91953]_  = \new_[91952]_  & \new_[91945]_ ;
  assign \new_[91956]_  = ~A266 & A265;
  assign \new_[91959]_  = ~A268 & ~A267;
  assign \new_[91960]_  = \new_[91959]_  & \new_[91956]_ ;
  assign \new_[91963]_  = A300 & ~A269;
  assign \new_[91966]_  = ~A302 & ~A301;
  assign \new_[91967]_  = \new_[91966]_  & \new_[91963]_ ;
  assign \new_[91968]_  = \new_[91967]_  & \new_[91960]_ ;
  assign \new_[91971]_  = A168 & A169;
  assign \new_[91974]_  = ~A166 & A167;
  assign \new_[91975]_  = \new_[91974]_  & \new_[91971]_ ;
  assign \new_[91978]_  = ~A200 & A199;
  assign \new_[91981]_  = A203 & A201;
  assign \new_[91982]_  = \new_[91981]_  & \new_[91978]_ ;
  assign \new_[91983]_  = \new_[91982]_  & \new_[91975]_ ;
  assign \new_[91986]_  = A266 & ~A265;
  assign \new_[91989]_  = ~A268 & ~A267;
  assign \new_[91990]_  = \new_[91989]_  & \new_[91986]_ ;
  assign \new_[91993]_  = A300 & ~A269;
  assign \new_[91996]_  = ~A302 & ~A301;
  assign \new_[91997]_  = \new_[91996]_  & \new_[91993]_ ;
  assign \new_[91998]_  = \new_[91997]_  & \new_[91990]_ ;
  assign \new_[92001]_  = A168 & A169;
  assign \new_[92004]_  = ~A166 & A167;
  assign \new_[92005]_  = \new_[92004]_  & \new_[92001]_ ;
  assign \new_[92008]_  = ~A200 & A199;
  assign \new_[92011]_  = A203 & A201;
  assign \new_[92012]_  = \new_[92011]_  & \new_[92008]_ ;
  assign \new_[92013]_  = \new_[92012]_  & \new_[92005]_ ;
  assign \new_[92016]_  = ~A266 & A265;
  assign \new_[92019]_  = ~A268 & ~A267;
  assign \new_[92020]_  = \new_[92019]_  & \new_[92016]_ ;
  assign \new_[92023]_  = A300 & ~A269;
  assign \new_[92026]_  = ~A302 & ~A301;
  assign \new_[92027]_  = \new_[92026]_  & \new_[92023]_ ;
  assign \new_[92028]_  = \new_[92027]_  & \new_[92020]_ ;
  assign \new_[92031]_  = A168 & A169;
  assign \new_[92034]_  = ~A166 & A167;
  assign \new_[92035]_  = \new_[92034]_  & \new_[92031]_ ;
  assign \new_[92038]_  = ~A200 & A199;
  assign \new_[92041]_  = ~A202 & ~A201;
  assign \new_[92042]_  = \new_[92041]_  & \new_[92038]_ ;
  assign \new_[92043]_  = \new_[92042]_  & \new_[92035]_ ;
  assign \new_[92046]_  = ~A265 & ~A203;
  assign \new_[92049]_  = A267 & A266;
  assign \new_[92050]_  = \new_[92049]_  & \new_[92046]_ ;
  assign \new_[92053]_  = A300 & A268;
  assign \new_[92056]_  = ~A302 & ~A301;
  assign \new_[92057]_  = \new_[92056]_  & \new_[92053]_ ;
  assign \new_[92058]_  = \new_[92057]_  & \new_[92050]_ ;
  assign \new_[92061]_  = A168 & A169;
  assign \new_[92064]_  = ~A166 & A167;
  assign \new_[92065]_  = \new_[92064]_  & \new_[92061]_ ;
  assign \new_[92068]_  = ~A200 & A199;
  assign \new_[92071]_  = ~A202 & ~A201;
  assign \new_[92072]_  = \new_[92071]_  & \new_[92068]_ ;
  assign \new_[92073]_  = \new_[92072]_  & \new_[92065]_ ;
  assign \new_[92076]_  = ~A265 & ~A203;
  assign \new_[92079]_  = A267 & A266;
  assign \new_[92080]_  = \new_[92079]_  & \new_[92076]_ ;
  assign \new_[92083]_  = A300 & A269;
  assign \new_[92086]_  = ~A302 & ~A301;
  assign \new_[92087]_  = \new_[92086]_  & \new_[92083]_ ;
  assign \new_[92088]_  = \new_[92087]_  & \new_[92080]_ ;
  assign \new_[92091]_  = A168 & A169;
  assign \new_[92094]_  = ~A166 & A167;
  assign \new_[92095]_  = \new_[92094]_  & \new_[92091]_ ;
  assign \new_[92098]_  = ~A200 & A199;
  assign \new_[92101]_  = ~A202 & ~A201;
  assign \new_[92102]_  = \new_[92101]_  & \new_[92098]_ ;
  assign \new_[92103]_  = \new_[92102]_  & \new_[92095]_ ;
  assign \new_[92106]_  = ~A265 & ~A203;
  assign \new_[92109]_  = ~A267 & A266;
  assign \new_[92110]_  = \new_[92109]_  & \new_[92106]_ ;
  assign \new_[92113]_  = ~A269 & ~A268;
  assign \new_[92116]_  = A301 & ~A300;
  assign \new_[92117]_  = \new_[92116]_  & \new_[92113]_ ;
  assign \new_[92118]_  = \new_[92117]_  & \new_[92110]_ ;
  assign \new_[92121]_  = A168 & A169;
  assign \new_[92124]_  = ~A166 & A167;
  assign \new_[92125]_  = \new_[92124]_  & \new_[92121]_ ;
  assign \new_[92128]_  = ~A200 & A199;
  assign \new_[92131]_  = ~A202 & ~A201;
  assign \new_[92132]_  = \new_[92131]_  & \new_[92128]_ ;
  assign \new_[92133]_  = \new_[92132]_  & \new_[92125]_ ;
  assign \new_[92136]_  = ~A265 & ~A203;
  assign \new_[92139]_  = ~A267 & A266;
  assign \new_[92140]_  = \new_[92139]_  & \new_[92136]_ ;
  assign \new_[92143]_  = ~A269 & ~A268;
  assign \new_[92146]_  = A302 & ~A300;
  assign \new_[92147]_  = \new_[92146]_  & \new_[92143]_ ;
  assign \new_[92148]_  = \new_[92147]_  & \new_[92140]_ ;
  assign \new_[92151]_  = A168 & A169;
  assign \new_[92154]_  = ~A166 & A167;
  assign \new_[92155]_  = \new_[92154]_  & \new_[92151]_ ;
  assign \new_[92158]_  = ~A200 & A199;
  assign \new_[92161]_  = ~A202 & ~A201;
  assign \new_[92162]_  = \new_[92161]_  & \new_[92158]_ ;
  assign \new_[92163]_  = \new_[92162]_  & \new_[92155]_ ;
  assign \new_[92166]_  = ~A265 & ~A203;
  assign \new_[92169]_  = ~A267 & A266;
  assign \new_[92170]_  = \new_[92169]_  & \new_[92166]_ ;
  assign \new_[92173]_  = ~A269 & ~A268;
  assign \new_[92176]_  = A299 & A298;
  assign \new_[92177]_  = \new_[92176]_  & \new_[92173]_ ;
  assign \new_[92178]_  = \new_[92177]_  & \new_[92170]_ ;
  assign \new_[92181]_  = A168 & A169;
  assign \new_[92184]_  = ~A166 & A167;
  assign \new_[92185]_  = \new_[92184]_  & \new_[92181]_ ;
  assign \new_[92188]_  = ~A200 & A199;
  assign \new_[92191]_  = ~A202 & ~A201;
  assign \new_[92192]_  = \new_[92191]_  & \new_[92188]_ ;
  assign \new_[92193]_  = \new_[92192]_  & \new_[92185]_ ;
  assign \new_[92196]_  = ~A265 & ~A203;
  assign \new_[92199]_  = ~A267 & A266;
  assign \new_[92200]_  = \new_[92199]_  & \new_[92196]_ ;
  assign \new_[92203]_  = ~A269 & ~A268;
  assign \new_[92206]_  = ~A299 & ~A298;
  assign \new_[92207]_  = \new_[92206]_  & \new_[92203]_ ;
  assign \new_[92208]_  = \new_[92207]_  & \new_[92200]_ ;
  assign \new_[92211]_  = A168 & A169;
  assign \new_[92214]_  = ~A166 & A167;
  assign \new_[92215]_  = \new_[92214]_  & \new_[92211]_ ;
  assign \new_[92218]_  = ~A200 & A199;
  assign \new_[92221]_  = ~A202 & ~A201;
  assign \new_[92222]_  = \new_[92221]_  & \new_[92218]_ ;
  assign \new_[92223]_  = \new_[92222]_  & \new_[92215]_ ;
  assign \new_[92226]_  = A265 & ~A203;
  assign \new_[92229]_  = A267 & ~A266;
  assign \new_[92230]_  = \new_[92229]_  & \new_[92226]_ ;
  assign \new_[92233]_  = A300 & A268;
  assign \new_[92236]_  = ~A302 & ~A301;
  assign \new_[92237]_  = \new_[92236]_  & \new_[92233]_ ;
  assign \new_[92238]_  = \new_[92237]_  & \new_[92230]_ ;
  assign \new_[92241]_  = A168 & A169;
  assign \new_[92244]_  = ~A166 & A167;
  assign \new_[92245]_  = \new_[92244]_  & \new_[92241]_ ;
  assign \new_[92248]_  = ~A200 & A199;
  assign \new_[92251]_  = ~A202 & ~A201;
  assign \new_[92252]_  = \new_[92251]_  & \new_[92248]_ ;
  assign \new_[92253]_  = \new_[92252]_  & \new_[92245]_ ;
  assign \new_[92256]_  = A265 & ~A203;
  assign \new_[92259]_  = A267 & ~A266;
  assign \new_[92260]_  = \new_[92259]_  & \new_[92256]_ ;
  assign \new_[92263]_  = A300 & A269;
  assign \new_[92266]_  = ~A302 & ~A301;
  assign \new_[92267]_  = \new_[92266]_  & \new_[92263]_ ;
  assign \new_[92268]_  = \new_[92267]_  & \new_[92260]_ ;
  assign \new_[92271]_  = A168 & A169;
  assign \new_[92274]_  = ~A166 & A167;
  assign \new_[92275]_  = \new_[92274]_  & \new_[92271]_ ;
  assign \new_[92278]_  = ~A200 & A199;
  assign \new_[92281]_  = ~A202 & ~A201;
  assign \new_[92282]_  = \new_[92281]_  & \new_[92278]_ ;
  assign \new_[92283]_  = \new_[92282]_  & \new_[92275]_ ;
  assign \new_[92286]_  = A265 & ~A203;
  assign \new_[92289]_  = ~A267 & ~A266;
  assign \new_[92290]_  = \new_[92289]_  & \new_[92286]_ ;
  assign \new_[92293]_  = ~A269 & ~A268;
  assign \new_[92296]_  = A301 & ~A300;
  assign \new_[92297]_  = \new_[92296]_  & \new_[92293]_ ;
  assign \new_[92298]_  = \new_[92297]_  & \new_[92290]_ ;
  assign \new_[92301]_  = A168 & A169;
  assign \new_[92304]_  = ~A166 & A167;
  assign \new_[92305]_  = \new_[92304]_  & \new_[92301]_ ;
  assign \new_[92308]_  = ~A200 & A199;
  assign \new_[92311]_  = ~A202 & ~A201;
  assign \new_[92312]_  = \new_[92311]_  & \new_[92308]_ ;
  assign \new_[92313]_  = \new_[92312]_  & \new_[92305]_ ;
  assign \new_[92316]_  = A265 & ~A203;
  assign \new_[92319]_  = ~A267 & ~A266;
  assign \new_[92320]_  = \new_[92319]_  & \new_[92316]_ ;
  assign \new_[92323]_  = ~A269 & ~A268;
  assign \new_[92326]_  = A302 & ~A300;
  assign \new_[92327]_  = \new_[92326]_  & \new_[92323]_ ;
  assign \new_[92328]_  = \new_[92327]_  & \new_[92320]_ ;
  assign \new_[92331]_  = A168 & A169;
  assign \new_[92334]_  = ~A166 & A167;
  assign \new_[92335]_  = \new_[92334]_  & \new_[92331]_ ;
  assign \new_[92338]_  = ~A200 & A199;
  assign \new_[92341]_  = ~A202 & ~A201;
  assign \new_[92342]_  = \new_[92341]_  & \new_[92338]_ ;
  assign \new_[92343]_  = \new_[92342]_  & \new_[92335]_ ;
  assign \new_[92346]_  = A265 & ~A203;
  assign \new_[92349]_  = ~A267 & ~A266;
  assign \new_[92350]_  = \new_[92349]_  & \new_[92346]_ ;
  assign \new_[92353]_  = ~A269 & ~A268;
  assign \new_[92356]_  = A299 & A298;
  assign \new_[92357]_  = \new_[92356]_  & \new_[92353]_ ;
  assign \new_[92358]_  = \new_[92357]_  & \new_[92350]_ ;
  assign \new_[92361]_  = A168 & A169;
  assign \new_[92364]_  = ~A166 & A167;
  assign \new_[92365]_  = \new_[92364]_  & \new_[92361]_ ;
  assign \new_[92368]_  = ~A200 & A199;
  assign \new_[92371]_  = ~A202 & ~A201;
  assign \new_[92372]_  = \new_[92371]_  & \new_[92368]_ ;
  assign \new_[92373]_  = \new_[92372]_  & \new_[92365]_ ;
  assign \new_[92376]_  = A265 & ~A203;
  assign \new_[92379]_  = ~A267 & ~A266;
  assign \new_[92380]_  = \new_[92379]_  & \new_[92376]_ ;
  assign \new_[92383]_  = ~A269 & ~A268;
  assign \new_[92386]_  = ~A299 & ~A298;
  assign \new_[92387]_  = \new_[92386]_  & \new_[92383]_ ;
  assign \new_[92388]_  = \new_[92387]_  & \new_[92380]_ ;
  assign \new_[92391]_  = A168 & A169;
  assign \new_[92394]_  = A166 & ~A167;
  assign \new_[92395]_  = \new_[92394]_  & \new_[92391]_ ;
  assign \new_[92398]_  = A200 & ~A199;
  assign \new_[92401]_  = A202 & A201;
  assign \new_[92402]_  = \new_[92401]_  & \new_[92398]_ ;
  assign \new_[92403]_  = \new_[92402]_  & \new_[92395]_ ;
  assign \new_[92406]_  = A266 & ~A265;
  assign \new_[92409]_  = ~A268 & ~A267;
  assign \new_[92410]_  = \new_[92409]_  & \new_[92406]_ ;
  assign \new_[92413]_  = A300 & ~A269;
  assign \new_[92416]_  = ~A302 & ~A301;
  assign \new_[92417]_  = \new_[92416]_  & \new_[92413]_ ;
  assign \new_[92418]_  = \new_[92417]_  & \new_[92410]_ ;
  assign \new_[92421]_  = A168 & A169;
  assign \new_[92424]_  = A166 & ~A167;
  assign \new_[92425]_  = \new_[92424]_  & \new_[92421]_ ;
  assign \new_[92428]_  = A200 & ~A199;
  assign \new_[92431]_  = A202 & A201;
  assign \new_[92432]_  = \new_[92431]_  & \new_[92428]_ ;
  assign \new_[92433]_  = \new_[92432]_  & \new_[92425]_ ;
  assign \new_[92436]_  = ~A266 & A265;
  assign \new_[92439]_  = ~A268 & ~A267;
  assign \new_[92440]_  = \new_[92439]_  & \new_[92436]_ ;
  assign \new_[92443]_  = A300 & ~A269;
  assign \new_[92446]_  = ~A302 & ~A301;
  assign \new_[92447]_  = \new_[92446]_  & \new_[92443]_ ;
  assign \new_[92448]_  = \new_[92447]_  & \new_[92440]_ ;
  assign \new_[92451]_  = A168 & A169;
  assign \new_[92454]_  = A166 & ~A167;
  assign \new_[92455]_  = \new_[92454]_  & \new_[92451]_ ;
  assign \new_[92458]_  = A200 & ~A199;
  assign \new_[92461]_  = A203 & A201;
  assign \new_[92462]_  = \new_[92461]_  & \new_[92458]_ ;
  assign \new_[92463]_  = \new_[92462]_  & \new_[92455]_ ;
  assign \new_[92466]_  = A266 & ~A265;
  assign \new_[92469]_  = ~A268 & ~A267;
  assign \new_[92470]_  = \new_[92469]_  & \new_[92466]_ ;
  assign \new_[92473]_  = A300 & ~A269;
  assign \new_[92476]_  = ~A302 & ~A301;
  assign \new_[92477]_  = \new_[92476]_  & \new_[92473]_ ;
  assign \new_[92478]_  = \new_[92477]_  & \new_[92470]_ ;
  assign \new_[92481]_  = A168 & A169;
  assign \new_[92484]_  = A166 & ~A167;
  assign \new_[92485]_  = \new_[92484]_  & \new_[92481]_ ;
  assign \new_[92488]_  = A200 & ~A199;
  assign \new_[92491]_  = A203 & A201;
  assign \new_[92492]_  = \new_[92491]_  & \new_[92488]_ ;
  assign \new_[92493]_  = \new_[92492]_  & \new_[92485]_ ;
  assign \new_[92496]_  = ~A266 & A265;
  assign \new_[92499]_  = ~A268 & ~A267;
  assign \new_[92500]_  = \new_[92499]_  & \new_[92496]_ ;
  assign \new_[92503]_  = A300 & ~A269;
  assign \new_[92506]_  = ~A302 & ~A301;
  assign \new_[92507]_  = \new_[92506]_  & \new_[92503]_ ;
  assign \new_[92508]_  = \new_[92507]_  & \new_[92500]_ ;
  assign \new_[92511]_  = A168 & A169;
  assign \new_[92514]_  = A166 & ~A167;
  assign \new_[92515]_  = \new_[92514]_  & \new_[92511]_ ;
  assign \new_[92518]_  = A200 & ~A199;
  assign \new_[92521]_  = ~A202 & ~A201;
  assign \new_[92522]_  = \new_[92521]_  & \new_[92518]_ ;
  assign \new_[92523]_  = \new_[92522]_  & \new_[92515]_ ;
  assign \new_[92526]_  = ~A265 & ~A203;
  assign \new_[92529]_  = A267 & A266;
  assign \new_[92530]_  = \new_[92529]_  & \new_[92526]_ ;
  assign \new_[92533]_  = A300 & A268;
  assign \new_[92536]_  = ~A302 & ~A301;
  assign \new_[92537]_  = \new_[92536]_  & \new_[92533]_ ;
  assign \new_[92538]_  = \new_[92537]_  & \new_[92530]_ ;
  assign \new_[92541]_  = A168 & A169;
  assign \new_[92544]_  = A166 & ~A167;
  assign \new_[92545]_  = \new_[92544]_  & \new_[92541]_ ;
  assign \new_[92548]_  = A200 & ~A199;
  assign \new_[92551]_  = ~A202 & ~A201;
  assign \new_[92552]_  = \new_[92551]_  & \new_[92548]_ ;
  assign \new_[92553]_  = \new_[92552]_  & \new_[92545]_ ;
  assign \new_[92556]_  = ~A265 & ~A203;
  assign \new_[92559]_  = A267 & A266;
  assign \new_[92560]_  = \new_[92559]_  & \new_[92556]_ ;
  assign \new_[92563]_  = A300 & A269;
  assign \new_[92566]_  = ~A302 & ~A301;
  assign \new_[92567]_  = \new_[92566]_  & \new_[92563]_ ;
  assign \new_[92568]_  = \new_[92567]_  & \new_[92560]_ ;
  assign \new_[92571]_  = A168 & A169;
  assign \new_[92574]_  = A166 & ~A167;
  assign \new_[92575]_  = \new_[92574]_  & \new_[92571]_ ;
  assign \new_[92578]_  = A200 & ~A199;
  assign \new_[92581]_  = ~A202 & ~A201;
  assign \new_[92582]_  = \new_[92581]_  & \new_[92578]_ ;
  assign \new_[92583]_  = \new_[92582]_  & \new_[92575]_ ;
  assign \new_[92586]_  = ~A265 & ~A203;
  assign \new_[92589]_  = ~A267 & A266;
  assign \new_[92590]_  = \new_[92589]_  & \new_[92586]_ ;
  assign \new_[92593]_  = ~A269 & ~A268;
  assign \new_[92596]_  = A301 & ~A300;
  assign \new_[92597]_  = \new_[92596]_  & \new_[92593]_ ;
  assign \new_[92598]_  = \new_[92597]_  & \new_[92590]_ ;
  assign \new_[92601]_  = A168 & A169;
  assign \new_[92604]_  = A166 & ~A167;
  assign \new_[92605]_  = \new_[92604]_  & \new_[92601]_ ;
  assign \new_[92608]_  = A200 & ~A199;
  assign \new_[92611]_  = ~A202 & ~A201;
  assign \new_[92612]_  = \new_[92611]_  & \new_[92608]_ ;
  assign \new_[92613]_  = \new_[92612]_  & \new_[92605]_ ;
  assign \new_[92616]_  = ~A265 & ~A203;
  assign \new_[92619]_  = ~A267 & A266;
  assign \new_[92620]_  = \new_[92619]_  & \new_[92616]_ ;
  assign \new_[92623]_  = ~A269 & ~A268;
  assign \new_[92626]_  = A302 & ~A300;
  assign \new_[92627]_  = \new_[92626]_  & \new_[92623]_ ;
  assign \new_[92628]_  = \new_[92627]_  & \new_[92620]_ ;
  assign \new_[92631]_  = A168 & A169;
  assign \new_[92634]_  = A166 & ~A167;
  assign \new_[92635]_  = \new_[92634]_  & \new_[92631]_ ;
  assign \new_[92638]_  = A200 & ~A199;
  assign \new_[92641]_  = ~A202 & ~A201;
  assign \new_[92642]_  = \new_[92641]_  & \new_[92638]_ ;
  assign \new_[92643]_  = \new_[92642]_  & \new_[92635]_ ;
  assign \new_[92646]_  = ~A265 & ~A203;
  assign \new_[92649]_  = ~A267 & A266;
  assign \new_[92650]_  = \new_[92649]_  & \new_[92646]_ ;
  assign \new_[92653]_  = ~A269 & ~A268;
  assign \new_[92656]_  = A299 & A298;
  assign \new_[92657]_  = \new_[92656]_  & \new_[92653]_ ;
  assign \new_[92658]_  = \new_[92657]_  & \new_[92650]_ ;
  assign \new_[92661]_  = A168 & A169;
  assign \new_[92664]_  = A166 & ~A167;
  assign \new_[92665]_  = \new_[92664]_  & \new_[92661]_ ;
  assign \new_[92668]_  = A200 & ~A199;
  assign \new_[92671]_  = ~A202 & ~A201;
  assign \new_[92672]_  = \new_[92671]_  & \new_[92668]_ ;
  assign \new_[92673]_  = \new_[92672]_  & \new_[92665]_ ;
  assign \new_[92676]_  = ~A265 & ~A203;
  assign \new_[92679]_  = ~A267 & A266;
  assign \new_[92680]_  = \new_[92679]_  & \new_[92676]_ ;
  assign \new_[92683]_  = ~A269 & ~A268;
  assign \new_[92686]_  = ~A299 & ~A298;
  assign \new_[92687]_  = \new_[92686]_  & \new_[92683]_ ;
  assign \new_[92688]_  = \new_[92687]_  & \new_[92680]_ ;
  assign \new_[92691]_  = A168 & A169;
  assign \new_[92694]_  = A166 & ~A167;
  assign \new_[92695]_  = \new_[92694]_  & \new_[92691]_ ;
  assign \new_[92698]_  = A200 & ~A199;
  assign \new_[92701]_  = ~A202 & ~A201;
  assign \new_[92702]_  = \new_[92701]_  & \new_[92698]_ ;
  assign \new_[92703]_  = \new_[92702]_  & \new_[92695]_ ;
  assign \new_[92706]_  = A265 & ~A203;
  assign \new_[92709]_  = A267 & ~A266;
  assign \new_[92710]_  = \new_[92709]_  & \new_[92706]_ ;
  assign \new_[92713]_  = A300 & A268;
  assign \new_[92716]_  = ~A302 & ~A301;
  assign \new_[92717]_  = \new_[92716]_  & \new_[92713]_ ;
  assign \new_[92718]_  = \new_[92717]_  & \new_[92710]_ ;
  assign \new_[92721]_  = A168 & A169;
  assign \new_[92724]_  = A166 & ~A167;
  assign \new_[92725]_  = \new_[92724]_  & \new_[92721]_ ;
  assign \new_[92728]_  = A200 & ~A199;
  assign \new_[92731]_  = ~A202 & ~A201;
  assign \new_[92732]_  = \new_[92731]_  & \new_[92728]_ ;
  assign \new_[92733]_  = \new_[92732]_  & \new_[92725]_ ;
  assign \new_[92736]_  = A265 & ~A203;
  assign \new_[92739]_  = A267 & ~A266;
  assign \new_[92740]_  = \new_[92739]_  & \new_[92736]_ ;
  assign \new_[92743]_  = A300 & A269;
  assign \new_[92746]_  = ~A302 & ~A301;
  assign \new_[92747]_  = \new_[92746]_  & \new_[92743]_ ;
  assign \new_[92748]_  = \new_[92747]_  & \new_[92740]_ ;
  assign \new_[92751]_  = A168 & A169;
  assign \new_[92754]_  = A166 & ~A167;
  assign \new_[92755]_  = \new_[92754]_  & \new_[92751]_ ;
  assign \new_[92758]_  = A200 & ~A199;
  assign \new_[92761]_  = ~A202 & ~A201;
  assign \new_[92762]_  = \new_[92761]_  & \new_[92758]_ ;
  assign \new_[92763]_  = \new_[92762]_  & \new_[92755]_ ;
  assign \new_[92766]_  = A265 & ~A203;
  assign \new_[92769]_  = ~A267 & ~A266;
  assign \new_[92770]_  = \new_[92769]_  & \new_[92766]_ ;
  assign \new_[92773]_  = ~A269 & ~A268;
  assign \new_[92776]_  = A301 & ~A300;
  assign \new_[92777]_  = \new_[92776]_  & \new_[92773]_ ;
  assign \new_[92778]_  = \new_[92777]_  & \new_[92770]_ ;
  assign \new_[92781]_  = A168 & A169;
  assign \new_[92784]_  = A166 & ~A167;
  assign \new_[92785]_  = \new_[92784]_  & \new_[92781]_ ;
  assign \new_[92788]_  = A200 & ~A199;
  assign \new_[92791]_  = ~A202 & ~A201;
  assign \new_[92792]_  = \new_[92791]_  & \new_[92788]_ ;
  assign \new_[92793]_  = \new_[92792]_  & \new_[92785]_ ;
  assign \new_[92796]_  = A265 & ~A203;
  assign \new_[92799]_  = ~A267 & ~A266;
  assign \new_[92800]_  = \new_[92799]_  & \new_[92796]_ ;
  assign \new_[92803]_  = ~A269 & ~A268;
  assign \new_[92806]_  = A302 & ~A300;
  assign \new_[92807]_  = \new_[92806]_  & \new_[92803]_ ;
  assign \new_[92808]_  = \new_[92807]_  & \new_[92800]_ ;
  assign \new_[92811]_  = A168 & A169;
  assign \new_[92814]_  = A166 & ~A167;
  assign \new_[92815]_  = \new_[92814]_  & \new_[92811]_ ;
  assign \new_[92818]_  = A200 & ~A199;
  assign \new_[92821]_  = ~A202 & ~A201;
  assign \new_[92822]_  = \new_[92821]_  & \new_[92818]_ ;
  assign \new_[92823]_  = \new_[92822]_  & \new_[92815]_ ;
  assign \new_[92826]_  = A265 & ~A203;
  assign \new_[92829]_  = ~A267 & ~A266;
  assign \new_[92830]_  = \new_[92829]_  & \new_[92826]_ ;
  assign \new_[92833]_  = ~A269 & ~A268;
  assign \new_[92836]_  = A299 & A298;
  assign \new_[92837]_  = \new_[92836]_  & \new_[92833]_ ;
  assign \new_[92838]_  = \new_[92837]_  & \new_[92830]_ ;
  assign \new_[92841]_  = A168 & A169;
  assign \new_[92844]_  = A166 & ~A167;
  assign \new_[92845]_  = \new_[92844]_  & \new_[92841]_ ;
  assign \new_[92848]_  = A200 & ~A199;
  assign \new_[92851]_  = ~A202 & ~A201;
  assign \new_[92852]_  = \new_[92851]_  & \new_[92848]_ ;
  assign \new_[92853]_  = \new_[92852]_  & \new_[92845]_ ;
  assign \new_[92856]_  = A265 & ~A203;
  assign \new_[92859]_  = ~A267 & ~A266;
  assign \new_[92860]_  = \new_[92859]_  & \new_[92856]_ ;
  assign \new_[92863]_  = ~A269 & ~A268;
  assign \new_[92866]_  = ~A299 & ~A298;
  assign \new_[92867]_  = \new_[92866]_  & \new_[92863]_ ;
  assign \new_[92868]_  = \new_[92867]_  & \new_[92860]_ ;
  assign \new_[92871]_  = A168 & A169;
  assign \new_[92874]_  = A166 & ~A167;
  assign \new_[92875]_  = \new_[92874]_  & \new_[92871]_ ;
  assign \new_[92878]_  = ~A200 & A199;
  assign \new_[92881]_  = A202 & A201;
  assign \new_[92882]_  = \new_[92881]_  & \new_[92878]_ ;
  assign \new_[92883]_  = \new_[92882]_  & \new_[92875]_ ;
  assign \new_[92886]_  = A266 & ~A265;
  assign \new_[92889]_  = ~A268 & ~A267;
  assign \new_[92890]_  = \new_[92889]_  & \new_[92886]_ ;
  assign \new_[92893]_  = A300 & ~A269;
  assign \new_[92896]_  = ~A302 & ~A301;
  assign \new_[92897]_  = \new_[92896]_  & \new_[92893]_ ;
  assign \new_[92898]_  = \new_[92897]_  & \new_[92890]_ ;
  assign \new_[92901]_  = A168 & A169;
  assign \new_[92904]_  = A166 & ~A167;
  assign \new_[92905]_  = \new_[92904]_  & \new_[92901]_ ;
  assign \new_[92908]_  = ~A200 & A199;
  assign \new_[92911]_  = A202 & A201;
  assign \new_[92912]_  = \new_[92911]_  & \new_[92908]_ ;
  assign \new_[92913]_  = \new_[92912]_  & \new_[92905]_ ;
  assign \new_[92916]_  = ~A266 & A265;
  assign \new_[92919]_  = ~A268 & ~A267;
  assign \new_[92920]_  = \new_[92919]_  & \new_[92916]_ ;
  assign \new_[92923]_  = A300 & ~A269;
  assign \new_[92926]_  = ~A302 & ~A301;
  assign \new_[92927]_  = \new_[92926]_  & \new_[92923]_ ;
  assign \new_[92928]_  = \new_[92927]_  & \new_[92920]_ ;
  assign \new_[92931]_  = A168 & A169;
  assign \new_[92934]_  = A166 & ~A167;
  assign \new_[92935]_  = \new_[92934]_  & \new_[92931]_ ;
  assign \new_[92938]_  = ~A200 & A199;
  assign \new_[92941]_  = A203 & A201;
  assign \new_[92942]_  = \new_[92941]_  & \new_[92938]_ ;
  assign \new_[92943]_  = \new_[92942]_  & \new_[92935]_ ;
  assign \new_[92946]_  = A266 & ~A265;
  assign \new_[92949]_  = ~A268 & ~A267;
  assign \new_[92950]_  = \new_[92949]_  & \new_[92946]_ ;
  assign \new_[92953]_  = A300 & ~A269;
  assign \new_[92956]_  = ~A302 & ~A301;
  assign \new_[92957]_  = \new_[92956]_  & \new_[92953]_ ;
  assign \new_[92958]_  = \new_[92957]_  & \new_[92950]_ ;
  assign \new_[92961]_  = A168 & A169;
  assign \new_[92964]_  = A166 & ~A167;
  assign \new_[92965]_  = \new_[92964]_  & \new_[92961]_ ;
  assign \new_[92968]_  = ~A200 & A199;
  assign \new_[92971]_  = A203 & A201;
  assign \new_[92972]_  = \new_[92971]_  & \new_[92968]_ ;
  assign \new_[92973]_  = \new_[92972]_  & \new_[92965]_ ;
  assign \new_[92976]_  = ~A266 & A265;
  assign \new_[92979]_  = ~A268 & ~A267;
  assign \new_[92980]_  = \new_[92979]_  & \new_[92976]_ ;
  assign \new_[92983]_  = A300 & ~A269;
  assign \new_[92986]_  = ~A302 & ~A301;
  assign \new_[92987]_  = \new_[92986]_  & \new_[92983]_ ;
  assign \new_[92988]_  = \new_[92987]_  & \new_[92980]_ ;
  assign \new_[92991]_  = A168 & A169;
  assign \new_[92994]_  = A166 & ~A167;
  assign \new_[92995]_  = \new_[92994]_  & \new_[92991]_ ;
  assign \new_[92998]_  = ~A200 & A199;
  assign \new_[93001]_  = ~A202 & ~A201;
  assign \new_[93002]_  = \new_[93001]_  & \new_[92998]_ ;
  assign \new_[93003]_  = \new_[93002]_  & \new_[92995]_ ;
  assign \new_[93006]_  = ~A265 & ~A203;
  assign \new_[93009]_  = A267 & A266;
  assign \new_[93010]_  = \new_[93009]_  & \new_[93006]_ ;
  assign \new_[93013]_  = A300 & A268;
  assign \new_[93016]_  = ~A302 & ~A301;
  assign \new_[93017]_  = \new_[93016]_  & \new_[93013]_ ;
  assign \new_[93018]_  = \new_[93017]_  & \new_[93010]_ ;
  assign \new_[93021]_  = A168 & A169;
  assign \new_[93024]_  = A166 & ~A167;
  assign \new_[93025]_  = \new_[93024]_  & \new_[93021]_ ;
  assign \new_[93028]_  = ~A200 & A199;
  assign \new_[93031]_  = ~A202 & ~A201;
  assign \new_[93032]_  = \new_[93031]_  & \new_[93028]_ ;
  assign \new_[93033]_  = \new_[93032]_  & \new_[93025]_ ;
  assign \new_[93036]_  = ~A265 & ~A203;
  assign \new_[93039]_  = A267 & A266;
  assign \new_[93040]_  = \new_[93039]_  & \new_[93036]_ ;
  assign \new_[93043]_  = A300 & A269;
  assign \new_[93046]_  = ~A302 & ~A301;
  assign \new_[93047]_  = \new_[93046]_  & \new_[93043]_ ;
  assign \new_[93048]_  = \new_[93047]_  & \new_[93040]_ ;
  assign \new_[93051]_  = A168 & A169;
  assign \new_[93054]_  = A166 & ~A167;
  assign \new_[93055]_  = \new_[93054]_  & \new_[93051]_ ;
  assign \new_[93058]_  = ~A200 & A199;
  assign \new_[93061]_  = ~A202 & ~A201;
  assign \new_[93062]_  = \new_[93061]_  & \new_[93058]_ ;
  assign \new_[93063]_  = \new_[93062]_  & \new_[93055]_ ;
  assign \new_[93066]_  = ~A265 & ~A203;
  assign \new_[93069]_  = ~A267 & A266;
  assign \new_[93070]_  = \new_[93069]_  & \new_[93066]_ ;
  assign \new_[93073]_  = ~A269 & ~A268;
  assign \new_[93076]_  = A301 & ~A300;
  assign \new_[93077]_  = \new_[93076]_  & \new_[93073]_ ;
  assign \new_[93078]_  = \new_[93077]_  & \new_[93070]_ ;
  assign \new_[93081]_  = A168 & A169;
  assign \new_[93084]_  = A166 & ~A167;
  assign \new_[93085]_  = \new_[93084]_  & \new_[93081]_ ;
  assign \new_[93088]_  = ~A200 & A199;
  assign \new_[93091]_  = ~A202 & ~A201;
  assign \new_[93092]_  = \new_[93091]_  & \new_[93088]_ ;
  assign \new_[93093]_  = \new_[93092]_  & \new_[93085]_ ;
  assign \new_[93096]_  = ~A265 & ~A203;
  assign \new_[93099]_  = ~A267 & A266;
  assign \new_[93100]_  = \new_[93099]_  & \new_[93096]_ ;
  assign \new_[93103]_  = ~A269 & ~A268;
  assign \new_[93106]_  = A302 & ~A300;
  assign \new_[93107]_  = \new_[93106]_  & \new_[93103]_ ;
  assign \new_[93108]_  = \new_[93107]_  & \new_[93100]_ ;
  assign \new_[93111]_  = A168 & A169;
  assign \new_[93114]_  = A166 & ~A167;
  assign \new_[93115]_  = \new_[93114]_  & \new_[93111]_ ;
  assign \new_[93118]_  = ~A200 & A199;
  assign \new_[93121]_  = ~A202 & ~A201;
  assign \new_[93122]_  = \new_[93121]_  & \new_[93118]_ ;
  assign \new_[93123]_  = \new_[93122]_  & \new_[93115]_ ;
  assign \new_[93126]_  = ~A265 & ~A203;
  assign \new_[93129]_  = ~A267 & A266;
  assign \new_[93130]_  = \new_[93129]_  & \new_[93126]_ ;
  assign \new_[93133]_  = ~A269 & ~A268;
  assign \new_[93136]_  = A299 & A298;
  assign \new_[93137]_  = \new_[93136]_  & \new_[93133]_ ;
  assign \new_[93138]_  = \new_[93137]_  & \new_[93130]_ ;
  assign \new_[93141]_  = A168 & A169;
  assign \new_[93144]_  = A166 & ~A167;
  assign \new_[93145]_  = \new_[93144]_  & \new_[93141]_ ;
  assign \new_[93148]_  = ~A200 & A199;
  assign \new_[93151]_  = ~A202 & ~A201;
  assign \new_[93152]_  = \new_[93151]_  & \new_[93148]_ ;
  assign \new_[93153]_  = \new_[93152]_  & \new_[93145]_ ;
  assign \new_[93156]_  = ~A265 & ~A203;
  assign \new_[93159]_  = ~A267 & A266;
  assign \new_[93160]_  = \new_[93159]_  & \new_[93156]_ ;
  assign \new_[93163]_  = ~A269 & ~A268;
  assign \new_[93166]_  = ~A299 & ~A298;
  assign \new_[93167]_  = \new_[93166]_  & \new_[93163]_ ;
  assign \new_[93168]_  = \new_[93167]_  & \new_[93160]_ ;
  assign \new_[93171]_  = A168 & A169;
  assign \new_[93174]_  = A166 & ~A167;
  assign \new_[93175]_  = \new_[93174]_  & \new_[93171]_ ;
  assign \new_[93178]_  = ~A200 & A199;
  assign \new_[93181]_  = ~A202 & ~A201;
  assign \new_[93182]_  = \new_[93181]_  & \new_[93178]_ ;
  assign \new_[93183]_  = \new_[93182]_  & \new_[93175]_ ;
  assign \new_[93186]_  = A265 & ~A203;
  assign \new_[93189]_  = A267 & ~A266;
  assign \new_[93190]_  = \new_[93189]_  & \new_[93186]_ ;
  assign \new_[93193]_  = A300 & A268;
  assign \new_[93196]_  = ~A302 & ~A301;
  assign \new_[93197]_  = \new_[93196]_  & \new_[93193]_ ;
  assign \new_[93198]_  = \new_[93197]_  & \new_[93190]_ ;
  assign \new_[93201]_  = A168 & A169;
  assign \new_[93204]_  = A166 & ~A167;
  assign \new_[93205]_  = \new_[93204]_  & \new_[93201]_ ;
  assign \new_[93208]_  = ~A200 & A199;
  assign \new_[93211]_  = ~A202 & ~A201;
  assign \new_[93212]_  = \new_[93211]_  & \new_[93208]_ ;
  assign \new_[93213]_  = \new_[93212]_  & \new_[93205]_ ;
  assign \new_[93216]_  = A265 & ~A203;
  assign \new_[93219]_  = A267 & ~A266;
  assign \new_[93220]_  = \new_[93219]_  & \new_[93216]_ ;
  assign \new_[93223]_  = A300 & A269;
  assign \new_[93226]_  = ~A302 & ~A301;
  assign \new_[93227]_  = \new_[93226]_  & \new_[93223]_ ;
  assign \new_[93228]_  = \new_[93227]_  & \new_[93220]_ ;
  assign \new_[93231]_  = A168 & A169;
  assign \new_[93234]_  = A166 & ~A167;
  assign \new_[93235]_  = \new_[93234]_  & \new_[93231]_ ;
  assign \new_[93238]_  = ~A200 & A199;
  assign \new_[93241]_  = ~A202 & ~A201;
  assign \new_[93242]_  = \new_[93241]_  & \new_[93238]_ ;
  assign \new_[93243]_  = \new_[93242]_  & \new_[93235]_ ;
  assign \new_[93246]_  = A265 & ~A203;
  assign \new_[93249]_  = ~A267 & ~A266;
  assign \new_[93250]_  = \new_[93249]_  & \new_[93246]_ ;
  assign \new_[93253]_  = ~A269 & ~A268;
  assign \new_[93256]_  = A301 & ~A300;
  assign \new_[93257]_  = \new_[93256]_  & \new_[93253]_ ;
  assign \new_[93258]_  = \new_[93257]_  & \new_[93250]_ ;
  assign \new_[93261]_  = A168 & A169;
  assign \new_[93264]_  = A166 & ~A167;
  assign \new_[93265]_  = \new_[93264]_  & \new_[93261]_ ;
  assign \new_[93268]_  = ~A200 & A199;
  assign \new_[93271]_  = ~A202 & ~A201;
  assign \new_[93272]_  = \new_[93271]_  & \new_[93268]_ ;
  assign \new_[93273]_  = \new_[93272]_  & \new_[93265]_ ;
  assign \new_[93276]_  = A265 & ~A203;
  assign \new_[93279]_  = ~A267 & ~A266;
  assign \new_[93280]_  = \new_[93279]_  & \new_[93276]_ ;
  assign \new_[93283]_  = ~A269 & ~A268;
  assign \new_[93286]_  = A302 & ~A300;
  assign \new_[93287]_  = \new_[93286]_  & \new_[93283]_ ;
  assign \new_[93288]_  = \new_[93287]_  & \new_[93280]_ ;
  assign \new_[93291]_  = A168 & A169;
  assign \new_[93294]_  = A166 & ~A167;
  assign \new_[93295]_  = \new_[93294]_  & \new_[93291]_ ;
  assign \new_[93298]_  = ~A200 & A199;
  assign \new_[93301]_  = ~A202 & ~A201;
  assign \new_[93302]_  = \new_[93301]_  & \new_[93298]_ ;
  assign \new_[93303]_  = \new_[93302]_  & \new_[93295]_ ;
  assign \new_[93306]_  = A265 & ~A203;
  assign \new_[93309]_  = ~A267 & ~A266;
  assign \new_[93310]_  = \new_[93309]_  & \new_[93306]_ ;
  assign \new_[93313]_  = ~A269 & ~A268;
  assign \new_[93316]_  = A299 & A298;
  assign \new_[93317]_  = \new_[93316]_  & \new_[93313]_ ;
  assign \new_[93318]_  = \new_[93317]_  & \new_[93310]_ ;
  assign \new_[93321]_  = A168 & A169;
  assign \new_[93324]_  = A166 & ~A167;
  assign \new_[93325]_  = \new_[93324]_  & \new_[93321]_ ;
  assign \new_[93328]_  = ~A200 & A199;
  assign \new_[93331]_  = ~A202 & ~A201;
  assign \new_[93332]_  = \new_[93331]_  & \new_[93328]_ ;
  assign \new_[93333]_  = \new_[93332]_  & \new_[93325]_ ;
  assign \new_[93336]_  = A265 & ~A203;
  assign \new_[93339]_  = ~A267 & ~A266;
  assign \new_[93340]_  = \new_[93339]_  & \new_[93336]_ ;
  assign \new_[93343]_  = ~A269 & ~A268;
  assign \new_[93346]_  = ~A299 & ~A298;
  assign \new_[93347]_  = \new_[93346]_  & \new_[93343]_ ;
  assign \new_[93348]_  = \new_[93347]_  & \new_[93340]_ ;
  assign \new_[93351]_  = ~A169 & A170;
  assign \new_[93354]_  = ~A199 & A168;
  assign \new_[93355]_  = \new_[93354]_  & \new_[93351]_ ;
  assign \new_[93358]_  = ~A201 & A200;
  assign \new_[93361]_  = ~A203 & ~A202;
  assign \new_[93362]_  = \new_[93361]_  & \new_[93358]_ ;
  assign \new_[93363]_  = \new_[93362]_  & \new_[93355]_ ;
  assign \new_[93366]_  = ~A268 & A267;
  assign \new_[93369]_  = A298 & ~A269;
  assign \new_[93370]_  = \new_[93369]_  & \new_[93366]_ ;
  assign \new_[93373]_  = ~A300 & ~A299;
  assign \new_[93376]_  = ~A302 & ~A301;
  assign \new_[93377]_  = \new_[93376]_  & \new_[93373]_ ;
  assign \new_[93378]_  = \new_[93377]_  & \new_[93370]_ ;
  assign \new_[93381]_  = ~A169 & A170;
  assign \new_[93384]_  = ~A199 & A168;
  assign \new_[93385]_  = \new_[93384]_  & \new_[93381]_ ;
  assign \new_[93388]_  = ~A201 & A200;
  assign \new_[93391]_  = ~A203 & ~A202;
  assign \new_[93392]_  = \new_[93391]_  & \new_[93388]_ ;
  assign \new_[93393]_  = \new_[93392]_  & \new_[93385]_ ;
  assign \new_[93396]_  = ~A268 & A267;
  assign \new_[93399]_  = ~A298 & ~A269;
  assign \new_[93400]_  = \new_[93399]_  & \new_[93396]_ ;
  assign \new_[93403]_  = ~A300 & A299;
  assign \new_[93406]_  = ~A302 & ~A301;
  assign \new_[93407]_  = \new_[93406]_  & \new_[93403]_ ;
  assign \new_[93408]_  = \new_[93407]_  & \new_[93400]_ ;
  assign \new_[93411]_  = ~A169 & A170;
  assign \new_[93414]_  = A199 & A168;
  assign \new_[93415]_  = \new_[93414]_  & \new_[93411]_ ;
  assign \new_[93418]_  = ~A201 & ~A200;
  assign \new_[93421]_  = ~A203 & ~A202;
  assign \new_[93422]_  = \new_[93421]_  & \new_[93418]_ ;
  assign \new_[93423]_  = \new_[93422]_  & \new_[93415]_ ;
  assign \new_[93426]_  = ~A268 & A267;
  assign \new_[93429]_  = A298 & ~A269;
  assign \new_[93430]_  = \new_[93429]_  & \new_[93426]_ ;
  assign \new_[93433]_  = ~A300 & ~A299;
  assign \new_[93436]_  = ~A302 & ~A301;
  assign \new_[93437]_  = \new_[93436]_  & \new_[93433]_ ;
  assign \new_[93438]_  = \new_[93437]_  & \new_[93430]_ ;
  assign \new_[93441]_  = ~A169 & A170;
  assign \new_[93444]_  = A199 & A168;
  assign \new_[93445]_  = \new_[93444]_  & \new_[93441]_ ;
  assign \new_[93448]_  = ~A201 & ~A200;
  assign \new_[93451]_  = ~A203 & ~A202;
  assign \new_[93452]_  = \new_[93451]_  & \new_[93448]_ ;
  assign \new_[93453]_  = \new_[93452]_  & \new_[93445]_ ;
  assign \new_[93456]_  = ~A268 & A267;
  assign \new_[93459]_  = ~A298 & ~A269;
  assign \new_[93460]_  = \new_[93459]_  & \new_[93456]_ ;
  assign \new_[93463]_  = ~A300 & A299;
  assign \new_[93466]_  = ~A302 & ~A301;
  assign \new_[93467]_  = \new_[93466]_  & \new_[93463]_ ;
  assign \new_[93468]_  = \new_[93467]_  & \new_[93460]_ ;
  assign \new_[93471]_  = ~A169 & A170;
  assign \new_[93474]_  = A167 & ~A168;
  assign \new_[93475]_  = \new_[93474]_  & \new_[93471]_ ;
  assign \new_[93478]_  = A201 & ~A166;
  assign \new_[93481]_  = ~A203 & ~A202;
  assign \new_[93482]_  = \new_[93481]_  & \new_[93478]_ ;
  assign \new_[93483]_  = \new_[93482]_  & \new_[93475]_ ;
  assign \new_[93486]_  = ~A268 & A267;
  assign \new_[93489]_  = A298 & ~A269;
  assign \new_[93490]_  = \new_[93489]_  & \new_[93486]_ ;
  assign \new_[93493]_  = ~A300 & ~A299;
  assign \new_[93496]_  = ~A302 & ~A301;
  assign \new_[93497]_  = \new_[93496]_  & \new_[93493]_ ;
  assign \new_[93498]_  = \new_[93497]_  & \new_[93490]_ ;
  assign \new_[93501]_  = ~A169 & A170;
  assign \new_[93504]_  = A167 & ~A168;
  assign \new_[93505]_  = \new_[93504]_  & \new_[93501]_ ;
  assign \new_[93508]_  = A201 & ~A166;
  assign \new_[93511]_  = ~A203 & ~A202;
  assign \new_[93512]_  = \new_[93511]_  & \new_[93508]_ ;
  assign \new_[93513]_  = \new_[93512]_  & \new_[93505]_ ;
  assign \new_[93516]_  = ~A268 & A267;
  assign \new_[93519]_  = ~A298 & ~A269;
  assign \new_[93520]_  = \new_[93519]_  & \new_[93516]_ ;
  assign \new_[93523]_  = ~A300 & A299;
  assign \new_[93526]_  = ~A302 & ~A301;
  assign \new_[93527]_  = \new_[93526]_  & \new_[93523]_ ;
  assign \new_[93528]_  = \new_[93527]_  & \new_[93520]_ ;
  assign \new_[93531]_  = ~A169 & A170;
  assign \new_[93534]_  = A167 & ~A168;
  assign \new_[93535]_  = \new_[93534]_  & \new_[93531]_ ;
  assign \new_[93538]_  = ~A199 & ~A166;
  assign \new_[93541]_  = A201 & A200;
  assign \new_[93542]_  = \new_[93541]_  & \new_[93538]_ ;
  assign \new_[93543]_  = \new_[93542]_  & \new_[93535]_ ;
  assign \new_[93546]_  = ~A265 & A202;
  assign \new_[93549]_  = A267 & A266;
  assign \new_[93550]_  = \new_[93549]_  & \new_[93546]_ ;
  assign \new_[93553]_  = A300 & A268;
  assign \new_[93556]_  = ~A302 & ~A301;
  assign \new_[93557]_  = \new_[93556]_  & \new_[93553]_ ;
  assign \new_[93558]_  = \new_[93557]_  & \new_[93550]_ ;
  assign \new_[93561]_  = ~A169 & A170;
  assign \new_[93564]_  = A167 & ~A168;
  assign \new_[93565]_  = \new_[93564]_  & \new_[93561]_ ;
  assign \new_[93568]_  = ~A199 & ~A166;
  assign \new_[93571]_  = A201 & A200;
  assign \new_[93572]_  = \new_[93571]_  & \new_[93568]_ ;
  assign \new_[93573]_  = \new_[93572]_  & \new_[93565]_ ;
  assign \new_[93576]_  = ~A265 & A202;
  assign \new_[93579]_  = A267 & A266;
  assign \new_[93580]_  = \new_[93579]_  & \new_[93576]_ ;
  assign \new_[93583]_  = A300 & A269;
  assign \new_[93586]_  = ~A302 & ~A301;
  assign \new_[93587]_  = \new_[93586]_  & \new_[93583]_ ;
  assign \new_[93588]_  = \new_[93587]_  & \new_[93580]_ ;
  assign \new_[93591]_  = ~A169 & A170;
  assign \new_[93594]_  = A167 & ~A168;
  assign \new_[93595]_  = \new_[93594]_  & \new_[93591]_ ;
  assign \new_[93598]_  = ~A199 & ~A166;
  assign \new_[93601]_  = A201 & A200;
  assign \new_[93602]_  = \new_[93601]_  & \new_[93598]_ ;
  assign \new_[93603]_  = \new_[93602]_  & \new_[93595]_ ;
  assign \new_[93606]_  = ~A265 & A202;
  assign \new_[93609]_  = ~A267 & A266;
  assign \new_[93610]_  = \new_[93609]_  & \new_[93606]_ ;
  assign \new_[93613]_  = ~A269 & ~A268;
  assign \new_[93616]_  = A301 & ~A300;
  assign \new_[93617]_  = \new_[93616]_  & \new_[93613]_ ;
  assign \new_[93618]_  = \new_[93617]_  & \new_[93610]_ ;
  assign \new_[93621]_  = ~A169 & A170;
  assign \new_[93624]_  = A167 & ~A168;
  assign \new_[93625]_  = \new_[93624]_  & \new_[93621]_ ;
  assign \new_[93628]_  = ~A199 & ~A166;
  assign \new_[93631]_  = A201 & A200;
  assign \new_[93632]_  = \new_[93631]_  & \new_[93628]_ ;
  assign \new_[93633]_  = \new_[93632]_  & \new_[93625]_ ;
  assign \new_[93636]_  = ~A265 & A202;
  assign \new_[93639]_  = ~A267 & A266;
  assign \new_[93640]_  = \new_[93639]_  & \new_[93636]_ ;
  assign \new_[93643]_  = ~A269 & ~A268;
  assign \new_[93646]_  = A302 & ~A300;
  assign \new_[93647]_  = \new_[93646]_  & \new_[93643]_ ;
  assign \new_[93648]_  = \new_[93647]_  & \new_[93640]_ ;
  assign \new_[93651]_  = ~A169 & A170;
  assign \new_[93654]_  = A167 & ~A168;
  assign \new_[93655]_  = \new_[93654]_  & \new_[93651]_ ;
  assign \new_[93658]_  = ~A199 & ~A166;
  assign \new_[93661]_  = A201 & A200;
  assign \new_[93662]_  = \new_[93661]_  & \new_[93658]_ ;
  assign \new_[93663]_  = \new_[93662]_  & \new_[93655]_ ;
  assign \new_[93666]_  = ~A265 & A202;
  assign \new_[93669]_  = ~A267 & A266;
  assign \new_[93670]_  = \new_[93669]_  & \new_[93666]_ ;
  assign \new_[93673]_  = ~A269 & ~A268;
  assign \new_[93676]_  = A299 & A298;
  assign \new_[93677]_  = \new_[93676]_  & \new_[93673]_ ;
  assign \new_[93678]_  = \new_[93677]_  & \new_[93670]_ ;
  assign \new_[93681]_  = ~A169 & A170;
  assign \new_[93684]_  = A167 & ~A168;
  assign \new_[93685]_  = \new_[93684]_  & \new_[93681]_ ;
  assign \new_[93688]_  = ~A199 & ~A166;
  assign \new_[93691]_  = A201 & A200;
  assign \new_[93692]_  = \new_[93691]_  & \new_[93688]_ ;
  assign \new_[93693]_  = \new_[93692]_  & \new_[93685]_ ;
  assign \new_[93696]_  = ~A265 & A202;
  assign \new_[93699]_  = ~A267 & A266;
  assign \new_[93700]_  = \new_[93699]_  & \new_[93696]_ ;
  assign \new_[93703]_  = ~A269 & ~A268;
  assign \new_[93706]_  = ~A299 & ~A298;
  assign \new_[93707]_  = \new_[93706]_  & \new_[93703]_ ;
  assign \new_[93708]_  = \new_[93707]_  & \new_[93700]_ ;
  assign \new_[93711]_  = ~A169 & A170;
  assign \new_[93714]_  = A167 & ~A168;
  assign \new_[93715]_  = \new_[93714]_  & \new_[93711]_ ;
  assign \new_[93718]_  = ~A199 & ~A166;
  assign \new_[93721]_  = A201 & A200;
  assign \new_[93722]_  = \new_[93721]_  & \new_[93718]_ ;
  assign \new_[93723]_  = \new_[93722]_  & \new_[93715]_ ;
  assign \new_[93726]_  = A265 & A202;
  assign \new_[93729]_  = A267 & ~A266;
  assign \new_[93730]_  = \new_[93729]_  & \new_[93726]_ ;
  assign \new_[93733]_  = A300 & A268;
  assign \new_[93736]_  = ~A302 & ~A301;
  assign \new_[93737]_  = \new_[93736]_  & \new_[93733]_ ;
  assign \new_[93738]_  = \new_[93737]_  & \new_[93730]_ ;
  assign \new_[93741]_  = ~A169 & A170;
  assign \new_[93744]_  = A167 & ~A168;
  assign \new_[93745]_  = \new_[93744]_  & \new_[93741]_ ;
  assign \new_[93748]_  = ~A199 & ~A166;
  assign \new_[93751]_  = A201 & A200;
  assign \new_[93752]_  = \new_[93751]_  & \new_[93748]_ ;
  assign \new_[93753]_  = \new_[93752]_  & \new_[93745]_ ;
  assign \new_[93756]_  = A265 & A202;
  assign \new_[93759]_  = A267 & ~A266;
  assign \new_[93760]_  = \new_[93759]_  & \new_[93756]_ ;
  assign \new_[93763]_  = A300 & A269;
  assign \new_[93766]_  = ~A302 & ~A301;
  assign \new_[93767]_  = \new_[93766]_  & \new_[93763]_ ;
  assign \new_[93768]_  = \new_[93767]_  & \new_[93760]_ ;
  assign \new_[93771]_  = ~A169 & A170;
  assign \new_[93774]_  = A167 & ~A168;
  assign \new_[93775]_  = \new_[93774]_  & \new_[93771]_ ;
  assign \new_[93778]_  = ~A199 & ~A166;
  assign \new_[93781]_  = A201 & A200;
  assign \new_[93782]_  = \new_[93781]_  & \new_[93778]_ ;
  assign \new_[93783]_  = \new_[93782]_  & \new_[93775]_ ;
  assign \new_[93786]_  = A265 & A202;
  assign \new_[93789]_  = ~A267 & ~A266;
  assign \new_[93790]_  = \new_[93789]_  & \new_[93786]_ ;
  assign \new_[93793]_  = ~A269 & ~A268;
  assign \new_[93796]_  = A301 & ~A300;
  assign \new_[93797]_  = \new_[93796]_  & \new_[93793]_ ;
  assign \new_[93798]_  = \new_[93797]_  & \new_[93790]_ ;
  assign \new_[93801]_  = ~A169 & A170;
  assign \new_[93804]_  = A167 & ~A168;
  assign \new_[93805]_  = \new_[93804]_  & \new_[93801]_ ;
  assign \new_[93808]_  = ~A199 & ~A166;
  assign \new_[93811]_  = A201 & A200;
  assign \new_[93812]_  = \new_[93811]_  & \new_[93808]_ ;
  assign \new_[93813]_  = \new_[93812]_  & \new_[93805]_ ;
  assign \new_[93816]_  = A265 & A202;
  assign \new_[93819]_  = ~A267 & ~A266;
  assign \new_[93820]_  = \new_[93819]_  & \new_[93816]_ ;
  assign \new_[93823]_  = ~A269 & ~A268;
  assign \new_[93826]_  = A302 & ~A300;
  assign \new_[93827]_  = \new_[93826]_  & \new_[93823]_ ;
  assign \new_[93828]_  = \new_[93827]_  & \new_[93820]_ ;
  assign \new_[93831]_  = ~A169 & A170;
  assign \new_[93834]_  = A167 & ~A168;
  assign \new_[93835]_  = \new_[93834]_  & \new_[93831]_ ;
  assign \new_[93838]_  = ~A199 & ~A166;
  assign \new_[93841]_  = A201 & A200;
  assign \new_[93842]_  = \new_[93841]_  & \new_[93838]_ ;
  assign \new_[93843]_  = \new_[93842]_  & \new_[93835]_ ;
  assign \new_[93846]_  = A265 & A202;
  assign \new_[93849]_  = ~A267 & ~A266;
  assign \new_[93850]_  = \new_[93849]_  & \new_[93846]_ ;
  assign \new_[93853]_  = ~A269 & ~A268;
  assign \new_[93856]_  = A299 & A298;
  assign \new_[93857]_  = \new_[93856]_  & \new_[93853]_ ;
  assign \new_[93858]_  = \new_[93857]_  & \new_[93850]_ ;
  assign \new_[93861]_  = ~A169 & A170;
  assign \new_[93864]_  = A167 & ~A168;
  assign \new_[93865]_  = \new_[93864]_  & \new_[93861]_ ;
  assign \new_[93868]_  = ~A199 & ~A166;
  assign \new_[93871]_  = A201 & A200;
  assign \new_[93872]_  = \new_[93871]_  & \new_[93868]_ ;
  assign \new_[93873]_  = \new_[93872]_  & \new_[93865]_ ;
  assign \new_[93876]_  = A265 & A202;
  assign \new_[93879]_  = ~A267 & ~A266;
  assign \new_[93880]_  = \new_[93879]_  & \new_[93876]_ ;
  assign \new_[93883]_  = ~A269 & ~A268;
  assign \new_[93886]_  = ~A299 & ~A298;
  assign \new_[93887]_  = \new_[93886]_  & \new_[93883]_ ;
  assign \new_[93888]_  = \new_[93887]_  & \new_[93880]_ ;
  assign \new_[93891]_  = ~A169 & A170;
  assign \new_[93894]_  = A167 & ~A168;
  assign \new_[93895]_  = \new_[93894]_  & \new_[93891]_ ;
  assign \new_[93898]_  = ~A199 & ~A166;
  assign \new_[93901]_  = A201 & A200;
  assign \new_[93902]_  = \new_[93901]_  & \new_[93898]_ ;
  assign \new_[93903]_  = \new_[93902]_  & \new_[93895]_ ;
  assign \new_[93906]_  = ~A265 & A203;
  assign \new_[93909]_  = A267 & A266;
  assign \new_[93910]_  = \new_[93909]_  & \new_[93906]_ ;
  assign \new_[93913]_  = A300 & A268;
  assign \new_[93916]_  = ~A302 & ~A301;
  assign \new_[93917]_  = \new_[93916]_  & \new_[93913]_ ;
  assign \new_[93918]_  = \new_[93917]_  & \new_[93910]_ ;
  assign \new_[93921]_  = ~A169 & A170;
  assign \new_[93924]_  = A167 & ~A168;
  assign \new_[93925]_  = \new_[93924]_  & \new_[93921]_ ;
  assign \new_[93928]_  = ~A199 & ~A166;
  assign \new_[93931]_  = A201 & A200;
  assign \new_[93932]_  = \new_[93931]_  & \new_[93928]_ ;
  assign \new_[93933]_  = \new_[93932]_  & \new_[93925]_ ;
  assign \new_[93936]_  = ~A265 & A203;
  assign \new_[93939]_  = A267 & A266;
  assign \new_[93940]_  = \new_[93939]_  & \new_[93936]_ ;
  assign \new_[93943]_  = A300 & A269;
  assign \new_[93946]_  = ~A302 & ~A301;
  assign \new_[93947]_  = \new_[93946]_  & \new_[93943]_ ;
  assign \new_[93948]_  = \new_[93947]_  & \new_[93940]_ ;
  assign \new_[93951]_  = ~A169 & A170;
  assign \new_[93954]_  = A167 & ~A168;
  assign \new_[93955]_  = \new_[93954]_  & \new_[93951]_ ;
  assign \new_[93958]_  = ~A199 & ~A166;
  assign \new_[93961]_  = A201 & A200;
  assign \new_[93962]_  = \new_[93961]_  & \new_[93958]_ ;
  assign \new_[93963]_  = \new_[93962]_  & \new_[93955]_ ;
  assign \new_[93966]_  = ~A265 & A203;
  assign \new_[93969]_  = ~A267 & A266;
  assign \new_[93970]_  = \new_[93969]_  & \new_[93966]_ ;
  assign \new_[93973]_  = ~A269 & ~A268;
  assign \new_[93976]_  = A301 & ~A300;
  assign \new_[93977]_  = \new_[93976]_  & \new_[93973]_ ;
  assign \new_[93978]_  = \new_[93977]_  & \new_[93970]_ ;
  assign \new_[93981]_  = ~A169 & A170;
  assign \new_[93984]_  = A167 & ~A168;
  assign \new_[93985]_  = \new_[93984]_  & \new_[93981]_ ;
  assign \new_[93988]_  = ~A199 & ~A166;
  assign \new_[93991]_  = A201 & A200;
  assign \new_[93992]_  = \new_[93991]_  & \new_[93988]_ ;
  assign \new_[93993]_  = \new_[93992]_  & \new_[93985]_ ;
  assign \new_[93996]_  = ~A265 & A203;
  assign \new_[93999]_  = ~A267 & A266;
  assign \new_[94000]_  = \new_[93999]_  & \new_[93996]_ ;
  assign \new_[94003]_  = ~A269 & ~A268;
  assign \new_[94006]_  = A302 & ~A300;
  assign \new_[94007]_  = \new_[94006]_  & \new_[94003]_ ;
  assign \new_[94008]_  = \new_[94007]_  & \new_[94000]_ ;
  assign \new_[94011]_  = ~A169 & A170;
  assign \new_[94014]_  = A167 & ~A168;
  assign \new_[94015]_  = \new_[94014]_  & \new_[94011]_ ;
  assign \new_[94018]_  = ~A199 & ~A166;
  assign \new_[94021]_  = A201 & A200;
  assign \new_[94022]_  = \new_[94021]_  & \new_[94018]_ ;
  assign \new_[94023]_  = \new_[94022]_  & \new_[94015]_ ;
  assign \new_[94026]_  = ~A265 & A203;
  assign \new_[94029]_  = ~A267 & A266;
  assign \new_[94030]_  = \new_[94029]_  & \new_[94026]_ ;
  assign \new_[94033]_  = ~A269 & ~A268;
  assign \new_[94036]_  = A299 & A298;
  assign \new_[94037]_  = \new_[94036]_  & \new_[94033]_ ;
  assign \new_[94038]_  = \new_[94037]_  & \new_[94030]_ ;
  assign \new_[94041]_  = ~A169 & A170;
  assign \new_[94044]_  = A167 & ~A168;
  assign \new_[94045]_  = \new_[94044]_  & \new_[94041]_ ;
  assign \new_[94048]_  = ~A199 & ~A166;
  assign \new_[94051]_  = A201 & A200;
  assign \new_[94052]_  = \new_[94051]_  & \new_[94048]_ ;
  assign \new_[94053]_  = \new_[94052]_  & \new_[94045]_ ;
  assign \new_[94056]_  = ~A265 & A203;
  assign \new_[94059]_  = ~A267 & A266;
  assign \new_[94060]_  = \new_[94059]_  & \new_[94056]_ ;
  assign \new_[94063]_  = ~A269 & ~A268;
  assign \new_[94066]_  = ~A299 & ~A298;
  assign \new_[94067]_  = \new_[94066]_  & \new_[94063]_ ;
  assign \new_[94068]_  = \new_[94067]_  & \new_[94060]_ ;
  assign \new_[94071]_  = ~A169 & A170;
  assign \new_[94074]_  = A167 & ~A168;
  assign \new_[94075]_  = \new_[94074]_  & \new_[94071]_ ;
  assign \new_[94078]_  = ~A199 & ~A166;
  assign \new_[94081]_  = A201 & A200;
  assign \new_[94082]_  = \new_[94081]_  & \new_[94078]_ ;
  assign \new_[94083]_  = \new_[94082]_  & \new_[94075]_ ;
  assign \new_[94086]_  = A265 & A203;
  assign \new_[94089]_  = A267 & ~A266;
  assign \new_[94090]_  = \new_[94089]_  & \new_[94086]_ ;
  assign \new_[94093]_  = A300 & A268;
  assign \new_[94096]_  = ~A302 & ~A301;
  assign \new_[94097]_  = \new_[94096]_  & \new_[94093]_ ;
  assign \new_[94098]_  = \new_[94097]_  & \new_[94090]_ ;
  assign \new_[94101]_  = ~A169 & A170;
  assign \new_[94104]_  = A167 & ~A168;
  assign \new_[94105]_  = \new_[94104]_  & \new_[94101]_ ;
  assign \new_[94108]_  = ~A199 & ~A166;
  assign \new_[94111]_  = A201 & A200;
  assign \new_[94112]_  = \new_[94111]_  & \new_[94108]_ ;
  assign \new_[94113]_  = \new_[94112]_  & \new_[94105]_ ;
  assign \new_[94116]_  = A265 & A203;
  assign \new_[94119]_  = A267 & ~A266;
  assign \new_[94120]_  = \new_[94119]_  & \new_[94116]_ ;
  assign \new_[94123]_  = A300 & A269;
  assign \new_[94126]_  = ~A302 & ~A301;
  assign \new_[94127]_  = \new_[94126]_  & \new_[94123]_ ;
  assign \new_[94128]_  = \new_[94127]_  & \new_[94120]_ ;
  assign \new_[94131]_  = ~A169 & A170;
  assign \new_[94134]_  = A167 & ~A168;
  assign \new_[94135]_  = \new_[94134]_  & \new_[94131]_ ;
  assign \new_[94138]_  = ~A199 & ~A166;
  assign \new_[94141]_  = A201 & A200;
  assign \new_[94142]_  = \new_[94141]_  & \new_[94138]_ ;
  assign \new_[94143]_  = \new_[94142]_  & \new_[94135]_ ;
  assign \new_[94146]_  = A265 & A203;
  assign \new_[94149]_  = ~A267 & ~A266;
  assign \new_[94150]_  = \new_[94149]_  & \new_[94146]_ ;
  assign \new_[94153]_  = ~A269 & ~A268;
  assign \new_[94156]_  = A301 & ~A300;
  assign \new_[94157]_  = \new_[94156]_  & \new_[94153]_ ;
  assign \new_[94158]_  = \new_[94157]_  & \new_[94150]_ ;
  assign \new_[94161]_  = ~A169 & A170;
  assign \new_[94164]_  = A167 & ~A168;
  assign \new_[94165]_  = \new_[94164]_  & \new_[94161]_ ;
  assign \new_[94168]_  = ~A199 & ~A166;
  assign \new_[94171]_  = A201 & A200;
  assign \new_[94172]_  = \new_[94171]_  & \new_[94168]_ ;
  assign \new_[94173]_  = \new_[94172]_  & \new_[94165]_ ;
  assign \new_[94176]_  = A265 & A203;
  assign \new_[94179]_  = ~A267 & ~A266;
  assign \new_[94180]_  = \new_[94179]_  & \new_[94176]_ ;
  assign \new_[94183]_  = ~A269 & ~A268;
  assign \new_[94186]_  = A302 & ~A300;
  assign \new_[94187]_  = \new_[94186]_  & \new_[94183]_ ;
  assign \new_[94188]_  = \new_[94187]_  & \new_[94180]_ ;
  assign \new_[94191]_  = ~A169 & A170;
  assign \new_[94194]_  = A167 & ~A168;
  assign \new_[94195]_  = \new_[94194]_  & \new_[94191]_ ;
  assign \new_[94198]_  = ~A199 & ~A166;
  assign \new_[94201]_  = A201 & A200;
  assign \new_[94202]_  = \new_[94201]_  & \new_[94198]_ ;
  assign \new_[94203]_  = \new_[94202]_  & \new_[94195]_ ;
  assign \new_[94206]_  = A265 & A203;
  assign \new_[94209]_  = ~A267 & ~A266;
  assign \new_[94210]_  = \new_[94209]_  & \new_[94206]_ ;
  assign \new_[94213]_  = ~A269 & ~A268;
  assign \new_[94216]_  = A299 & A298;
  assign \new_[94217]_  = \new_[94216]_  & \new_[94213]_ ;
  assign \new_[94218]_  = \new_[94217]_  & \new_[94210]_ ;
  assign \new_[94221]_  = ~A169 & A170;
  assign \new_[94224]_  = A167 & ~A168;
  assign \new_[94225]_  = \new_[94224]_  & \new_[94221]_ ;
  assign \new_[94228]_  = ~A199 & ~A166;
  assign \new_[94231]_  = A201 & A200;
  assign \new_[94232]_  = \new_[94231]_  & \new_[94228]_ ;
  assign \new_[94233]_  = \new_[94232]_  & \new_[94225]_ ;
  assign \new_[94236]_  = A265 & A203;
  assign \new_[94239]_  = ~A267 & ~A266;
  assign \new_[94240]_  = \new_[94239]_  & \new_[94236]_ ;
  assign \new_[94243]_  = ~A269 & ~A268;
  assign \new_[94246]_  = ~A299 & ~A298;
  assign \new_[94247]_  = \new_[94246]_  & \new_[94243]_ ;
  assign \new_[94248]_  = \new_[94247]_  & \new_[94240]_ ;
  assign \new_[94251]_  = ~A169 & A170;
  assign \new_[94254]_  = A167 & ~A168;
  assign \new_[94255]_  = \new_[94254]_  & \new_[94251]_ ;
  assign \new_[94258]_  = ~A199 & ~A166;
  assign \new_[94261]_  = ~A201 & A200;
  assign \new_[94262]_  = \new_[94261]_  & \new_[94258]_ ;
  assign \new_[94263]_  = \new_[94262]_  & \new_[94255]_ ;
  assign \new_[94266]_  = ~A203 & ~A202;
  assign \new_[94269]_  = A266 & ~A265;
  assign \new_[94270]_  = \new_[94269]_  & \new_[94266]_ ;
  assign \new_[94273]_  = A268 & A267;
  assign \new_[94276]_  = A301 & ~A300;
  assign \new_[94277]_  = \new_[94276]_  & \new_[94273]_ ;
  assign \new_[94278]_  = \new_[94277]_  & \new_[94270]_ ;
  assign \new_[94281]_  = ~A169 & A170;
  assign \new_[94284]_  = A167 & ~A168;
  assign \new_[94285]_  = \new_[94284]_  & \new_[94281]_ ;
  assign \new_[94288]_  = ~A199 & ~A166;
  assign \new_[94291]_  = ~A201 & A200;
  assign \new_[94292]_  = \new_[94291]_  & \new_[94288]_ ;
  assign \new_[94293]_  = \new_[94292]_  & \new_[94285]_ ;
  assign \new_[94296]_  = ~A203 & ~A202;
  assign \new_[94299]_  = A266 & ~A265;
  assign \new_[94300]_  = \new_[94299]_  & \new_[94296]_ ;
  assign \new_[94303]_  = A268 & A267;
  assign \new_[94306]_  = A302 & ~A300;
  assign \new_[94307]_  = \new_[94306]_  & \new_[94303]_ ;
  assign \new_[94308]_  = \new_[94307]_  & \new_[94300]_ ;
  assign \new_[94311]_  = ~A169 & A170;
  assign \new_[94314]_  = A167 & ~A168;
  assign \new_[94315]_  = \new_[94314]_  & \new_[94311]_ ;
  assign \new_[94318]_  = ~A199 & ~A166;
  assign \new_[94321]_  = ~A201 & A200;
  assign \new_[94322]_  = \new_[94321]_  & \new_[94318]_ ;
  assign \new_[94323]_  = \new_[94322]_  & \new_[94315]_ ;
  assign \new_[94326]_  = ~A203 & ~A202;
  assign \new_[94329]_  = A266 & ~A265;
  assign \new_[94330]_  = \new_[94329]_  & \new_[94326]_ ;
  assign \new_[94333]_  = A268 & A267;
  assign \new_[94336]_  = A299 & A298;
  assign \new_[94337]_  = \new_[94336]_  & \new_[94333]_ ;
  assign \new_[94338]_  = \new_[94337]_  & \new_[94330]_ ;
  assign \new_[94341]_  = ~A169 & A170;
  assign \new_[94344]_  = A167 & ~A168;
  assign \new_[94345]_  = \new_[94344]_  & \new_[94341]_ ;
  assign \new_[94348]_  = ~A199 & ~A166;
  assign \new_[94351]_  = ~A201 & A200;
  assign \new_[94352]_  = \new_[94351]_  & \new_[94348]_ ;
  assign \new_[94353]_  = \new_[94352]_  & \new_[94345]_ ;
  assign \new_[94356]_  = ~A203 & ~A202;
  assign \new_[94359]_  = A266 & ~A265;
  assign \new_[94360]_  = \new_[94359]_  & \new_[94356]_ ;
  assign \new_[94363]_  = A268 & A267;
  assign \new_[94366]_  = ~A299 & ~A298;
  assign \new_[94367]_  = \new_[94366]_  & \new_[94363]_ ;
  assign \new_[94368]_  = \new_[94367]_  & \new_[94360]_ ;
  assign \new_[94371]_  = ~A169 & A170;
  assign \new_[94374]_  = A167 & ~A168;
  assign \new_[94375]_  = \new_[94374]_  & \new_[94371]_ ;
  assign \new_[94378]_  = ~A199 & ~A166;
  assign \new_[94381]_  = ~A201 & A200;
  assign \new_[94382]_  = \new_[94381]_  & \new_[94378]_ ;
  assign \new_[94383]_  = \new_[94382]_  & \new_[94375]_ ;
  assign \new_[94386]_  = ~A203 & ~A202;
  assign \new_[94389]_  = A266 & ~A265;
  assign \new_[94390]_  = \new_[94389]_  & \new_[94386]_ ;
  assign \new_[94393]_  = A269 & A267;
  assign \new_[94396]_  = A301 & ~A300;
  assign \new_[94397]_  = \new_[94396]_  & \new_[94393]_ ;
  assign \new_[94398]_  = \new_[94397]_  & \new_[94390]_ ;
  assign \new_[94401]_  = ~A169 & A170;
  assign \new_[94404]_  = A167 & ~A168;
  assign \new_[94405]_  = \new_[94404]_  & \new_[94401]_ ;
  assign \new_[94408]_  = ~A199 & ~A166;
  assign \new_[94411]_  = ~A201 & A200;
  assign \new_[94412]_  = \new_[94411]_  & \new_[94408]_ ;
  assign \new_[94413]_  = \new_[94412]_  & \new_[94405]_ ;
  assign \new_[94416]_  = ~A203 & ~A202;
  assign \new_[94419]_  = A266 & ~A265;
  assign \new_[94420]_  = \new_[94419]_  & \new_[94416]_ ;
  assign \new_[94423]_  = A269 & A267;
  assign \new_[94426]_  = A302 & ~A300;
  assign \new_[94427]_  = \new_[94426]_  & \new_[94423]_ ;
  assign \new_[94428]_  = \new_[94427]_  & \new_[94420]_ ;
  assign \new_[94431]_  = ~A169 & A170;
  assign \new_[94434]_  = A167 & ~A168;
  assign \new_[94435]_  = \new_[94434]_  & \new_[94431]_ ;
  assign \new_[94438]_  = ~A199 & ~A166;
  assign \new_[94441]_  = ~A201 & A200;
  assign \new_[94442]_  = \new_[94441]_  & \new_[94438]_ ;
  assign \new_[94443]_  = \new_[94442]_  & \new_[94435]_ ;
  assign \new_[94446]_  = ~A203 & ~A202;
  assign \new_[94449]_  = A266 & ~A265;
  assign \new_[94450]_  = \new_[94449]_  & \new_[94446]_ ;
  assign \new_[94453]_  = A269 & A267;
  assign \new_[94456]_  = A299 & A298;
  assign \new_[94457]_  = \new_[94456]_  & \new_[94453]_ ;
  assign \new_[94458]_  = \new_[94457]_  & \new_[94450]_ ;
  assign \new_[94461]_  = ~A169 & A170;
  assign \new_[94464]_  = A167 & ~A168;
  assign \new_[94465]_  = \new_[94464]_  & \new_[94461]_ ;
  assign \new_[94468]_  = ~A199 & ~A166;
  assign \new_[94471]_  = ~A201 & A200;
  assign \new_[94472]_  = \new_[94471]_  & \new_[94468]_ ;
  assign \new_[94473]_  = \new_[94472]_  & \new_[94465]_ ;
  assign \new_[94476]_  = ~A203 & ~A202;
  assign \new_[94479]_  = A266 & ~A265;
  assign \new_[94480]_  = \new_[94479]_  & \new_[94476]_ ;
  assign \new_[94483]_  = A269 & A267;
  assign \new_[94486]_  = ~A299 & ~A298;
  assign \new_[94487]_  = \new_[94486]_  & \new_[94483]_ ;
  assign \new_[94488]_  = \new_[94487]_  & \new_[94480]_ ;
  assign \new_[94491]_  = ~A169 & A170;
  assign \new_[94494]_  = A167 & ~A168;
  assign \new_[94495]_  = \new_[94494]_  & \new_[94491]_ ;
  assign \new_[94498]_  = ~A199 & ~A166;
  assign \new_[94501]_  = ~A201 & A200;
  assign \new_[94502]_  = \new_[94501]_  & \new_[94498]_ ;
  assign \new_[94503]_  = \new_[94502]_  & \new_[94495]_ ;
  assign \new_[94506]_  = ~A203 & ~A202;
  assign \new_[94509]_  = ~A266 & A265;
  assign \new_[94510]_  = \new_[94509]_  & \new_[94506]_ ;
  assign \new_[94513]_  = A268 & A267;
  assign \new_[94516]_  = A301 & ~A300;
  assign \new_[94517]_  = \new_[94516]_  & \new_[94513]_ ;
  assign \new_[94518]_  = \new_[94517]_  & \new_[94510]_ ;
  assign \new_[94521]_  = ~A169 & A170;
  assign \new_[94524]_  = A167 & ~A168;
  assign \new_[94525]_  = \new_[94524]_  & \new_[94521]_ ;
  assign \new_[94528]_  = ~A199 & ~A166;
  assign \new_[94531]_  = ~A201 & A200;
  assign \new_[94532]_  = \new_[94531]_  & \new_[94528]_ ;
  assign \new_[94533]_  = \new_[94532]_  & \new_[94525]_ ;
  assign \new_[94536]_  = ~A203 & ~A202;
  assign \new_[94539]_  = ~A266 & A265;
  assign \new_[94540]_  = \new_[94539]_  & \new_[94536]_ ;
  assign \new_[94543]_  = A268 & A267;
  assign \new_[94546]_  = A302 & ~A300;
  assign \new_[94547]_  = \new_[94546]_  & \new_[94543]_ ;
  assign \new_[94548]_  = \new_[94547]_  & \new_[94540]_ ;
  assign \new_[94551]_  = ~A169 & A170;
  assign \new_[94554]_  = A167 & ~A168;
  assign \new_[94555]_  = \new_[94554]_  & \new_[94551]_ ;
  assign \new_[94558]_  = ~A199 & ~A166;
  assign \new_[94561]_  = ~A201 & A200;
  assign \new_[94562]_  = \new_[94561]_  & \new_[94558]_ ;
  assign \new_[94563]_  = \new_[94562]_  & \new_[94555]_ ;
  assign \new_[94566]_  = ~A203 & ~A202;
  assign \new_[94569]_  = ~A266 & A265;
  assign \new_[94570]_  = \new_[94569]_  & \new_[94566]_ ;
  assign \new_[94573]_  = A268 & A267;
  assign \new_[94576]_  = A299 & A298;
  assign \new_[94577]_  = \new_[94576]_  & \new_[94573]_ ;
  assign \new_[94578]_  = \new_[94577]_  & \new_[94570]_ ;
  assign \new_[94581]_  = ~A169 & A170;
  assign \new_[94584]_  = A167 & ~A168;
  assign \new_[94585]_  = \new_[94584]_  & \new_[94581]_ ;
  assign \new_[94588]_  = ~A199 & ~A166;
  assign \new_[94591]_  = ~A201 & A200;
  assign \new_[94592]_  = \new_[94591]_  & \new_[94588]_ ;
  assign \new_[94593]_  = \new_[94592]_  & \new_[94585]_ ;
  assign \new_[94596]_  = ~A203 & ~A202;
  assign \new_[94599]_  = ~A266 & A265;
  assign \new_[94600]_  = \new_[94599]_  & \new_[94596]_ ;
  assign \new_[94603]_  = A268 & A267;
  assign \new_[94606]_  = ~A299 & ~A298;
  assign \new_[94607]_  = \new_[94606]_  & \new_[94603]_ ;
  assign \new_[94608]_  = \new_[94607]_  & \new_[94600]_ ;
  assign \new_[94611]_  = ~A169 & A170;
  assign \new_[94614]_  = A167 & ~A168;
  assign \new_[94615]_  = \new_[94614]_  & \new_[94611]_ ;
  assign \new_[94618]_  = ~A199 & ~A166;
  assign \new_[94621]_  = ~A201 & A200;
  assign \new_[94622]_  = \new_[94621]_  & \new_[94618]_ ;
  assign \new_[94623]_  = \new_[94622]_  & \new_[94615]_ ;
  assign \new_[94626]_  = ~A203 & ~A202;
  assign \new_[94629]_  = ~A266 & A265;
  assign \new_[94630]_  = \new_[94629]_  & \new_[94626]_ ;
  assign \new_[94633]_  = A269 & A267;
  assign \new_[94636]_  = A301 & ~A300;
  assign \new_[94637]_  = \new_[94636]_  & \new_[94633]_ ;
  assign \new_[94638]_  = \new_[94637]_  & \new_[94630]_ ;
  assign \new_[94641]_  = ~A169 & A170;
  assign \new_[94644]_  = A167 & ~A168;
  assign \new_[94645]_  = \new_[94644]_  & \new_[94641]_ ;
  assign \new_[94648]_  = ~A199 & ~A166;
  assign \new_[94651]_  = ~A201 & A200;
  assign \new_[94652]_  = \new_[94651]_  & \new_[94648]_ ;
  assign \new_[94653]_  = \new_[94652]_  & \new_[94645]_ ;
  assign \new_[94656]_  = ~A203 & ~A202;
  assign \new_[94659]_  = ~A266 & A265;
  assign \new_[94660]_  = \new_[94659]_  & \new_[94656]_ ;
  assign \new_[94663]_  = A269 & A267;
  assign \new_[94666]_  = A302 & ~A300;
  assign \new_[94667]_  = \new_[94666]_  & \new_[94663]_ ;
  assign \new_[94668]_  = \new_[94667]_  & \new_[94660]_ ;
  assign \new_[94671]_  = ~A169 & A170;
  assign \new_[94674]_  = A167 & ~A168;
  assign \new_[94675]_  = \new_[94674]_  & \new_[94671]_ ;
  assign \new_[94678]_  = ~A199 & ~A166;
  assign \new_[94681]_  = ~A201 & A200;
  assign \new_[94682]_  = \new_[94681]_  & \new_[94678]_ ;
  assign \new_[94683]_  = \new_[94682]_  & \new_[94675]_ ;
  assign \new_[94686]_  = ~A203 & ~A202;
  assign \new_[94689]_  = ~A266 & A265;
  assign \new_[94690]_  = \new_[94689]_  & \new_[94686]_ ;
  assign \new_[94693]_  = A269 & A267;
  assign \new_[94696]_  = A299 & A298;
  assign \new_[94697]_  = \new_[94696]_  & \new_[94693]_ ;
  assign \new_[94698]_  = \new_[94697]_  & \new_[94690]_ ;
  assign \new_[94701]_  = ~A169 & A170;
  assign \new_[94704]_  = A167 & ~A168;
  assign \new_[94705]_  = \new_[94704]_  & \new_[94701]_ ;
  assign \new_[94708]_  = ~A199 & ~A166;
  assign \new_[94711]_  = ~A201 & A200;
  assign \new_[94712]_  = \new_[94711]_  & \new_[94708]_ ;
  assign \new_[94713]_  = \new_[94712]_  & \new_[94705]_ ;
  assign \new_[94716]_  = ~A203 & ~A202;
  assign \new_[94719]_  = ~A266 & A265;
  assign \new_[94720]_  = \new_[94719]_  & \new_[94716]_ ;
  assign \new_[94723]_  = A269 & A267;
  assign \new_[94726]_  = ~A299 & ~A298;
  assign \new_[94727]_  = \new_[94726]_  & \new_[94723]_ ;
  assign \new_[94728]_  = \new_[94727]_  & \new_[94720]_ ;
  assign \new_[94731]_  = ~A169 & A170;
  assign \new_[94734]_  = A167 & ~A168;
  assign \new_[94735]_  = \new_[94734]_  & \new_[94731]_ ;
  assign \new_[94738]_  = A199 & ~A166;
  assign \new_[94741]_  = A201 & ~A200;
  assign \new_[94742]_  = \new_[94741]_  & \new_[94738]_ ;
  assign \new_[94743]_  = \new_[94742]_  & \new_[94735]_ ;
  assign \new_[94746]_  = ~A265 & A202;
  assign \new_[94749]_  = A267 & A266;
  assign \new_[94750]_  = \new_[94749]_  & \new_[94746]_ ;
  assign \new_[94753]_  = A300 & A268;
  assign \new_[94756]_  = ~A302 & ~A301;
  assign \new_[94757]_  = \new_[94756]_  & \new_[94753]_ ;
  assign \new_[94758]_  = \new_[94757]_  & \new_[94750]_ ;
  assign \new_[94761]_  = ~A169 & A170;
  assign \new_[94764]_  = A167 & ~A168;
  assign \new_[94765]_  = \new_[94764]_  & \new_[94761]_ ;
  assign \new_[94768]_  = A199 & ~A166;
  assign \new_[94771]_  = A201 & ~A200;
  assign \new_[94772]_  = \new_[94771]_  & \new_[94768]_ ;
  assign \new_[94773]_  = \new_[94772]_  & \new_[94765]_ ;
  assign \new_[94776]_  = ~A265 & A202;
  assign \new_[94779]_  = A267 & A266;
  assign \new_[94780]_  = \new_[94779]_  & \new_[94776]_ ;
  assign \new_[94783]_  = A300 & A269;
  assign \new_[94786]_  = ~A302 & ~A301;
  assign \new_[94787]_  = \new_[94786]_  & \new_[94783]_ ;
  assign \new_[94788]_  = \new_[94787]_  & \new_[94780]_ ;
  assign \new_[94791]_  = ~A169 & A170;
  assign \new_[94794]_  = A167 & ~A168;
  assign \new_[94795]_  = \new_[94794]_  & \new_[94791]_ ;
  assign \new_[94798]_  = A199 & ~A166;
  assign \new_[94801]_  = A201 & ~A200;
  assign \new_[94802]_  = \new_[94801]_  & \new_[94798]_ ;
  assign \new_[94803]_  = \new_[94802]_  & \new_[94795]_ ;
  assign \new_[94806]_  = ~A265 & A202;
  assign \new_[94809]_  = ~A267 & A266;
  assign \new_[94810]_  = \new_[94809]_  & \new_[94806]_ ;
  assign \new_[94813]_  = ~A269 & ~A268;
  assign \new_[94816]_  = A301 & ~A300;
  assign \new_[94817]_  = \new_[94816]_  & \new_[94813]_ ;
  assign \new_[94818]_  = \new_[94817]_  & \new_[94810]_ ;
  assign \new_[94821]_  = ~A169 & A170;
  assign \new_[94824]_  = A167 & ~A168;
  assign \new_[94825]_  = \new_[94824]_  & \new_[94821]_ ;
  assign \new_[94828]_  = A199 & ~A166;
  assign \new_[94831]_  = A201 & ~A200;
  assign \new_[94832]_  = \new_[94831]_  & \new_[94828]_ ;
  assign \new_[94833]_  = \new_[94832]_  & \new_[94825]_ ;
  assign \new_[94836]_  = ~A265 & A202;
  assign \new_[94839]_  = ~A267 & A266;
  assign \new_[94840]_  = \new_[94839]_  & \new_[94836]_ ;
  assign \new_[94843]_  = ~A269 & ~A268;
  assign \new_[94846]_  = A302 & ~A300;
  assign \new_[94847]_  = \new_[94846]_  & \new_[94843]_ ;
  assign \new_[94848]_  = \new_[94847]_  & \new_[94840]_ ;
  assign \new_[94851]_  = ~A169 & A170;
  assign \new_[94854]_  = A167 & ~A168;
  assign \new_[94855]_  = \new_[94854]_  & \new_[94851]_ ;
  assign \new_[94858]_  = A199 & ~A166;
  assign \new_[94861]_  = A201 & ~A200;
  assign \new_[94862]_  = \new_[94861]_  & \new_[94858]_ ;
  assign \new_[94863]_  = \new_[94862]_  & \new_[94855]_ ;
  assign \new_[94866]_  = ~A265 & A202;
  assign \new_[94869]_  = ~A267 & A266;
  assign \new_[94870]_  = \new_[94869]_  & \new_[94866]_ ;
  assign \new_[94873]_  = ~A269 & ~A268;
  assign \new_[94876]_  = A299 & A298;
  assign \new_[94877]_  = \new_[94876]_  & \new_[94873]_ ;
  assign \new_[94878]_  = \new_[94877]_  & \new_[94870]_ ;
  assign \new_[94881]_  = ~A169 & A170;
  assign \new_[94884]_  = A167 & ~A168;
  assign \new_[94885]_  = \new_[94884]_  & \new_[94881]_ ;
  assign \new_[94888]_  = A199 & ~A166;
  assign \new_[94891]_  = A201 & ~A200;
  assign \new_[94892]_  = \new_[94891]_  & \new_[94888]_ ;
  assign \new_[94893]_  = \new_[94892]_  & \new_[94885]_ ;
  assign \new_[94896]_  = ~A265 & A202;
  assign \new_[94899]_  = ~A267 & A266;
  assign \new_[94900]_  = \new_[94899]_  & \new_[94896]_ ;
  assign \new_[94903]_  = ~A269 & ~A268;
  assign \new_[94906]_  = ~A299 & ~A298;
  assign \new_[94907]_  = \new_[94906]_  & \new_[94903]_ ;
  assign \new_[94908]_  = \new_[94907]_  & \new_[94900]_ ;
  assign \new_[94911]_  = ~A169 & A170;
  assign \new_[94914]_  = A167 & ~A168;
  assign \new_[94915]_  = \new_[94914]_  & \new_[94911]_ ;
  assign \new_[94918]_  = A199 & ~A166;
  assign \new_[94921]_  = A201 & ~A200;
  assign \new_[94922]_  = \new_[94921]_  & \new_[94918]_ ;
  assign \new_[94923]_  = \new_[94922]_  & \new_[94915]_ ;
  assign \new_[94926]_  = A265 & A202;
  assign \new_[94929]_  = A267 & ~A266;
  assign \new_[94930]_  = \new_[94929]_  & \new_[94926]_ ;
  assign \new_[94933]_  = A300 & A268;
  assign \new_[94936]_  = ~A302 & ~A301;
  assign \new_[94937]_  = \new_[94936]_  & \new_[94933]_ ;
  assign \new_[94938]_  = \new_[94937]_  & \new_[94930]_ ;
  assign \new_[94941]_  = ~A169 & A170;
  assign \new_[94944]_  = A167 & ~A168;
  assign \new_[94945]_  = \new_[94944]_  & \new_[94941]_ ;
  assign \new_[94948]_  = A199 & ~A166;
  assign \new_[94951]_  = A201 & ~A200;
  assign \new_[94952]_  = \new_[94951]_  & \new_[94948]_ ;
  assign \new_[94953]_  = \new_[94952]_  & \new_[94945]_ ;
  assign \new_[94956]_  = A265 & A202;
  assign \new_[94959]_  = A267 & ~A266;
  assign \new_[94960]_  = \new_[94959]_  & \new_[94956]_ ;
  assign \new_[94963]_  = A300 & A269;
  assign \new_[94966]_  = ~A302 & ~A301;
  assign \new_[94967]_  = \new_[94966]_  & \new_[94963]_ ;
  assign \new_[94968]_  = \new_[94967]_  & \new_[94960]_ ;
  assign \new_[94971]_  = ~A169 & A170;
  assign \new_[94974]_  = A167 & ~A168;
  assign \new_[94975]_  = \new_[94974]_  & \new_[94971]_ ;
  assign \new_[94978]_  = A199 & ~A166;
  assign \new_[94981]_  = A201 & ~A200;
  assign \new_[94982]_  = \new_[94981]_  & \new_[94978]_ ;
  assign \new_[94983]_  = \new_[94982]_  & \new_[94975]_ ;
  assign \new_[94986]_  = A265 & A202;
  assign \new_[94989]_  = ~A267 & ~A266;
  assign \new_[94990]_  = \new_[94989]_  & \new_[94986]_ ;
  assign \new_[94993]_  = ~A269 & ~A268;
  assign \new_[94996]_  = A301 & ~A300;
  assign \new_[94997]_  = \new_[94996]_  & \new_[94993]_ ;
  assign \new_[94998]_  = \new_[94997]_  & \new_[94990]_ ;
  assign \new_[95001]_  = ~A169 & A170;
  assign \new_[95004]_  = A167 & ~A168;
  assign \new_[95005]_  = \new_[95004]_  & \new_[95001]_ ;
  assign \new_[95008]_  = A199 & ~A166;
  assign \new_[95011]_  = A201 & ~A200;
  assign \new_[95012]_  = \new_[95011]_  & \new_[95008]_ ;
  assign \new_[95013]_  = \new_[95012]_  & \new_[95005]_ ;
  assign \new_[95016]_  = A265 & A202;
  assign \new_[95019]_  = ~A267 & ~A266;
  assign \new_[95020]_  = \new_[95019]_  & \new_[95016]_ ;
  assign \new_[95023]_  = ~A269 & ~A268;
  assign \new_[95026]_  = A302 & ~A300;
  assign \new_[95027]_  = \new_[95026]_  & \new_[95023]_ ;
  assign \new_[95028]_  = \new_[95027]_  & \new_[95020]_ ;
  assign \new_[95031]_  = ~A169 & A170;
  assign \new_[95034]_  = A167 & ~A168;
  assign \new_[95035]_  = \new_[95034]_  & \new_[95031]_ ;
  assign \new_[95038]_  = A199 & ~A166;
  assign \new_[95041]_  = A201 & ~A200;
  assign \new_[95042]_  = \new_[95041]_  & \new_[95038]_ ;
  assign \new_[95043]_  = \new_[95042]_  & \new_[95035]_ ;
  assign \new_[95046]_  = A265 & A202;
  assign \new_[95049]_  = ~A267 & ~A266;
  assign \new_[95050]_  = \new_[95049]_  & \new_[95046]_ ;
  assign \new_[95053]_  = ~A269 & ~A268;
  assign \new_[95056]_  = A299 & A298;
  assign \new_[95057]_  = \new_[95056]_  & \new_[95053]_ ;
  assign \new_[95058]_  = \new_[95057]_  & \new_[95050]_ ;
  assign \new_[95061]_  = ~A169 & A170;
  assign \new_[95064]_  = A167 & ~A168;
  assign \new_[95065]_  = \new_[95064]_  & \new_[95061]_ ;
  assign \new_[95068]_  = A199 & ~A166;
  assign \new_[95071]_  = A201 & ~A200;
  assign \new_[95072]_  = \new_[95071]_  & \new_[95068]_ ;
  assign \new_[95073]_  = \new_[95072]_  & \new_[95065]_ ;
  assign \new_[95076]_  = A265 & A202;
  assign \new_[95079]_  = ~A267 & ~A266;
  assign \new_[95080]_  = \new_[95079]_  & \new_[95076]_ ;
  assign \new_[95083]_  = ~A269 & ~A268;
  assign \new_[95086]_  = ~A299 & ~A298;
  assign \new_[95087]_  = \new_[95086]_  & \new_[95083]_ ;
  assign \new_[95088]_  = \new_[95087]_  & \new_[95080]_ ;
  assign \new_[95091]_  = ~A169 & A170;
  assign \new_[95094]_  = A167 & ~A168;
  assign \new_[95095]_  = \new_[95094]_  & \new_[95091]_ ;
  assign \new_[95098]_  = A199 & ~A166;
  assign \new_[95101]_  = A201 & ~A200;
  assign \new_[95102]_  = \new_[95101]_  & \new_[95098]_ ;
  assign \new_[95103]_  = \new_[95102]_  & \new_[95095]_ ;
  assign \new_[95106]_  = ~A265 & A203;
  assign \new_[95109]_  = A267 & A266;
  assign \new_[95110]_  = \new_[95109]_  & \new_[95106]_ ;
  assign \new_[95113]_  = A300 & A268;
  assign \new_[95116]_  = ~A302 & ~A301;
  assign \new_[95117]_  = \new_[95116]_  & \new_[95113]_ ;
  assign \new_[95118]_  = \new_[95117]_  & \new_[95110]_ ;
  assign \new_[95121]_  = ~A169 & A170;
  assign \new_[95124]_  = A167 & ~A168;
  assign \new_[95125]_  = \new_[95124]_  & \new_[95121]_ ;
  assign \new_[95128]_  = A199 & ~A166;
  assign \new_[95131]_  = A201 & ~A200;
  assign \new_[95132]_  = \new_[95131]_  & \new_[95128]_ ;
  assign \new_[95133]_  = \new_[95132]_  & \new_[95125]_ ;
  assign \new_[95136]_  = ~A265 & A203;
  assign \new_[95139]_  = A267 & A266;
  assign \new_[95140]_  = \new_[95139]_  & \new_[95136]_ ;
  assign \new_[95143]_  = A300 & A269;
  assign \new_[95146]_  = ~A302 & ~A301;
  assign \new_[95147]_  = \new_[95146]_  & \new_[95143]_ ;
  assign \new_[95148]_  = \new_[95147]_  & \new_[95140]_ ;
  assign \new_[95151]_  = ~A169 & A170;
  assign \new_[95154]_  = A167 & ~A168;
  assign \new_[95155]_  = \new_[95154]_  & \new_[95151]_ ;
  assign \new_[95158]_  = A199 & ~A166;
  assign \new_[95161]_  = A201 & ~A200;
  assign \new_[95162]_  = \new_[95161]_  & \new_[95158]_ ;
  assign \new_[95163]_  = \new_[95162]_  & \new_[95155]_ ;
  assign \new_[95166]_  = ~A265 & A203;
  assign \new_[95169]_  = ~A267 & A266;
  assign \new_[95170]_  = \new_[95169]_  & \new_[95166]_ ;
  assign \new_[95173]_  = ~A269 & ~A268;
  assign \new_[95176]_  = A301 & ~A300;
  assign \new_[95177]_  = \new_[95176]_  & \new_[95173]_ ;
  assign \new_[95178]_  = \new_[95177]_  & \new_[95170]_ ;
  assign \new_[95181]_  = ~A169 & A170;
  assign \new_[95184]_  = A167 & ~A168;
  assign \new_[95185]_  = \new_[95184]_  & \new_[95181]_ ;
  assign \new_[95188]_  = A199 & ~A166;
  assign \new_[95191]_  = A201 & ~A200;
  assign \new_[95192]_  = \new_[95191]_  & \new_[95188]_ ;
  assign \new_[95193]_  = \new_[95192]_  & \new_[95185]_ ;
  assign \new_[95196]_  = ~A265 & A203;
  assign \new_[95199]_  = ~A267 & A266;
  assign \new_[95200]_  = \new_[95199]_  & \new_[95196]_ ;
  assign \new_[95203]_  = ~A269 & ~A268;
  assign \new_[95206]_  = A302 & ~A300;
  assign \new_[95207]_  = \new_[95206]_  & \new_[95203]_ ;
  assign \new_[95208]_  = \new_[95207]_  & \new_[95200]_ ;
  assign \new_[95211]_  = ~A169 & A170;
  assign \new_[95214]_  = A167 & ~A168;
  assign \new_[95215]_  = \new_[95214]_  & \new_[95211]_ ;
  assign \new_[95218]_  = A199 & ~A166;
  assign \new_[95221]_  = A201 & ~A200;
  assign \new_[95222]_  = \new_[95221]_  & \new_[95218]_ ;
  assign \new_[95223]_  = \new_[95222]_  & \new_[95215]_ ;
  assign \new_[95226]_  = ~A265 & A203;
  assign \new_[95229]_  = ~A267 & A266;
  assign \new_[95230]_  = \new_[95229]_  & \new_[95226]_ ;
  assign \new_[95233]_  = ~A269 & ~A268;
  assign \new_[95236]_  = A299 & A298;
  assign \new_[95237]_  = \new_[95236]_  & \new_[95233]_ ;
  assign \new_[95238]_  = \new_[95237]_  & \new_[95230]_ ;
  assign \new_[95241]_  = ~A169 & A170;
  assign \new_[95244]_  = A167 & ~A168;
  assign \new_[95245]_  = \new_[95244]_  & \new_[95241]_ ;
  assign \new_[95248]_  = A199 & ~A166;
  assign \new_[95251]_  = A201 & ~A200;
  assign \new_[95252]_  = \new_[95251]_  & \new_[95248]_ ;
  assign \new_[95253]_  = \new_[95252]_  & \new_[95245]_ ;
  assign \new_[95256]_  = ~A265 & A203;
  assign \new_[95259]_  = ~A267 & A266;
  assign \new_[95260]_  = \new_[95259]_  & \new_[95256]_ ;
  assign \new_[95263]_  = ~A269 & ~A268;
  assign \new_[95266]_  = ~A299 & ~A298;
  assign \new_[95267]_  = \new_[95266]_  & \new_[95263]_ ;
  assign \new_[95268]_  = \new_[95267]_  & \new_[95260]_ ;
  assign \new_[95271]_  = ~A169 & A170;
  assign \new_[95274]_  = A167 & ~A168;
  assign \new_[95275]_  = \new_[95274]_  & \new_[95271]_ ;
  assign \new_[95278]_  = A199 & ~A166;
  assign \new_[95281]_  = A201 & ~A200;
  assign \new_[95282]_  = \new_[95281]_  & \new_[95278]_ ;
  assign \new_[95283]_  = \new_[95282]_  & \new_[95275]_ ;
  assign \new_[95286]_  = A265 & A203;
  assign \new_[95289]_  = A267 & ~A266;
  assign \new_[95290]_  = \new_[95289]_  & \new_[95286]_ ;
  assign \new_[95293]_  = A300 & A268;
  assign \new_[95296]_  = ~A302 & ~A301;
  assign \new_[95297]_  = \new_[95296]_  & \new_[95293]_ ;
  assign \new_[95298]_  = \new_[95297]_  & \new_[95290]_ ;
  assign \new_[95301]_  = ~A169 & A170;
  assign \new_[95304]_  = A167 & ~A168;
  assign \new_[95305]_  = \new_[95304]_  & \new_[95301]_ ;
  assign \new_[95308]_  = A199 & ~A166;
  assign \new_[95311]_  = A201 & ~A200;
  assign \new_[95312]_  = \new_[95311]_  & \new_[95308]_ ;
  assign \new_[95313]_  = \new_[95312]_  & \new_[95305]_ ;
  assign \new_[95316]_  = A265 & A203;
  assign \new_[95319]_  = A267 & ~A266;
  assign \new_[95320]_  = \new_[95319]_  & \new_[95316]_ ;
  assign \new_[95323]_  = A300 & A269;
  assign \new_[95326]_  = ~A302 & ~A301;
  assign \new_[95327]_  = \new_[95326]_  & \new_[95323]_ ;
  assign \new_[95328]_  = \new_[95327]_  & \new_[95320]_ ;
  assign \new_[95331]_  = ~A169 & A170;
  assign \new_[95334]_  = A167 & ~A168;
  assign \new_[95335]_  = \new_[95334]_  & \new_[95331]_ ;
  assign \new_[95338]_  = A199 & ~A166;
  assign \new_[95341]_  = A201 & ~A200;
  assign \new_[95342]_  = \new_[95341]_  & \new_[95338]_ ;
  assign \new_[95343]_  = \new_[95342]_  & \new_[95335]_ ;
  assign \new_[95346]_  = A265 & A203;
  assign \new_[95349]_  = ~A267 & ~A266;
  assign \new_[95350]_  = \new_[95349]_  & \new_[95346]_ ;
  assign \new_[95353]_  = ~A269 & ~A268;
  assign \new_[95356]_  = A301 & ~A300;
  assign \new_[95357]_  = \new_[95356]_  & \new_[95353]_ ;
  assign \new_[95358]_  = \new_[95357]_  & \new_[95350]_ ;
  assign \new_[95361]_  = ~A169 & A170;
  assign \new_[95364]_  = A167 & ~A168;
  assign \new_[95365]_  = \new_[95364]_  & \new_[95361]_ ;
  assign \new_[95368]_  = A199 & ~A166;
  assign \new_[95371]_  = A201 & ~A200;
  assign \new_[95372]_  = \new_[95371]_  & \new_[95368]_ ;
  assign \new_[95373]_  = \new_[95372]_  & \new_[95365]_ ;
  assign \new_[95376]_  = A265 & A203;
  assign \new_[95379]_  = ~A267 & ~A266;
  assign \new_[95380]_  = \new_[95379]_  & \new_[95376]_ ;
  assign \new_[95383]_  = ~A269 & ~A268;
  assign \new_[95386]_  = A302 & ~A300;
  assign \new_[95387]_  = \new_[95386]_  & \new_[95383]_ ;
  assign \new_[95388]_  = \new_[95387]_  & \new_[95380]_ ;
  assign \new_[95391]_  = ~A169 & A170;
  assign \new_[95394]_  = A167 & ~A168;
  assign \new_[95395]_  = \new_[95394]_  & \new_[95391]_ ;
  assign \new_[95398]_  = A199 & ~A166;
  assign \new_[95401]_  = A201 & ~A200;
  assign \new_[95402]_  = \new_[95401]_  & \new_[95398]_ ;
  assign \new_[95403]_  = \new_[95402]_  & \new_[95395]_ ;
  assign \new_[95406]_  = A265 & A203;
  assign \new_[95409]_  = ~A267 & ~A266;
  assign \new_[95410]_  = \new_[95409]_  & \new_[95406]_ ;
  assign \new_[95413]_  = ~A269 & ~A268;
  assign \new_[95416]_  = A299 & A298;
  assign \new_[95417]_  = \new_[95416]_  & \new_[95413]_ ;
  assign \new_[95418]_  = \new_[95417]_  & \new_[95410]_ ;
  assign \new_[95421]_  = ~A169 & A170;
  assign \new_[95424]_  = A167 & ~A168;
  assign \new_[95425]_  = \new_[95424]_  & \new_[95421]_ ;
  assign \new_[95428]_  = A199 & ~A166;
  assign \new_[95431]_  = A201 & ~A200;
  assign \new_[95432]_  = \new_[95431]_  & \new_[95428]_ ;
  assign \new_[95433]_  = \new_[95432]_  & \new_[95425]_ ;
  assign \new_[95436]_  = A265 & A203;
  assign \new_[95439]_  = ~A267 & ~A266;
  assign \new_[95440]_  = \new_[95439]_  & \new_[95436]_ ;
  assign \new_[95443]_  = ~A269 & ~A268;
  assign \new_[95446]_  = ~A299 & ~A298;
  assign \new_[95447]_  = \new_[95446]_  & \new_[95443]_ ;
  assign \new_[95448]_  = \new_[95447]_  & \new_[95440]_ ;
  assign \new_[95451]_  = ~A169 & A170;
  assign \new_[95454]_  = A167 & ~A168;
  assign \new_[95455]_  = \new_[95454]_  & \new_[95451]_ ;
  assign \new_[95458]_  = A199 & ~A166;
  assign \new_[95461]_  = ~A201 & ~A200;
  assign \new_[95462]_  = \new_[95461]_  & \new_[95458]_ ;
  assign \new_[95463]_  = \new_[95462]_  & \new_[95455]_ ;
  assign \new_[95466]_  = ~A203 & ~A202;
  assign \new_[95469]_  = A266 & ~A265;
  assign \new_[95470]_  = \new_[95469]_  & \new_[95466]_ ;
  assign \new_[95473]_  = A268 & A267;
  assign \new_[95476]_  = A301 & ~A300;
  assign \new_[95477]_  = \new_[95476]_  & \new_[95473]_ ;
  assign \new_[95478]_  = \new_[95477]_  & \new_[95470]_ ;
  assign \new_[95481]_  = ~A169 & A170;
  assign \new_[95484]_  = A167 & ~A168;
  assign \new_[95485]_  = \new_[95484]_  & \new_[95481]_ ;
  assign \new_[95488]_  = A199 & ~A166;
  assign \new_[95491]_  = ~A201 & ~A200;
  assign \new_[95492]_  = \new_[95491]_  & \new_[95488]_ ;
  assign \new_[95493]_  = \new_[95492]_  & \new_[95485]_ ;
  assign \new_[95496]_  = ~A203 & ~A202;
  assign \new_[95499]_  = A266 & ~A265;
  assign \new_[95500]_  = \new_[95499]_  & \new_[95496]_ ;
  assign \new_[95503]_  = A268 & A267;
  assign \new_[95506]_  = A302 & ~A300;
  assign \new_[95507]_  = \new_[95506]_  & \new_[95503]_ ;
  assign \new_[95508]_  = \new_[95507]_  & \new_[95500]_ ;
  assign \new_[95511]_  = ~A169 & A170;
  assign \new_[95514]_  = A167 & ~A168;
  assign \new_[95515]_  = \new_[95514]_  & \new_[95511]_ ;
  assign \new_[95518]_  = A199 & ~A166;
  assign \new_[95521]_  = ~A201 & ~A200;
  assign \new_[95522]_  = \new_[95521]_  & \new_[95518]_ ;
  assign \new_[95523]_  = \new_[95522]_  & \new_[95515]_ ;
  assign \new_[95526]_  = ~A203 & ~A202;
  assign \new_[95529]_  = A266 & ~A265;
  assign \new_[95530]_  = \new_[95529]_  & \new_[95526]_ ;
  assign \new_[95533]_  = A268 & A267;
  assign \new_[95536]_  = A299 & A298;
  assign \new_[95537]_  = \new_[95536]_  & \new_[95533]_ ;
  assign \new_[95538]_  = \new_[95537]_  & \new_[95530]_ ;
  assign \new_[95541]_  = ~A169 & A170;
  assign \new_[95544]_  = A167 & ~A168;
  assign \new_[95545]_  = \new_[95544]_  & \new_[95541]_ ;
  assign \new_[95548]_  = A199 & ~A166;
  assign \new_[95551]_  = ~A201 & ~A200;
  assign \new_[95552]_  = \new_[95551]_  & \new_[95548]_ ;
  assign \new_[95553]_  = \new_[95552]_  & \new_[95545]_ ;
  assign \new_[95556]_  = ~A203 & ~A202;
  assign \new_[95559]_  = A266 & ~A265;
  assign \new_[95560]_  = \new_[95559]_  & \new_[95556]_ ;
  assign \new_[95563]_  = A268 & A267;
  assign \new_[95566]_  = ~A299 & ~A298;
  assign \new_[95567]_  = \new_[95566]_  & \new_[95563]_ ;
  assign \new_[95568]_  = \new_[95567]_  & \new_[95560]_ ;
  assign \new_[95571]_  = ~A169 & A170;
  assign \new_[95574]_  = A167 & ~A168;
  assign \new_[95575]_  = \new_[95574]_  & \new_[95571]_ ;
  assign \new_[95578]_  = A199 & ~A166;
  assign \new_[95581]_  = ~A201 & ~A200;
  assign \new_[95582]_  = \new_[95581]_  & \new_[95578]_ ;
  assign \new_[95583]_  = \new_[95582]_  & \new_[95575]_ ;
  assign \new_[95586]_  = ~A203 & ~A202;
  assign \new_[95589]_  = A266 & ~A265;
  assign \new_[95590]_  = \new_[95589]_  & \new_[95586]_ ;
  assign \new_[95593]_  = A269 & A267;
  assign \new_[95596]_  = A301 & ~A300;
  assign \new_[95597]_  = \new_[95596]_  & \new_[95593]_ ;
  assign \new_[95598]_  = \new_[95597]_  & \new_[95590]_ ;
  assign \new_[95601]_  = ~A169 & A170;
  assign \new_[95604]_  = A167 & ~A168;
  assign \new_[95605]_  = \new_[95604]_  & \new_[95601]_ ;
  assign \new_[95608]_  = A199 & ~A166;
  assign \new_[95611]_  = ~A201 & ~A200;
  assign \new_[95612]_  = \new_[95611]_  & \new_[95608]_ ;
  assign \new_[95613]_  = \new_[95612]_  & \new_[95605]_ ;
  assign \new_[95616]_  = ~A203 & ~A202;
  assign \new_[95619]_  = A266 & ~A265;
  assign \new_[95620]_  = \new_[95619]_  & \new_[95616]_ ;
  assign \new_[95623]_  = A269 & A267;
  assign \new_[95626]_  = A302 & ~A300;
  assign \new_[95627]_  = \new_[95626]_  & \new_[95623]_ ;
  assign \new_[95628]_  = \new_[95627]_  & \new_[95620]_ ;
  assign \new_[95631]_  = ~A169 & A170;
  assign \new_[95634]_  = A167 & ~A168;
  assign \new_[95635]_  = \new_[95634]_  & \new_[95631]_ ;
  assign \new_[95638]_  = A199 & ~A166;
  assign \new_[95641]_  = ~A201 & ~A200;
  assign \new_[95642]_  = \new_[95641]_  & \new_[95638]_ ;
  assign \new_[95643]_  = \new_[95642]_  & \new_[95635]_ ;
  assign \new_[95646]_  = ~A203 & ~A202;
  assign \new_[95649]_  = A266 & ~A265;
  assign \new_[95650]_  = \new_[95649]_  & \new_[95646]_ ;
  assign \new_[95653]_  = A269 & A267;
  assign \new_[95656]_  = A299 & A298;
  assign \new_[95657]_  = \new_[95656]_  & \new_[95653]_ ;
  assign \new_[95658]_  = \new_[95657]_  & \new_[95650]_ ;
  assign \new_[95661]_  = ~A169 & A170;
  assign \new_[95664]_  = A167 & ~A168;
  assign \new_[95665]_  = \new_[95664]_  & \new_[95661]_ ;
  assign \new_[95668]_  = A199 & ~A166;
  assign \new_[95671]_  = ~A201 & ~A200;
  assign \new_[95672]_  = \new_[95671]_  & \new_[95668]_ ;
  assign \new_[95673]_  = \new_[95672]_  & \new_[95665]_ ;
  assign \new_[95676]_  = ~A203 & ~A202;
  assign \new_[95679]_  = A266 & ~A265;
  assign \new_[95680]_  = \new_[95679]_  & \new_[95676]_ ;
  assign \new_[95683]_  = A269 & A267;
  assign \new_[95686]_  = ~A299 & ~A298;
  assign \new_[95687]_  = \new_[95686]_  & \new_[95683]_ ;
  assign \new_[95688]_  = \new_[95687]_  & \new_[95680]_ ;
  assign \new_[95691]_  = ~A169 & A170;
  assign \new_[95694]_  = A167 & ~A168;
  assign \new_[95695]_  = \new_[95694]_  & \new_[95691]_ ;
  assign \new_[95698]_  = A199 & ~A166;
  assign \new_[95701]_  = ~A201 & ~A200;
  assign \new_[95702]_  = \new_[95701]_  & \new_[95698]_ ;
  assign \new_[95703]_  = \new_[95702]_  & \new_[95695]_ ;
  assign \new_[95706]_  = ~A203 & ~A202;
  assign \new_[95709]_  = ~A266 & A265;
  assign \new_[95710]_  = \new_[95709]_  & \new_[95706]_ ;
  assign \new_[95713]_  = A268 & A267;
  assign \new_[95716]_  = A301 & ~A300;
  assign \new_[95717]_  = \new_[95716]_  & \new_[95713]_ ;
  assign \new_[95718]_  = \new_[95717]_  & \new_[95710]_ ;
  assign \new_[95721]_  = ~A169 & A170;
  assign \new_[95724]_  = A167 & ~A168;
  assign \new_[95725]_  = \new_[95724]_  & \new_[95721]_ ;
  assign \new_[95728]_  = A199 & ~A166;
  assign \new_[95731]_  = ~A201 & ~A200;
  assign \new_[95732]_  = \new_[95731]_  & \new_[95728]_ ;
  assign \new_[95733]_  = \new_[95732]_  & \new_[95725]_ ;
  assign \new_[95736]_  = ~A203 & ~A202;
  assign \new_[95739]_  = ~A266 & A265;
  assign \new_[95740]_  = \new_[95739]_  & \new_[95736]_ ;
  assign \new_[95743]_  = A268 & A267;
  assign \new_[95746]_  = A302 & ~A300;
  assign \new_[95747]_  = \new_[95746]_  & \new_[95743]_ ;
  assign \new_[95748]_  = \new_[95747]_  & \new_[95740]_ ;
  assign \new_[95751]_  = ~A169 & A170;
  assign \new_[95754]_  = A167 & ~A168;
  assign \new_[95755]_  = \new_[95754]_  & \new_[95751]_ ;
  assign \new_[95758]_  = A199 & ~A166;
  assign \new_[95761]_  = ~A201 & ~A200;
  assign \new_[95762]_  = \new_[95761]_  & \new_[95758]_ ;
  assign \new_[95763]_  = \new_[95762]_  & \new_[95755]_ ;
  assign \new_[95766]_  = ~A203 & ~A202;
  assign \new_[95769]_  = ~A266 & A265;
  assign \new_[95770]_  = \new_[95769]_  & \new_[95766]_ ;
  assign \new_[95773]_  = A268 & A267;
  assign \new_[95776]_  = A299 & A298;
  assign \new_[95777]_  = \new_[95776]_  & \new_[95773]_ ;
  assign \new_[95778]_  = \new_[95777]_  & \new_[95770]_ ;
  assign \new_[95781]_  = ~A169 & A170;
  assign \new_[95784]_  = A167 & ~A168;
  assign \new_[95785]_  = \new_[95784]_  & \new_[95781]_ ;
  assign \new_[95788]_  = A199 & ~A166;
  assign \new_[95791]_  = ~A201 & ~A200;
  assign \new_[95792]_  = \new_[95791]_  & \new_[95788]_ ;
  assign \new_[95793]_  = \new_[95792]_  & \new_[95785]_ ;
  assign \new_[95796]_  = ~A203 & ~A202;
  assign \new_[95799]_  = ~A266 & A265;
  assign \new_[95800]_  = \new_[95799]_  & \new_[95796]_ ;
  assign \new_[95803]_  = A268 & A267;
  assign \new_[95806]_  = ~A299 & ~A298;
  assign \new_[95807]_  = \new_[95806]_  & \new_[95803]_ ;
  assign \new_[95808]_  = \new_[95807]_  & \new_[95800]_ ;
  assign \new_[95811]_  = ~A169 & A170;
  assign \new_[95814]_  = A167 & ~A168;
  assign \new_[95815]_  = \new_[95814]_  & \new_[95811]_ ;
  assign \new_[95818]_  = A199 & ~A166;
  assign \new_[95821]_  = ~A201 & ~A200;
  assign \new_[95822]_  = \new_[95821]_  & \new_[95818]_ ;
  assign \new_[95823]_  = \new_[95822]_  & \new_[95815]_ ;
  assign \new_[95826]_  = ~A203 & ~A202;
  assign \new_[95829]_  = ~A266 & A265;
  assign \new_[95830]_  = \new_[95829]_  & \new_[95826]_ ;
  assign \new_[95833]_  = A269 & A267;
  assign \new_[95836]_  = A301 & ~A300;
  assign \new_[95837]_  = \new_[95836]_  & \new_[95833]_ ;
  assign \new_[95838]_  = \new_[95837]_  & \new_[95830]_ ;
  assign \new_[95841]_  = ~A169 & A170;
  assign \new_[95844]_  = A167 & ~A168;
  assign \new_[95845]_  = \new_[95844]_  & \new_[95841]_ ;
  assign \new_[95848]_  = A199 & ~A166;
  assign \new_[95851]_  = ~A201 & ~A200;
  assign \new_[95852]_  = \new_[95851]_  & \new_[95848]_ ;
  assign \new_[95853]_  = \new_[95852]_  & \new_[95845]_ ;
  assign \new_[95856]_  = ~A203 & ~A202;
  assign \new_[95859]_  = ~A266 & A265;
  assign \new_[95860]_  = \new_[95859]_  & \new_[95856]_ ;
  assign \new_[95863]_  = A269 & A267;
  assign \new_[95866]_  = A302 & ~A300;
  assign \new_[95867]_  = \new_[95866]_  & \new_[95863]_ ;
  assign \new_[95868]_  = \new_[95867]_  & \new_[95860]_ ;
  assign \new_[95871]_  = ~A169 & A170;
  assign \new_[95874]_  = A167 & ~A168;
  assign \new_[95875]_  = \new_[95874]_  & \new_[95871]_ ;
  assign \new_[95878]_  = A199 & ~A166;
  assign \new_[95881]_  = ~A201 & ~A200;
  assign \new_[95882]_  = \new_[95881]_  & \new_[95878]_ ;
  assign \new_[95883]_  = \new_[95882]_  & \new_[95875]_ ;
  assign \new_[95886]_  = ~A203 & ~A202;
  assign \new_[95889]_  = ~A266 & A265;
  assign \new_[95890]_  = \new_[95889]_  & \new_[95886]_ ;
  assign \new_[95893]_  = A269 & A267;
  assign \new_[95896]_  = A299 & A298;
  assign \new_[95897]_  = \new_[95896]_  & \new_[95893]_ ;
  assign \new_[95898]_  = \new_[95897]_  & \new_[95890]_ ;
  assign \new_[95901]_  = ~A169 & A170;
  assign \new_[95904]_  = A167 & ~A168;
  assign \new_[95905]_  = \new_[95904]_  & \new_[95901]_ ;
  assign \new_[95908]_  = A199 & ~A166;
  assign \new_[95911]_  = ~A201 & ~A200;
  assign \new_[95912]_  = \new_[95911]_  & \new_[95908]_ ;
  assign \new_[95913]_  = \new_[95912]_  & \new_[95905]_ ;
  assign \new_[95916]_  = ~A203 & ~A202;
  assign \new_[95919]_  = ~A266 & A265;
  assign \new_[95920]_  = \new_[95919]_  & \new_[95916]_ ;
  assign \new_[95923]_  = A269 & A267;
  assign \new_[95926]_  = ~A299 & ~A298;
  assign \new_[95927]_  = \new_[95926]_  & \new_[95923]_ ;
  assign \new_[95928]_  = \new_[95927]_  & \new_[95920]_ ;
  assign \new_[95931]_  = ~A169 & A170;
  assign \new_[95934]_  = ~A167 & ~A168;
  assign \new_[95935]_  = \new_[95934]_  & \new_[95931]_ ;
  assign \new_[95938]_  = A201 & A166;
  assign \new_[95941]_  = ~A203 & ~A202;
  assign \new_[95942]_  = \new_[95941]_  & \new_[95938]_ ;
  assign \new_[95943]_  = \new_[95942]_  & \new_[95935]_ ;
  assign \new_[95946]_  = ~A268 & A267;
  assign \new_[95949]_  = A298 & ~A269;
  assign \new_[95950]_  = \new_[95949]_  & \new_[95946]_ ;
  assign \new_[95953]_  = ~A300 & ~A299;
  assign \new_[95956]_  = ~A302 & ~A301;
  assign \new_[95957]_  = \new_[95956]_  & \new_[95953]_ ;
  assign \new_[95958]_  = \new_[95957]_  & \new_[95950]_ ;
  assign \new_[95961]_  = ~A169 & A170;
  assign \new_[95964]_  = ~A167 & ~A168;
  assign \new_[95965]_  = \new_[95964]_  & \new_[95961]_ ;
  assign \new_[95968]_  = A201 & A166;
  assign \new_[95971]_  = ~A203 & ~A202;
  assign \new_[95972]_  = \new_[95971]_  & \new_[95968]_ ;
  assign \new_[95973]_  = \new_[95972]_  & \new_[95965]_ ;
  assign \new_[95976]_  = ~A268 & A267;
  assign \new_[95979]_  = ~A298 & ~A269;
  assign \new_[95980]_  = \new_[95979]_  & \new_[95976]_ ;
  assign \new_[95983]_  = ~A300 & A299;
  assign \new_[95986]_  = ~A302 & ~A301;
  assign \new_[95987]_  = \new_[95986]_  & \new_[95983]_ ;
  assign \new_[95988]_  = \new_[95987]_  & \new_[95980]_ ;
  assign \new_[95991]_  = ~A169 & A170;
  assign \new_[95994]_  = ~A167 & ~A168;
  assign \new_[95995]_  = \new_[95994]_  & \new_[95991]_ ;
  assign \new_[95998]_  = ~A199 & A166;
  assign \new_[96001]_  = A201 & A200;
  assign \new_[96002]_  = \new_[96001]_  & \new_[95998]_ ;
  assign \new_[96003]_  = \new_[96002]_  & \new_[95995]_ ;
  assign \new_[96006]_  = ~A265 & A202;
  assign \new_[96009]_  = A267 & A266;
  assign \new_[96010]_  = \new_[96009]_  & \new_[96006]_ ;
  assign \new_[96013]_  = A300 & A268;
  assign \new_[96016]_  = ~A302 & ~A301;
  assign \new_[96017]_  = \new_[96016]_  & \new_[96013]_ ;
  assign \new_[96018]_  = \new_[96017]_  & \new_[96010]_ ;
  assign \new_[96021]_  = ~A169 & A170;
  assign \new_[96024]_  = ~A167 & ~A168;
  assign \new_[96025]_  = \new_[96024]_  & \new_[96021]_ ;
  assign \new_[96028]_  = ~A199 & A166;
  assign \new_[96031]_  = A201 & A200;
  assign \new_[96032]_  = \new_[96031]_  & \new_[96028]_ ;
  assign \new_[96033]_  = \new_[96032]_  & \new_[96025]_ ;
  assign \new_[96036]_  = ~A265 & A202;
  assign \new_[96039]_  = A267 & A266;
  assign \new_[96040]_  = \new_[96039]_  & \new_[96036]_ ;
  assign \new_[96043]_  = A300 & A269;
  assign \new_[96046]_  = ~A302 & ~A301;
  assign \new_[96047]_  = \new_[96046]_  & \new_[96043]_ ;
  assign \new_[96048]_  = \new_[96047]_  & \new_[96040]_ ;
  assign \new_[96051]_  = ~A169 & A170;
  assign \new_[96054]_  = ~A167 & ~A168;
  assign \new_[96055]_  = \new_[96054]_  & \new_[96051]_ ;
  assign \new_[96058]_  = ~A199 & A166;
  assign \new_[96061]_  = A201 & A200;
  assign \new_[96062]_  = \new_[96061]_  & \new_[96058]_ ;
  assign \new_[96063]_  = \new_[96062]_  & \new_[96055]_ ;
  assign \new_[96066]_  = ~A265 & A202;
  assign \new_[96069]_  = ~A267 & A266;
  assign \new_[96070]_  = \new_[96069]_  & \new_[96066]_ ;
  assign \new_[96073]_  = ~A269 & ~A268;
  assign \new_[96076]_  = A301 & ~A300;
  assign \new_[96077]_  = \new_[96076]_  & \new_[96073]_ ;
  assign \new_[96078]_  = \new_[96077]_  & \new_[96070]_ ;
  assign \new_[96081]_  = ~A169 & A170;
  assign \new_[96084]_  = ~A167 & ~A168;
  assign \new_[96085]_  = \new_[96084]_  & \new_[96081]_ ;
  assign \new_[96088]_  = ~A199 & A166;
  assign \new_[96091]_  = A201 & A200;
  assign \new_[96092]_  = \new_[96091]_  & \new_[96088]_ ;
  assign \new_[96093]_  = \new_[96092]_  & \new_[96085]_ ;
  assign \new_[96096]_  = ~A265 & A202;
  assign \new_[96099]_  = ~A267 & A266;
  assign \new_[96100]_  = \new_[96099]_  & \new_[96096]_ ;
  assign \new_[96103]_  = ~A269 & ~A268;
  assign \new_[96106]_  = A302 & ~A300;
  assign \new_[96107]_  = \new_[96106]_  & \new_[96103]_ ;
  assign \new_[96108]_  = \new_[96107]_  & \new_[96100]_ ;
  assign \new_[96111]_  = ~A169 & A170;
  assign \new_[96114]_  = ~A167 & ~A168;
  assign \new_[96115]_  = \new_[96114]_  & \new_[96111]_ ;
  assign \new_[96118]_  = ~A199 & A166;
  assign \new_[96121]_  = A201 & A200;
  assign \new_[96122]_  = \new_[96121]_  & \new_[96118]_ ;
  assign \new_[96123]_  = \new_[96122]_  & \new_[96115]_ ;
  assign \new_[96126]_  = ~A265 & A202;
  assign \new_[96129]_  = ~A267 & A266;
  assign \new_[96130]_  = \new_[96129]_  & \new_[96126]_ ;
  assign \new_[96133]_  = ~A269 & ~A268;
  assign \new_[96136]_  = A299 & A298;
  assign \new_[96137]_  = \new_[96136]_  & \new_[96133]_ ;
  assign \new_[96138]_  = \new_[96137]_  & \new_[96130]_ ;
  assign \new_[96141]_  = ~A169 & A170;
  assign \new_[96144]_  = ~A167 & ~A168;
  assign \new_[96145]_  = \new_[96144]_  & \new_[96141]_ ;
  assign \new_[96148]_  = ~A199 & A166;
  assign \new_[96151]_  = A201 & A200;
  assign \new_[96152]_  = \new_[96151]_  & \new_[96148]_ ;
  assign \new_[96153]_  = \new_[96152]_  & \new_[96145]_ ;
  assign \new_[96156]_  = ~A265 & A202;
  assign \new_[96159]_  = ~A267 & A266;
  assign \new_[96160]_  = \new_[96159]_  & \new_[96156]_ ;
  assign \new_[96163]_  = ~A269 & ~A268;
  assign \new_[96166]_  = ~A299 & ~A298;
  assign \new_[96167]_  = \new_[96166]_  & \new_[96163]_ ;
  assign \new_[96168]_  = \new_[96167]_  & \new_[96160]_ ;
  assign \new_[96171]_  = ~A169 & A170;
  assign \new_[96174]_  = ~A167 & ~A168;
  assign \new_[96175]_  = \new_[96174]_  & \new_[96171]_ ;
  assign \new_[96178]_  = ~A199 & A166;
  assign \new_[96181]_  = A201 & A200;
  assign \new_[96182]_  = \new_[96181]_  & \new_[96178]_ ;
  assign \new_[96183]_  = \new_[96182]_  & \new_[96175]_ ;
  assign \new_[96186]_  = A265 & A202;
  assign \new_[96189]_  = A267 & ~A266;
  assign \new_[96190]_  = \new_[96189]_  & \new_[96186]_ ;
  assign \new_[96193]_  = A300 & A268;
  assign \new_[96196]_  = ~A302 & ~A301;
  assign \new_[96197]_  = \new_[96196]_  & \new_[96193]_ ;
  assign \new_[96198]_  = \new_[96197]_  & \new_[96190]_ ;
  assign \new_[96201]_  = ~A169 & A170;
  assign \new_[96204]_  = ~A167 & ~A168;
  assign \new_[96205]_  = \new_[96204]_  & \new_[96201]_ ;
  assign \new_[96208]_  = ~A199 & A166;
  assign \new_[96211]_  = A201 & A200;
  assign \new_[96212]_  = \new_[96211]_  & \new_[96208]_ ;
  assign \new_[96213]_  = \new_[96212]_  & \new_[96205]_ ;
  assign \new_[96216]_  = A265 & A202;
  assign \new_[96219]_  = A267 & ~A266;
  assign \new_[96220]_  = \new_[96219]_  & \new_[96216]_ ;
  assign \new_[96223]_  = A300 & A269;
  assign \new_[96226]_  = ~A302 & ~A301;
  assign \new_[96227]_  = \new_[96226]_  & \new_[96223]_ ;
  assign \new_[96228]_  = \new_[96227]_  & \new_[96220]_ ;
  assign \new_[96231]_  = ~A169 & A170;
  assign \new_[96234]_  = ~A167 & ~A168;
  assign \new_[96235]_  = \new_[96234]_  & \new_[96231]_ ;
  assign \new_[96238]_  = ~A199 & A166;
  assign \new_[96241]_  = A201 & A200;
  assign \new_[96242]_  = \new_[96241]_  & \new_[96238]_ ;
  assign \new_[96243]_  = \new_[96242]_  & \new_[96235]_ ;
  assign \new_[96246]_  = A265 & A202;
  assign \new_[96249]_  = ~A267 & ~A266;
  assign \new_[96250]_  = \new_[96249]_  & \new_[96246]_ ;
  assign \new_[96253]_  = ~A269 & ~A268;
  assign \new_[96256]_  = A301 & ~A300;
  assign \new_[96257]_  = \new_[96256]_  & \new_[96253]_ ;
  assign \new_[96258]_  = \new_[96257]_  & \new_[96250]_ ;
  assign \new_[96261]_  = ~A169 & A170;
  assign \new_[96264]_  = ~A167 & ~A168;
  assign \new_[96265]_  = \new_[96264]_  & \new_[96261]_ ;
  assign \new_[96268]_  = ~A199 & A166;
  assign \new_[96271]_  = A201 & A200;
  assign \new_[96272]_  = \new_[96271]_  & \new_[96268]_ ;
  assign \new_[96273]_  = \new_[96272]_  & \new_[96265]_ ;
  assign \new_[96276]_  = A265 & A202;
  assign \new_[96279]_  = ~A267 & ~A266;
  assign \new_[96280]_  = \new_[96279]_  & \new_[96276]_ ;
  assign \new_[96283]_  = ~A269 & ~A268;
  assign \new_[96286]_  = A302 & ~A300;
  assign \new_[96287]_  = \new_[96286]_  & \new_[96283]_ ;
  assign \new_[96288]_  = \new_[96287]_  & \new_[96280]_ ;
  assign \new_[96291]_  = ~A169 & A170;
  assign \new_[96294]_  = ~A167 & ~A168;
  assign \new_[96295]_  = \new_[96294]_  & \new_[96291]_ ;
  assign \new_[96298]_  = ~A199 & A166;
  assign \new_[96301]_  = A201 & A200;
  assign \new_[96302]_  = \new_[96301]_  & \new_[96298]_ ;
  assign \new_[96303]_  = \new_[96302]_  & \new_[96295]_ ;
  assign \new_[96306]_  = A265 & A202;
  assign \new_[96309]_  = ~A267 & ~A266;
  assign \new_[96310]_  = \new_[96309]_  & \new_[96306]_ ;
  assign \new_[96313]_  = ~A269 & ~A268;
  assign \new_[96316]_  = A299 & A298;
  assign \new_[96317]_  = \new_[96316]_  & \new_[96313]_ ;
  assign \new_[96318]_  = \new_[96317]_  & \new_[96310]_ ;
  assign \new_[96321]_  = ~A169 & A170;
  assign \new_[96324]_  = ~A167 & ~A168;
  assign \new_[96325]_  = \new_[96324]_  & \new_[96321]_ ;
  assign \new_[96328]_  = ~A199 & A166;
  assign \new_[96331]_  = A201 & A200;
  assign \new_[96332]_  = \new_[96331]_  & \new_[96328]_ ;
  assign \new_[96333]_  = \new_[96332]_  & \new_[96325]_ ;
  assign \new_[96336]_  = A265 & A202;
  assign \new_[96339]_  = ~A267 & ~A266;
  assign \new_[96340]_  = \new_[96339]_  & \new_[96336]_ ;
  assign \new_[96343]_  = ~A269 & ~A268;
  assign \new_[96346]_  = ~A299 & ~A298;
  assign \new_[96347]_  = \new_[96346]_  & \new_[96343]_ ;
  assign \new_[96348]_  = \new_[96347]_  & \new_[96340]_ ;
  assign \new_[96351]_  = ~A169 & A170;
  assign \new_[96354]_  = ~A167 & ~A168;
  assign \new_[96355]_  = \new_[96354]_  & \new_[96351]_ ;
  assign \new_[96358]_  = ~A199 & A166;
  assign \new_[96361]_  = A201 & A200;
  assign \new_[96362]_  = \new_[96361]_  & \new_[96358]_ ;
  assign \new_[96363]_  = \new_[96362]_  & \new_[96355]_ ;
  assign \new_[96366]_  = ~A265 & A203;
  assign \new_[96369]_  = A267 & A266;
  assign \new_[96370]_  = \new_[96369]_  & \new_[96366]_ ;
  assign \new_[96373]_  = A300 & A268;
  assign \new_[96376]_  = ~A302 & ~A301;
  assign \new_[96377]_  = \new_[96376]_  & \new_[96373]_ ;
  assign \new_[96378]_  = \new_[96377]_  & \new_[96370]_ ;
  assign \new_[96381]_  = ~A169 & A170;
  assign \new_[96384]_  = ~A167 & ~A168;
  assign \new_[96385]_  = \new_[96384]_  & \new_[96381]_ ;
  assign \new_[96388]_  = ~A199 & A166;
  assign \new_[96391]_  = A201 & A200;
  assign \new_[96392]_  = \new_[96391]_  & \new_[96388]_ ;
  assign \new_[96393]_  = \new_[96392]_  & \new_[96385]_ ;
  assign \new_[96396]_  = ~A265 & A203;
  assign \new_[96399]_  = A267 & A266;
  assign \new_[96400]_  = \new_[96399]_  & \new_[96396]_ ;
  assign \new_[96403]_  = A300 & A269;
  assign \new_[96406]_  = ~A302 & ~A301;
  assign \new_[96407]_  = \new_[96406]_  & \new_[96403]_ ;
  assign \new_[96408]_  = \new_[96407]_  & \new_[96400]_ ;
  assign \new_[96411]_  = ~A169 & A170;
  assign \new_[96414]_  = ~A167 & ~A168;
  assign \new_[96415]_  = \new_[96414]_  & \new_[96411]_ ;
  assign \new_[96418]_  = ~A199 & A166;
  assign \new_[96421]_  = A201 & A200;
  assign \new_[96422]_  = \new_[96421]_  & \new_[96418]_ ;
  assign \new_[96423]_  = \new_[96422]_  & \new_[96415]_ ;
  assign \new_[96426]_  = ~A265 & A203;
  assign \new_[96429]_  = ~A267 & A266;
  assign \new_[96430]_  = \new_[96429]_  & \new_[96426]_ ;
  assign \new_[96433]_  = ~A269 & ~A268;
  assign \new_[96436]_  = A301 & ~A300;
  assign \new_[96437]_  = \new_[96436]_  & \new_[96433]_ ;
  assign \new_[96438]_  = \new_[96437]_  & \new_[96430]_ ;
  assign \new_[96441]_  = ~A169 & A170;
  assign \new_[96444]_  = ~A167 & ~A168;
  assign \new_[96445]_  = \new_[96444]_  & \new_[96441]_ ;
  assign \new_[96448]_  = ~A199 & A166;
  assign \new_[96451]_  = A201 & A200;
  assign \new_[96452]_  = \new_[96451]_  & \new_[96448]_ ;
  assign \new_[96453]_  = \new_[96452]_  & \new_[96445]_ ;
  assign \new_[96456]_  = ~A265 & A203;
  assign \new_[96459]_  = ~A267 & A266;
  assign \new_[96460]_  = \new_[96459]_  & \new_[96456]_ ;
  assign \new_[96463]_  = ~A269 & ~A268;
  assign \new_[96466]_  = A302 & ~A300;
  assign \new_[96467]_  = \new_[96466]_  & \new_[96463]_ ;
  assign \new_[96468]_  = \new_[96467]_  & \new_[96460]_ ;
  assign \new_[96471]_  = ~A169 & A170;
  assign \new_[96474]_  = ~A167 & ~A168;
  assign \new_[96475]_  = \new_[96474]_  & \new_[96471]_ ;
  assign \new_[96478]_  = ~A199 & A166;
  assign \new_[96481]_  = A201 & A200;
  assign \new_[96482]_  = \new_[96481]_  & \new_[96478]_ ;
  assign \new_[96483]_  = \new_[96482]_  & \new_[96475]_ ;
  assign \new_[96486]_  = ~A265 & A203;
  assign \new_[96489]_  = ~A267 & A266;
  assign \new_[96490]_  = \new_[96489]_  & \new_[96486]_ ;
  assign \new_[96493]_  = ~A269 & ~A268;
  assign \new_[96496]_  = A299 & A298;
  assign \new_[96497]_  = \new_[96496]_  & \new_[96493]_ ;
  assign \new_[96498]_  = \new_[96497]_  & \new_[96490]_ ;
  assign \new_[96501]_  = ~A169 & A170;
  assign \new_[96504]_  = ~A167 & ~A168;
  assign \new_[96505]_  = \new_[96504]_  & \new_[96501]_ ;
  assign \new_[96508]_  = ~A199 & A166;
  assign \new_[96511]_  = A201 & A200;
  assign \new_[96512]_  = \new_[96511]_  & \new_[96508]_ ;
  assign \new_[96513]_  = \new_[96512]_  & \new_[96505]_ ;
  assign \new_[96516]_  = ~A265 & A203;
  assign \new_[96519]_  = ~A267 & A266;
  assign \new_[96520]_  = \new_[96519]_  & \new_[96516]_ ;
  assign \new_[96523]_  = ~A269 & ~A268;
  assign \new_[96526]_  = ~A299 & ~A298;
  assign \new_[96527]_  = \new_[96526]_  & \new_[96523]_ ;
  assign \new_[96528]_  = \new_[96527]_  & \new_[96520]_ ;
  assign \new_[96531]_  = ~A169 & A170;
  assign \new_[96534]_  = ~A167 & ~A168;
  assign \new_[96535]_  = \new_[96534]_  & \new_[96531]_ ;
  assign \new_[96538]_  = ~A199 & A166;
  assign \new_[96541]_  = A201 & A200;
  assign \new_[96542]_  = \new_[96541]_  & \new_[96538]_ ;
  assign \new_[96543]_  = \new_[96542]_  & \new_[96535]_ ;
  assign \new_[96546]_  = A265 & A203;
  assign \new_[96549]_  = A267 & ~A266;
  assign \new_[96550]_  = \new_[96549]_  & \new_[96546]_ ;
  assign \new_[96553]_  = A300 & A268;
  assign \new_[96556]_  = ~A302 & ~A301;
  assign \new_[96557]_  = \new_[96556]_  & \new_[96553]_ ;
  assign \new_[96558]_  = \new_[96557]_  & \new_[96550]_ ;
  assign \new_[96561]_  = ~A169 & A170;
  assign \new_[96564]_  = ~A167 & ~A168;
  assign \new_[96565]_  = \new_[96564]_  & \new_[96561]_ ;
  assign \new_[96568]_  = ~A199 & A166;
  assign \new_[96571]_  = A201 & A200;
  assign \new_[96572]_  = \new_[96571]_  & \new_[96568]_ ;
  assign \new_[96573]_  = \new_[96572]_  & \new_[96565]_ ;
  assign \new_[96576]_  = A265 & A203;
  assign \new_[96579]_  = A267 & ~A266;
  assign \new_[96580]_  = \new_[96579]_  & \new_[96576]_ ;
  assign \new_[96583]_  = A300 & A269;
  assign \new_[96586]_  = ~A302 & ~A301;
  assign \new_[96587]_  = \new_[96586]_  & \new_[96583]_ ;
  assign \new_[96588]_  = \new_[96587]_  & \new_[96580]_ ;
  assign \new_[96591]_  = ~A169 & A170;
  assign \new_[96594]_  = ~A167 & ~A168;
  assign \new_[96595]_  = \new_[96594]_  & \new_[96591]_ ;
  assign \new_[96598]_  = ~A199 & A166;
  assign \new_[96601]_  = A201 & A200;
  assign \new_[96602]_  = \new_[96601]_  & \new_[96598]_ ;
  assign \new_[96603]_  = \new_[96602]_  & \new_[96595]_ ;
  assign \new_[96606]_  = A265 & A203;
  assign \new_[96609]_  = ~A267 & ~A266;
  assign \new_[96610]_  = \new_[96609]_  & \new_[96606]_ ;
  assign \new_[96613]_  = ~A269 & ~A268;
  assign \new_[96616]_  = A301 & ~A300;
  assign \new_[96617]_  = \new_[96616]_  & \new_[96613]_ ;
  assign \new_[96618]_  = \new_[96617]_  & \new_[96610]_ ;
  assign \new_[96621]_  = ~A169 & A170;
  assign \new_[96624]_  = ~A167 & ~A168;
  assign \new_[96625]_  = \new_[96624]_  & \new_[96621]_ ;
  assign \new_[96628]_  = ~A199 & A166;
  assign \new_[96631]_  = A201 & A200;
  assign \new_[96632]_  = \new_[96631]_  & \new_[96628]_ ;
  assign \new_[96633]_  = \new_[96632]_  & \new_[96625]_ ;
  assign \new_[96636]_  = A265 & A203;
  assign \new_[96639]_  = ~A267 & ~A266;
  assign \new_[96640]_  = \new_[96639]_  & \new_[96636]_ ;
  assign \new_[96643]_  = ~A269 & ~A268;
  assign \new_[96646]_  = A302 & ~A300;
  assign \new_[96647]_  = \new_[96646]_  & \new_[96643]_ ;
  assign \new_[96648]_  = \new_[96647]_  & \new_[96640]_ ;
  assign \new_[96651]_  = ~A169 & A170;
  assign \new_[96654]_  = ~A167 & ~A168;
  assign \new_[96655]_  = \new_[96654]_  & \new_[96651]_ ;
  assign \new_[96658]_  = ~A199 & A166;
  assign \new_[96661]_  = A201 & A200;
  assign \new_[96662]_  = \new_[96661]_  & \new_[96658]_ ;
  assign \new_[96663]_  = \new_[96662]_  & \new_[96655]_ ;
  assign \new_[96666]_  = A265 & A203;
  assign \new_[96669]_  = ~A267 & ~A266;
  assign \new_[96670]_  = \new_[96669]_  & \new_[96666]_ ;
  assign \new_[96673]_  = ~A269 & ~A268;
  assign \new_[96676]_  = A299 & A298;
  assign \new_[96677]_  = \new_[96676]_  & \new_[96673]_ ;
  assign \new_[96678]_  = \new_[96677]_  & \new_[96670]_ ;
  assign \new_[96681]_  = ~A169 & A170;
  assign \new_[96684]_  = ~A167 & ~A168;
  assign \new_[96685]_  = \new_[96684]_  & \new_[96681]_ ;
  assign \new_[96688]_  = ~A199 & A166;
  assign \new_[96691]_  = A201 & A200;
  assign \new_[96692]_  = \new_[96691]_  & \new_[96688]_ ;
  assign \new_[96693]_  = \new_[96692]_  & \new_[96685]_ ;
  assign \new_[96696]_  = A265 & A203;
  assign \new_[96699]_  = ~A267 & ~A266;
  assign \new_[96700]_  = \new_[96699]_  & \new_[96696]_ ;
  assign \new_[96703]_  = ~A269 & ~A268;
  assign \new_[96706]_  = ~A299 & ~A298;
  assign \new_[96707]_  = \new_[96706]_  & \new_[96703]_ ;
  assign \new_[96708]_  = \new_[96707]_  & \new_[96700]_ ;
  assign \new_[96711]_  = ~A169 & A170;
  assign \new_[96714]_  = ~A167 & ~A168;
  assign \new_[96715]_  = \new_[96714]_  & \new_[96711]_ ;
  assign \new_[96718]_  = ~A199 & A166;
  assign \new_[96721]_  = ~A201 & A200;
  assign \new_[96722]_  = \new_[96721]_  & \new_[96718]_ ;
  assign \new_[96723]_  = \new_[96722]_  & \new_[96715]_ ;
  assign \new_[96726]_  = ~A203 & ~A202;
  assign \new_[96729]_  = A266 & ~A265;
  assign \new_[96730]_  = \new_[96729]_  & \new_[96726]_ ;
  assign \new_[96733]_  = A268 & A267;
  assign \new_[96736]_  = A301 & ~A300;
  assign \new_[96737]_  = \new_[96736]_  & \new_[96733]_ ;
  assign \new_[96738]_  = \new_[96737]_  & \new_[96730]_ ;
  assign \new_[96741]_  = ~A169 & A170;
  assign \new_[96744]_  = ~A167 & ~A168;
  assign \new_[96745]_  = \new_[96744]_  & \new_[96741]_ ;
  assign \new_[96748]_  = ~A199 & A166;
  assign \new_[96751]_  = ~A201 & A200;
  assign \new_[96752]_  = \new_[96751]_  & \new_[96748]_ ;
  assign \new_[96753]_  = \new_[96752]_  & \new_[96745]_ ;
  assign \new_[96756]_  = ~A203 & ~A202;
  assign \new_[96759]_  = A266 & ~A265;
  assign \new_[96760]_  = \new_[96759]_  & \new_[96756]_ ;
  assign \new_[96763]_  = A268 & A267;
  assign \new_[96766]_  = A302 & ~A300;
  assign \new_[96767]_  = \new_[96766]_  & \new_[96763]_ ;
  assign \new_[96768]_  = \new_[96767]_  & \new_[96760]_ ;
  assign \new_[96771]_  = ~A169 & A170;
  assign \new_[96774]_  = ~A167 & ~A168;
  assign \new_[96775]_  = \new_[96774]_  & \new_[96771]_ ;
  assign \new_[96778]_  = ~A199 & A166;
  assign \new_[96781]_  = ~A201 & A200;
  assign \new_[96782]_  = \new_[96781]_  & \new_[96778]_ ;
  assign \new_[96783]_  = \new_[96782]_  & \new_[96775]_ ;
  assign \new_[96786]_  = ~A203 & ~A202;
  assign \new_[96789]_  = A266 & ~A265;
  assign \new_[96790]_  = \new_[96789]_  & \new_[96786]_ ;
  assign \new_[96793]_  = A268 & A267;
  assign \new_[96796]_  = A299 & A298;
  assign \new_[96797]_  = \new_[96796]_  & \new_[96793]_ ;
  assign \new_[96798]_  = \new_[96797]_  & \new_[96790]_ ;
  assign \new_[96801]_  = ~A169 & A170;
  assign \new_[96804]_  = ~A167 & ~A168;
  assign \new_[96805]_  = \new_[96804]_  & \new_[96801]_ ;
  assign \new_[96808]_  = ~A199 & A166;
  assign \new_[96811]_  = ~A201 & A200;
  assign \new_[96812]_  = \new_[96811]_  & \new_[96808]_ ;
  assign \new_[96813]_  = \new_[96812]_  & \new_[96805]_ ;
  assign \new_[96816]_  = ~A203 & ~A202;
  assign \new_[96819]_  = A266 & ~A265;
  assign \new_[96820]_  = \new_[96819]_  & \new_[96816]_ ;
  assign \new_[96823]_  = A268 & A267;
  assign \new_[96826]_  = ~A299 & ~A298;
  assign \new_[96827]_  = \new_[96826]_  & \new_[96823]_ ;
  assign \new_[96828]_  = \new_[96827]_  & \new_[96820]_ ;
  assign \new_[96831]_  = ~A169 & A170;
  assign \new_[96834]_  = ~A167 & ~A168;
  assign \new_[96835]_  = \new_[96834]_  & \new_[96831]_ ;
  assign \new_[96838]_  = ~A199 & A166;
  assign \new_[96841]_  = ~A201 & A200;
  assign \new_[96842]_  = \new_[96841]_  & \new_[96838]_ ;
  assign \new_[96843]_  = \new_[96842]_  & \new_[96835]_ ;
  assign \new_[96846]_  = ~A203 & ~A202;
  assign \new_[96849]_  = A266 & ~A265;
  assign \new_[96850]_  = \new_[96849]_  & \new_[96846]_ ;
  assign \new_[96853]_  = A269 & A267;
  assign \new_[96856]_  = A301 & ~A300;
  assign \new_[96857]_  = \new_[96856]_  & \new_[96853]_ ;
  assign \new_[96858]_  = \new_[96857]_  & \new_[96850]_ ;
  assign \new_[96861]_  = ~A169 & A170;
  assign \new_[96864]_  = ~A167 & ~A168;
  assign \new_[96865]_  = \new_[96864]_  & \new_[96861]_ ;
  assign \new_[96868]_  = ~A199 & A166;
  assign \new_[96871]_  = ~A201 & A200;
  assign \new_[96872]_  = \new_[96871]_  & \new_[96868]_ ;
  assign \new_[96873]_  = \new_[96872]_  & \new_[96865]_ ;
  assign \new_[96876]_  = ~A203 & ~A202;
  assign \new_[96879]_  = A266 & ~A265;
  assign \new_[96880]_  = \new_[96879]_  & \new_[96876]_ ;
  assign \new_[96883]_  = A269 & A267;
  assign \new_[96886]_  = A302 & ~A300;
  assign \new_[96887]_  = \new_[96886]_  & \new_[96883]_ ;
  assign \new_[96888]_  = \new_[96887]_  & \new_[96880]_ ;
  assign \new_[96891]_  = ~A169 & A170;
  assign \new_[96894]_  = ~A167 & ~A168;
  assign \new_[96895]_  = \new_[96894]_  & \new_[96891]_ ;
  assign \new_[96898]_  = ~A199 & A166;
  assign \new_[96901]_  = ~A201 & A200;
  assign \new_[96902]_  = \new_[96901]_  & \new_[96898]_ ;
  assign \new_[96903]_  = \new_[96902]_  & \new_[96895]_ ;
  assign \new_[96906]_  = ~A203 & ~A202;
  assign \new_[96909]_  = A266 & ~A265;
  assign \new_[96910]_  = \new_[96909]_  & \new_[96906]_ ;
  assign \new_[96913]_  = A269 & A267;
  assign \new_[96916]_  = A299 & A298;
  assign \new_[96917]_  = \new_[96916]_  & \new_[96913]_ ;
  assign \new_[96918]_  = \new_[96917]_  & \new_[96910]_ ;
  assign \new_[96921]_  = ~A169 & A170;
  assign \new_[96924]_  = ~A167 & ~A168;
  assign \new_[96925]_  = \new_[96924]_  & \new_[96921]_ ;
  assign \new_[96928]_  = ~A199 & A166;
  assign \new_[96931]_  = ~A201 & A200;
  assign \new_[96932]_  = \new_[96931]_  & \new_[96928]_ ;
  assign \new_[96933]_  = \new_[96932]_  & \new_[96925]_ ;
  assign \new_[96936]_  = ~A203 & ~A202;
  assign \new_[96939]_  = A266 & ~A265;
  assign \new_[96940]_  = \new_[96939]_  & \new_[96936]_ ;
  assign \new_[96943]_  = A269 & A267;
  assign \new_[96946]_  = ~A299 & ~A298;
  assign \new_[96947]_  = \new_[96946]_  & \new_[96943]_ ;
  assign \new_[96948]_  = \new_[96947]_  & \new_[96940]_ ;
  assign \new_[96951]_  = ~A169 & A170;
  assign \new_[96954]_  = ~A167 & ~A168;
  assign \new_[96955]_  = \new_[96954]_  & \new_[96951]_ ;
  assign \new_[96958]_  = ~A199 & A166;
  assign \new_[96961]_  = ~A201 & A200;
  assign \new_[96962]_  = \new_[96961]_  & \new_[96958]_ ;
  assign \new_[96963]_  = \new_[96962]_  & \new_[96955]_ ;
  assign \new_[96966]_  = ~A203 & ~A202;
  assign \new_[96969]_  = ~A266 & A265;
  assign \new_[96970]_  = \new_[96969]_  & \new_[96966]_ ;
  assign \new_[96973]_  = A268 & A267;
  assign \new_[96976]_  = A301 & ~A300;
  assign \new_[96977]_  = \new_[96976]_  & \new_[96973]_ ;
  assign \new_[96978]_  = \new_[96977]_  & \new_[96970]_ ;
  assign \new_[96981]_  = ~A169 & A170;
  assign \new_[96984]_  = ~A167 & ~A168;
  assign \new_[96985]_  = \new_[96984]_  & \new_[96981]_ ;
  assign \new_[96988]_  = ~A199 & A166;
  assign \new_[96991]_  = ~A201 & A200;
  assign \new_[96992]_  = \new_[96991]_  & \new_[96988]_ ;
  assign \new_[96993]_  = \new_[96992]_  & \new_[96985]_ ;
  assign \new_[96996]_  = ~A203 & ~A202;
  assign \new_[96999]_  = ~A266 & A265;
  assign \new_[97000]_  = \new_[96999]_  & \new_[96996]_ ;
  assign \new_[97003]_  = A268 & A267;
  assign \new_[97006]_  = A302 & ~A300;
  assign \new_[97007]_  = \new_[97006]_  & \new_[97003]_ ;
  assign \new_[97008]_  = \new_[97007]_  & \new_[97000]_ ;
  assign \new_[97011]_  = ~A169 & A170;
  assign \new_[97014]_  = ~A167 & ~A168;
  assign \new_[97015]_  = \new_[97014]_  & \new_[97011]_ ;
  assign \new_[97018]_  = ~A199 & A166;
  assign \new_[97021]_  = ~A201 & A200;
  assign \new_[97022]_  = \new_[97021]_  & \new_[97018]_ ;
  assign \new_[97023]_  = \new_[97022]_  & \new_[97015]_ ;
  assign \new_[97026]_  = ~A203 & ~A202;
  assign \new_[97029]_  = ~A266 & A265;
  assign \new_[97030]_  = \new_[97029]_  & \new_[97026]_ ;
  assign \new_[97033]_  = A268 & A267;
  assign \new_[97036]_  = A299 & A298;
  assign \new_[97037]_  = \new_[97036]_  & \new_[97033]_ ;
  assign \new_[97038]_  = \new_[97037]_  & \new_[97030]_ ;
  assign \new_[97041]_  = ~A169 & A170;
  assign \new_[97044]_  = ~A167 & ~A168;
  assign \new_[97045]_  = \new_[97044]_  & \new_[97041]_ ;
  assign \new_[97048]_  = ~A199 & A166;
  assign \new_[97051]_  = ~A201 & A200;
  assign \new_[97052]_  = \new_[97051]_  & \new_[97048]_ ;
  assign \new_[97053]_  = \new_[97052]_  & \new_[97045]_ ;
  assign \new_[97056]_  = ~A203 & ~A202;
  assign \new_[97059]_  = ~A266 & A265;
  assign \new_[97060]_  = \new_[97059]_  & \new_[97056]_ ;
  assign \new_[97063]_  = A268 & A267;
  assign \new_[97066]_  = ~A299 & ~A298;
  assign \new_[97067]_  = \new_[97066]_  & \new_[97063]_ ;
  assign \new_[97068]_  = \new_[97067]_  & \new_[97060]_ ;
  assign \new_[97071]_  = ~A169 & A170;
  assign \new_[97074]_  = ~A167 & ~A168;
  assign \new_[97075]_  = \new_[97074]_  & \new_[97071]_ ;
  assign \new_[97078]_  = ~A199 & A166;
  assign \new_[97081]_  = ~A201 & A200;
  assign \new_[97082]_  = \new_[97081]_  & \new_[97078]_ ;
  assign \new_[97083]_  = \new_[97082]_  & \new_[97075]_ ;
  assign \new_[97086]_  = ~A203 & ~A202;
  assign \new_[97089]_  = ~A266 & A265;
  assign \new_[97090]_  = \new_[97089]_  & \new_[97086]_ ;
  assign \new_[97093]_  = A269 & A267;
  assign \new_[97096]_  = A301 & ~A300;
  assign \new_[97097]_  = \new_[97096]_  & \new_[97093]_ ;
  assign \new_[97098]_  = \new_[97097]_  & \new_[97090]_ ;
  assign \new_[97101]_  = ~A169 & A170;
  assign \new_[97104]_  = ~A167 & ~A168;
  assign \new_[97105]_  = \new_[97104]_  & \new_[97101]_ ;
  assign \new_[97108]_  = ~A199 & A166;
  assign \new_[97111]_  = ~A201 & A200;
  assign \new_[97112]_  = \new_[97111]_  & \new_[97108]_ ;
  assign \new_[97113]_  = \new_[97112]_  & \new_[97105]_ ;
  assign \new_[97116]_  = ~A203 & ~A202;
  assign \new_[97119]_  = ~A266 & A265;
  assign \new_[97120]_  = \new_[97119]_  & \new_[97116]_ ;
  assign \new_[97123]_  = A269 & A267;
  assign \new_[97126]_  = A302 & ~A300;
  assign \new_[97127]_  = \new_[97126]_  & \new_[97123]_ ;
  assign \new_[97128]_  = \new_[97127]_  & \new_[97120]_ ;
  assign \new_[97131]_  = ~A169 & A170;
  assign \new_[97134]_  = ~A167 & ~A168;
  assign \new_[97135]_  = \new_[97134]_  & \new_[97131]_ ;
  assign \new_[97138]_  = ~A199 & A166;
  assign \new_[97141]_  = ~A201 & A200;
  assign \new_[97142]_  = \new_[97141]_  & \new_[97138]_ ;
  assign \new_[97143]_  = \new_[97142]_  & \new_[97135]_ ;
  assign \new_[97146]_  = ~A203 & ~A202;
  assign \new_[97149]_  = ~A266 & A265;
  assign \new_[97150]_  = \new_[97149]_  & \new_[97146]_ ;
  assign \new_[97153]_  = A269 & A267;
  assign \new_[97156]_  = A299 & A298;
  assign \new_[97157]_  = \new_[97156]_  & \new_[97153]_ ;
  assign \new_[97158]_  = \new_[97157]_  & \new_[97150]_ ;
  assign \new_[97161]_  = ~A169 & A170;
  assign \new_[97164]_  = ~A167 & ~A168;
  assign \new_[97165]_  = \new_[97164]_  & \new_[97161]_ ;
  assign \new_[97168]_  = ~A199 & A166;
  assign \new_[97171]_  = ~A201 & A200;
  assign \new_[97172]_  = \new_[97171]_  & \new_[97168]_ ;
  assign \new_[97173]_  = \new_[97172]_  & \new_[97165]_ ;
  assign \new_[97176]_  = ~A203 & ~A202;
  assign \new_[97179]_  = ~A266 & A265;
  assign \new_[97180]_  = \new_[97179]_  & \new_[97176]_ ;
  assign \new_[97183]_  = A269 & A267;
  assign \new_[97186]_  = ~A299 & ~A298;
  assign \new_[97187]_  = \new_[97186]_  & \new_[97183]_ ;
  assign \new_[97188]_  = \new_[97187]_  & \new_[97180]_ ;
  assign \new_[97191]_  = ~A169 & A170;
  assign \new_[97194]_  = ~A167 & ~A168;
  assign \new_[97195]_  = \new_[97194]_  & \new_[97191]_ ;
  assign \new_[97198]_  = A199 & A166;
  assign \new_[97201]_  = A201 & ~A200;
  assign \new_[97202]_  = \new_[97201]_  & \new_[97198]_ ;
  assign \new_[97203]_  = \new_[97202]_  & \new_[97195]_ ;
  assign \new_[97206]_  = ~A265 & A202;
  assign \new_[97209]_  = A267 & A266;
  assign \new_[97210]_  = \new_[97209]_  & \new_[97206]_ ;
  assign \new_[97213]_  = A300 & A268;
  assign \new_[97216]_  = ~A302 & ~A301;
  assign \new_[97217]_  = \new_[97216]_  & \new_[97213]_ ;
  assign \new_[97218]_  = \new_[97217]_  & \new_[97210]_ ;
  assign \new_[97221]_  = ~A169 & A170;
  assign \new_[97224]_  = ~A167 & ~A168;
  assign \new_[97225]_  = \new_[97224]_  & \new_[97221]_ ;
  assign \new_[97228]_  = A199 & A166;
  assign \new_[97231]_  = A201 & ~A200;
  assign \new_[97232]_  = \new_[97231]_  & \new_[97228]_ ;
  assign \new_[97233]_  = \new_[97232]_  & \new_[97225]_ ;
  assign \new_[97236]_  = ~A265 & A202;
  assign \new_[97239]_  = A267 & A266;
  assign \new_[97240]_  = \new_[97239]_  & \new_[97236]_ ;
  assign \new_[97243]_  = A300 & A269;
  assign \new_[97246]_  = ~A302 & ~A301;
  assign \new_[97247]_  = \new_[97246]_  & \new_[97243]_ ;
  assign \new_[97248]_  = \new_[97247]_  & \new_[97240]_ ;
  assign \new_[97251]_  = ~A169 & A170;
  assign \new_[97254]_  = ~A167 & ~A168;
  assign \new_[97255]_  = \new_[97254]_  & \new_[97251]_ ;
  assign \new_[97258]_  = A199 & A166;
  assign \new_[97261]_  = A201 & ~A200;
  assign \new_[97262]_  = \new_[97261]_  & \new_[97258]_ ;
  assign \new_[97263]_  = \new_[97262]_  & \new_[97255]_ ;
  assign \new_[97266]_  = ~A265 & A202;
  assign \new_[97269]_  = ~A267 & A266;
  assign \new_[97270]_  = \new_[97269]_  & \new_[97266]_ ;
  assign \new_[97273]_  = ~A269 & ~A268;
  assign \new_[97276]_  = A301 & ~A300;
  assign \new_[97277]_  = \new_[97276]_  & \new_[97273]_ ;
  assign \new_[97278]_  = \new_[97277]_  & \new_[97270]_ ;
  assign \new_[97281]_  = ~A169 & A170;
  assign \new_[97284]_  = ~A167 & ~A168;
  assign \new_[97285]_  = \new_[97284]_  & \new_[97281]_ ;
  assign \new_[97288]_  = A199 & A166;
  assign \new_[97291]_  = A201 & ~A200;
  assign \new_[97292]_  = \new_[97291]_  & \new_[97288]_ ;
  assign \new_[97293]_  = \new_[97292]_  & \new_[97285]_ ;
  assign \new_[97296]_  = ~A265 & A202;
  assign \new_[97299]_  = ~A267 & A266;
  assign \new_[97300]_  = \new_[97299]_  & \new_[97296]_ ;
  assign \new_[97303]_  = ~A269 & ~A268;
  assign \new_[97306]_  = A302 & ~A300;
  assign \new_[97307]_  = \new_[97306]_  & \new_[97303]_ ;
  assign \new_[97308]_  = \new_[97307]_  & \new_[97300]_ ;
  assign \new_[97311]_  = ~A169 & A170;
  assign \new_[97314]_  = ~A167 & ~A168;
  assign \new_[97315]_  = \new_[97314]_  & \new_[97311]_ ;
  assign \new_[97318]_  = A199 & A166;
  assign \new_[97321]_  = A201 & ~A200;
  assign \new_[97322]_  = \new_[97321]_  & \new_[97318]_ ;
  assign \new_[97323]_  = \new_[97322]_  & \new_[97315]_ ;
  assign \new_[97326]_  = ~A265 & A202;
  assign \new_[97329]_  = ~A267 & A266;
  assign \new_[97330]_  = \new_[97329]_  & \new_[97326]_ ;
  assign \new_[97333]_  = ~A269 & ~A268;
  assign \new_[97336]_  = A299 & A298;
  assign \new_[97337]_  = \new_[97336]_  & \new_[97333]_ ;
  assign \new_[97338]_  = \new_[97337]_  & \new_[97330]_ ;
  assign \new_[97341]_  = ~A169 & A170;
  assign \new_[97344]_  = ~A167 & ~A168;
  assign \new_[97345]_  = \new_[97344]_  & \new_[97341]_ ;
  assign \new_[97348]_  = A199 & A166;
  assign \new_[97351]_  = A201 & ~A200;
  assign \new_[97352]_  = \new_[97351]_  & \new_[97348]_ ;
  assign \new_[97353]_  = \new_[97352]_  & \new_[97345]_ ;
  assign \new_[97356]_  = ~A265 & A202;
  assign \new_[97359]_  = ~A267 & A266;
  assign \new_[97360]_  = \new_[97359]_  & \new_[97356]_ ;
  assign \new_[97363]_  = ~A269 & ~A268;
  assign \new_[97366]_  = ~A299 & ~A298;
  assign \new_[97367]_  = \new_[97366]_  & \new_[97363]_ ;
  assign \new_[97368]_  = \new_[97367]_  & \new_[97360]_ ;
  assign \new_[97371]_  = ~A169 & A170;
  assign \new_[97374]_  = ~A167 & ~A168;
  assign \new_[97375]_  = \new_[97374]_  & \new_[97371]_ ;
  assign \new_[97378]_  = A199 & A166;
  assign \new_[97381]_  = A201 & ~A200;
  assign \new_[97382]_  = \new_[97381]_  & \new_[97378]_ ;
  assign \new_[97383]_  = \new_[97382]_  & \new_[97375]_ ;
  assign \new_[97386]_  = A265 & A202;
  assign \new_[97389]_  = A267 & ~A266;
  assign \new_[97390]_  = \new_[97389]_  & \new_[97386]_ ;
  assign \new_[97393]_  = A300 & A268;
  assign \new_[97396]_  = ~A302 & ~A301;
  assign \new_[97397]_  = \new_[97396]_  & \new_[97393]_ ;
  assign \new_[97398]_  = \new_[97397]_  & \new_[97390]_ ;
  assign \new_[97401]_  = ~A169 & A170;
  assign \new_[97404]_  = ~A167 & ~A168;
  assign \new_[97405]_  = \new_[97404]_  & \new_[97401]_ ;
  assign \new_[97408]_  = A199 & A166;
  assign \new_[97411]_  = A201 & ~A200;
  assign \new_[97412]_  = \new_[97411]_  & \new_[97408]_ ;
  assign \new_[97413]_  = \new_[97412]_  & \new_[97405]_ ;
  assign \new_[97416]_  = A265 & A202;
  assign \new_[97419]_  = A267 & ~A266;
  assign \new_[97420]_  = \new_[97419]_  & \new_[97416]_ ;
  assign \new_[97423]_  = A300 & A269;
  assign \new_[97426]_  = ~A302 & ~A301;
  assign \new_[97427]_  = \new_[97426]_  & \new_[97423]_ ;
  assign \new_[97428]_  = \new_[97427]_  & \new_[97420]_ ;
  assign \new_[97431]_  = ~A169 & A170;
  assign \new_[97434]_  = ~A167 & ~A168;
  assign \new_[97435]_  = \new_[97434]_  & \new_[97431]_ ;
  assign \new_[97438]_  = A199 & A166;
  assign \new_[97441]_  = A201 & ~A200;
  assign \new_[97442]_  = \new_[97441]_  & \new_[97438]_ ;
  assign \new_[97443]_  = \new_[97442]_  & \new_[97435]_ ;
  assign \new_[97446]_  = A265 & A202;
  assign \new_[97449]_  = ~A267 & ~A266;
  assign \new_[97450]_  = \new_[97449]_  & \new_[97446]_ ;
  assign \new_[97453]_  = ~A269 & ~A268;
  assign \new_[97456]_  = A301 & ~A300;
  assign \new_[97457]_  = \new_[97456]_  & \new_[97453]_ ;
  assign \new_[97458]_  = \new_[97457]_  & \new_[97450]_ ;
  assign \new_[97461]_  = ~A169 & A170;
  assign \new_[97464]_  = ~A167 & ~A168;
  assign \new_[97465]_  = \new_[97464]_  & \new_[97461]_ ;
  assign \new_[97468]_  = A199 & A166;
  assign \new_[97471]_  = A201 & ~A200;
  assign \new_[97472]_  = \new_[97471]_  & \new_[97468]_ ;
  assign \new_[97473]_  = \new_[97472]_  & \new_[97465]_ ;
  assign \new_[97476]_  = A265 & A202;
  assign \new_[97479]_  = ~A267 & ~A266;
  assign \new_[97480]_  = \new_[97479]_  & \new_[97476]_ ;
  assign \new_[97483]_  = ~A269 & ~A268;
  assign \new_[97486]_  = A302 & ~A300;
  assign \new_[97487]_  = \new_[97486]_  & \new_[97483]_ ;
  assign \new_[97488]_  = \new_[97487]_  & \new_[97480]_ ;
  assign \new_[97491]_  = ~A169 & A170;
  assign \new_[97494]_  = ~A167 & ~A168;
  assign \new_[97495]_  = \new_[97494]_  & \new_[97491]_ ;
  assign \new_[97498]_  = A199 & A166;
  assign \new_[97501]_  = A201 & ~A200;
  assign \new_[97502]_  = \new_[97501]_  & \new_[97498]_ ;
  assign \new_[97503]_  = \new_[97502]_  & \new_[97495]_ ;
  assign \new_[97506]_  = A265 & A202;
  assign \new_[97509]_  = ~A267 & ~A266;
  assign \new_[97510]_  = \new_[97509]_  & \new_[97506]_ ;
  assign \new_[97513]_  = ~A269 & ~A268;
  assign \new_[97516]_  = A299 & A298;
  assign \new_[97517]_  = \new_[97516]_  & \new_[97513]_ ;
  assign \new_[97518]_  = \new_[97517]_  & \new_[97510]_ ;
  assign \new_[97521]_  = ~A169 & A170;
  assign \new_[97524]_  = ~A167 & ~A168;
  assign \new_[97525]_  = \new_[97524]_  & \new_[97521]_ ;
  assign \new_[97528]_  = A199 & A166;
  assign \new_[97531]_  = A201 & ~A200;
  assign \new_[97532]_  = \new_[97531]_  & \new_[97528]_ ;
  assign \new_[97533]_  = \new_[97532]_  & \new_[97525]_ ;
  assign \new_[97536]_  = A265 & A202;
  assign \new_[97539]_  = ~A267 & ~A266;
  assign \new_[97540]_  = \new_[97539]_  & \new_[97536]_ ;
  assign \new_[97543]_  = ~A269 & ~A268;
  assign \new_[97546]_  = ~A299 & ~A298;
  assign \new_[97547]_  = \new_[97546]_  & \new_[97543]_ ;
  assign \new_[97548]_  = \new_[97547]_  & \new_[97540]_ ;
  assign \new_[97551]_  = ~A169 & A170;
  assign \new_[97554]_  = ~A167 & ~A168;
  assign \new_[97555]_  = \new_[97554]_  & \new_[97551]_ ;
  assign \new_[97558]_  = A199 & A166;
  assign \new_[97561]_  = A201 & ~A200;
  assign \new_[97562]_  = \new_[97561]_  & \new_[97558]_ ;
  assign \new_[97563]_  = \new_[97562]_  & \new_[97555]_ ;
  assign \new_[97566]_  = ~A265 & A203;
  assign \new_[97569]_  = A267 & A266;
  assign \new_[97570]_  = \new_[97569]_  & \new_[97566]_ ;
  assign \new_[97573]_  = A300 & A268;
  assign \new_[97576]_  = ~A302 & ~A301;
  assign \new_[97577]_  = \new_[97576]_  & \new_[97573]_ ;
  assign \new_[97578]_  = \new_[97577]_  & \new_[97570]_ ;
  assign \new_[97581]_  = ~A169 & A170;
  assign \new_[97584]_  = ~A167 & ~A168;
  assign \new_[97585]_  = \new_[97584]_  & \new_[97581]_ ;
  assign \new_[97588]_  = A199 & A166;
  assign \new_[97591]_  = A201 & ~A200;
  assign \new_[97592]_  = \new_[97591]_  & \new_[97588]_ ;
  assign \new_[97593]_  = \new_[97592]_  & \new_[97585]_ ;
  assign \new_[97596]_  = ~A265 & A203;
  assign \new_[97599]_  = A267 & A266;
  assign \new_[97600]_  = \new_[97599]_  & \new_[97596]_ ;
  assign \new_[97603]_  = A300 & A269;
  assign \new_[97606]_  = ~A302 & ~A301;
  assign \new_[97607]_  = \new_[97606]_  & \new_[97603]_ ;
  assign \new_[97608]_  = \new_[97607]_  & \new_[97600]_ ;
  assign \new_[97611]_  = ~A169 & A170;
  assign \new_[97614]_  = ~A167 & ~A168;
  assign \new_[97615]_  = \new_[97614]_  & \new_[97611]_ ;
  assign \new_[97618]_  = A199 & A166;
  assign \new_[97621]_  = A201 & ~A200;
  assign \new_[97622]_  = \new_[97621]_  & \new_[97618]_ ;
  assign \new_[97623]_  = \new_[97622]_  & \new_[97615]_ ;
  assign \new_[97626]_  = ~A265 & A203;
  assign \new_[97629]_  = ~A267 & A266;
  assign \new_[97630]_  = \new_[97629]_  & \new_[97626]_ ;
  assign \new_[97633]_  = ~A269 & ~A268;
  assign \new_[97636]_  = A301 & ~A300;
  assign \new_[97637]_  = \new_[97636]_  & \new_[97633]_ ;
  assign \new_[97638]_  = \new_[97637]_  & \new_[97630]_ ;
  assign \new_[97641]_  = ~A169 & A170;
  assign \new_[97644]_  = ~A167 & ~A168;
  assign \new_[97645]_  = \new_[97644]_  & \new_[97641]_ ;
  assign \new_[97648]_  = A199 & A166;
  assign \new_[97651]_  = A201 & ~A200;
  assign \new_[97652]_  = \new_[97651]_  & \new_[97648]_ ;
  assign \new_[97653]_  = \new_[97652]_  & \new_[97645]_ ;
  assign \new_[97656]_  = ~A265 & A203;
  assign \new_[97659]_  = ~A267 & A266;
  assign \new_[97660]_  = \new_[97659]_  & \new_[97656]_ ;
  assign \new_[97663]_  = ~A269 & ~A268;
  assign \new_[97666]_  = A302 & ~A300;
  assign \new_[97667]_  = \new_[97666]_  & \new_[97663]_ ;
  assign \new_[97668]_  = \new_[97667]_  & \new_[97660]_ ;
  assign \new_[97671]_  = ~A169 & A170;
  assign \new_[97674]_  = ~A167 & ~A168;
  assign \new_[97675]_  = \new_[97674]_  & \new_[97671]_ ;
  assign \new_[97678]_  = A199 & A166;
  assign \new_[97681]_  = A201 & ~A200;
  assign \new_[97682]_  = \new_[97681]_  & \new_[97678]_ ;
  assign \new_[97683]_  = \new_[97682]_  & \new_[97675]_ ;
  assign \new_[97686]_  = ~A265 & A203;
  assign \new_[97689]_  = ~A267 & A266;
  assign \new_[97690]_  = \new_[97689]_  & \new_[97686]_ ;
  assign \new_[97693]_  = ~A269 & ~A268;
  assign \new_[97696]_  = A299 & A298;
  assign \new_[97697]_  = \new_[97696]_  & \new_[97693]_ ;
  assign \new_[97698]_  = \new_[97697]_  & \new_[97690]_ ;
  assign \new_[97701]_  = ~A169 & A170;
  assign \new_[97704]_  = ~A167 & ~A168;
  assign \new_[97705]_  = \new_[97704]_  & \new_[97701]_ ;
  assign \new_[97708]_  = A199 & A166;
  assign \new_[97711]_  = A201 & ~A200;
  assign \new_[97712]_  = \new_[97711]_  & \new_[97708]_ ;
  assign \new_[97713]_  = \new_[97712]_  & \new_[97705]_ ;
  assign \new_[97716]_  = ~A265 & A203;
  assign \new_[97719]_  = ~A267 & A266;
  assign \new_[97720]_  = \new_[97719]_  & \new_[97716]_ ;
  assign \new_[97723]_  = ~A269 & ~A268;
  assign \new_[97726]_  = ~A299 & ~A298;
  assign \new_[97727]_  = \new_[97726]_  & \new_[97723]_ ;
  assign \new_[97728]_  = \new_[97727]_  & \new_[97720]_ ;
  assign \new_[97731]_  = ~A169 & A170;
  assign \new_[97734]_  = ~A167 & ~A168;
  assign \new_[97735]_  = \new_[97734]_  & \new_[97731]_ ;
  assign \new_[97738]_  = A199 & A166;
  assign \new_[97741]_  = A201 & ~A200;
  assign \new_[97742]_  = \new_[97741]_  & \new_[97738]_ ;
  assign \new_[97743]_  = \new_[97742]_  & \new_[97735]_ ;
  assign \new_[97746]_  = A265 & A203;
  assign \new_[97749]_  = A267 & ~A266;
  assign \new_[97750]_  = \new_[97749]_  & \new_[97746]_ ;
  assign \new_[97753]_  = A300 & A268;
  assign \new_[97756]_  = ~A302 & ~A301;
  assign \new_[97757]_  = \new_[97756]_  & \new_[97753]_ ;
  assign \new_[97758]_  = \new_[97757]_  & \new_[97750]_ ;
  assign \new_[97761]_  = ~A169 & A170;
  assign \new_[97764]_  = ~A167 & ~A168;
  assign \new_[97765]_  = \new_[97764]_  & \new_[97761]_ ;
  assign \new_[97768]_  = A199 & A166;
  assign \new_[97771]_  = A201 & ~A200;
  assign \new_[97772]_  = \new_[97771]_  & \new_[97768]_ ;
  assign \new_[97773]_  = \new_[97772]_  & \new_[97765]_ ;
  assign \new_[97776]_  = A265 & A203;
  assign \new_[97779]_  = A267 & ~A266;
  assign \new_[97780]_  = \new_[97779]_  & \new_[97776]_ ;
  assign \new_[97783]_  = A300 & A269;
  assign \new_[97786]_  = ~A302 & ~A301;
  assign \new_[97787]_  = \new_[97786]_  & \new_[97783]_ ;
  assign \new_[97788]_  = \new_[97787]_  & \new_[97780]_ ;
  assign \new_[97791]_  = ~A169 & A170;
  assign \new_[97794]_  = ~A167 & ~A168;
  assign \new_[97795]_  = \new_[97794]_  & \new_[97791]_ ;
  assign \new_[97798]_  = A199 & A166;
  assign \new_[97801]_  = A201 & ~A200;
  assign \new_[97802]_  = \new_[97801]_  & \new_[97798]_ ;
  assign \new_[97803]_  = \new_[97802]_  & \new_[97795]_ ;
  assign \new_[97806]_  = A265 & A203;
  assign \new_[97809]_  = ~A267 & ~A266;
  assign \new_[97810]_  = \new_[97809]_  & \new_[97806]_ ;
  assign \new_[97813]_  = ~A269 & ~A268;
  assign \new_[97816]_  = A301 & ~A300;
  assign \new_[97817]_  = \new_[97816]_  & \new_[97813]_ ;
  assign \new_[97818]_  = \new_[97817]_  & \new_[97810]_ ;
  assign \new_[97821]_  = ~A169 & A170;
  assign \new_[97824]_  = ~A167 & ~A168;
  assign \new_[97825]_  = \new_[97824]_  & \new_[97821]_ ;
  assign \new_[97828]_  = A199 & A166;
  assign \new_[97831]_  = A201 & ~A200;
  assign \new_[97832]_  = \new_[97831]_  & \new_[97828]_ ;
  assign \new_[97833]_  = \new_[97832]_  & \new_[97825]_ ;
  assign \new_[97836]_  = A265 & A203;
  assign \new_[97839]_  = ~A267 & ~A266;
  assign \new_[97840]_  = \new_[97839]_  & \new_[97836]_ ;
  assign \new_[97843]_  = ~A269 & ~A268;
  assign \new_[97846]_  = A302 & ~A300;
  assign \new_[97847]_  = \new_[97846]_  & \new_[97843]_ ;
  assign \new_[97848]_  = \new_[97847]_  & \new_[97840]_ ;
  assign \new_[97851]_  = ~A169 & A170;
  assign \new_[97854]_  = ~A167 & ~A168;
  assign \new_[97855]_  = \new_[97854]_  & \new_[97851]_ ;
  assign \new_[97858]_  = A199 & A166;
  assign \new_[97861]_  = A201 & ~A200;
  assign \new_[97862]_  = \new_[97861]_  & \new_[97858]_ ;
  assign \new_[97863]_  = \new_[97862]_  & \new_[97855]_ ;
  assign \new_[97866]_  = A265 & A203;
  assign \new_[97869]_  = ~A267 & ~A266;
  assign \new_[97870]_  = \new_[97869]_  & \new_[97866]_ ;
  assign \new_[97873]_  = ~A269 & ~A268;
  assign \new_[97876]_  = A299 & A298;
  assign \new_[97877]_  = \new_[97876]_  & \new_[97873]_ ;
  assign \new_[97878]_  = \new_[97877]_  & \new_[97870]_ ;
  assign \new_[97881]_  = ~A169 & A170;
  assign \new_[97884]_  = ~A167 & ~A168;
  assign \new_[97885]_  = \new_[97884]_  & \new_[97881]_ ;
  assign \new_[97888]_  = A199 & A166;
  assign \new_[97891]_  = A201 & ~A200;
  assign \new_[97892]_  = \new_[97891]_  & \new_[97888]_ ;
  assign \new_[97893]_  = \new_[97892]_  & \new_[97885]_ ;
  assign \new_[97896]_  = A265 & A203;
  assign \new_[97899]_  = ~A267 & ~A266;
  assign \new_[97900]_  = \new_[97899]_  & \new_[97896]_ ;
  assign \new_[97903]_  = ~A269 & ~A268;
  assign \new_[97906]_  = ~A299 & ~A298;
  assign \new_[97907]_  = \new_[97906]_  & \new_[97903]_ ;
  assign \new_[97908]_  = \new_[97907]_  & \new_[97900]_ ;
  assign \new_[97911]_  = ~A169 & A170;
  assign \new_[97914]_  = ~A167 & ~A168;
  assign \new_[97915]_  = \new_[97914]_  & \new_[97911]_ ;
  assign \new_[97918]_  = A199 & A166;
  assign \new_[97921]_  = ~A201 & ~A200;
  assign \new_[97922]_  = \new_[97921]_  & \new_[97918]_ ;
  assign \new_[97923]_  = \new_[97922]_  & \new_[97915]_ ;
  assign \new_[97926]_  = ~A203 & ~A202;
  assign \new_[97929]_  = A266 & ~A265;
  assign \new_[97930]_  = \new_[97929]_  & \new_[97926]_ ;
  assign \new_[97933]_  = A268 & A267;
  assign \new_[97936]_  = A301 & ~A300;
  assign \new_[97937]_  = \new_[97936]_  & \new_[97933]_ ;
  assign \new_[97938]_  = \new_[97937]_  & \new_[97930]_ ;
  assign \new_[97941]_  = ~A169 & A170;
  assign \new_[97944]_  = ~A167 & ~A168;
  assign \new_[97945]_  = \new_[97944]_  & \new_[97941]_ ;
  assign \new_[97948]_  = A199 & A166;
  assign \new_[97951]_  = ~A201 & ~A200;
  assign \new_[97952]_  = \new_[97951]_  & \new_[97948]_ ;
  assign \new_[97953]_  = \new_[97952]_  & \new_[97945]_ ;
  assign \new_[97956]_  = ~A203 & ~A202;
  assign \new_[97959]_  = A266 & ~A265;
  assign \new_[97960]_  = \new_[97959]_  & \new_[97956]_ ;
  assign \new_[97963]_  = A268 & A267;
  assign \new_[97966]_  = A302 & ~A300;
  assign \new_[97967]_  = \new_[97966]_  & \new_[97963]_ ;
  assign \new_[97968]_  = \new_[97967]_  & \new_[97960]_ ;
  assign \new_[97971]_  = ~A169 & A170;
  assign \new_[97974]_  = ~A167 & ~A168;
  assign \new_[97975]_  = \new_[97974]_  & \new_[97971]_ ;
  assign \new_[97978]_  = A199 & A166;
  assign \new_[97981]_  = ~A201 & ~A200;
  assign \new_[97982]_  = \new_[97981]_  & \new_[97978]_ ;
  assign \new_[97983]_  = \new_[97982]_  & \new_[97975]_ ;
  assign \new_[97986]_  = ~A203 & ~A202;
  assign \new_[97989]_  = A266 & ~A265;
  assign \new_[97990]_  = \new_[97989]_  & \new_[97986]_ ;
  assign \new_[97993]_  = A268 & A267;
  assign \new_[97996]_  = A299 & A298;
  assign \new_[97997]_  = \new_[97996]_  & \new_[97993]_ ;
  assign \new_[97998]_  = \new_[97997]_  & \new_[97990]_ ;
  assign \new_[98001]_  = ~A169 & A170;
  assign \new_[98004]_  = ~A167 & ~A168;
  assign \new_[98005]_  = \new_[98004]_  & \new_[98001]_ ;
  assign \new_[98008]_  = A199 & A166;
  assign \new_[98011]_  = ~A201 & ~A200;
  assign \new_[98012]_  = \new_[98011]_  & \new_[98008]_ ;
  assign \new_[98013]_  = \new_[98012]_  & \new_[98005]_ ;
  assign \new_[98016]_  = ~A203 & ~A202;
  assign \new_[98019]_  = A266 & ~A265;
  assign \new_[98020]_  = \new_[98019]_  & \new_[98016]_ ;
  assign \new_[98023]_  = A268 & A267;
  assign \new_[98026]_  = ~A299 & ~A298;
  assign \new_[98027]_  = \new_[98026]_  & \new_[98023]_ ;
  assign \new_[98028]_  = \new_[98027]_  & \new_[98020]_ ;
  assign \new_[98031]_  = ~A169 & A170;
  assign \new_[98034]_  = ~A167 & ~A168;
  assign \new_[98035]_  = \new_[98034]_  & \new_[98031]_ ;
  assign \new_[98038]_  = A199 & A166;
  assign \new_[98041]_  = ~A201 & ~A200;
  assign \new_[98042]_  = \new_[98041]_  & \new_[98038]_ ;
  assign \new_[98043]_  = \new_[98042]_  & \new_[98035]_ ;
  assign \new_[98046]_  = ~A203 & ~A202;
  assign \new_[98049]_  = A266 & ~A265;
  assign \new_[98050]_  = \new_[98049]_  & \new_[98046]_ ;
  assign \new_[98053]_  = A269 & A267;
  assign \new_[98056]_  = A301 & ~A300;
  assign \new_[98057]_  = \new_[98056]_  & \new_[98053]_ ;
  assign \new_[98058]_  = \new_[98057]_  & \new_[98050]_ ;
  assign \new_[98061]_  = ~A169 & A170;
  assign \new_[98064]_  = ~A167 & ~A168;
  assign \new_[98065]_  = \new_[98064]_  & \new_[98061]_ ;
  assign \new_[98068]_  = A199 & A166;
  assign \new_[98071]_  = ~A201 & ~A200;
  assign \new_[98072]_  = \new_[98071]_  & \new_[98068]_ ;
  assign \new_[98073]_  = \new_[98072]_  & \new_[98065]_ ;
  assign \new_[98076]_  = ~A203 & ~A202;
  assign \new_[98079]_  = A266 & ~A265;
  assign \new_[98080]_  = \new_[98079]_  & \new_[98076]_ ;
  assign \new_[98083]_  = A269 & A267;
  assign \new_[98086]_  = A302 & ~A300;
  assign \new_[98087]_  = \new_[98086]_  & \new_[98083]_ ;
  assign \new_[98088]_  = \new_[98087]_  & \new_[98080]_ ;
  assign \new_[98091]_  = ~A169 & A170;
  assign \new_[98094]_  = ~A167 & ~A168;
  assign \new_[98095]_  = \new_[98094]_  & \new_[98091]_ ;
  assign \new_[98098]_  = A199 & A166;
  assign \new_[98101]_  = ~A201 & ~A200;
  assign \new_[98102]_  = \new_[98101]_  & \new_[98098]_ ;
  assign \new_[98103]_  = \new_[98102]_  & \new_[98095]_ ;
  assign \new_[98106]_  = ~A203 & ~A202;
  assign \new_[98109]_  = A266 & ~A265;
  assign \new_[98110]_  = \new_[98109]_  & \new_[98106]_ ;
  assign \new_[98113]_  = A269 & A267;
  assign \new_[98116]_  = A299 & A298;
  assign \new_[98117]_  = \new_[98116]_  & \new_[98113]_ ;
  assign \new_[98118]_  = \new_[98117]_  & \new_[98110]_ ;
  assign \new_[98121]_  = ~A169 & A170;
  assign \new_[98124]_  = ~A167 & ~A168;
  assign \new_[98125]_  = \new_[98124]_  & \new_[98121]_ ;
  assign \new_[98128]_  = A199 & A166;
  assign \new_[98131]_  = ~A201 & ~A200;
  assign \new_[98132]_  = \new_[98131]_  & \new_[98128]_ ;
  assign \new_[98133]_  = \new_[98132]_  & \new_[98125]_ ;
  assign \new_[98136]_  = ~A203 & ~A202;
  assign \new_[98139]_  = A266 & ~A265;
  assign \new_[98140]_  = \new_[98139]_  & \new_[98136]_ ;
  assign \new_[98143]_  = A269 & A267;
  assign \new_[98146]_  = ~A299 & ~A298;
  assign \new_[98147]_  = \new_[98146]_  & \new_[98143]_ ;
  assign \new_[98148]_  = \new_[98147]_  & \new_[98140]_ ;
  assign \new_[98151]_  = ~A169 & A170;
  assign \new_[98154]_  = ~A167 & ~A168;
  assign \new_[98155]_  = \new_[98154]_  & \new_[98151]_ ;
  assign \new_[98158]_  = A199 & A166;
  assign \new_[98161]_  = ~A201 & ~A200;
  assign \new_[98162]_  = \new_[98161]_  & \new_[98158]_ ;
  assign \new_[98163]_  = \new_[98162]_  & \new_[98155]_ ;
  assign \new_[98166]_  = ~A203 & ~A202;
  assign \new_[98169]_  = ~A266 & A265;
  assign \new_[98170]_  = \new_[98169]_  & \new_[98166]_ ;
  assign \new_[98173]_  = A268 & A267;
  assign \new_[98176]_  = A301 & ~A300;
  assign \new_[98177]_  = \new_[98176]_  & \new_[98173]_ ;
  assign \new_[98178]_  = \new_[98177]_  & \new_[98170]_ ;
  assign \new_[98181]_  = ~A169 & A170;
  assign \new_[98184]_  = ~A167 & ~A168;
  assign \new_[98185]_  = \new_[98184]_  & \new_[98181]_ ;
  assign \new_[98188]_  = A199 & A166;
  assign \new_[98191]_  = ~A201 & ~A200;
  assign \new_[98192]_  = \new_[98191]_  & \new_[98188]_ ;
  assign \new_[98193]_  = \new_[98192]_  & \new_[98185]_ ;
  assign \new_[98196]_  = ~A203 & ~A202;
  assign \new_[98199]_  = ~A266 & A265;
  assign \new_[98200]_  = \new_[98199]_  & \new_[98196]_ ;
  assign \new_[98203]_  = A268 & A267;
  assign \new_[98206]_  = A302 & ~A300;
  assign \new_[98207]_  = \new_[98206]_  & \new_[98203]_ ;
  assign \new_[98208]_  = \new_[98207]_  & \new_[98200]_ ;
  assign \new_[98211]_  = ~A169 & A170;
  assign \new_[98214]_  = ~A167 & ~A168;
  assign \new_[98215]_  = \new_[98214]_  & \new_[98211]_ ;
  assign \new_[98218]_  = A199 & A166;
  assign \new_[98221]_  = ~A201 & ~A200;
  assign \new_[98222]_  = \new_[98221]_  & \new_[98218]_ ;
  assign \new_[98223]_  = \new_[98222]_  & \new_[98215]_ ;
  assign \new_[98226]_  = ~A203 & ~A202;
  assign \new_[98229]_  = ~A266 & A265;
  assign \new_[98230]_  = \new_[98229]_  & \new_[98226]_ ;
  assign \new_[98233]_  = A268 & A267;
  assign \new_[98236]_  = A299 & A298;
  assign \new_[98237]_  = \new_[98236]_  & \new_[98233]_ ;
  assign \new_[98238]_  = \new_[98237]_  & \new_[98230]_ ;
  assign \new_[98241]_  = ~A169 & A170;
  assign \new_[98244]_  = ~A167 & ~A168;
  assign \new_[98245]_  = \new_[98244]_  & \new_[98241]_ ;
  assign \new_[98248]_  = A199 & A166;
  assign \new_[98251]_  = ~A201 & ~A200;
  assign \new_[98252]_  = \new_[98251]_  & \new_[98248]_ ;
  assign \new_[98253]_  = \new_[98252]_  & \new_[98245]_ ;
  assign \new_[98256]_  = ~A203 & ~A202;
  assign \new_[98259]_  = ~A266 & A265;
  assign \new_[98260]_  = \new_[98259]_  & \new_[98256]_ ;
  assign \new_[98263]_  = A268 & A267;
  assign \new_[98266]_  = ~A299 & ~A298;
  assign \new_[98267]_  = \new_[98266]_  & \new_[98263]_ ;
  assign \new_[98268]_  = \new_[98267]_  & \new_[98260]_ ;
  assign \new_[98271]_  = ~A169 & A170;
  assign \new_[98274]_  = ~A167 & ~A168;
  assign \new_[98275]_  = \new_[98274]_  & \new_[98271]_ ;
  assign \new_[98278]_  = A199 & A166;
  assign \new_[98281]_  = ~A201 & ~A200;
  assign \new_[98282]_  = \new_[98281]_  & \new_[98278]_ ;
  assign \new_[98283]_  = \new_[98282]_  & \new_[98275]_ ;
  assign \new_[98286]_  = ~A203 & ~A202;
  assign \new_[98289]_  = ~A266 & A265;
  assign \new_[98290]_  = \new_[98289]_  & \new_[98286]_ ;
  assign \new_[98293]_  = A269 & A267;
  assign \new_[98296]_  = A301 & ~A300;
  assign \new_[98297]_  = \new_[98296]_  & \new_[98293]_ ;
  assign \new_[98298]_  = \new_[98297]_  & \new_[98290]_ ;
  assign \new_[98301]_  = ~A169 & A170;
  assign \new_[98304]_  = ~A167 & ~A168;
  assign \new_[98305]_  = \new_[98304]_  & \new_[98301]_ ;
  assign \new_[98308]_  = A199 & A166;
  assign \new_[98311]_  = ~A201 & ~A200;
  assign \new_[98312]_  = \new_[98311]_  & \new_[98308]_ ;
  assign \new_[98313]_  = \new_[98312]_  & \new_[98305]_ ;
  assign \new_[98316]_  = ~A203 & ~A202;
  assign \new_[98319]_  = ~A266 & A265;
  assign \new_[98320]_  = \new_[98319]_  & \new_[98316]_ ;
  assign \new_[98323]_  = A269 & A267;
  assign \new_[98326]_  = A302 & ~A300;
  assign \new_[98327]_  = \new_[98326]_  & \new_[98323]_ ;
  assign \new_[98328]_  = \new_[98327]_  & \new_[98320]_ ;
  assign \new_[98331]_  = ~A169 & A170;
  assign \new_[98334]_  = ~A167 & ~A168;
  assign \new_[98335]_  = \new_[98334]_  & \new_[98331]_ ;
  assign \new_[98338]_  = A199 & A166;
  assign \new_[98341]_  = ~A201 & ~A200;
  assign \new_[98342]_  = \new_[98341]_  & \new_[98338]_ ;
  assign \new_[98343]_  = \new_[98342]_  & \new_[98335]_ ;
  assign \new_[98346]_  = ~A203 & ~A202;
  assign \new_[98349]_  = ~A266 & A265;
  assign \new_[98350]_  = \new_[98349]_  & \new_[98346]_ ;
  assign \new_[98353]_  = A269 & A267;
  assign \new_[98356]_  = A299 & A298;
  assign \new_[98357]_  = \new_[98356]_  & \new_[98353]_ ;
  assign \new_[98358]_  = \new_[98357]_  & \new_[98350]_ ;
  assign \new_[98361]_  = ~A169 & A170;
  assign \new_[98364]_  = ~A167 & ~A168;
  assign \new_[98365]_  = \new_[98364]_  & \new_[98361]_ ;
  assign \new_[98368]_  = A199 & A166;
  assign \new_[98371]_  = ~A201 & ~A200;
  assign \new_[98372]_  = \new_[98371]_  & \new_[98368]_ ;
  assign \new_[98373]_  = \new_[98372]_  & \new_[98365]_ ;
  assign \new_[98376]_  = ~A203 & ~A202;
  assign \new_[98379]_  = ~A266 & A265;
  assign \new_[98380]_  = \new_[98379]_  & \new_[98376]_ ;
  assign \new_[98383]_  = A269 & A267;
  assign \new_[98386]_  = ~A299 & ~A298;
  assign \new_[98387]_  = \new_[98386]_  & \new_[98383]_ ;
  assign \new_[98388]_  = \new_[98387]_  & \new_[98380]_ ;
  assign \new_[98391]_  = A168 & ~A170;
  assign \new_[98394]_  = ~A166 & A167;
  assign \new_[98395]_  = \new_[98394]_  & \new_[98391]_ ;
  assign \new_[98398]_  = A200 & ~A199;
  assign \new_[98401]_  = ~A202 & ~A201;
  assign \new_[98402]_  = \new_[98401]_  & \new_[98398]_ ;
  assign \new_[98403]_  = \new_[98402]_  & \new_[98395]_ ;
  assign \new_[98406]_  = ~A265 & ~A203;
  assign \new_[98409]_  = ~A267 & A266;
  assign \new_[98410]_  = \new_[98409]_  & \new_[98406]_ ;
  assign \new_[98413]_  = ~A269 & ~A268;
  assign \new_[98417]_  = ~A302 & ~A301;
  assign \new_[98418]_  = A300 & \new_[98417]_ ;
  assign \new_[98419]_  = \new_[98418]_  & \new_[98413]_ ;
  assign \new_[98420]_  = \new_[98419]_  & \new_[98410]_ ;
  assign \new_[98423]_  = A168 & ~A170;
  assign \new_[98426]_  = ~A166 & A167;
  assign \new_[98427]_  = \new_[98426]_  & \new_[98423]_ ;
  assign \new_[98430]_  = A200 & ~A199;
  assign \new_[98433]_  = ~A202 & ~A201;
  assign \new_[98434]_  = \new_[98433]_  & \new_[98430]_ ;
  assign \new_[98435]_  = \new_[98434]_  & \new_[98427]_ ;
  assign \new_[98438]_  = A265 & ~A203;
  assign \new_[98441]_  = ~A267 & ~A266;
  assign \new_[98442]_  = \new_[98441]_  & \new_[98438]_ ;
  assign \new_[98445]_  = ~A269 & ~A268;
  assign \new_[98449]_  = ~A302 & ~A301;
  assign \new_[98450]_  = A300 & \new_[98449]_ ;
  assign \new_[98451]_  = \new_[98450]_  & \new_[98445]_ ;
  assign \new_[98452]_  = \new_[98451]_  & \new_[98442]_ ;
  assign \new_[98455]_  = A168 & ~A170;
  assign \new_[98458]_  = ~A166 & A167;
  assign \new_[98459]_  = \new_[98458]_  & \new_[98455]_ ;
  assign \new_[98462]_  = ~A200 & A199;
  assign \new_[98465]_  = ~A202 & ~A201;
  assign \new_[98466]_  = \new_[98465]_  & \new_[98462]_ ;
  assign \new_[98467]_  = \new_[98466]_  & \new_[98459]_ ;
  assign \new_[98470]_  = ~A265 & ~A203;
  assign \new_[98473]_  = ~A267 & A266;
  assign \new_[98474]_  = \new_[98473]_  & \new_[98470]_ ;
  assign \new_[98477]_  = ~A269 & ~A268;
  assign \new_[98481]_  = ~A302 & ~A301;
  assign \new_[98482]_  = A300 & \new_[98481]_ ;
  assign \new_[98483]_  = \new_[98482]_  & \new_[98477]_ ;
  assign \new_[98484]_  = \new_[98483]_  & \new_[98474]_ ;
  assign \new_[98487]_  = A168 & ~A170;
  assign \new_[98490]_  = ~A166 & A167;
  assign \new_[98491]_  = \new_[98490]_  & \new_[98487]_ ;
  assign \new_[98494]_  = ~A200 & A199;
  assign \new_[98497]_  = ~A202 & ~A201;
  assign \new_[98498]_  = \new_[98497]_  & \new_[98494]_ ;
  assign \new_[98499]_  = \new_[98498]_  & \new_[98491]_ ;
  assign \new_[98502]_  = A265 & ~A203;
  assign \new_[98505]_  = ~A267 & ~A266;
  assign \new_[98506]_  = \new_[98505]_  & \new_[98502]_ ;
  assign \new_[98509]_  = ~A269 & ~A268;
  assign \new_[98513]_  = ~A302 & ~A301;
  assign \new_[98514]_  = A300 & \new_[98513]_ ;
  assign \new_[98515]_  = \new_[98514]_  & \new_[98509]_ ;
  assign \new_[98516]_  = \new_[98515]_  & \new_[98506]_ ;
  assign \new_[98519]_  = A168 & ~A170;
  assign \new_[98522]_  = A166 & ~A167;
  assign \new_[98523]_  = \new_[98522]_  & \new_[98519]_ ;
  assign \new_[98526]_  = A200 & ~A199;
  assign \new_[98529]_  = ~A202 & ~A201;
  assign \new_[98530]_  = \new_[98529]_  & \new_[98526]_ ;
  assign \new_[98531]_  = \new_[98530]_  & \new_[98523]_ ;
  assign \new_[98534]_  = ~A265 & ~A203;
  assign \new_[98537]_  = ~A267 & A266;
  assign \new_[98538]_  = \new_[98537]_  & \new_[98534]_ ;
  assign \new_[98541]_  = ~A269 & ~A268;
  assign \new_[98545]_  = ~A302 & ~A301;
  assign \new_[98546]_  = A300 & \new_[98545]_ ;
  assign \new_[98547]_  = \new_[98546]_  & \new_[98541]_ ;
  assign \new_[98548]_  = \new_[98547]_  & \new_[98538]_ ;
  assign \new_[98551]_  = A168 & ~A170;
  assign \new_[98554]_  = A166 & ~A167;
  assign \new_[98555]_  = \new_[98554]_  & \new_[98551]_ ;
  assign \new_[98558]_  = A200 & ~A199;
  assign \new_[98561]_  = ~A202 & ~A201;
  assign \new_[98562]_  = \new_[98561]_  & \new_[98558]_ ;
  assign \new_[98563]_  = \new_[98562]_  & \new_[98555]_ ;
  assign \new_[98566]_  = A265 & ~A203;
  assign \new_[98569]_  = ~A267 & ~A266;
  assign \new_[98570]_  = \new_[98569]_  & \new_[98566]_ ;
  assign \new_[98573]_  = ~A269 & ~A268;
  assign \new_[98577]_  = ~A302 & ~A301;
  assign \new_[98578]_  = A300 & \new_[98577]_ ;
  assign \new_[98579]_  = \new_[98578]_  & \new_[98573]_ ;
  assign \new_[98580]_  = \new_[98579]_  & \new_[98570]_ ;
  assign \new_[98583]_  = A168 & ~A170;
  assign \new_[98586]_  = A166 & ~A167;
  assign \new_[98587]_  = \new_[98586]_  & \new_[98583]_ ;
  assign \new_[98590]_  = ~A200 & A199;
  assign \new_[98593]_  = ~A202 & ~A201;
  assign \new_[98594]_  = \new_[98593]_  & \new_[98590]_ ;
  assign \new_[98595]_  = \new_[98594]_  & \new_[98587]_ ;
  assign \new_[98598]_  = ~A265 & ~A203;
  assign \new_[98601]_  = ~A267 & A266;
  assign \new_[98602]_  = \new_[98601]_  & \new_[98598]_ ;
  assign \new_[98605]_  = ~A269 & ~A268;
  assign \new_[98609]_  = ~A302 & ~A301;
  assign \new_[98610]_  = A300 & \new_[98609]_ ;
  assign \new_[98611]_  = \new_[98610]_  & \new_[98605]_ ;
  assign \new_[98612]_  = \new_[98611]_  & \new_[98602]_ ;
  assign \new_[98615]_  = A168 & ~A170;
  assign \new_[98618]_  = A166 & ~A167;
  assign \new_[98619]_  = \new_[98618]_  & \new_[98615]_ ;
  assign \new_[98622]_  = ~A200 & A199;
  assign \new_[98625]_  = ~A202 & ~A201;
  assign \new_[98626]_  = \new_[98625]_  & \new_[98622]_ ;
  assign \new_[98627]_  = \new_[98626]_  & \new_[98619]_ ;
  assign \new_[98630]_  = A265 & ~A203;
  assign \new_[98633]_  = ~A267 & ~A266;
  assign \new_[98634]_  = \new_[98633]_  & \new_[98630]_ ;
  assign \new_[98637]_  = ~A269 & ~A268;
  assign \new_[98641]_  = ~A302 & ~A301;
  assign \new_[98642]_  = A300 & \new_[98641]_ ;
  assign \new_[98643]_  = \new_[98642]_  & \new_[98637]_ ;
  assign \new_[98644]_  = \new_[98643]_  & \new_[98634]_ ;
  assign \new_[98647]_  = A168 & A169;
  assign \new_[98650]_  = ~A166 & A167;
  assign \new_[98651]_  = \new_[98650]_  & \new_[98647]_ ;
  assign \new_[98654]_  = A200 & ~A199;
  assign \new_[98657]_  = ~A202 & ~A201;
  assign \new_[98658]_  = \new_[98657]_  & \new_[98654]_ ;
  assign \new_[98659]_  = \new_[98658]_  & \new_[98651]_ ;
  assign \new_[98662]_  = ~A265 & ~A203;
  assign \new_[98665]_  = ~A267 & A266;
  assign \new_[98666]_  = \new_[98665]_  & \new_[98662]_ ;
  assign \new_[98669]_  = ~A269 & ~A268;
  assign \new_[98673]_  = ~A302 & ~A301;
  assign \new_[98674]_  = A300 & \new_[98673]_ ;
  assign \new_[98675]_  = \new_[98674]_  & \new_[98669]_ ;
  assign \new_[98676]_  = \new_[98675]_  & \new_[98666]_ ;
  assign \new_[98679]_  = A168 & A169;
  assign \new_[98682]_  = ~A166 & A167;
  assign \new_[98683]_  = \new_[98682]_  & \new_[98679]_ ;
  assign \new_[98686]_  = A200 & ~A199;
  assign \new_[98689]_  = ~A202 & ~A201;
  assign \new_[98690]_  = \new_[98689]_  & \new_[98686]_ ;
  assign \new_[98691]_  = \new_[98690]_  & \new_[98683]_ ;
  assign \new_[98694]_  = A265 & ~A203;
  assign \new_[98697]_  = ~A267 & ~A266;
  assign \new_[98698]_  = \new_[98697]_  & \new_[98694]_ ;
  assign \new_[98701]_  = ~A269 & ~A268;
  assign \new_[98705]_  = ~A302 & ~A301;
  assign \new_[98706]_  = A300 & \new_[98705]_ ;
  assign \new_[98707]_  = \new_[98706]_  & \new_[98701]_ ;
  assign \new_[98708]_  = \new_[98707]_  & \new_[98698]_ ;
  assign \new_[98711]_  = A168 & A169;
  assign \new_[98714]_  = ~A166 & A167;
  assign \new_[98715]_  = \new_[98714]_  & \new_[98711]_ ;
  assign \new_[98718]_  = ~A200 & A199;
  assign \new_[98721]_  = ~A202 & ~A201;
  assign \new_[98722]_  = \new_[98721]_  & \new_[98718]_ ;
  assign \new_[98723]_  = \new_[98722]_  & \new_[98715]_ ;
  assign \new_[98726]_  = ~A265 & ~A203;
  assign \new_[98729]_  = ~A267 & A266;
  assign \new_[98730]_  = \new_[98729]_  & \new_[98726]_ ;
  assign \new_[98733]_  = ~A269 & ~A268;
  assign \new_[98737]_  = ~A302 & ~A301;
  assign \new_[98738]_  = A300 & \new_[98737]_ ;
  assign \new_[98739]_  = \new_[98738]_  & \new_[98733]_ ;
  assign \new_[98740]_  = \new_[98739]_  & \new_[98730]_ ;
  assign \new_[98743]_  = A168 & A169;
  assign \new_[98746]_  = ~A166 & A167;
  assign \new_[98747]_  = \new_[98746]_  & \new_[98743]_ ;
  assign \new_[98750]_  = ~A200 & A199;
  assign \new_[98753]_  = ~A202 & ~A201;
  assign \new_[98754]_  = \new_[98753]_  & \new_[98750]_ ;
  assign \new_[98755]_  = \new_[98754]_  & \new_[98747]_ ;
  assign \new_[98758]_  = A265 & ~A203;
  assign \new_[98761]_  = ~A267 & ~A266;
  assign \new_[98762]_  = \new_[98761]_  & \new_[98758]_ ;
  assign \new_[98765]_  = ~A269 & ~A268;
  assign \new_[98769]_  = ~A302 & ~A301;
  assign \new_[98770]_  = A300 & \new_[98769]_ ;
  assign \new_[98771]_  = \new_[98770]_  & \new_[98765]_ ;
  assign \new_[98772]_  = \new_[98771]_  & \new_[98762]_ ;
  assign \new_[98775]_  = A168 & A169;
  assign \new_[98778]_  = A166 & ~A167;
  assign \new_[98779]_  = \new_[98778]_  & \new_[98775]_ ;
  assign \new_[98782]_  = A200 & ~A199;
  assign \new_[98785]_  = ~A202 & ~A201;
  assign \new_[98786]_  = \new_[98785]_  & \new_[98782]_ ;
  assign \new_[98787]_  = \new_[98786]_  & \new_[98779]_ ;
  assign \new_[98790]_  = ~A265 & ~A203;
  assign \new_[98793]_  = ~A267 & A266;
  assign \new_[98794]_  = \new_[98793]_  & \new_[98790]_ ;
  assign \new_[98797]_  = ~A269 & ~A268;
  assign \new_[98801]_  = ~A302 & ~A301;
  assign \new_[98802]_  = A300 & \new_[98801]_ ;
  assign \new_[98803]_  = \new_[98802]_  & \new_[98797]_ ;
  assign \new_[98804]_  = \new_[98803]_  & \new_[98794]_ ;
  assign \new_[98807]_  = A168 & A169;
  assign \new_[98810]_  = A166 & ~A167;
  assign \new_[98811]_  = \new_[98810]_  & \new_[98807]_ ;
  assign \new_[98814]_  = A200 & ~A199;
  assign \new_[98817]_  = ~A202 & ~A201;
  assign \new_[98818]_  = \new_[98817]_  & \new_[98814]_ ;
  assign \new_[98819]_  = \new_[98818]_  & \new_[98811]_ ;
  assign \new_[98822]_  = A265 & ~A203;
  assign \new_[98825]_  = ~A267 & ~A266;
  assign \new_[98826]_  = \new_[98825]_  & \new_[98822]_ ;
  assign \new_[98829]_  = ~A269 & ~A268;
  assign \new_[98833]_  = ~A302 & ~A301;
  assign \new_[98834]_  = A300 & \new_[98833]_ ;
  assign \new_[98835]_  = \new_[98834]_  & \new_[98829]_ ;
  assign \new_[98836]_  = \new_[98835]_  & \new_[98826]_ ;
  assign \new_[98839]_  = A168 & A169;
  assign \new_[98842]_  = A166 & ~A167;
  assign \new_[98843]_  = \new_[98842]_  & \new_[98839]_ ;
  assign \new_[98846]_  = ~A200 & A199;
  assign \new_[98849]_  = ~A202 & ~A201;
  assign \new_[98850]_  = \new_[98849]_  & \new_[98846]_ ;
  assign \new_[98851]_  = \new_[98850]_  & \new_[98843]_ ;
  assign \new_[98854]_  = ~A265 & ~A203;
  assign \new_[98857]_  = ~A267 & A266;
  assign \new_[98858]_  = \new_[98857]_  & \new_[98854]_ ;
  assign \new_[98861]_  = ~A269 & ~A268;
  assign \new_[98865]_  = ~A302 & ~A301;
  assign \new_[98866]_  = A300 & \new_[98865]_ ;
  assign \new_[98867]_  = \new_[98866]_  & \new_[98861]_ ;
  assign \new_[98868]_  = \new_[98867]_  & \new_[98858]_ ;
  assign \new_[98871]_  = A168 & A169;
  assign \new_[98874]_  = A166 & ~A167;
  assign \new_[98875]_  = \new_[98874]_  & \new_[98871]_ ;
  assign \new_[98878]_  = ~A200 & A199;
  assign \new_[98881]_  = ~A202 & ~A201;
  assign \new_[98882]_  = \new_[98881]_  & \new_[98878]_ ;
  assign \new_[98883]_  = \new_[98882]_  & \new_[98875]_ ;
  assign \new_[98886]_  = A265 & ~A203;
  assign \new_[98889]_  = ~A267 & ~A266;
  assign \new_[98890]_  = \new_[98889]_  & \new_[98886]_ ;
  assign \new_[98893]_  = ~A269 & ~A268;
  assign \new_[98897]_  = ~A302 & ~A301;
  assign \new_[98898]_  = A300 & \new_[98897]_ ;
  assign \new_[98899]_  = \new_[98898]_  & \new_[98893]_ ;
  assign \new_[98900]_  = \new_[98899]_  & \new_[98890]_ ;
  assign \new_[98903]_  = ~A169 & A170;
  assign \new_[98906]_  = A167 & ~A168;
  assign \new_[98907]_  = \new_[98906]_  & \new_[98903]_ ;
  assign \new_[98910]_  = ~A199 & ~A166;
  assign \new_[98913]_  = A201 & A200;
  assign \new_[98914]_  = \new_[98913]_  & \new_[98910]_ ;
  assign \new_[98915]_  = \new_[98914]_  & \new_[98907]_ ;
  assign \new_[98918]_  = ~A265 & A202;
  assign \new_[98921]_  = ~A267 & A266;
  assign \new_[98922]_  = \new_[98921]_  & \new_[98918]_ ;
  assign \new_[98925]_  = ~A269 & ~A268;
  assign \new_[98929]_  = ~A302 & ~A301;
  assign \new_[98930]_  = A300 & \new_[98929]_ ;
  assign \new_[98931]_  = \new_[98930]_  & \new_[98925]_ ;
  assign \new_[98932]_  = \new_[98931]_  & \new_[98922]_ ;
  assign \new_[98935]_  = ~A169 & A170;
  assign \new_[98938]_  = A167 & ~A168;
  assign \new_[98939]_  = \new_[98938]_  & \new_[98935]_ ;
  assign \new_[98942]_  = ~A199 & ~A166;
  assign \new_[98945]_  = A201 & A200;
  assign \new_[98946]_  = \new_[98945]_  & \new_[98942]_ ;
  assign \new_[98947]_  = \new_[98946]_  & \new_[98939]_ ;
  assign \new_[98950]_  = A265 & A202;
  assign \new_[98953]_  = ~A267 & ~A266;
  assign \new_[98954]_  = \new_[98953]_  & \new_[98950]_ ;
  assign \new_[98957]_  = ~A269 & ~A268;
  assign \new_[98961]_  = ~A302 & ~A301;
  assign \new_[98962]_  = A300 & \new_[98961]_ ;
  assign \new_[98963]_  = \new_[98962]_  & \new_[98957]_ ;
  assign \new_[98964]_  = \new_[98963]_  & \new_[98954]_ ;
  assign \new_[98967]_  = ~A169 & A170;
  assign \new_[98970]_  = A167 & ~A168;
  assign \new_[98971]_  = \new_[98970]_  & \new_[98967]_ ;
  assign \new_[98974]_  = ~A199 & ~A166;
  assign \new_[98977]_  = A201 & A200;
  assign \new_[98978]_  = \new_[98977]_  & \new_[98974]_ ;
  assign \new_[98979]_  = \new_[98978]_  & \new_[98971]_ ;
  assign \new_[98982]_  = ~A265 & A203;
  assign \new_[98985]_  = ~A267 & A266;
  assign \new_[98986]_  = \new_[98985]_  & \new_[98982]_ ;
  assign \new_[98989]_  = ~A269 & ~A268;
  assign \new_[98993]_  = ~A302 & ~A301;
  assign \new_[98994]_  = A300 & \new_[98993]_ ;
  assign \new_[98995]_  = \new_[98994]_  & \new_[98989]_ ;
  assign \new_[98996]_  = \new_[98995]_  & \new_[98986]_ ;
  assign \new_[98999]_  = ~A169 & A170;
  assign \new_[99002]_  = A167 & ~A168;
  assign \new_[99003]_  = \new_[99002]_  & \new_[98999]_ ;
  assign \new_[99006]_  = ~A199 & ~A166;
  assign \new_[99009]_  = A201 & A200;
  assign \new_[99010]_  = \new_[99009]_  & \new_[99006]_ ;
  assign \new_[99011]_  = \new_[99010]_  & \new_[99003]_ ;
  assign \new_[99014]_  = A265 & A203;
  assign \new_[99017]_  = ~A267 & ~A266;
  assign \new_[99018]_  = \new_[99017]_  & \new_[99014]_ ;
  assign \new_[99021]_  = ~A269 & ~A268;
  assign \new_[99025]_  = ~A302 & ~A301;
  assign \new_[99026]_  = A300 & \new_[99025]_ ;
  assign \new_[99027]_  = \new_[99026]_  & \new_[99021]_ ;
  assign \new_[99028]_  = \new_[99027]_  & \new_[99018]_ ;
  assign \new_[99031]_  = ~A169 & A170;
  assign \new_[99034]_  = A167 & ~A168;
  assign \new_[99035]_  = \new_[99034]_  & \new_[99031]_ ;
  assign \new_[99038]_  = ~A199 & ~A166;
  assign \new_[99041]_  = ~A201 & A200;
  assign \new_[99042]_  = \new_[99041]_  & \new_[99038]_ ;
  assign \new_[99043]_  = \new_[99042]_  & \new_[99035]_ ;
  assign \new_[99046]_  = ~A203 & ~A202;
  assign \new_[99049]_  = A266 & ~A265;
  assign \new_[99050]_  = \new_[99049]_  & \new_[99046]_ ;
  assign \new_[99053]_  = A268 & A267;
  assign \new_[99057]_  = ~A302 & ~A301;
  assign \new_[99058]_  = A300 & \new_[99057]_ ;
  assign \new_[99059]_  = \new_[99058]_  & \new_[99053]_ ;
  assign \new_[99060]_  = \new_[99059]_  & \new_[99050]_ ;
  assign \new_[99063]_  = ~A169 & A170;
  assign \new_[99066]_  = A167 & ~A168;
  assign \new_[99067]_  = \new_[99066]_  & \new_[99063]_ ;
  assign \new_[99070]_  = ~A199 & ~A166;
  assign \new_[99073]_  = ~A201 & A200;
  assign \new_[99074]_  = \new_[99073]_  & \new_[99070]_ ;
  assign \new_[99075]_  = \new_[99074]_  & \new_[99067]_ ;
  assign \new_[99078]_  = ~A203 & ~A202;
  assign \new_[99081]_  = A266 & ~A265;
  assign \new_[99082]_  = \new_[99081]_  & \new_[99078]_ ;
  assign \new_[99085]_  = A269 & A267;
  assign \new_[99089]_  = ~A302 & ~A301;
  assign \new_[99090]_  = A300 & \new_[99089]_ ;
  assign \new_[99091]_  = \new_[99090]_  & \new_[99085]_ ;
  assign \new_[99092]_  = \new_[99091]_  & \new_[99082]_ ;
  assign \new_[99095]_  = ~A169 & A170;
  assign \new_[99098]_  = A167 & ~A168;
  assign \new_[99099]_  = \new_[99098]_  & \new_[99095]_ ;
  assign \new_[99102]_  = ~A199 & ~A166;
  assign \new_[99105]_  = ~A201 & A200;
  assign \new_[99106]_  = \new_[99105]_  & \new_[99102]_ ;
  assign \new_[99107]_  = \new_[99106]_  & \new_[99099]_ ;
  assign \new_[99110]_  = ~A203 & ~A202;
  assign \new_[99113]_  = A266 & ~A265;
  assign \new_[99114]_  = \new_[99113]_  & \new_[99110]_ ;
  assign \new_[99117]_  = ~A268 & ~A267;
  assign \new_[99121]_  = A301 & ~A300;
  assign \new_[99122]_  = ~A269 & \new_[99121]_ ;
  assign \new_[99123]_  = \new_[99122]_  & \new_[99117]_ ;
  assign \new_[99124]_  = \new_[99123]_  & \new_[99114]_ ;
  assign \new_[99127]_  = ~A169 & A170;
  assign \new_[99130]_  = A167 & ~A168;
  assign \new_[99131]_  = \new_[99130]_  & \new_[99127]_ ;
  assign \new_[99134]_  = ~A199 & ~A166;
  assign \new_[99137]_  = ~A201 & A200;
  assign \new_[99138]_  = \new_[99137]_  & \new_[99134]_ ;
  assign \new_[99139]_  = \new_[99138]_  & \new_[99131]_ ;
  assign \new_[99142]_  = ~A203 & ~A202;
  assign \new_[99145]_  = A266 & ~A265;
  assign \new_[99146]_  = \new_[99145]_  & \new_[99142]_ ;
  assign \new_[99149]_  = ~A268 & ~A267;
  assign \new_[99153]_  = A302 & ~A300;
  assign \new_[99154]_  = ~A269 & \new_[99153]_ ;
  assign \new_[99155]_  = \new_[99154]_  & \new_[99149]_ ;
  assign \new_[99156]_  = \new_[99155]_  & \new_[99146]_ ;
  assign \new_[99159]_  = ~A169 & A170;
  assign \new_[99162]_  = A167 & ~A168;
  assign \new_[99163]_  = \new_[99162]_  & \new_[99159]_ ;
  assign \new_[99166]_  = ~A199 & ~A166;
  assign \new_[99169]_  = ~A201 & A200;
  assign \new_[99170]_  = \new_[99169]_  & \new_[99166]_ ;
  assign \new_[99171]_  = \new_[99170]_  & \new_[99163]_ ;
  assign \new_[99174]_  = ~A203 & ~A202;
  assign \new_[99177]_  = A266 & ~A265;
  assign \new_[99178]_  = \new_[99177]_  & \new_[99174]_ ;
  assign \new_[99181]_  = ~A268 & ~A267;
  assign \new_[99185]_  = A299 & A298;
  assign \new_[99186]_  = ~A269 & \new_[99185]_ ;
  assign \new_[99187]_  = \new_[99186]_  & \new_[99181]_ ;
  assign \new_[99188]_  = \new_[99187]_  & \new_[99178]_ ;
  assign \new_[99191]_  = ~A169 & A170;
  assign \new_[99194]_  = A167 & ~A168;
  assign \new_[99195]_  = \new_[99194]_  & \new_[99191]_ ;
  assign \new_[99198]_  = ~A199 & ~A166;
  assign \new_[99201]_  = ~A201 & A200;
  assign \new_[99202]_  = \new_[99201]_  & \new_[99198]_ ;
  assign \new_[99203]_  = \new_[99202]_  & \new_[99195]_ ;
  assign \new_[99206]_  = ~A203 & ~A202;
  assign \new_[99209]_  = A266 & ~A265;
  assign \new_[99210]_  = \new_[99209]_  & \new_[99206]_ ;
  assign \new_[99213]_  = ~A268 & ~A267;
  assign \new_[99217]_  = ~A299 & ~A298;
  assign \new_[99218]_  = ~A269 & \new_[99217]_ ;
  assign \new_[99219]_  = \new_[99218]_  & \new_[99213]_ ;
  assign \new_[99220]_  = \new_[99219]_  & \new_[99210]_ ;
  assign \new_[99223]_  = ~A169 & A170;
  assign \new_[99226]_  = A167 & ~A168;
  assign \new_[99227]_  = \new_[99226]_  & \new_[99223]_ ;
  assign \new_[99230]_  = ~A199 & ~A166;
  assign \new_[99233]_  = ~A201 & A200;
  assign \new_[99234]_  = \new_[99233]_  & \new_[99230]_ ;
  assign \new_[99235]_  = \new_[99234]_  & \new_[99227]_ ;
  assign \new_[99238]_  = ~A203 & ~A202;
  assign \new_[99241]_  = ~A266 & A265;
  assign \new_[99242]_  = \new_[99241]_  & \new_[99238]_ ;
  assign \new_[99245]_  = A268 & A267;
  assign \new_[99249]_  = ~A302 & ~A301;
  assign \new_[99250]_  = A300 & \new_[99249]_ ;
  assign \new_[99251]_  = \new_[99250]_  & \new_[99245]_ ;
  assign \new_[99252]_  = \new_[99251]_  & \new_[99242]_ ;
  assign \new_[99255]_  = ~A169 & A170;
  assign \new_[99258]_  = A167 & ~A168;
  assign \new_[99259]_  = \new_[99258]_  & \new_[99255]_ ;
  assign \new_[99262]_  = ~A199 & ~A166;
  assign \new_[99265]_  = ~A201 & A200;
  assign \new_[99266]_  = \new_[99265]_  & \new_[99262]_ ;
  assign \new_[99267]_  = \new_[99266]_  & \new_[99259]_ ;
  assign \new_[99270]_  = ~A203 & ~A202;
  assign \new_[99273]_  = ~A266 & A265;
  assign \new_[99274]_  = \new_[99273]_  & \new_[99270]_ ;
  assign \new_[99277]_  = A269 & A267;
  assign \new_[99281]_  = ~A302 & ~A301;
  assign \new_[99282]_  = A300 & \new_[99281]_ ;
  assign \new_[99283]_  = \new_[99282]_  & \new_[99277]_ ;
  assign \new_[99284]_  = \new_[99283]_  & \new_[99274]_ ;
  assign \new_[99287]_  = ~A169 & A170;
  assign \new_[99290]_  = A167 & ~A168;
  assign \new_[99291]_  = \new_[99290]_  & \new_[99287]_ ;
  assign \new_[99294]_  = ~A199 & ~A166;
  assign \new_[99297]_  = ~A201 & A200;
  assign \new_[99298]_  = \new_[99297]_  & \new_[99294]_ ;
  assign \new_[99299]_  = \new_[99298]_  & \new_[99291]_ ;
  assign \new_[99302]_  = ~A203 & ~A202;
  assign \new_[99305]_  = ~A266 & A265;
  assign \new_[99306]_  = \new_[99305]_  & \new_[99302]_ ;
  assign \new_[99309]_  = ~A268 & ~A267;
  assign \new_[99313]_  = A301 & ~A300;
  assign \new_[99314]_  = ~A269 & \new_[99313]_ ;
  assign \new_[99315]_  = \new_[99314]_  & \new_[99309]_ ;
  assign \new_[99316]_  = \new_[99315]_  & \new_[99306]_ ;
  assign \new_[99319]_  = ~A169 & A170;
  assign \new_[99322]_  = A167 & ~A168;
  assign \new_[99323]_  = \new_[99322]_  & \new_[99319]_ ;
  assign \new_[99326]_  = ~A199 & ~A166;
  assign \new_[99329]_  = ~A201 & A200;
  assign \new_[99330]_  = \new_[99329]_  & \new_[99326]_ ;
  assign \new_[99331]_  = \new_[99330]_  & \new_[99323]_ ;
  assign \new_[99334]_  = ~A203 & ~A202;
  assign \new_[99337]_  = ~A266 & A265;
  assign \new_[99338]_  = \new_[99337]_  & \new_[99334]_ ;
  assign \new_[99341]_  = ~A268 & ~A267;
  assign \new_[99345]_  = A302 & ~A300;
  assign \new_[99346]_  = ~A269 & \new_[99345]_ ;
  assign \new_[99347]_  = \new_[99346]_  & \new_[99341]_ ;
  assign \new_[99348]_  = \new_[99347]_  & \new_[99338]_ ;
  assign \new_[99351]_  = ~A169 & A170;
  assign \new_[99354]_  = A167 & ~A168;
  assign \new_[99355]_  = \new_[99354]_  & \new_[99351]_ ;
  assign \new_[99358]_  = ~A199 & ~A166;
  assign \new_[99361]_  = ~A201 & A200;
  assign \new_[99362]_  = \new_[99361]_  & \new_[99358]_ ;
  assign \new_[99363]_  = \new_[99362]_  & \new_[99355]_ ;
  assign \new_[99366]_  = ~A203 & ~A202;
  assign \new_[99369]_  = ~A266 & A265;
  assign \new_[99370]_  = \new_[99369]_  & \new_[99366]_ ;
  assign \new_[99373]_  = ~A268 & ~A267;
  assign \new_[99377]_  = A299 & A298;
  assign \new_[99378]_  = ~A269 & \new_[99377]_ ;
  assign \new_[99379]_  = \new_[99378]_  & \new_[99373]_ ;
  assign \new_[99380]_  = \new_[99379]_  & \new_[99370]_ ;
  assign \new_[99383]_  = ~A169 & A170;
  assign \new_[99386]_  = A167 & ~A168;
  assign \new_[99387]_  = \new_[99386]_  & \new_[99383]_ ;
  assign \new_[99390]_  = ~A199 & ~A166;
  assign \new_[99393]_  = ~A201 & A200;
  assign \new_[99394]_  = \new_[99393]_  & \new_[99390]_ ;
  assign \new_[99395]_  = \new_[99394]_  & \new_[99387]_ ;
  assign \new_[99398]_  = ~A203 & ~A202;
  assign \new_[99401]_  = ~A266 & A265;
  assign \new_[99402]_  = \new_[99401]_  & \new_[99398]_ ;
  assign \new_[99405]_  = ~A268 & ~A267;
  assign \new_[99409]_  = ~A299 & ~A298;
  assign \new_[99410]_  = ~A269 & \new_[99409]_ ;
  assign \new_[99411]_  = \new_[99410]_  & \new_[99405]_ ;
  assign \new_[99412]_  = \new_[99411]_  & \new_[99402]_ ;
  assign \new_[99415]_  = ~A169 & A170;
  assign \new_[99418]_  = A167 & ~A168;
  assign \new_[99419]_  = \new_[99418]_  & \new_[99415]_ ;
  assign \new_[99422]_  = A199 & ~A166;
  assign \new_[99425]_  = A201 & ~A200;
  assign \new_[99426]_  = \new_[99425]_  & \new_[99422]_ ;
  assign \new_[99427]_  = \new_[99426]_  & \new_[99419]_ ;
  assign \new_[99430]_  = ~A265 & A202;
  assign \new_[99433]_  = ~A267 & A266;
  assign \new_[99434]_  = \new_[99433]_  & \new_[99430]_ ;
  assign \new_[99437]_  = ~A269 & ~A268;
  assign \new_[99441]_  = ~A302 & ~A301;
  assign \new_[99442]_  = A300 & \new_[99441]_ ;
  assign \new_[99443]_  = \new_[99442]_  & \new_[99437]_ ;
  assign \new_[99444]_  = \new_[99443]_  & \new_[99434]_ ;
  assign \new_[99447]_  = ~A169 & A170;
  assign \new_[99450]_  = A167 & ~A168;
  assign \new_[99451]_  = \new_[99450]_  & \new_[99447]_ ;
  assign \new_[99454]_  = A199 & ~A166;
  assign \new_[99457]_  = A201 & ~A200;
  assign \new_[99458]_  = \new_[99457]_  & \new_[99454]_ ;
  assign \new_[99459]_  = \new_[99458]_  & \new_[99451]_ ;
  assign \new_[99462]_  = A265 & A202;
  assign \new_[99465]_  = ~A267 & ~A266;
  assign \new_[99466]_  = \new_[99465]_  & \new_[99462]_ ;
  assign \new_[99469]_  = ~A269 & ~A268;
  assign \new_[99473]_  = ~A302 & ~A301;
  assign \new_[99474]_  = A300 & \new_[99473]_ ;
  assign \new_[99475]_  = \new_[99474]_  & \new_[99469]_ ;
  assign \new_[99476]_  = \new_[99475]_  & \new_[99466]_ ;
  assign \new_[99479]_  = ~A169 & A170;
  assign \new_[99482]_  = A167 & ~A168;
  assign \new_[99483]_  = \new_[99482]_  & \new_[99479]_ ;
  assign \new_[99486]_  = A199 & ~A166;
  assign \new_[99489]_  = A201 & ~A200;
  assign \new_[99490]_  = \new_[99489]_  & \new_[99486]_ ;
  assign \new_[99491]_  = \new_[99490]_  & \new_[99483]_ ;
  assign \new_[99494]_  = ~A265 & A203;
  assign \new_[99497]_  = ~A267 & A266;
  assign \new_[99498]_  = \new_[99497]_  & \new_[99494]_ ;
  assign \new_[99501]_  = ~A269 & ~A268;
  assign \new_[99505]_  = ~A302 & ~A301;
  assign \new_[99506]_  = A300 & \new_[99505]_ ;
  assign \new_[99507]_  = \new_[99506]_  & \new_[99501]_ ;
  assign \new_[99508]_  = \new_[99507]_  & \new_[99498]_ ;
  assign \new_[99511]_  = ~A169 & A170;
  assign \new_[99514]_  = A167 & ~A168;
  assign \new_[99515]_  = \new_[99514]_  & \new_[99511]_ ;
  assign \new_[99518]_  = A199 & ~A166;
  assign \new_[99521]_  = A201 & ~A200;
  assign \new_[99522]_  = \new_[99521]_  & \new_[99518]_ ;
  assign \new_[99523]_  = \new_[99522]_  & \new_[99515]_ ;
  assign \new_[99526]_  = A265 & A203;
  assign \new_[99529]_  = ~A267 & ~A266;
  assign \new_[99530]_  = \new_[99529]_  & \new_[99526]_ ;
  assign \new_[99533]_  = ~A269 & ~A268;
  assign \new_[99537]_  = ~A302 & ~A301;
  assign \new_[99538]_  = A300 & \new_[99537]_ ;
  assign \new_[99539]_  = \new_[99538]_  & \new_[99533]_ ;
  assign \new_[99540]_  = \new_[99539]_  & \new_[99530]_ ;
  assign \new_[99543]_  = ~A169 & A170;
  assign \new_[99546]_  = A167 & ~A168;
  assign \new_[99547]_  = \new_[99546]_  & \new_[99543]_ ;
  assign \new_[99550]_  = A199 & ~A166;
  assign \new_[99553]_  = ~A201 & ~A200;
  assign \new_[99554]_  = \new_[99553]_  & \new_[99550]_ ;
  assign \new_[99555]_  = \new_[99554]_  & \new_[99547]_ ;
  assign \new_[99558]_  = ~A203 & ~A202;
  assign \new_[99561]_  = A266 & ~A265;
  assign \new_[99562]_  = \new_[99561]_  & \new_[99558]_ ;
  assign \new_[99565]_  = A268 & A267;
  assign \new_[99569]_  = ~A302 & ~A301;
  assign \new_[99570]_  = A300 & \new_[99569]_ ;
  assign \new_[99571]_  = \new_[99570]_  & \new_[99565]_ ;
  assign \new_[99572]_  = \new_[99571]_  & \new_[99562]_ ;
  assign \new_[99575]_  = ~A169 & A170;
  assign \new_[99578]_  = A167 & ~A168;
  assign \new_[99579]_  = \new_[99578]_  & \new_[99575]_ ;
  assign \new_[99582]_  = A199 & ~A166;
  assign \new_[99585]_  = ~A201 & ~A200;
  assign \new_[99586]_  = \new_[99585]_  & \new_[99582]_ ;
  assign \new_[99587]_  = \new_[99586]_  & \new_[99579]_ ;
  assign \new_[99590]_  = ~A203 & ~A202;
  assign \new_[99593]_  = A266 & ~A265;
  assign \new_[99594]_  = \new_[99593]_  & \new_[99590]_ ;
  assign \new_[99597]_  = A269 & A267;
  assign \new_[99601]_  = ~A302 & ~A301;
  assign \new_[99602]_  = A300 & \new_[99601]_ ;
  assign \new_[99603]_  = \new_[99602]_  & \new_[99597]_ ;
  assign \new_[99604]_  = \new_[99603]_  & \new_[99594]_ ;
  assign \new_[99607]_  = ~A169 & A170;
  assign \new_[99610]_  = A167 & ~A168;
  assign \new_[99611]_  = \new_[99610]_  & \new_[99607]_ ;
  assign \new_[99614]_  = A199 & ~A166;
  assign \new_[99617]_  = ~A201 & ~A200;
  assign \new_[99618]_  = \new_[99617]_  & \new_[99614]_ ;
  assign \new_[99619]_  = \new_[99618]_  & \new_[99611]_ ;
  assign \new_[99622]_  = ~A203 & ~A202;
  assign \new_[99625]_  = A266 & ~A265;
  assign \new_[99626]_  = \new_[99625]_  & \new_[99622]_ ;
  assign \new_[99629]_  = ~A268 & ~A267;
  assign \new_[99633]_  = A301 & ~A300;
  assign \new_[99634]_  = ~A269 & \new_[99633]_ ;
  assign \new_[99635]_  = \new_[99634]_  & \new_[99629]_ ;
  assign \new_[99636]_  = \new_[99635]_  & \new_[99626]_ ;
  assign \new_[99639]_  = ~A169 & A170;
  assign \new_[99642]_  = A167 & ~A168;
  assign \new_[99643]_  = \new_[99642]_  & \new_[99639]_ ;
  assign \new_[99646]_  = A199 & ~A166;
  assign \new_[99649]_  = ~A201 & ~A200;
  assign \new_[99650]_  = \new_[99649]_  & \new_[99646]_ ;
  assign \new_[99651]_  = \new_[99650]_  & \new_[99643]_ ;
  assign \new_[99654]_  = ~A203 & ~A202;
  assign \new_[99657]_  = A266 & ~A265;
  assign \new_[99658]_  = \new_[99657]_  & \new_[99654]_ ;
  assign \new_[99661]_  = ~A268 & ~A267;
  assign \new_[99665]_  = A302 & ~A300;
  assign \new_[99666]_  = ~A269 & \new_[99665]_ ;
  assign \new_[99667]_  = \new_[99666]_  & \new_[99661]_ ;
  assign \new_[99668]_  = \new_[99667]_  & \new_[99658]_ ;
  assign \new_[99671]_  = ~A169 & A170;
  assign \new_[99674]_  = A167 & ~A168;
  assign \new_[99675]_  = \new_[99674]_  & \new_[99671]_ ;
  assign \new_[99678]_  = A199 & ~A166;
  assign \new_[99681]_  = ~A201 & ~A200;
  assign \new_[99682]_  = \new_[99681]_  & \new_[99678]_ ;
  assign \new_[99683]_  = \new_[99682]_  & \new_[99675]_ ;
  assign \new_[99686]_  = ~A203 & ~A202;
  assign \new_[99689]_  = A266 & ~A265;
  assign \new_[99690]_  = \new_[99689]_  & \new_[99686]_ ;
  assign \new_[99693]_  = ~A268 & ~A267;
  assign \new_[99697]_  = A299 & A298;
  assign \new_[99698]_  = ~A269 & \new_[99697]_ ;
  assign \new_[99699]_  = \new_[99698]_  & \new_[99693]_ ;
  assign \new_[99700]_  = \new_[99699]_  & \new_[99690]_ ;
  assign \new_[99703]_  = ~A169 & A170;
  assign \new_[99706]_  = A167 & ~A168;
  assign \new_[99707]_  = \new_[99706]_  & \new_[99703]_ ;
  assign \new_[99710]_  = A199 & ~A166;
  assign \new_[99713]_  = ~A201 & ~A200;
  assign \new_[99714]_  = \new_[99713]_  & \new_[99710]_ ;
  assign \new_[99715]_  = \new_[99714]_  & \new_[99707]_ ;
  assign \new_[99718]_  = ~A203 & ~A202;
  assign \new_[99721]_  = A266 & ~A265;
  assign \new_[99722]_  = \new_[99721]_  & \new_[99718]_ ;
  assign \new_[99725]_  = ~A268 & ~A267;
  assign \new_[99729]_  = ~A299 & ~A298;
  assign \new_[99730]_  = ~A269 & \new_[99729]_ ;
  assign \new_[99731]_  = \new_[99730]_  & \new_[99725]_ ;
  assign \new_[99732]_  = \new_[99731]_  & \new_[99722]_ ;
  assign \new_[99735]_  = ~A169 & A170;
  assign \new_[99738]_  = A167 & ~A168;
  assign \new_[99739]_  = \new_[99738]_  & \new_[99735]_ ;
  assign \new_[99742]_  = A199 & ~A166;
  assign \new_[99745]_  = ~A201 & ~A200;
  assign \new_[99746]_  = \new_[99745]_  & \new_[99742]_ ;
  assign \new_[99747]_  = \new_[99746]_  & \new_[99739]_ ;
  assign \new_[99750]_  = ~A203 & ~A202;
  assign \new_[99753]_  = ~A266 & A265;
  assign \new_[99754]_  = \new_[99753]_  & \new_[99750]_ ;
  assign \new_[99757]_  = A268 & A267;
  assign \new_[99761]_  = ~A302 & ~A301;
  assign \new_[99762]_  = A300 & \new_[99761]_ ;
  assign \new_[99763]_  = \new_[99762]_  & \new_[99757]_ ;
  assign \new_[99764]_  = \new_[99763]_  & \new_[99754]_ ;
  assign \new_[99767]_  = ~A169 & A170;
  assign \new_[99770]_  = A167 & ~A168;
  assign \new_[99771]_  = \new_[99770]_  & \new_[99767]_ ;
  assign \new_[99774]_  = A199 & ~A166;
  assign \new_[99777]_  = ~A201 & ~A200;
  assign \new_[99778]_  = \new_[99777]_  & \new_[99774]_ ;
  assign \new_[99779]_  = \new_[99778]_  & \new_[99771]_ ;
  assign \new_[99782]_  = ~A203 & ~A202;
  assign \new_[99785]_  = ~A266 & A265;
  assign \new_[99786]_  = \new_[99785]_  & \new_[99782]_ ;
  assign \new_[99789]_  = A269 & A267;
  assign \new_[99793]_  = ~A302 & ~A301;
  assign \new_[99794]_  = A300 & \new_[99793]_ ;
  assign \new_[99795]_  = \new_[99794]_  & \new_[99789]_ ;
  assign \new_[99796]_  = \new_[99795]_  & \new_[99786]_ ;
  assign \new_[99799]_  = ~A169 & A170;
  assign \new_[99802]_  = A167 & ~A168;
  assign \new_[99803]_  = \new_[99802]_  & \new_[99799]_ ;
  assign \new_[99806]_  = A199 & ~A166;
  assign \new_[99809]_  = ~A201 & ~A200;
  assign \new_[99810]_  = \new_[99809]_  & \new_[99806]_ ;
  assign \new_[99811]_  = \new_[99810]_  & \new_[99803]_ ;
  assign \new_[99814]_  = ~A203 & ~A202;
  assign \new_[99817]_  = ~A266 & A265;
  assign \new_[99818]_  = \new_[99817]_  & \new_[99814]_ ;
  assign \new_[99821]_  = ~A268 & ~A267;
  assign \new_[99825]_  = A301 & ~A300;
  assign \new_[99826]_  = ~A269 & \new_[99825]_ ;
  assign \new_[99827]_  = \new_[99826]_  & \new_[99821]_ ;
  assign \new_[99828]_  = \new_[99827]_  & \new_[99818]_ ;
  assign \new_[99831]_  = ~A169 & A170;
  assign \new_[99834]_  = A167 & ~A168;
  assign \new_[99835]_  = \new_[99834]_  & \new_[99831]_ ;
  assign \new_[99838]_  = A199 & ~A166;
  assign \new_[99841]_  = ~A201 & ~A200;
  assign \new_[99842]_  = \new_[99841]_  & \new_[99838]_ ;
  assign \new_[99843]_  = \new_[99842]_  & \new_[99835]_ ;
  assign \new_[99846]_  = ~A203 & ~A202;
  assign \new_[99849]_  = ~A266 & A265;
  assign \new_[99850]_  = \new_[99849]_  & \new_[99846]_ ;
  assign \new_[99853]_  = ~A268 & ~A267;
  assign \new_[99857]_  = A302 & ~A300;
  assign \new_[99858]_  = ~A269 & \new_[99857]_ ;
  assign \new_[99859]_  = \new_[99858]_  & \new_[99853]_ ;
  assign \new_[99860]_  = \new_[99859]_  & \new_[99850]_ ;
  assign \new_[99863]_  = ~A169 & A170;
  assign \new_[99866]_  = A167 & ~A168;
  assign \new_[99867]_  = \new_[99866]_  & \new_[99863]_ ;
  assign \new_[99870]_  = A199 & ~A166;
  assign \new_[99873]_  = ~A201 & ~A200;
  assign \new_[99874]_  = \new_[99873]_  & \new_[99870]_ ;
  assign \new_[99875]_  = \new_[99874]_  & \new_[99867]_ ;
  assign \new_[99878]_  = ~A203 & ~A202;
  assign \new_[99881]_  = ~A266 & A265;
  assign \new_[99882]_  = \new_[99881]_  & \new_[99878]_ ;
  assign \new_[99885]_  = ~A268 & ~A267;
  assign \new_[99889]_  = A299 & A298;
  assign \new_[99890]_  = ~A269 & \new_[99889]_ ;
  assign \new_[99891]_  = \new_[99890]_  & \new_[99885]_ ;
  assign \new_[99892]_  = \new_[99891]_  & \new_[99882]_ ;
  assign \new_[99895]_  = ~A169 & A170;
  assign \new_[99898]_  = A167 & ~A168;
  assign \new_[99899]_  = \new_[99898]_  & \new_[99895]_ ;
  assign \new_[99902]_  = A199 & ~A166;
  assign \new_[99905]_  = ~A201 & ~A200;
  assign \new_[99906]_  = \new_[99905]_  & \new_[99902]_ ;
  assign \new_[99907]_  = \new_[99906]_  & \new_[99899]_ ;
  assign \new_[99910]_  = ~A203 & ~A202;
  assign \new_[99913]_  = ~A266 & A265;
  assign \new_[99914]_  = \new_[99913]_  & \new_[99910]_ ;
  assign \new_[99917]_  = ~A268 & ~A267;
  assign \new_[99921]_  = ~A299 & ~A298;
  assign \new_[99922]_  = ~A269 & \new_[99921]_ ;
  assign \new_[99923]_  = \new_[99922]_  & \new_[99917]_ ;
  assign \new_[99924]_  = \new_[99923]_  & \new_[99914]_ ;
  assign \new_[99927]_  = ~A169 & A170;
  assign \new_[99930]_  = ~A167 & ~A168;
  assign \new_[99931]_  = \new_[99930]_  & \new_[99927]_ ;
  assign \new_[99934]_  = ~A199 & A166;
  assign \new_[99937]_  = A201 & A200;
  assign \new_[99938]_  = \new_[99937]_  & \new_[99934]_ ;
  assign \new_[99939]_  = \new_[99938]_  & \new_[99931]_ ;
  assign \new_[99942]_  = ~A265 & A202;
  assign \new_[99945]_  = ~A267 & A266;
  assign \new_[99946]_  = \new_[99945]_  & \new_[99942]_ ;
  assign \new_[99949]_  = ~A269 & ~A268;
  assign \new_[99953]_  = ~A302 & ~A301;
  assign \new_[99954]_  = A300 & \new_[99953]_ ;
  assign \new_[99955]_  = \new_[99954]_  & \new_[99949]_ ;
  assign \new_[99956]_  = \new_[99955]_  & \new_[99946]_ ;
  assign \new_[99959]_  = ~A169 & A170;
  assign \new_[99962]_  = ~A167 & ~A168;
  assign \new_[99963]_  = \new_[99962]_  & \new_[99959]_ ;
  assign \new_[99966]_  = ~A199 & A166;
  assign \new_[99969]_  = A201 & A200;
  assign \new_[99970]_  = \new_[99969]_  & \new_[99966]_ ;
  assign \new_[99971]_  = \new_[99970]_  & \new_[99963]_ ;
  assign \new_[99974]_  = A265 & A202;
  assign \new_[99977]_  = ~A267 & ~A266;
  assign \new_[99978]_  = \new_[99977]_  & \new_[99974]_ ;
  assign \new_[99981]_  = ~A269 & ~A268;
  assign \new_[99985]_  = ~A302 & ~A301;
  assign \new_[99986]_  = A300 & \new_[99985]_ ;
  assign \new_[99987]_  = \new_[99986]_  & \new_[99981]_ ;
  assign \new_[99988]_  = \new_[99987]_  & \new_[99978]_ ;
  assign \new_[99991]_  = ~A169 & A170;
  assign \new_[99994]_  = ~A167 & ~A168;
  assign \new_[99995]_  = \new_[99994]_  & \new_[99991]_ ;
  assign \new_[99998]_  = ~A199 & A166;
  assign \new_[100001]_  = A201 & A200;
  assign \new_[100002]_  = \new_[100001]_  & \new_[99998]_ ;
  assign \new_[100003]_  = \new_[100002]_  & \new_[99995]_ ;
  assign \new_[100006]_  = ~A265 & A203;
  assign \new_[100009]_  = ~A267 & A266;
  assign \new_[100010]_  = \new_[100009]_  & \new_[100006]_ ;
  assign \new_[100013]_  = ~A269 & ~A268;
  assign \new_[100017]_  = ~A302 & ~A301;
  assign \new_[100018]_  = A300 & \new_[100017]_ ;
  assign \new_[100019]_  = \new_[100018]_  & \new_[100013]_ ;
  assign \new_[100020]_  = \new_[100019]_  & \new_[100010]_ ;
  assign \new_[100023]_  = ~A169 & A170;
  assign \new_[100026]_  = ~A167 & ~A168;
  assign \new_[100027]_  = \new_[100026]_  & \new_[100023]_ ;
  assign \new_[100030]_  = ~A199 & A166;
  assign \new_[100033]_  = A201 & A200;
  assign \new_[100034]_  = \new_[100033]_  & \new_[100030]_ ;
  assign \new_[100035]_  = \new_[100034]_  & \new_[100027]_ ;
  assign \new_[100038]_  = A265 & A203;
  assign \new_[100041]_  = ~A267 & ~A266;
  assign \new_[100042]_  = \new_[100041]_  & \new_[100038]_ ;
  assign \new_[100045]_  = ~A269 & ~A268;
  assign \new_[100049]_  = ~A302 & ~A301;
  assign \new_[100050]_  = A300 & \new_[100049]_ ;
  assign \new_[100051]_  = \new_[100050]_  & \new_[100045]_ ;
  assign \new_[100052]_  = \new_[100051]_  & \new_[100042]_ ;
  assign \new_[100055]_  = ~A169 & A170;
  assign \new_[100058]_  = ~A167 & ~A168;
  assign \new_[100059]_  = \new_[100058]_  & \new_[100055]_ ;
  assign \new_[100062]_  = ~A199 & A166;
  assign \new_[100065]_  = ~A201 & A200;
  assign \new_[100066]_  = \new_[100065]_  & \new_[100062]_ ;
  assign \new_[100067]_  = \new_[100066]_  & \new_[100059]_ ;
  assign \new_[100070]_  = ~A203 & ~A202;
  assign \new_[100073]_  = A266 & ~A265;
  assign \new_[100074]_  = \new_[100073]_  & \new_[100070]_ ;
  assign \new_[100077]_  = A268 & A267;
  assign \new_[100081]_  = ~A302 & ~A301;
  assign \new_[100082]_  = A300 & \new_[100081]_ ;
  assign \new_[100083]_  = \new_[100082]_  & \new_[100077]_ ;
  assign \new_[100084]_  = \new_[100083]_  & \new_[100074]_ ;
  assign \new_[100087]_  = ~A169 & A170;
  assign \new_[100090]_  = ~A167 & ~A168;
  assign \new_[100091]_  = \new_[100090]_  & \new_[100087]_ ;
  assign \new_[100094]_  = ~A199 & A166;
  assign \new_[100097]_  = ~A201 & A200;
  assign \new_[100098]_  = \new_[100097]_  & \new_[100094]_ ;
  assign \new_[100099]_  = \new_[100098]_  & \new_[100091]_ ;
  assign \new_[100102]_  = ~A203 & ~A202;
  assign \new_[100105]_  = A266 & ~A265;
  assign \new_[100106]_  = \new_[100105]_  & \new_[100102]_ ;
  assign \new_[100109]_  = A269 & A267;
  assign \new_[100113]_  = ~A302 & ~A301;
  assign \new_[100114]_  = A300 & \new_[100113]_ ;
  assign \new_[100115]_  = \new_[100114]_  & \new_[100109]_ ;
  assign \new_[100116]_  = \new_[100115]_  & \new_[100106]_ ;
  assign \new_[100119]_  = ~A169 & A170;
  assign \new_[100122]_  = ~A167 & ~A168;
  assign \new_[100123]_  = \new_[100122]_  & \new_[100119]_ ;
  assign \new_[100126]_  = ~A199 & A166;
  assign \new_[100129]_  = ~A201 & A200;
  assign \new_[100130]_  = \new_[100129]_  & \new_[100126]_ ;
  assign \new_[100131]_  = \new_[100130]_  & \new_[100123]_ ;
  assign \new_[100134]_  = ~A203 & ~A202;
  assign \new_[100137]_  = A266 & ~A265;
  assign \new_[100138]_  = \new_[100137]_  & \new_[100134]_ ;
  assign \new_[100141]_  = ~A268 & ~A267;
  assign \new_[100145]_  = A301 & ~A300;
  assign \new_[100146]_  = ~A269 & \new_[100145]_ ;
  assign \new_[100147]_  = \new_[100146]_  & \new_[100141]_ ;
  assign \new_[100148]_  = \new_[100147]_  & \new_[100138]_ ;
  assign \new_[100151]_  = ~A169 & A170;
  assign \new_[100154]_  = ~A167 & ~A168;
  assign \new_[100155]_  = \new_[100154]_  & \new_[100151]_ ;
  assign \new_[100158]_  = ~A199 & A166;
  assign \new_[100161]_  = ~A201 & A200;
  assign \new_[100162]_  = \new_[100161]_  & \new_[100158]_ ;
  assign \new_[100163]_  = \new_[100162]_  & \new_[100155]_ ;
  assign \new_[100166]_  = ~A203 & ~A202;
  assign \new_[100169]_  = A266 & ~A265;
  assign \new_[100170]_  = \new_[100169]_  & \new_[100166]_ ;
  assign \new_[100173]_  = ~A268 & ~A267;
  assign \new_[100177]_  = A302 & ~A300;
  assign \new_[100178]_  = ~A269 & \new_[100177]_ ;
  assign \new_[100179]_  = \new_[100178]_  & \new_[100173]_ ;
  assign \new_[100180]_  = \new_[100179]_  & \new_[100170]_ ;
  assign \new_[100183]_  = ~A169 & A170;
  assign \new_[100186]_  = ~A167 & ~A168;
  assign \new_[100187]_  = \new_[100186]_  & \new_[100183]_ ;
  assign \new_[100190]_  = ~A199 & A166;
  assign \new_[100193]_  = ~A201 & A200;
  assign \new_[100194]_  = \new_[100193]_  & \new_[100190]_ ;
  assign \new_[100195]_  = \new_[100194]_  & \new_[100187]_ ;
  assign \new_[100198]_  = ~A203 & ~A202;
  assign \new_[100201]_  = A266 & ~A265;
  assign \new_[100202]_  = \new_[100201]_  & \new_[100198]_ ;
  assign \new_[100205]_  = ~A268 & ~A267;
  assign \new_[100209]_  = A299 & A298;
  assign \new_[100210]_  = ~A269 & \new_[100209]_ ;
  assign \new_[100211]_  = \new_[100210]_  & \new_[100205]_ ;
  assign \new_[100212]_  = \new_[100211]_  & \new_[100202]_ ;
  assign \new_[100215]_  = ~A169 & A170;
  assign \new_[100218]_  = ~A167 & ~A168;
  assign \new_[100219]_  = \new_[100218]_  & \new_[100215]_ ;
  assign \new_[100222]_  = ~A199 & A166;
  assign \new_[100225]_  = ~A201 & A200;
  assign \new_[100226]_  = \new_[100225]_  & \new_[100222]_ ;
  assign \new_[100227]_  = \new_[100226]_  & \new_[100219]_ ;
  assign \new_[100230]_  = ~A203 & ~A202;
  assign \new_[100233]_  = A266 & ~A265;
  assign \new_[100234]_  = \new_[100233]_  & \new_[100230]_ ;
  assign \new_[100237]_  = ~A268 & ~A267;
  assign \new_[100241]_  = ~A299 & ~A298;
  assign \new_[100242]_  = ~A269 & \new_[100241]_ ;
  assign \new_[100243]_  = \new_[100242]_  & \new_[100237]_ ;
  assign \new_[100244]_  = \new_[100243]_  & \new_[100234]_ ;
  assign \new_[100247]_  = ~A169 & A170;
  assign \new_[100250]_  = ~A167 & ~A168;
  assign \new_[100251]_  = \new_[100250]_  & \new_[100247]_ ;
  assign \new_[100254]_  = ~A199 & A166;
  assign \new_[100257]_  = ~A201 & A200;
  assign \new_[100258]_  = \new_[100257]_  & \new_[100254]_ ;
  assign \new_[100259]_  = \new_[100258]_  & \new_[100251]_ ;
  assign \new_[100262]_  = ~A203 & ~A202;
  assign \new_[100265]_  = ~A266 & A265;
  assign \new_[100266]_  = \new_[100265]_  & \new_[100262]_ ;
  assign \new_[100269]_  = A268 & A267;
  assign \new_[100273]_  = ~A302 & ~A301;
  assign \new_[100274]_  = A300 & \new_[100273]_ ;
  assign \new_[100275]_  = \new_[100274]_  & \new_[100269]_ ;
  assign \new_[100276]_  = \new_[100275]_  & \new_[100266]_ ;
  assign \new_[100279]_  = ~A169 & A170;
  assign \new_[100282]_  = ~A167 & ~A168;
  assign \new_[100283]_  = \new_[100282]_  & \new_[100279]_ ;
  assign \new_[100286]_  = ~A199 & A166;
  assign \new_[100289]_  = ~A201 & A200;
  assign \new_[100290]_  = \new_[100289]_  & \new_[100286]_ ;
  assign \new_[100291]_  = \new_[100290]_  & \new_[100283]_ ;
  assign \new_[100294]_  = ~A203 & ~A202;
  assign \new_[100297]_  = ~A266 & A265;
  assign \new_[100298]_  = \new_[100297]_  & \new_[100294]_ ;
  assign \new_[100301]_  = A269 & A267;
  assign \new_[100305]_  = ~A302 & ~A301;
  assign \new_[100306]_  = A300 & \new_[100305]_ ;
  assign \new_[100307]_  = \new_[100306]_  & \new_[100301]_ ;
  assign \new_[100308]_  = \new_[100307]_  & \new_[100298]_ ;
  assign \new_[100311]_  = ~A169 & A170;
  assign \new_[100314]_  = ~A167 & ~A168;
  assign \new_[100315]_  = \new_[100314]_  & \new_[100311]_ ;
  assign \new_[100318]_  = ~A199 & A166;
  assign \new_[100321]_  = ~A201 & A200;
  assign \new_[100322]_  = \new_[100321]_  & \new_[100318]_ ;
  assign \new_[100323]_  = \new_[100322]_  & \new_[100315]_ ;
  assign \new_[100326]_  = ~A203 & ~A202;
  assign \new_[100329]_  = ~A266 & A265;
  assign \new_[100330]_  = \new_[100329]_  & \new_[100326]_ ;
  assign \new_[100333]_  = ~A268 & ~A267;
  assign \new_[100337]_  = A301 & ~A300;
  assign \new_[100338]_  = ~A269 & \new_[100337]_ ;
  assign \new_[100339]_  = \new_[100338]_  & \new_[100333]_ ;
  assign \new_[100340]_  = \new_[100339]_  & \new_[100330]_ ;
  assign \new_[100343]_  = ~A169 & A170;
  assign \new_[100346]_  = ~A167 & ~A168;
  assign \new_[100347]_  = \new_[100346]_  & \new_[100343]_ ;
  assign \new_[100350]_  = ~A199 & A166;
  assign \new_[100353]_  = ~A201 & A200;
  assign \new_[100354]_  = \new_[100353]_  & \new_[100350]_ ;
  assign \new_[100355]_  = \new_[100354]_  & \new_[100347]_ ;
  assign \new_[100358]_  = ~A203 & ~A202;
  assign \new_[100361]_  = ~A266 & A265;
  assign \new_[100362]_  = \new_[100361]_  & \new_[100358]_ ;
  assign \new_[100365]_  = ~A268 & ~A267;
  assign \new_[100369]_  = A302 & ~A300;
  assign \new_[100370]_  = ~A269 & \new_[100369]_ ;
  assign \new_[100371]_  = \new_[100370]_  & \new_[100365]_ ;
  assign \new_[100372]_  = \new_[100371]_  & \new_[100362]_ ;
  assign \new_[100375]_  = ~A169 & A170;
  assign \new_[100378]_  = ~A167 & ~A168;
  assign \new_[100379]_  = \new_[100378]_  & \new_[100375]_ ;
  assign \new_[100382]_  = ~A199 & A166;
  assign \new_[100385]_  = ~A201 & A200;
  assign \new_[100386]_  = \new_[100385]_  & \new_[100382]_ ;
  assign \new_[100387]_  = \new_[100386]_  & \new_[100379]_ ;
  assign \new_[100390]_  = ~A203 & ~A202;
  assign \new_[100393]_  = ~A266 & A265;
  assign \new_[100394]_  = \new_[100393]_  & \new_[100390]_ ;
  assign \new_[100397]_  = ~A268 & ~A267;
  assign \new_[100401]_  = A299 & A298;
  assign \new_[100402]_  = ~A269 & \new_[100401]_ ;
  assign \new_[100403]_  = \new_[100402]_  & \new_[100397]_ ;
  assign \new_[100404]_  = \new_[100403]_  & \new_[100394]_ ;
  assign \new_[100407]_  = ~A169 & A170;
  assign \new_[100410]_  = ~A167 & ~A168;
  assign \new_[100411]_  = \new_[100410]_  & \new_[100407]_ ;
  assign \new_[100414]_  = ~A199 & A166;
  assign \new_[100417]_  = ~A201 & A200;
  assign \new_[100418]_  = \new_[100417]_  & \new_[100414]_ ;
  assign \new_[100419]_  = \new_[100418]_  & \new_[100411]_ ;
  assign \new_[100422]_  = ~A203 & ~A202;
  assign \new_[100425]_  = ~A266 & A265;
  assign \new_[100426]_  = \new_[100425]_  & \new_[100422]_ ;
  assign \new_[100429]_  = ~A268 & ~A267;
  assign \new_[100433]_  = ~A299 & ~A298;
  assign \new_[100434]_  = ~A269 & \new_[100433]_ ;
  assign \new_[100435]_  = \new_[100434]_  & \new_[100429]_ ;
  assign \new_[100436]_  = \new_[100435]_  & \new_[100426]_ ;
  assign \new_[100439]_  = ~A169 & A170;
  assign \new_[100442]_  = ~A167 & ~A168;
  assign \new_[100443]_  = \new_[100442]_  & \new_[100439]_ ;
  assign \new_[100446]_  = A199 & A166;
  assign \new_[100449]_  = A201 & ~A200;
  assign \new_[100450]_  = \new_[100449]_  & \new_[100446]_ ;
  assign \new_[100451]_  = \new_[100450]_  & \new_[100443]_ ;
  assign \new_[100454]_  = ~A265 & A202;
  assign \new_[100457]_  = ~A267 & A266;
  assign \new_[100458]_  = \new_[100457]_  & \new_[100454]_ ;
  assign \new_[100461]_  = ~A269 & ~A268;
  assign \new_[100465]_  = ~A302 & ~A301;
  assign \new_[100466]_  = A300 & \new_[100465]_ ;
  assign \new_[100467]_  = \new_[100466]_  & \new_[100461]_ ;
  assign \new_[100468]_  = \new_[100467]_  & \new_[100458]_ ;
  assign \new_[100471]_  = ~A169 & A170;
  assign \new_[100474]_  = ~A167 & ~A168;
  assign \new_[100475]_  = \new_[100474]_  & \new_[100471]_ ;
  assign \new_[100478]_  = A199 & A166;
  assign \new_[100481]_  = A201 & ~A200;
  assign \new_[100482]_  = \new_[100481]_  & \new_[100478]_ ;
  assign \new_[100483]_  = \new_[100482]_  & \new_[100475]_ ;
  assign \new_[100486]_  = A265 & A202;
  assign \new_[100489]_  = ~A267 & ~A266;
  assign \new_[100490]_  = \new_[100489]_  & \new_[100486]_ ;
  assign \new_[100493]_  = ~A269 & ~A268;
  assign \new_[100497]_  = ~A302 & ~A301;
  assign \new_[100498]_  = A300 & \new_[100497]_ ;
  assign \new_[100499]_  = \new_[100498]_  & \new_[100493]_ ;
  assign \new_[100500]_  = \new_[100499]_  & \new_[100490]_ ;
  assign \new_[100503]_  = ~A169 & A170;
  assign \new_[100506]_  = ~A167 & ~A168;
  assign \new_[100507]_  = \new_[100506]_  & \new_[100503]_ ;
  assign \new_[100510]_  = A199 & A166;
  assign \new_[100513]_  = A201 & ~A200;
  assign \new_[100514]_  = \new_[100513]_  & \new_[100510]_ ;
  assign \new_[100515]_  = \new_[100514]_  & \new_[100507]_ ;
  assign \new_[100518]_  = ~A265 & A203;
  assign \new_[100521]_  = ~A267 & A266;
  assign \new_[100522]_  = \new_[100521]_  & \new_[100518]_ ;
  assign \new_[100525]_  = ~A269 & ~A268;
  assign \new_[100529]_  = ~A302 & ~A301;
  assign \new_[100530]_  = A300 & \new_[100529]_ ;
  assign \new_[100531]_  = \new_[100530]_  & \new_[100525]_ ;
  assign \new_[100532]_  = \new_[100531]_  & \new_[100522]_ ;
  assign \new_[100535]_  = ~A169 & A170;
  assign \new_[100538]_  = ~A167 & ~A168;
  assign \new_[100539]_  = \new_[100538]_  & \new_[100535]_ ;
  assign \new_[100542]_  = A199 & A166;
  assign \new_[100545]_  = A201 & ~A200;
  assign \new_[100546]_  = \new_[100545]_  & \new_[100542]_ ;
  assign \new_[100547]_  = \new_[100546]_  & \new_[100539]_ ;
  assign \new_[100550]_  = A265 & A203;
  assign \new_[100553]_  = ~A267 & ~A266;
  assign \new_[100554]_  = \new_[100553]_  & \new_[100550]_ ;
  assign \new_[100557]_  = ~A269 & ~A268;
  assign \new_[100561]_  = ~A302 & ~A301;
  assign \new_[100562]_  = A300 & \new_[100561]_ ;
  assign \new_[100563]_  = \new_[100562]_  & \new_[100557]_ ;
  assign \new_[100564]_  = \new_[100563]_  & \new_[100554]_ ;
  assign \new_[100567]_  = ~A169 & A170;
  assign \new_[100570]_  = ~A167 & ~A168;
  assign \new_[100571]_  = \new_[100570]_  & \new_[100567]_ ;
  assign \new_[100574]_  = A199 & A166;
  assign \new_[100577]_  = ~A201 & ~A200;
  assign \new_[100578]_  = \new_[100577]_  & \new_[100574]_ ;
  assign \new_[100579]_  = \new_[100578]_  & \new_[100571]_ ;
  assign \new_[100582]_  = ~A203 & ~A202;
  assign \new_[100585]_  = A266 & ~A265;
  assign \new_[100586]_  = \new_[100585]_  & \new_[100582]_ ;
  assign \new_[100589]_  = A268 & A267;
  assign \new_[100593]_  = ~A302 & ~A301;
  assign \new_[100594]_  = A300 & \new_[100593]_ ;
  assign \new_[100595]_  = \new_[100594]_  & \new_[100589]_ ;
  assign \new_[100596]_  = \new_[100595]_  & \new_[100586]_ ;
  assign \new_[100599]_  = ~A169 & A170;
  assign \new_[100602]_  = ~A167 & ~A168;
  assign \new_[100603]_  = \new_[100602]_  & \new_[100599]_ ;
  assign \new_[100606]_  = A199 & A166;
  assign \new_[100609]_  = ~A201 & ~A200;
  assign \new_[100610]_  = \new_[100609]_  & \new_[100606]_ ;
  assign \new_[100611]_  = \new_[100610]_  & \new_[100603]_ ;
  assign \new_[100614]_  = ~A203 & ~A202;
  assign \new_[100617]_  = A266 & ~A265;
  assign \new_[100618]_  = \new_[100617]_  & \new_[100614]_ ;
  assign \new_[100621]_  = A269 & A267;
  assign \new_[100625]_  = ~A302 & ~A301;
  assign \new_[100626]_  = A300 & \new_[100625]_ ;
  assign \new_[100627]_  = \new_[100626]_  & \new_[100621]_ ;
  assign \new_[100628]_  = \new_[100627]_  & \new_[100618]_ ;
  assign \new_[100631]_  = ~A169 & A170;
  assign \new_[100634]_  = ~A167 & ~A168;
  assign \new_[100635]_  = \new_[100634]_  & \new_[100631]_ ;
  assign \new_[100638]_  = A199 & A166;
  assign \new_[100641]_  = ~A201 & ~A200;
  assign \new_[100642]_  = \new_[100641]_  & \new_[100638]_ ;
  assign \new_[100643]_  = \new_[100642]_  & \new_[100635]_ ;
  assign \new_[100646]_  = ~A203 & ~A202;
  assign \new_[100649]_  = A266 & ~A265;
  assign \new_[100650]_  = \new_[100649]_  & \new_[100646]_ ;
  assign \new_[100653]_  = ~A268 & ~A267;
  assign \new_[100657]_  = A301 & ~A300;
  assign \new_[100658]_  = ~A269 & \new_[100657]_ ;
  assign \new_[100659]_  = \new_[100658]_  & \new_[100653]_ ;
  assign \new_[100660]_  = \new_[100659]_  & \new_[100650]_ ;
  assign \new_[100663]_  = ~A169 & A170;
  assign \new_[100666]_  = ~A167 & ~A168;
  assign \new_[100667]_  = \new_[100666]_  & \new_[100663]_ ;
  assign \new_[100670]_  = A199 & A166;
  assign \new_[100673]_  = ~A201 & ~A200;
  assign \new_[100674]_  = \new_[100673]_  & \new_[100670]_ ;
  assign \new_[100675]_  = \new_[100674]_  & \new_[100667]_ ;
  assign \new_[100678]_  = ~A203 & ~A202;
  assign \new_[100681]_  = A266 & ~A265;
  assign \new_[100682]_  = \new_[100681]_  & \new_[100678]_ ;
  assign \new_[100685]_  = ~A268 & ~A267;
  assign \new_[100689]_  = A302 & ~A300;
  assign \new_[100690]_  = ~A269 & \new_[100689]_ ;
  assign \new_[100691]_  = \new_[100690]_  & \new_[100685]_ ;
  assign \new_[100692]_  = \new_[100691]_  & \new_[100682]_ ;
  assign \new_[100695]_  = ~A169 & A170;
  assign \new_[100698]_  = ~A167 & ~A168;
  assign \new_[100699]_  = \new_[100698]_  & \new_[100695]_ ;
  assign \new_[100702]_  = A199 & A166;
  assign \new_[100705]_  = ~A201 & ~A200;
  assign \new_[100706]_  = \new_[100705]_  & \new_[100702]_ ;
  assign \new_[100707]_  = \new_[100706]_  & \new_[100699]_ ;
  assign \new_[100710]_  = ~A203 & ~A202;
  assign \new_[100713]_  = A266 & ~A265;
  assign \new_[100714]_  = \new_[100713]_  & \new_[100710]_ ;
  assign \new_[100717]_  = ~A268 & ~A267;
  assign \new_[100721]_  = A299 & A298;
  assign \new_[100722]_  = ~A269 & \new_[100721]_ ;
  assign \new_[100723]_  = \new_[100722]_  & \new_[100717]_ ;
  assign \new_[100724]_  = \new_[100723]_  & \new_[100714]_ ;
  assign \new_[100727]_  = ~A169 & A170;
  assign \new_[100730]_  = ~A167 & ~A168;
  assign \new_[100731]_  = \new_[100730]_  & \new_[100727]_ ;
  assign \new_[100734]_  = A199 & A166;
  assign \new_[100737]_  = ~A201 & ~A200;
  assign \new_[100738]_  = \new_[100737]_  & \new_[100734]_ ;
  assign \new_[100739]_  = \new_[100738]_  & \new_[100731]_ ;
  assign \new_[100742]_  = ~A203 & ~A202;
  assign \new_[100745]_  = A266 & ~A265;
  assign \new_[100746]_  = \new_[100745]_  & \new_[100742]_ ;
  assign \new_[100749]_  = ~A268 & ~A267;
  assign \new_[100753]_  = ~A299 & ~A298;
  assign \new_[100754]_  = ~A269 & \new_[100753]_ ;
  assign \new_[100755]_  = \new_[100754]_  & \new_[100749]_ ;
  assign \new_[100756]_  = \new_[100755]_  & \new_[100746]_ ;
  assign \new_[100759]_  = ~A169 & A170;
  assign \new_[100762]_  = ~A167 & ~A168;
  assign \new_[100763]_  = \new_[100762]_  & \new_[100759]_ ;
  assign \new_[100766]_  = A199 & A166;
  assign \new_[100769]_  = ~A201 & ~A200;
  assign \new_[100770]_  = \new_[100769]_  & \new_[100766]_ ;
  assign \new_[100771]_  = \new_[100770]_  & \new_[100763]_ ;
  assign \new_[100774]_  = ~A203 & ~A202;
  assign \new_[100777]_  = ~A266 & A265;
  assign \new_[100778]_  = \new_[100777]_  & \new_[100774]_ ;
  assign \new_[100781]_  = A268 & A267;
  assign \new_[100785]_  = ~A302 & ~A301;
  assign \new_[100786]_  = A300 & \new_[100785]_ ;
  assign \new_[100787]_  = \new_[100786]_  & \new_[100781]_ ;
  assign \new_[100788]_  = \new_[100787]_  & \new_[100778]_ ;
  assign \new_[100791]_  = ~A169 & A170;
  assign \new_[100794]_  = ~A167 & ~A168;
  assign \new_[100795]_  = \new_[100794]_  & \new_[100791]_ ;
  assign \new_[100798]_  = A199 & A166;
  assign \new_[100801]_  = ~A201 & ~A200;
  assign \new_[100802]_  = \new_[100801]_  & \new_[100798]_ ;
  assign \new_[100803]_  = \new_[100802]_  & \new_[100795]_ ;
  assign \new_[100806]_  = ~A203 & ~A202;
  assign \new_[100809]_  = ~A266 & A265;
  assign \new_[100810]_  = \new_[100809]_  & \new_[100806]_ ;
  assign \new_[100813]_  = A269 & A267;
  assign \new_[100817]_  = ~A302 & ~A301;
  assign \new_[100818]_  = A300 & \new_[100817]_ ;
  assign \new_[100819]_  = \new_[100818]_  & \new_[100813]_ ;
  assign \new_[100820]_  = \new_[100819]_  & \new_[100810]_ ;
  assign \new_[100823]_  = ~A169 & A170;
  assign \new_[100826]_  = ~A167 & ~A168;
  assign \new_[100827]_  = \new_[100826]_  & \new_[100823]_ ;
  assign \new_[100830]_  = A199 & A166;
  assign \new_[100833]_  = ~A201 & ~A200;
  assign \new_[100834]_  = \new_[100833]_  & \new_[100830]_ ;
  assign \new_[100835]_  = \new_[100834]_  & \new_[100827]_ ;
  assign \new_[100838]_  = ~A203 & ~A202;
  assign \new_[100841]_  = ~A266 & A265;
  assign \new_[100842]_  = \new_[100841]_  & \new_[100838]_ ;
  assign \new_[100845]_  = ~A268 & ~A267;
  assign \new_[100849]_  = A301 & ~A300;
  assign \new_[100850]_  = ~A269 & \new_[100849]_ ;
  assign \new_[100851]_  = \new_[100850]_  & \new_[100845]_ ;
  assign \new_[100852]_  = \new_[100851]_  & \new_[100842]_ ;
  assign \new_[100855]_  = ~A169 & A170;
  assign \new_[100858]_  = ~A167 & ~A168;
  assign \new_[100859]_  = \new_[100858]_  & \new_[100855]_ ;
  assign \new_[100862]_  = A199 & A166;
  assign \new_[100865]_  = ~A201 & ~A200;
  assign \new_[100866]_  = \new_[100865]_  & \new_[100862]_ ;
  assign \new_[100867]_  = \new_[100866]_  & \new_[100859]_ ;
  assign \new_[100870]_  = ~A203 & ~A202;
  assign \new_[100873]_  = ~A266 & A265;
  assign \new_[100874]_  = \new_[100873]_  & \new_[100870]_ ;
  assign \new_[100877]_  = ~A268 & ~A267;
  assign \new_[100881]_  = A302 & ~A300;
  assign \new_[100882]_  = ~A269 & \new_[100881]_ ;
  assign \new_[100883]_  = \new_[100882]_  & \new_[100877]_ ;
  assign \new_[100884]_  = \new_[100883]_  & \new_[100874]_ ;
  assign \new_[100887]_  = ~A169 & A170;
  assign \new_[100890]_  = ~A167 & ~A168;
  assign \new_[100891]_  = \new_[100890]_  & \new_[100887]_ ;
  assign \new_[100894]_  = A199 & A166;
  assign \new_[100897]_  = ~A201 & ~A200;
  assign \new_[100898]_  = \new_[100897]_  & \new_[100894]_ ;
  assign \new_[100899]_  = \new_[100898]_  & \new_[100891]_ ;
  assign \new_[100902]_  = ~A203 & ~A202;
  assign \new_[100905]_  = ~A266 & A265;
  assign \new_[100906]_  = \new_[100905]_  & \new_[100902]_ ;
  assign \new_[100909]_  = ~A268 & ~A267;
  assign \new_[100913]_  = A299 & A298;
  assign \new_[100914]_  = ~A269 & \new_[100913]_ ;
  assign \new_[100915]_  = \new_[100914]_  & \new_[100909]_ ;
  assign \new_[100916]_  = \new_[100915]_  & \new_[100906]_ ;
  assign \new_[100919]_  = ~A169 & A170;
  assign \new_[100922]_  = ~A167 & ~A168;
  assign \new_[100923]_  = \new_[100922]_  & \new_[100919]_ ;
  assign \new_[100926]_  = A199 & A166;
  assign \new_[100929]_  = ~A201 & ~A200;
  assign \new_[100930]_  = \new_[100929]_  & \new_[100926]_ ;
  assign \new_[100931]_  = \new_[100930]_  & \new_[100923]_ ;
  assign \new_[100934]_  = ~A203 & ~A202;
  assign \new_[100937]_  = ~A266 & A265;
  assign \new_[100938]_  = \new_[100937]_  & \new_[100934]_ ;
  assign \new_[100941]_  = ~A268 & ~A267;
  assign \new_[100945]_  = ~A299 & ~A298;
  assign \new_[100946]_  = ~A269 & \new_[100945]_ ;
  assign \new_[100947]_  = \new_[100946]_  & \new_[100941]_ ;
  assign \new_[100948]_  = \new_[100947]_  & \new_[100938]_ ;
  assign \new_[100951]_  = ~A169 & A170;
  assign \new_[100954]_  = A167 & ~A168;
  assign \new_[100955]_  = \new_[100954]_  & \new_[100951]_ ;
  assign \new_[100958]_  = ~A199 & ~A166;
  assign \new_[100962]_  = ~A202 & ~A201;
  assign \new_[100963]_  = A200 & \new_[100962]_ ;
  assign \new_[100964]_  = \new_[100963]_  & \new_[100958]_ ;
  assign \new_[100965]_  = \new_[100964]_  & \new_[100955]_ ;
  assign \new_[100968]_  = ~A265 & ~A203;
  assign \new_[100971]_  = ~A267 & A266;
  assign \new_[100972]_  = \new_[100971]_  & \new_[100968]_ ;
  assign \new_[100975]_  = ~A269 & ~A268;
  assign \new_[100979]_  = ~A302 & ~A301;
  assign \new_[100980]_  = A300 & \new_[100979]_ ;
  assign \new_[100981]_  = \new_[100980]_  & \new_[100975]_ ;
  assign \new_[100982]_  = \new_[100981]_  & \new_[100972]_ ;
  assign \new_[100985]_  = ~A169 & A170;
  assign \new_[100988]_  = A167 & ~A168;
  assign \new_[100989]_  = \new_[100988]_  & \new_[100985]_ ;
  assign \new_[100992]_  = ~A199 & ~A166;
  assign \new_[100996]_  = ~A202 & ~A201;
  assign \new_[100997]_  = A200 & \new_[100996]_ ;
  assign \new_[100998]_  = \new_[100997]_  & \new_[100992]_ ;
  assign \new_[100999]_  = \new_[100998]_  & \new_[100989]_ ;
  assign \new_[101002]_  = A265 & ~A203;
  assign \new_[101005]_  = ~A267 & ~A266;
  assign \new_[101006]_  = \new_[101005]_  & \new_[101002]_ ;
  assign \new_[101009]_  = ~A269 & ~A268;
  assign \new_[101013]_  = ~A302 & ~A301;
  assign \new_[101014]_  = A300 & \new_[101013]_ ;
  assign \new_[101015]_  = \new_[101014]_  & \new_[101009]_ ;
  assign \new_[101016]_  = \new_[101015]_  & \new_[101006]_ ;
  assign \new_[101019]_  = ~A169 & A170;
  assign \new_[101022]_  = A167 & ~A168;
  assign \new_[101023]_  = \new_[101022]_  & \new_[101019]_ ;
  assign \new_[101026]_  = A199 & ~A166;
  assign \new_[101030]_  = ~A202 & ~A201;
  assign \new_[101031]_  = ~A200 & \new_[101030]_ ;
  assign \new_[101032]_  = \new_[101031]_  & \new_[101026]_ ;
  assign \new_[101033]_  = \new_[101032]_  & \new_[101023]_ ;
  assign \new_[101036]_  = ~A265 & ~A203;
  assign \new_[101039]_  = ~A267 & A266;
  assign \new_[101040]_  = \new_[101039]_  & \new_[101036]_ ;
  assign \new_[101043]_  = ~A269 & ~A268;
  assign \new_[101047]_  = ~A302 & ~A301;
  assign \new_[101048]_  = A300 & \new_[101047]_ ;
  assign \new_[101049]_  = \new_[101048]_  & \new_[101043]_ ;
  assign \new_[101050]_  = \new_[101049]_  & \new_[101040]_ ;
  assign \new_[101053]_  = ~A169 & A170;
  assign \new_[101056]_  = A167 & ~A168;
  assign \new_[101057]_  = \new_[101056]_  & \new_[101053]_ ;
  assign \new_[101060]_  = A199 & ~A166;
  assign \new_[101064]_  = ~A202 & ~A201;
  assign \new_[101065]_  = ~A200 & \new_[101064]_ ;
  assign \new_[101066]_  = \new_[101065]_  & \new_[101060]_ ;
  assign \new_[101067]_  = \new_[101066]_  & \new_[101057]_ ;
  assign \new_[101070]_  = A265 & ~A203;
  assign \new_[101073]_  = ~A267 & ~A266;
  assign \new_[101074]_  = \new_[101073]_  & \new_[101070]_ ;
  assign \new_[101077]_  = ~A269 & ~A268;
  assign \new_[101081]_  = ~A302 & ~A301;
  assign \new_[101082]_  = A300 & \new_[101081]_ ;
  assign \new_[101083]_  = \new_[101082]_  & \new_[101077]_ ;
  assign \new_[101084]_  = \new_[101083]_  & \new_[101074]_ ;
  assign \new_[101087]_  = ~A169 & A170;
  assign \new_[101090]_  = ~A167 & ~A168;
  assign \new_[101091]_  = \new_[101090]_  & \new_[101087]_ ;
  assign \new_[101094]_  = ~A199 & A166;
  assign \new_[101098]_  = ~A202 & ~A201;
  assign \new_[101099]_  = A200 & \new_[101098]_ ;
  assign \new_[101100]_  = \new_[101099]_  & \new_[101094]_ ;
  assign \new_[101101]_  = \new_[101100]_  & \new_[101091]_ ;
  assign \new_[101104]_  = ~A265 & ~A203;
  assign \new_[101107]_  = ~A267 & A266;
  assign \new_[101108]_  = \new_[101107]_  & \new_[101104]_ ;
  assign \new_[101111]_  = ~A269 & ~A268;
  assign \new_[101115]_  = ~A302 & ~A301;
  assign \new_[101116]_  = A300 & \new_[101115]_ ;
  assign \new_[101117]_  = \new_[101116]_  & \new_[101111]_ ;
  assign \new_[101118]_  = \new_[101117]_  & \new_[101108]_ ;
  assign \new_[101121]_  = ~A169 & A170;
  assign \new_[101124]_  = ~A167 & ~A168;
  assign \new_[101125]_  = \new_[101124]_  & \new_[101121]_ ;
  assign \new_[101128]_  = ~A199 & A166;
  assign \new_[101132]_  = ~A202 & ~A201;
  assign \new_[101133]_  = A200 & \new_[101132]_ ;
  assign \new_[101134]_  = \new_[101133]_  & \new_[101128]_ ;
  assign \new_[101135]_  = \new_[101134]_  & \new_[101125]_ ;
  assign \new_[101138]_  = A265 & ~A203;
  assign \new_[101141]_  = ~A267 & ~A266;
  assign \new_[101142]_  = \new_[101141]_  & \new_[101138]_ ;
  assign \new_[101145]_  = ~A269 & ~A268;
  assign \new_[101149]_  = ~A302 & ~A301;
  assign \new_[101150]_  = A300 & \new_[101149]_ ;
  assign \new_[101151]_  = \new_[101150]_  & \new_[101145]_ ;
  assign \new_[101152]_  = \new_[101151]_  & \new_[101142]_ ;
  assign \new_[101155]_  = ~A169 & A170;
  assign \new_[101158]_  = ~A167 & ~A168;
  assign \new_[101159]_  = \new_[101158]_  & \new_[101155]_ ;
  assign \new_[101162]_  = A199 & A166;
  assign \new_[101166]_  = ~A202 & ~A201;
  assign \new_[101167]_  = ~A200 & \new_[101166]_ ;
  assign \new_[101168]_  = \new_[101167]_  & \new_[101162]_ ;
  assign \new_[101169]_  = \new_[101168]_  & \new_[101159]_ ;
  assign \new_[101172]_  = ~A265 & ~A203;
  assign \new_[101175]_  = ~A267 & A266;
  assign \new_[101176]_  = \new_[101175]_  & \new_[101172]_ ;
  assign \new_[101179]_  = ~A269 & ~A268;
  assign \new_[101183]_  = ~A302 & ~A301;
  assign \new_[101184]_  = A300 & \new_[101183]_ ;
  assign \new_[101185]_  = \new_[101184]_  & \new_[101179]_ ;
  assign \new_[101186]_  = \new_[101185]_  & \new_[101176]_ ;
  assign \new_[101189]_  = ~A169 & A170;
  assign \new_[101192]_  = ~A167 & ~A168;
  assign \new_[101193]_  = \new_[101192]_  & \new_[101189]_ ;
  assign \new_[101196]_  = A199 & A166;
  assign \new_[101200]_  = ~A202 & ~A201;
  assign \new_[101201]_  = ~A200 & \new_[101200]_ ;
  assign \new_[101202]_  = \new_[101201]_  & \new_[101196]_ ;
  assign \new_[101203]_  = \new_[101202]_  & \new_[101193]_ ;
  assign \new_[101206]_  = A265 & ~A203;
  assign \new_[101209]_  = ~A267 & ~A266;
  assign \new_[101210]_  = \new_[101209]_  & \new_[101206]_ ;
  assign \new_[101213]_  = ~A269 & ~A268;
  assign \new_[101217]_  = ~A302 & ~A301;
  assign \new_[101218]_  = A300 & \new_[101217]_ ;
  assign \new_[101219]_  = \new_[101218]_  & \new_[101213]_ ;
  assign \new_[101220]_  = \new_[101219]_  & \new_[101210]_ ;
endmodule


