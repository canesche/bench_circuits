// Benchmark "pci_conf_cyc_addr_dec" written by ABC on Thu Oct  8 22:04:25 2020

module pci_conf_cyc_addr_dec ( 
    \ccyc_addr_in[0] , \ccyc_addr_in[1] , \ccyc_addr_in[2] ,
    \ccyc_addr_in[3] , \ccyc_addr_in[4] , \ccyc_addr_in[5] ,
    \ccyc_addr_in[6] , \ccyc_addr_in[7] , \ccyc_addr_in[8] ,
    \ccyc_addr_in[9] , \ccyc_addr_in[10] , \ccyc_addr_in[11] ,
    \ccyc_addr_in[12] , \ccyc_addr_in[13] , \ccyc_addr_in[14] ,
    \ccyc_addr_in[15] , \ccyc_addr_in[16] , \ccyc_addr_in[17] ,
    \ccyc_addr_in[18] , \ccyc_addr_in[19] , \ccyc_addr_in[20] ,
    \ccyc_addr_in[21] , \ccyc_addr_in[22] , \ccyc_addr_in[23] ,
    \ccyc_addr_in[24] , \ccyc_addr_in[25] , \ccyc_addr_in[26] ,
    \ccyc_addr_in[27] , \ccyc_addr_in[28] , \ccyc_addr_in[29] ,
    \ccyc_addr_in[30] , \ccyc_addr_in[31] ,
    \ccyc_addr_out[0] , \ccyc_addr_out[1] , \ccyc_addr_out[2] ,
    \ccyc_addr_out[3] , \ccyc_addr_out[4] , \ccyc_addr_out[5] ,
    \ccyc_addr_out[6] , \ccyc_addr_out[7] , \ccyc_addr_out[8] ,
    \ccyc_addr_out[9] , \ccyc_addr_out[10] , \ccyc_addr_out[11] ,
    \ccyc_addr_out[12] , \ccyc_addr_out[13] , \ccyc_addr_out[14] ,
    \ccyc_addr_out[15] , \ccyc_addr_out[16] , \ccyc_addr_out[17] ,
    \ccyc_addr_out[18] , \ccyc_addr_out[19] , \ccyc_addr_out[20] ,
    \ccyc_addr_out[21] , \ccyc_addr_out[22] , \ccyc_addr_out[23] ,
    \ccyc_addr_out[24] , \ccyc_addr_out[25] , \ccyc_addr_out[26] ,
    \ccyc_addr_out[27] , \ccyc_addr_out[28] , \ccyc_addr_out[29] ,
    \ccyc_addr_out[30] , \ccyc_addr_out[31]   );
  input  \ccyc_addr_in[0] , \ccyc_addr_in[1] , \ccyc_addr_in[2] ,
    \ccyc_addr_in[3] , \ccyc_addr_in[4] , \ccyc_addr_in[5] ,
    \ccyc_addr_in[6] , \ccyc_addr_in[7] , \ccyc_addr_in[8] ,
    \ccyc_addr_in[9] , \ccyc_addr_in[10] , \ccyc_addr_in[11] ,
    \ccyc_addr_in[12] , \ccyc_addr_in[13] , \ccyc_addr_in[14] ,
    \ccyc_addr_in[15] , \ccyc_addr_in[16] , \ccyc_addr_in[17] ,
    \ccyc_addr_in[18] , \ccyc_addr_in[19] , \ccyc_addr_in[20] ,
    \ccyc_addr_in[21] , \ccyc_addr_in[22] , \ccyc_addr_in[23] ,
    \ccyc_addr_in[24] , \ccyc_addr_in[25] , \ccyc_addr_in[26] ,
    \ccyc_addr_in[27] , \ccyc_addr_in[28] , \ccyc_addr_in[29] ,
    \ccyc_addr_in[30] , \ccyc_addr_in[31] ;
  output \ccyc_addr_out[0] , \ccyc_addr_out[1] , \ccyc_addr_out[2] ,
    \ccyc_addr_out[3] , \ccyc_addr_out[4] , \ccyc_addr_out[5] ,
    \ccyc_addr_out[6] , \ccyc_addr_out[7] , \ccyc_addr_out[8] ,
    \ccyc_addr_out[9] , \ccyc_addr_out[10] , \ccyc_addr_out[11] ,
    \ccyc_addr_out[12] , \ccyc_addr_out[13] , \ccyc_addr_out[14] ,
    \ccyc_addr_out[15] , \ccyc_addr_out[16] , \ccyc_addr_out[17] ,
    \ccyc_addr_out[18] , \ccyc_addr_out[19] , \ccyc_addr_out[20] ,
    \ccyc_addr_out[21] , \ccyc_addr_out[22] , \ccyc_addr_out[23] ,
    \ccyc_addr_out[24] , \ccyc_addr_out[25] , \ccyc_addr_out[26] ,
    \ccyc_addr_out[27] , \ccyc_addr_out[28] , \ccyc_addr_out[29] ,
    \ccyc_addr_out[30] , \ccyc_addr_out[31] ;
  wire \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ , \new_[101]_ ,
    \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ , \new_[106]_ ,
    \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ , \new_[111]_ ,
    \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ , \new_[116]_ ,
    \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ , \new_[121]_ ,
    \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ , \new_[126]_ ,
    \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ , \new_[131]_ ,
    \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ , \new_[136]_ ,
    \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ , \new_[141]_ ,
    \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ , \new_[146]_ ,
    \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ , \new_[151]_ ,
    \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ , \new_[156]_ ,
    \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ , \new_[162]_ ,
    \new_[163]_ , \new_[164]_ , \new_[165]_ , \new_[166]_ , \new_[167]_ ,
    \new_[168]_ , \new_[169]_ , \new_[170]_ , \new_[171]_ , \new_[172]_ ;
  assign \ccyc_addr_out[1]  = \ccyc_addr_in[1] ;
  assign \ccyc_addr_out[2]  = \ccyc_addr_in[2] ;
  assign \ccyc_addr_out[3]  = \ccyc_addr_in[3] ;
  assign \ccyc_addr_out[4]  = \ccyc_addr_in[4] ;
  assign \ccyc_addr_out[5]  = \ccyc_addr_in[5] ;
  assign \ccyc_addr_out[6]  = \ccyc_addr_in[6] ;
  assign \ccyc_addr_out[7]  = \ccyc_addr_in[7] ;
  assign \ccyc_addr_out[8]  = \ccyc_addr_in[8] ;
  assign \ccyc_addr_out[9]  = \ccyc_addr_in[9] ;
  assign \ccyc_addr_out[10]  = \ccyc_addr_in[10] ;
  assign \ccyc_addr_out[30]  = ~\new_[115]_  | (~\new_[126]_  & ~\new_[98]_ );
  assign \ccyc_addr_out[29]  = ~\new_[151]_  | (~\new_[147]_  & ~\new_[98]_ );
  assign \ccyc_addr_out[28]  = ~\new_[123]_  | (~\new_[131]_  & ~\new_[97]_ );
  assign \ccyc_addr_out[27]  = ~\new_[116]_  | (~\new_[120]_  & ~\new_[97]_ );
  assign \ccyc_addr_out[31]  = ~\new_[143]_  | (~\new_[105]_  & ~\ccyc_addr_out[0] );
  assign \ccyc_addr_out[26]  = ~\new_[118]_  | (~\new_[134]_  & ~\new_[99]_ );
  assign \ccyc_addr_out[25]  = ~\new_[138]_  | (~\new_[142]_  & ~\new_[99]_ );
  assign \ccyc_addr_out[24]  = ~\new_[144]_  | (~\new_[145]_  & ~\new_[104]_ );
  assign \ccyc_addr_out[23]  = ~\new_[148]_  | (~\new_[122]_  & ~\new_[104]_ );
  assign \ccyc_addr_out[22]  = ~\new_[152]_  | (~\new_[121]_  & ~\new_[106]_ );
  assign \ccyc_addr_out[21]  = ~\new_[117]_  | (~\new_[119]_  & ~\new_[106]_ );
  assign \ccyc_addr_out[20]  = ~\new_[133]_  | (~\new_[128]_  & ~\new_[107]_ );
  assign \ccyc_addr_out[19]  = ~\new_[125]_  | (~\new_[130]_  & ~\new_[107]_ );
  assign \ccyc_addr_out[18]  = ~\new_[132]_  | (~\new_[137]_  & ~\new_[102]_ );
  assign \ccyc_addr_out[17]  = ~\new_[135]_  | (~\new_[139]_  & ~\new_[102]_ );
  assign \ccyc_addr_out[16]  = ~\new_[141]_  | (~\new_[140]_  & ~\new_[100]_ );
  assign \ccyc_addr_out[15]  = ~\new_[158]_  | (~\new_[129]_  & ~\new_[100]_ );
  assign \ccyc_addr_out[14]  = ~\new_[153]_  | (~\new_[146]_  & ~\new_[101]_ );
  assign \ccyc_addr_out[13]  = ~\new_[154]_  | (~\new_[149]_  & ~\new_[101]_ );
  assign \ccyc_addr_out[12]  = ~\new_[157]_  | (~\new_[150]_  & ~\new_[103]_ );
  assign \ccyc_addr_out[11]  = ~\new_[136]_  | (~\new_[124]_  & ~\new_[103]_ );
  assign \new_[97]_  = ~\new_[108]_  | ~\new_[168]_ ;
  assign \new_[98]_  = ~\new_[109]_  | ~\ccyc_addr_in[12] ;
  assign \new_[99]_  = ~\new_[111]_  | ~\ccyc_addr_in[12] ;
  assign \new_[100]_  = ~\new_[112]_  | ~\new_[168]_ ;
  assign \new_[101]_  = ~\new_[113]_  | ~\ccyc_addr_in[12] ;
  assign \new_[102]_  = ~\new_[112]_  | ~\ccyc_addr_in[12] ;
  assign \new_[103]_  = ~\new_[113]_  | ~\new_[168]_ ;
  assign \new_[104]_  = ~\new_[111]_  | ~\new_[168]_ ;
  assign \new_[105]_  = ~\ccyc_addr_in[13]  | ~\new_[155]_  | ~\new_[127]_ ;
  assign \new_[106]_  = ~\new_[114]_  | ~\ccyc_addr_in[12] ;
  assign \new_[107]_  = ~\new_[114]_  | ~\new_[168]_ ;
  assign \new_[108]_  = ~\new_[110]_ ;
  assign \new_[109]_  = ~\new_[110]_ ;
  assign \new_[110]_  = ~\new_[167]_  | ~\new_[171]_  | ~\new_[165]_ ;
  assign \new_[111]_  = ~\new_[156]_  & ~\new_[167]_ ;
  assign \new_[112]_  = ~\new_[159]_  & ~\new_[167]_ ;
  assign \new_[113]_  = ~\new_[159]_  & ~\ccyc_addr_in[13] ;
  assign \new_[114]_  = ~\new_[156]_  & ~\ccyc_addr_in[13] ;
  assign \new_[115]_  = ~\ccyc_addr_in[30]  | ~\ccyc_addr_out[0] ;
  assign \new_[116]_  = ~\ccyc_addr_in[27]  | ~\ccyc_addr_out[0] ;
  assign \new_[117]_  = ~\ccyc_addr_in[21]  | ~\ccyc_addr_out[0] ;
  assign \new_[118]_  = ~\ccyc_addr_in[26]  | ~\ccyc_addr_out[0] ;
  assign \new_[119]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[120]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[121]_  = ~\ccyc_addr_in[11]  | ~\new_[162]_ ;
  assign \new_[122]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[123]_  = ~\ccyc_addr_in[28]  | ~\ccyc_addr_out[0] ;
  assign \new_[124]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[125]_  = ~\ccyc_addr_in[19]  | ~\ccyc_addr_out[0] ;
  assign \new_[126]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[127]_  = \new_[165]_  & \new_[171]_ ;
  assign \new_[128]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[129]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[130]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[131]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[132]_  = ~\ccyc_addr_in[18]  | ~\ccyc_addr_out[0] ;
  assign \new_[133]_  = ~\ccyc_addr_in[20]  | ~\ccyc_addr_out[0] ;
  assign \new_[134]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[135]_  = ~\ccyc_addr_in[17]  | ~\ccyc_addr_out[0] ;
  assign \new_[136]_  = ~\new_[160]_  | ~\ccyc_addr_out[0] ;
  assign \new_[137]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[138]_  = ~\ccyc_addr_in[25]  | ~\ccyc_addr_out[0] ;
  assign \new_[139]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[140]_  = ~\ccyc_addr_in[11]  | ~\new_[162]_ ;
  assign \new_[141]_  = ~\ccyc_addr_in[16]  | ~\ccyc_addr_out[0] ;
  assign \new_[142]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[143]_  = ~\ccyc_addr_in[31]  | ~\ccyc_addr_out[0] ;
  assign \new_[144]_  = ~\ccyc_addr_in[24]  | ~\ccyc_addr_out[0] ;
  assign \new_[145]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[146]_  = ~\new_[160]_  | ~\new_[162]_ ;
  assign \new_[147]_  = \new_[163]_  | \ccyc_addr_out[0] ;
  assign \new_[148]_  = ~\ccyc_addr_in[23]  | ~\ccyc_addr_out[0] ;
  assign \new_[149]_  = \new_[163]_  | \ccyc_addr_in[0] ;
  assign \new_[150]_  = ~\ccyc_addr_in[11]  | ~\new_[162]_ ;
  assign \new_[151]_  = ~\ccyc_addr_in[29]  | ~\ccyc_addr_out[0] ;
  assign \new_[152]_  = ~\ccyc_addr_in[22]  | ~\ccyc_addr_out[0] ;
  assign \new_[153]_  = \new_[165]_  | \new_[166]_ ;
  assign \new_[154]_  = \new_[167]_  | \new_[166]_ ;
  assign \new_[155]_  = ~\new_[163]_  & ~\ccyc_addr_in[12] ;
  assign \new_[156]_  = ~\new_[172]_  | ~\ccyc_addr_in[14] ;
  assign \new_[157]_  = \new_[168]_  | \new_[166]_ ;
  assign \new_[158]_  = \new_[170]_  | \new_[166]_ ;
  assign \new_[159]_  = ~\new_[172]_  | ~\new_[169]_ ;
  assign \new_[160]_  = ~\new_[164]_ ;
  assign \ccyc_addr_out[0]  = ~\new_[166]_ ;
  assign \new_[162]_  = ~\ccyc_addr_in[0] ;
  assign \new_[163]_  = \ccyc_addr_in[11] ;
  assign \new_[164]_  = ~\ccyc_addr_in[11] ;
  assign \new_[165]_  = ~\ccyc_addr_in[14] ;
  assign \new_[166]_  = ~\ccyc_addr_in[0] ;
  assign \new_[167]_  = ~\ccyc_addr_in[13] ;
  assign \new_[168]_  = ~\ccyc_addr_in[12] ;
  assign \new_[169]_  = ~\ccyc_addr_in[14] ;
  assign \new_[170]_  = ~\new_[171]_ ;
  assign \new_[171]_  = ~\new_[172]_ ;
  assign \new_[172]_  = ~\ccyc_addr_in[15] ;
endmodule


