module top ( clock, 
    pg115, pg126, pg116, pg125, pg5, pg135, pg127, pg100, pg6751, pg99,
    pg6750, pg120, pg134, pg113, pg124, pg114, pg92, pg6748, pg91, pg6749,
    pclk, pg6746, pg84, pg6747, pg6744, pg6745, pg6753, pg6752, pg56, pg57,
    pg64, pg73, pg36, pg54, pg72, pg90, pg35, pg44, pg53,
    pg8342, pg8353, pg8870, pg9048, pg9741, pg13272, pg13906, pg28030,
    pg28041, pg33533, pg34437, pg8132, pg8783, pg9555, pg12184, pg13068,
    pg13099, pg31521, pg33435, pg34425, pg7260, pg8344, pg8784, pg14167,
    pg17320, pg18101, pg30327, pg31793, pg34435, pg8398, pg8785, pg18100,
    pg20899, pg34436, pg8786, pg14828, pg20557, pg20654, pg21727, pg24171,
    pg24182, pg26876, pg30329, pg33894, pg34239, pg7243, pg7540, pg8235,
    pg8787, pg12470, pg17819, pg19334, pg24172, pg24181, pg26877, pg32454,
    pg34597, pg8403, pg8788, pg9497, pg13926, pg14189, pg14451, pg23190,
    pg24151, pg24162, pg24180, pg26801, pg33874, pg34237, pg7245, pg8215,
    pg8789, pg10122, pg12919, pg16924, pg17291, pg20763, pg24161, pg24170,
    pg28042, pg34238, pg12833, pg14705, pg14738, pg14749, pg16693, pg16718,
    pg17423, pg18097, pg24164, pg24175, pg29211, pg34235, pg18098, pg20901,
    pg23652, pg24163, pg24176, pg24185, pg29210, pg34201, pg34236, pg11388,
    pg17577, pg17674, pg17760, pg18099, pg20652, pg24166, pg24173, pg24184,
    pg29213, pg29220, pg34233, pg34972, pg14597, pg14694, pg17813, pg21292,
    pg24165, pg24174, pg24183, pg29212, pg29221, pg32975, pg34234, pg34788,
    pg11678, pg12923, pg14518, pg14662, pg14673, pg17607, pg17715, pg19357,
    pg24168, pg24179, pg25219, pg29215, pg30332, pg34956, pg16627, pg23612,
    pg24167, pg29214, pg34232, pg14635, pg17519, pg17580, pg24177, pg25167,
    pg29217, pg30330, pg34240, pg12832, pg16722, pg24169, pg24178, pg29216,
    pg30331, pg34221, pg7916, pg8919, pg11447, pg13881, pg16624, pg17711,
    pg17722, pg20049, pg25259, pg25583, pg29219, pg33948, pg33959, pg34927,
    pg8918, pg11770, pg16874, pg17604, pg21245, pg25584, pg29218, pg33949,
    pg34917, pg25585, pg32185, pg33946, pg34839, pg8839, pg16603, pg16656,
    pg16744, pg17646, pg17743, pg17778, pg17787, pg18092, pg25586, pg33947,
    pg34919, pg11418, pg16686, pg17845, pg21176, pg25114, pg25590, pg34383,
    pg34923, pg12368, pg13895, pg14779, pg17639, pg17688, pg18094, pg18881,
    pg23683, pg33079, pg33945, pg34913, pg10527, pg13865, pg16659, pg17649,
    pg17678, pg17685, pg17739, pg17764, pg18095, pg33935, pg34925, pg11349,
    pg13259, pg16748, pg16775, pg17316, pg17404, pg17871, pg18096, pg21270,
    pg25582, pg34915, pg8416, pg9617, pg31863, pg33659, pg33950, pg7257,
    pg8920, pg9251, pg9817, pg13966, pg14217, pg27831, pg31861, pg34921,
    pg8291, pg12238, pg12300, pg14096, pg14201, pg14421, pg16955, pg17400,
    pg26875, pg31862, pg32429, pg8283, pg8915, pg9019, pg9682, pg12350,
    pg12422, pg13049, pg13085, pg14125, pg14147, pg25587, pg31665, pg8279,
    pg21698, pg25588, pg31860, pg8719, pg8917, pg9615, pg9680, pg9743,
    pg23002, pg25589, pg28753, pg31656, pg33636, pg7946, pg8178, pg8277,
    pg8358, pg8475, pg8916, pg9553, pg10306, pg10500, pg13039, pg23759  );
  input  clock;
  input  pg115, pg126, pg116, pg125, pg5, pg135, pg127, pg100, pg6751,
    pg99, pg6750, pg120, pg134, pg113, pg124, pg114, pg92, pg6748, pg91,
    pg6749, pclk, pg6746, pg84, pg6747, pg6744, pg6745, pg6753, pg6752,
    pg56, pg57, pg64, pg73, pg36, pg54, pg72, pg90, pg35, pg44, pg53;
  output pg8342, pg8353, pg8870, pg9048, pg9741, pg13272, pg13906, pg28030,
    pg28041, pg33533, pg34437, pg8132, pg8783, pg9555, pg12184, pg13068,
    pg13099, pg31521, pg33435, pg34425, pg7260, pg8344, pg8784, pg14167,
    pg17320, pg18101, pg30327, pg31793, pg34435, pg8398, pg8785, pg18100,
    pg20899, pg34436, pg8786, pg14828, pg20557, pg20654, pg21727, pg24171,
    pg24182, pg26876, pg30329, pg33894, pg34239, pg7243, pg7540, pg8235,
    pg8787, pg12470, pg17819, pg19334, pg24172, pg24181, pg26877, pg32454,
    pg34597, pg8403, pg8788, pg9497, pg13926, pg14189, pg14451, pg23190,
    pg24151, pg24162, pg24180, pg26801, pg33874, pg34237, pg7245, pg8215,
    pg8789, pg10122, pg12919, pg16924, pg17291, pg20763, pg24161, pg24170,
    pg28042, pg34238, pg12833, pg14705, pg14738, pg14749, pg16693, pg16718,
    pg17423, pg18097, pg24164, pg24175, pg29211, pg34235, pg18098, pg20901,
    pg23652, pg24163, pg24176, pg24185, pg29210, pg34201, pg34236, pg11388,
    pg17577, pg17674, pg17760, pg18099, pg20652, pg24166, pg24173, pg24184,
    pg29213, pg29220, pg34233, pg34972, pg14597, pg14694, pg17813, pg21292,
    pg24165, pg24174, pg24183, pg29212, pg29221, pg32975, pg34234, pg34788,
    pg11678, pg12923, pg14518, pg14662, pg14673, pg17607, pg17715, pg19357,
    pg24168, pg24179, pg25219, pg29215, pg30332, pg34956, pg16627, pg23612,
    pg24167, pg29214, pg34232, pg14635, pg17519, pg17580, pg24177, pg25167,
    pg29217, pg30330, pg34240, pg12832, pg16722, pg24169, pg24178, pg29216,
    pg30331, pg34221, pg7916, pg8919, pg11447, pg13881, pg16624, pg17711,
    pg17722, pg20049, pg25259, pg25583, pg29219, pg33948, pg33959, pg34927,
    pg8918, pg11770, pg16874, pg17604, pg21245, pg25584, pg29218, pg33949,
    pg34917, pg25585, pg32185, pg33946, pg34839, pg8839, pg16603, pg16656,
    pg16744, pg17646, pg17743, pg17778, pg17787, pg18092, pg25586, pg33947,
    pg34919, pg11418, pg16686, pg17845, pg21176, pg25114, pg25590, pg34383,
    pg34923, pg12368, pg13895, pg14779, pg17639, pg17688, pg18094, pg18881,
    pg23683, pg33079, pg33945, pg34913, pg10527, pg13865, pg16659, pg17649,
    pg17678, pg17685, pg17739, pg17764, pg18095, pg33935, pg34925, pg11349,
    pg13259, pg16748, pg16775, pg17316, pg17404, pg17871, pg18096, pg21270,
    pg25582, pg34915, pg8416, pg9617, pg31863, pg33659, pg33950, pg7257,
    pg8920, pg9251, pg9817, pg13966, pg14217, pg27831, pg31861, pg34921,
    pg8291, pg12238, pg12300, pg14096, pg14201, pg14421, pg16955, pg17400,
    pg26875, pg31862, pg32429, pg8283, pg8915, pg9019, pg9682, pg12350,
    pg12422, pg13049, pg13085, pg14125, pg14147, pg25587, pg31665, pg8279,
    pg21698, pg25588, pg31860, pg8719, pg8917, pg9615, pg9680, pg9743,
    pg23002, pg25589, pg28753, pg31656, pg33636, pg7946, pg8178, pg8277,
    pg8358, pg8475, pg8916, pg9553, pg10306, pg10500, pg13039, pg23759;
  reg ng6215, ng4332, ng2837, ng1135, ng2485, ng4375, ng4304, ng1171,
    ng3235, ng2852, ng4135, ng222, ng365, ng2815, ng4888, ng433, ng3736,
    ng246, ng102, ng1030, ng110, ng3983, ng4801, ng4045, ng4169, ng2145,
    ng5138, ng3873, ng3752, ng136, ng1772, ng990, ng3171, ng168, ng441,
    ng160, ng5283, ng1361, ng6621, ng5689, ng6593, ng55, ng5827, ng1079,
    ng74, ng5381, ng5723, ng4443, ng979, ng1484, ng6044, ng3817, ng316,
    ng887, ng3080, ng499, ng6012, ng3443, ng2269, ng2927, ng577, ng599,
    ng4222, ng781, ng6428, ng2759, ng2715, ng1870, ng1768, ng4031, ng6181,
    ng5731, ng2173, ng1783, ng6058, ng106, ng2711, ng2803, ng6303, ng3462,
    ng482, ng3085, ng1811, ng2890, ng1542, ng111, ng2161, ng947, ng546,
    ng3913, ng1570, ng4213, ng5599, ng3893, ng4141, ng3106, ng3841, ng2004,
    ng3586, ng4132, ng939, ng6195, ng925, ng6255, ng2177, ng5835, ng4543,
    ng5802, ng5092, ng3933, ng6027, ng911, ng3901, ng4297, ng1582, ng4049,
    ng3139, ng3672, ng6649, ng2599, ng4087, ng1467, ng6519, ng1700, ng1950,
    ng3632, ng46, ng2417, ng4741, ng475, ng3787, ng333, ng5105, ng6351,
    ng1779, ng2834, ng3470, ng5188, ng1116, ng504, ng3767, ng6541, ng6209,
    ng5685, ng1157, ng3466, ng3333, ng4922, ng6613, ng93, ng637, ng5327,
    ng1478, ng5413, ng63, ng2643, ng191, ng6052, ng1620, ng3668, ng2495,
    ng5583, ng2138, ng5244, ng936, ng429, ng4854, ng37, ng6381, ng347,
    ng4287, ng2767, ng4207, ng5921, ng6023, ng85, ng5069, ng1061, ng4401,
    ng3298, ng3431, ng3610, ng4975, ng4427, ng4145, ng1834, ng5703, ng4537,
    ng1141, ng6120, ng4512, ng4253, ng4570, ng1548, ng4284, ng385, ng291,
    ng5666, ng3111, ng718, ng6497, ng6267, ng3010, ng2399, ng2898, ng4414,
    ng4831, ng5889, ng822, ng43, ng6315, ng2112, ng5543, ng4449, ng142,
    ng5022, ng6148, ng1448, ng3961, ng1018, ng5029, ng513, ng5109, ng2016,
    ng5575, ng5052, ng3412, ng1992, ng2902, ng3808, ng5373, ng1608, ng5535,
    ng405, ng215, ng5448, ng3203, ng655, ng4423, ng4633, ng4116, ng298,
    ng1075, ng4501, ng6513, ng3368, ng5240, ng1002, ng896, ng3451, ng2712,
    ng5929, ng6486, ng837, ng2437, ng6373, ng3661, ng785, ng2575, ng6711,
    ng3925, ng4812, ng4765, ng1266, ng6605, ng2868, ng6573, ng5485, ng1211,
    ng1821, ng5124, ng5377, ng6434, ng6697, ng4932, ng5008, ng790, ng5142,
    ng3594, ng5953, ng5677, ng6561, ng2775, ng4366, ng5016, ng5654, ng5128,
    ng3763, ng5456, ng4674, ng4153, ng117, ng3239, ng1437, ng4809, ng52,
    ng4269, ng3343, ng2819, ng3050, ng4495, ng1070, ng4012, ng6251, ng1283,
    ng6537, ng2932, ng4584, ng4019, ng5798, ng881, ng2984, ng1418, ng1256,
    ng2841, ng2307, ng5759, ng3719, ng5452, ng31, ng3029, ng4455, ng9,
    ng5445, ng4197, ng4950, ng5216, ng2710, ng1936, ng1668, ng5290, ng3689,
    ng4146, ng4681, ng3774, ng827, ng287, ng1277, ng2799, ng1945, ng776,
    ng358, ng967, ng626, ng4340, ng2036, ng1249, ng2102, ng6173, ng2338,
    ng6741, ng65, ng6365, ng6509, ng2070, ng5563, ng4473, ng2445, ng2407,
    ng1677, ng86, ng2827, ng6451, ng1083, ng1306, ng1514, ng4727, ng3219,
    ng6597, ng5913, ng3259, ng2999, ng2472, ng3195, ng4417, ng2922, ng3401,
    ng3119, ng3211, ng3821, ng3191, ng2527, ng3243, ng5204, ng1862, ng6065,
    ng1178, ng6329, ng3530, ng4273, ng4572, ng2259, ng6191, ng6307, ng4281,
    ng4639, ng5037, ng6279, ng471, ng5297, ng4216, ng232, ng3759, ng3498,
    ng6555, ng1472, ng4760, ng2204, ng862, ng6736, ng6500, ng2724, ng2882,
    ng2541, ng6653, ng4894, ng2476, ng2729, ng3317, ng930, ng6682, ng2873,
    ng4899, ng4229, ng3484, ng604, ng1825, ng4392, ng4520, ng1395, ng714,
    ng79, ng6505, ng5462, ng3731, ng6423, ng5073, ng1636, ng5849, ng2197,
    ng4129, ng1858, ng6581, ng1902, ng2126, ng4200, ng582, ng3845, ng5747,
    ng2079, ng6082, ng5841, ng4239, ng5148, ng5630, ng5969, ng6322, ng128,
    ng2610, ng6727, ng4742, ng3143, ng4927, ng5077, ng2342, ng3574, ng4138,
    ng2319, ng5752, ng51, ng5791, ng1041, ng3770, ng4467, ng2279, ng859,
    ng2606, ng262, ng3502, ng5817, ng4944, ng3827, ng4704, ng336, ng2153,
    ng3480, ng5681, ng4646, ng5357, ng4907, ng3937, ng5949, ng1854, ng4064,
    ng6247, ng1259, ng6589, ng3004, ng5002, ng1322, ng1913, ng5489, ng182,
    ng1592, ng2689, ng3089, ng875, ng2509, ng3921, ng1756, ng6116, ng2950,
    ng446, ng4349, ng6163, ng5248, ng4446, ng4191, ng2116, ng2697, ng3676,
    ng49, ng2453, ng3391, ng4420, ng3606, ng843, ng3506, ng1036, ng4104,
    ng1706, ng6398, ng5523, ng6159, ng2960, ng5495, ng2975, ng6549, ng2315,
    ng2595, ng6545, ng2652, ng6235, ng3385, ng542, ng1840, ng703, ng5101,
    ng4072, ng3133, ng22, ng1906, ng4912, ng1959, ng3857, ng2375, ng4991,
    ng2946, ng2831, ng739, ng5084, ng4785, ng2791, ng6609, ng2098, ng6455,
    ng3546, ng2185, ng2491, ng1312, ng1129, ng1221, ng1624, ng1848, ng4859,
    ng4815, ng2994, ng956, ng2421, ng6533, ng370, ng1874, ng4125, ng5481,
    ng7, ng2361, ng2327, ng723, ng94, ng3703, ng4549, ng4180, ng1926,
    ng676, ng4558, ng4864, ng1532, ng1389, ng3618, ng3802, ng2255, ng5499,
    ng4185, ng5917, ng6167, ng3917, ng2537, ng5268, ng5459, ng3419, ng3881,
    ng6113, ng5256, ng5421, ng4732, ng344, ng5673, ng2878, ng933, ng4157,
    ng3863, ng3976, ng1657, ng6019, ng4035, ng667, ng5475, ng5603, ng2719,
    ng3949, ng209, ng4462, ng4249, ng5236, ng4219, ng4849, ng3310, ng2227,
    ng6411, ng5062, ng34, ng424, ng1280, ng650, ng2181, ng1046, ng1345,
    ng5694, ng2441, ng4821, ng3694, ng2779, ng376, ng907, ng699, ng3129,
    ng4698, ng6035, ng4507, ng4040, ng3380, ng5555, ng590, ng1752, ng4477,
    ng1296, ng4382, ng1052, ng1728, ng969, ng355, ng5335, ng6490, ng225,
    ng5869, ng153, ng2811, ng1585, ng3454, ng4108, ng5881, ng1146, ng518,
    ng4531, ng3045, ng468, ng5041, ng2988, ng1526, ng568, ng4294, ng3361,
    ng4546, ng3072, ng6098, ng6283, ng6415, ng5120, ng1399, ng4322, ng5252,
    ng1274, ng112, ng5033, ng4939, ng5097, ng5112, ng3408, ng3329, ng943,
    ng5200, ng2912, ng3352, ng3125, ng1988, ng5348, ng1, ng1878, ng2547,
    ng5343, ng48, ng6692, ng5567, ng1233, ng753, ng351, ng58, ng3179,
    ng2807, ng1682, ng5831, ng3231, ng4486, ng5579, ng6625, ng3798, ng4388,
    ng4564, ng4308, ng5385, ng2625, ng3897, ng2860, ng6641, ng5396, ng2151,
    ng3538, ng6523, ng3263, ng3562, ng6675, ng5937, ng1242, ng4771, ng6369,
    ng4966, ng5320, ng1199, ng5941, ng1152, ng6346, ng2856, ng4818, ng1056,
    ng1964, ng19, ng5401, ng5170, ng1559, ng4843, ng5637, ng6657, ng2894,
    ng4311, ng3223, ng3251, ng5619, ng559, ng554, ng1798, ng4871, ng1579,
    ng4643, ng2980, ng5901, ng479, ng4653, ng5424, ng1105, ng3889, ng4098,
    ng4504, ng1589, ng5990, ng3805, ng6275, ng6239, ng4571, ng5406, ng150,
    ng538, ng4743, ng5571, ng5196, ng2351, ng4434, ng301, ng854, ng2518,
    ng5976, ng6719, ng1236, ng4616, ng2523, ng2551, ng6715, ng2579, ng5276,
    ng3929, ng2012, ng4836, ng2108, ng2571, ng2093, ng6479, ng1554, ng3207,
    ng4027, ng1720, ng1193, ng3255, ng5893, ng4456, ng6140, ng1300, ng3747,
    ng4552, ng5417, ng3187, ng4931, ng1996, ng3654, ng3017, ng496, ng878,
    ng4722, ng6154, ng5264, ng3151, ng2886, ng6386, ng5736, ng4054, ng1087,
    ng3476, ng4575, ng5873, ng5719, ng4578, ng4459, ng6311, ng4826, ng3281,
    ng3338, ng1696, ng3025, ng6, ng3578, ng2380, ng2648, ng5441, ng341,
    ng4601, ng2567, ng890, ng2864, ng28, ng4561, ng3103, ng5156, ng2273,
    ng904, ng6459, ng6227, ng6203, ng66, ng6000, ng2165, ng4112, ng1982,
    ng4717, ng4483, ng3215, ng1367, ng2051, ng1691, ng1111, ng5821, ng411,
    ng4057, ng5763, ng3325, ng2661, ng3061, ng2970, ng4628, ng12, ng2771,
    ng3570, ng622, ng3853, ng2941, ng3100, ng4737, ng3440, ng5360, ng4754,
    ng4983, ng4961, ng3494, ng4749, ng2465, ng4917, ng3680, ng1748, ng3092,
    ng758, ng1227, ng1664, ng528, ng2848, ng1564, ng3712, ng962, ng457,
    ng5787, ng3831, ng4793, ng5808, ng6358, ng1890, ng799, ng5897, ng5331,
    ng3791, ng4093, ng2619, ng661, ng6494, ng1413, ng2311, ng5774, ng70,
    ng794, ng4999, ng2667, ng2555, ng4581, ng1616, ng305, ng255, ng3423,
    ng613, ng5390, ng3034, ng817, ng686, ng4489, ng4955, ng2675, ng25,
    ng391, ng329, ng6668, ng6704, ng5727, ng6439, ng2533, ng6404, ng2936,
    ng3267, ng6299, ng3068, ng319, ng1351, ng3274, ng728, ng2084, ng691,
    ng5698, ng4515, ng1882, ng640, ng6336, ng5134, ng4076, ng1495, ng3040,
    ng3969, ng5160, ng1189, ng3372, ng437, ng5511, ng3965, ng6483, ng6187,
    ng914, ng5551, ng1373, ng5712, ng632, ng1246, ng4498, ng5805, ng2241,
    ng2370, ng5770, ng2756, ng3436, ng2514, ng2763, ng6645, ng3869, ng2629,
    ng45, ng4165, ng3639, ng269, ng3957, ng1183, ng5767, ng4669, ng4411,
    ng3602, ng4688, ng3227, ng4023, ng2040, ng3396, ng6077, ng3021, ng5857,
    ng8, ng550, ng283, ng2795, ng194, ng6049, ng4082, ng1252, ng5527,
    ng5224, ng1287, ng1644, ng5176, ng1536, ng5228, ng3849, ng2303, ng3096,
    ng324, ng6527, ng5644, ng1311, ng1239, ng3953, ng164, ng1648, ng929,
    ng6295, ng1792, ng2583, ng3416, ng3447, ng6462, ng278, ng6395, ng1422,
    ng763, ng1632, ng744, ng1442, ng1454, ng2287, ng3566, ng681, ng3518,
    ng736, ng5623, ng3835, ng5339, ng174, ng5742, ng2783, ng5983, ng6243,
    ng6128, ng16, ng239, ng4452, ng884, ng2152, ng5164, ng4226, ng2461,
    ng4369, ng3288, ng1263, ng4664, ng2047, ng4430, ng572, ng3990, ng812,
    ng3684, ng401, ng6151, ng586, ng2393, ng5428, ng5308, ng2587, ng6271,
    ng2020, ng460, ng3247, ng4210, ng199, ng5080, ng2965, ng1404, ng617,
    ng3161, ng1844, ng6109, ng1955, ng6419, ng671, ng1270, ng5925, ng2787,
    ng6601, ng4119, ng5845, ng6661, ng3550, ng1687, ng1710, ng5152, ng2060,
    ng3727, ng5046, ng4232, ng4519, ng3614, ng5272, ng4358, ng3003, ng5366,
    ng5260, ng4300, ng71, ng2299, ng4492, ng6137, ng3794, ng3905, ng5313,
    ng1917, ng5965, ng5933, ng5611, ng4534, ng417, ng1604, ng2008, ng2122,
    ng2433, ng4164, ng6637, ng3558, ng157, ng1459, ng5961, ng6629, ng5436,
    ng1216, ng1430, ng3742, ng5208, ng1333, ng101, ng5706, ng1816, ng2403,
    ng952, ng2223, ng5957, ng4188, ng2130, ng3706, ng832, ng2823, ng6040,
    ng1760, ng869, ng2193, ng996, ng4474, ng4480, ng3582, ng4000, ng5467,
    ng4608, ng1894, ng5011, ng5863, ng6444, ng3723, ng5220, ng2384, ng4527,
    ng1489, ng4277, ng3347, ng2265, ng1974, ng1124, ng2429, ng1978, ng6390,
    ng3199, ng3065, ng1740, ng2681, ng2413, ng5352, ng6617, ng2704, ng2250,
    ng2357, ng5115, ng5595, ng2735, ng4659, ng1094, ng534, ng1521, ng4204,
    ng59, ng772, ng2563, ng3598, ng294, ng921, ng3522, ng1379, ng5587,
    ng1500, ng4264, ng6291, ng2955, ng3115, ng1724, ng6177, ng4593, ng1024,
    ng3625, ng203, ng5057, ng6377, ng4776, ng5591, ng5507, ng6088, ng452,
    ng807, ng1600, ng4621, ng1099, ng2024, ng901, ng4242, ng2741, ng2217,
    ng464, ng6219, ng1714, ng1968, ng4878, ng3303, ng4194, ng5503, ng802,
    ng595, ng3542, ng847, ng6005, ng1736, ng47, ng2389, ng3782, ng2638,
    ng2066, ng4258, ng5232, ng6031, ng4235, ng6073, ng3147, ng4438, ng5547,
    ng4122, ng1319, ng1612, ng5813, ng4172, ng3355, ng490, ng3457, ng2844,
    ng4709, ng1291, ng2449, ng5212, ng1830, ng6474, ng4408, ng3376, ng2907,
    ng976, ng2236, ng5659, ng6287, ng5180, ng918, ng5945, ng5517, ng4245,
    ng2246, ng1932, ng1576, ng3941, ng1744, ng3512, ng3649, ng2657, ng4933,
    ng608, ng5782, ng1886, ng1008, ng645, ng392, ng146, ng2671, ng6565,
    ng5909, ng4372, ng3155, ng5607, ng4521, ng562, ng6105, ng6466, ng6133,
    ng4291, ng3590, ng218, ng2028, ng2685, ng1802, ng3490, ng3167, ng2295,
    ng3321, ng3813, ng1205, ng2208, ng732, ng968, ng4176, ng6263, ng4540,
    ng121, ng6732, ng3554, ng749, ng5615, ng6199, ng2089, ng6144, ng3909,
    ng2917, ng2504, ng6093, ng4005, ng2331, ng6723, ng6585, ng6633, ng4555,
    ng6069, ng4567, ng1339, ng767, ng5794, ng6259, ng4405, ng3945, ng2748,
    ng2283, ng1426, ng3698, ng311, ng3057, ng1384, ng5853, ng5559, ng5905,
    ng872, ng50, ng5471, ng2169, ng5005;
  wire new_n4623_1_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_1_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_1_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_1_, new_n4639_, new_n4640_, new_n4641_, new_n4642_,
    new_n4643_1_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_1_, new_n4649_, new_n4650_, new_n4651_, new_n4652_,
    new_n4653_1_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_1_, new_n4659_, new_n4660_, new_n4661_, new_n4662_,
    new_n4663_1_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_1_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_1_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_1_, new_n4679_, new_n4680_, new_n4681_, new_n4682_1_,
    new_n4683_, new_n4685_, new_n4686_, new_n4687_1_, new_n4688_,
    new_n4689_, new_n4690_, new_n4691_1_, new_n4692_, new_n4693_,
    new_n4694_, new_n4696_1_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_1_, new_n4702_, new_n4705_, new_n4706_1_,
    new_n4707_, new_n4708_, new_n4709_, new_n4710_1_, new_n4711_,
    new_n4712_, new_n4714_1_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_1_, new_n4719_, new_n4720_, new_n4721_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_1_, new_n4728_,
    new_n4729_, new_n4730_, new_n4731_, new_n4732_1_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_1_, new_n4738_,
    new_n4739_, new_n4740_, new_n4742_1_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_1_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_1_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_1_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_1_, new_n4763_, new_n4764_,
    new_n4765_, new_n4766_, new_n4767_1_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_1_, new_n4772_, new_n4773_, new_n4774_,
    new_n4776_1_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_1_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_1_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_1_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_1_, new_n4797_, new_n4798_, new_n4799_, new_n4800_1_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_1_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_1_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_1_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_1_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_1_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_1_,
    new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_1_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_1_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_1_, new_n4848_1_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_1_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_1_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_1_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_1_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_1_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_1_, new_n4878_, new_n4879_,
    new_n4881_, new_n4882_1_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_1_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_1_, new_n4893_, new_n4894_, new_n4895_, new_n4896_1_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_1_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_1_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_1_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_1_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_1_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_1_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_1_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_1_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_1_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_1_, new_n4946_,
    new_n4947_, new_n4948_, new_n4949_, new_n4950_1_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_1_, new_n4956_,
    new_n4957_, new_n4958_, new_n4959_, new_n4960_1_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_1_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_1_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_1_, new_n4976_,
    new_n4977_, new_n4978_, new_n4979_, new_n4980_1_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_1_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_1_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_1_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_1_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_1_, new_n5006_,
    new_n5007_, new_n5008_, new_n5009_, new_n5010_1_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_1_, new_n5016_,
    new_n5018_, new_n5019_, new_n5020_1_, new_n5021_, new_n5022_,
    new_n5023_, new_n5024_, new_n5025_1_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_1_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_1_, new_n5036_, new_n5037_,
    new_n5039_, new_n5040_1_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_1_, new_n5046_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_1_, new_n5053_, new_n5055_, new_n5056_,
    new_n5058_1_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_1_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_1_, new_n5069_, new_n5070_, new_n5071_, new_n5072_,
    new_n5073_1_, new_n5074_, new_n5075_, new_n5076_, new_n5077_1_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_1_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_1_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_1_,
    new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_1_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_1_,
    new_n5103_, new_n5104_, new_n5105_, new_n5107_1_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_1_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_1_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_1_, new_n5123_, new_n5124_,
    new_n5125_, new_n5126_, new_n5127_1_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_1_, new_n5132_, new_n5133_, new_n5134_,
    new_n5135_, new_n5136_1_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_1_, new_n5142_, new_n5143_, new_n5144_,
    new_n5145_, new_n5146_1_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_1_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_1_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_1_, new_n5167_, new_n5168_, new_n5169_, new_n5170_,
    new_n5171_1_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_1_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_1_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_1_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_1_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_1_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_1_, new_n5203_, new_n5204_, new_n5205_, new_n5206_1_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_1_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_1_,
    new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_1_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5227_, new_n5228_,
    new_n5229_, new_n5230_, new_n5231_1_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_1_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_1_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_1_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_1_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_1_, new_n5255_, new_n5256_, new_n5257_, new_n5258_1_,
    new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_1_, new_n5269_, new_n5270_,
    new_n5271_, new_n5272_, new_n5273_1_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_1_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_1_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_1_, new_n5289_, new_n5290_,
    new_n5291_, new_n5292_, new_n5293_1_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_1_, new_n5299_, new_n5300_,
    new_n5302_, new_n5303_1_, new_n5304_, new_n5305_, new_n5306_,
    new_n5307_, new_n5308_1_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_1_, new_n5313_, new_n5314_, new_n5315_, new_n5316_1_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_1_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_1_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_1_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_1_, new_n5335_, new_n5336_,
    new_n5338_, new_n5339_1_, new_n5340_, new_n5341_, new_n5342_,
    new_n5343_, new_n5344_1_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_1_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_1_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_1_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_1_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_1_, new_n5369_, new_n5370_, new_n5371_, new_n5372_,
    new_n5373_1_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_1_, new_n5379_, new_n5380_, new_n5381_, new_n5383_1_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_1_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_1_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_1_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_1_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_1_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_1_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_1_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_1_, new_n5423_,
    new_n5425_, new_n5426_, new_n5427_1_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_1_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_1_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_1_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_1_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_1_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_1_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_1_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_1_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_1_, new_n5478_, new_n5479_, new_n5480_1_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_1_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_1_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_1_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_1_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_1_, new_n5506_,
    new_n5507_, new_n5508_, new_n5509_1_, new_n5510_, new_n5512_,
    new_n5513_, new_n5514_1_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_1_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_1_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_1_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_1_, new_n5534_, new_n5535_, new_n5536_, new_n5537_1_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_1_,
    new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_1_,
    new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_1_,
    new_n5553_, new_n5554_, new_n5555_, new_n5557_1_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_1_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_1_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_1_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_1_, new_n5576_, new_n5577_, new_n5578_,
    new_n5579_, new_n5580_1_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_1_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_1_, new_n5591_, new_n5593_, new_n5594_1_,
    new_n5595_, new_n5596_, new_n5597_, new_n5598_1_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_1_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5609_, new_n5611_, new_n5612_,
    new_n5613_1_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_1_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_1_, new_n5624_, new_n5625_, new_n5626_, new_n5628_1_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_1_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_1_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_1_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_1_,
    new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_1_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_1_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_1_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_1_,
    new_n5669_, new_n5670_, new_n5671_, new_n5672_1_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_1_, new_n5678_,
    new_n5679_, new_n5680_, new_n5681_, new_n5682_1_, new_n5683_,
    new_n5684_, new_n5687_1_, new_n5688_, new_n5689_, new_n5690_,
    new_n5691_, new_n5692_1_, new_n5693_, new_n5694_, new_n5696_,
    new_n5698_, new_n5700_, new_n5701_, new_n5702_1_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_1_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_1_, new_n5713_, new_n5714_,
    new_n5715_, new_n5716_, new_n5717_1_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_1_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_1_, new_n5729_, new_n5731_,
    new_n5732_1_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_1_, new_n5738_, new_n5740_, new_n5742_1_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_1_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_1_, new_n5754_,
    new_n5756_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_1_, new_n5763_, new_n5764_, new_n5765_, new_n5766_1_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_1_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_1_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_1_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_1_, new_n5786_,
    new_n5787_, new_n5788_, new_n5789_1_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_1_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_1_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_1_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_1_, new_n5810_, new_n5811_,
    new_n5812_, new_n5813_, new_n5814_1_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_1_, new_n5821_, new_n5823_,
    new_n5824_1_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_1_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_1_, new_n5836_, new_n5837_, new_n5838_1_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_1_, new_n5844_,
    new_n5845_, new_n5846_, new_n5848_1_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_1_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_1_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_1_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_1_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_1_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_1_, new_n5879_, new_n5880_, new_n5882_,
    new_n5883_1_, new_n5884_, new_n5886_, new_n5887_, new_n5888_1_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_1_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_1_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_1_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_1_, new_n5913_, new_n5914_, new_n5915_,
    new_n5917_1_, new_n5918_, new_n5920_, new_n5921_1_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_1_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_1_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_1_, new_n5936_, new_n5937_, new_n5938_,
    new_n5939_, new_n5940_1_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_1_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_1_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_1_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_1_, new_n5966_, new_n5967_, new_n5968_, new_n5969_1_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_1_, new_n5975_,
    new_n5976_, new_n5978_, new_n5979_1_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_1_, new_n5984_, new_n5985_, new_n5986_,
    new_n5988_1_, new_n5989_, new_n5990_, new_n5991_, new_n5992_,
    new_n5993_1_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_1_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_1_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_1_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_1_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_1_, new_n6019_, new_n6020_, new_n6021_, new_n6022_,
    new_n6023_1_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_1_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_1_, new_n6039_,
    new_n6040_, new_n6041_1_, new_n6042_, new_n6043_, new_n6044_,
    new_n6045_1_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_1_, new_n6052_, new_n6053_, new_n6054_, new_n6055_1_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_1_,
    new_n6061_, new_n6062_, new_n6063_, new_n6065_1_, new_n6066_,
    new_n6067_, new_n6068_, new_n6069_1_, new_n6070_, new_n6071_,
    new_n6073_, new_n6074_1_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_1_, new_n6080_, new_n6081_, new_n6082_,
    new_n6083_, new_n6084_1_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_1_, new_n6089_, new_n6090_, new_n6091_, new_n6092_1_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_1_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_1_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_1_, new_n6106_, new_n6107_,
    new_n6108_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_1_, new_n6115_, new_n6116_, new_n6118_, new_n6119_1_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_1_,
    new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_1_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_1_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_1_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_1_, new_n6151_, new_n6152_,
    new_n6154_1_, new_n6155_, new_n6156_, new_n6157_, new_n6158_,
    new_n6159_1_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_1_, new_n6165_, new_n6166_, new_n6167_, new_n6169_1_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_1_,
    new_n6175_, new_n6177_, new_n6178_, new_n6180_, new_n6181_, new_n6182_,
    new_n6183_, new_n6184_1_, new_n6185_, new_n6187_, new_n6188_1_,
    new_n6189_, new_n6190_, new_n6191_, new_n6192_1_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_1_, new_n6198_,
    new_n6199_, new_n6201_, new_n6202_1_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_1_, new_n6208_, new_n6209_,
    new_n6210_, new_n6212_1_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_1_, new_n6218_, new_n6219_, new_n6220_1_, new_n6221_,
    new_n6222_, new_n6223_, new_n6225_1_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_1_, new_n6231_, new_n6232_,
    new_n6233_, new_n6234_, new_n6235_1_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_1_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_1_, new_n6251_, new_n6252_, new_n6253_, new_n6254_,
    new_n6255_1_, new_n6257_, new_n6258_, new_n6259_, new_n6260_1_,
    new_n6261_, new_n6263_, new_n6264_, new_n6265_1_, new_n6266_,
    new_n6267_, new_n6269_, new_n6270_1_, new_n6271_, new_n6272_,
    new_n6273_, new_n6274_, new_n6275_1_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_1_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_1_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_1_, new_n6291_, new_n6293_,
    new_n6294_, new_n6295_1_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_1_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_1_, new_n6305_, new_n6306_, new_n6307_, new_n6308_1_,
    new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_1_,
    new_n6315_, new_n6316_, new_n6317_, new_n6318_1_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6324_, new_n6325_, new_n6326_,
    new_n6327_, new_n6328_1_, new_n6329_, new_n6330_, new_n6331_,
    new_n6333_1_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_1_, new_n6339_, new_n6340_, new_n6341_, new_n6343_,
    new_n6344_, new_n6346_, new_n6347_1_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_1_, new_n6353_, new_n6354_,
    new_n6355_, new_n6356_, new_n6357_1_, new_n6358_, new_n6360_,
    new_n6361_, new_n6362_1_, new_n6363_, new_n6364_, new_n6365_,
    new_n6367_1_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_1_, new_n6373_, new_n6374_, new_n6375_, new_n6376_,
    new_n6377_1_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_1_, new_n6383_, new_n6384_, new_n6385_, new_n6386_,
    new_n6387_1_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_1_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_1_, new_n6398_, new_n6400_, new_n6401_, new_n6402_1_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_1_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_1_, new_n6412_,
    new_n6413_, new_n6414_, new_n6415_, new_n6416_1_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_1_, new_n6421_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_1_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_1_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_1_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_1_, new_n6446_, new_n6447_, new_n6449_, new_n6450_1_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_1_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_1_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_1_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_1_, new_n6471_,
    new_n6472_, new_n6473_, new_n6474_, new_n6475_1_, new_n6476_,
    new_n6478_, new_n6479_, new_n6480_1_, new_n6481_, new_n6482_,
    new_n6484_, new_n6485_1_, new_n6486_, new_n6487_, new_n6488_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_1_, new_n6494_,
    new_n6495_, new_n6496_, new_n6497_, new_n6498_1_, new_n6499_,
    new_n6500_, new_n6501_, new_n6503_1_, new_n6504_, new_n6505_,
    new_n6507_, new_n6508_1_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_1_, new_n6514_, new_n6515_, new_n6516_,
    new_n6517_, new_n6518_1_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_1_, new_n6524_, new_n6525_, new_n6526_,
    new_n6527_1_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_1_, new_n6534_, new_n6535_, new_n6536_, new_n6537_1_,
    new_n6538_, new_n6539_, new_n6540_, new_n6542_1_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_1_, new_n6548_,
    new_n6549_, new_n6550_, new_n6551_, new_n6552_1_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_1_, new_n6558_,
    new_n6560_, new_n6561_, new_n6562_1_, new_n6563_, new_n6564_,
    new_n6565_, new_n6566_1_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_1_, new_n6572_, new_n6573_, new_n6575_,
    new_n6576_1_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_1_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_1_, new_n6587_, new_n6588_, new_n6589_, new_n6590_,
    new_n6591_1_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_1_, new_n6597_, new_n6598_, new_n6599_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_1_, new_n6605_, new_n6606_,
    new_n6607_, new_n6608_, new_n6609_1_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_1_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_1_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_1_, new_n6625_, new_n6626_,
    new_n6627_, new_n6628_1_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_1_, new_n6633_, new_n6634_, new_n6635_, new_n6636_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_1_,
    new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_1_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_1_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_1_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_1_, new_n6673_, new_n6674_, new_n6675_, new_n6676_,
    new_n6677_1_, new_n6679_, new_n6680_, new_n6681_, new_n6682_1_,
    new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_1_,
    new_n6688_, new_n6689_, new_n6691_1_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_1_, new_n6697_, new_n6698_,
    new_n6699_, new_n6700_, new_n6701_1_, new_n6702_, new_n6703_,
    new_n6704_, new_n6706_1_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_1_, new_n6712_, new_n6713_, new_n6714_,
    new_n6715_, new_n6716_1_, new_n6718_, new_n6719_, new_n6720_,
    new_n6721_1_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_1_, new_n6727_, new_n6728_, new_n6730_, new_n6731_1_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_1_,
    new_n6737_, new_n6739_, new_n6740_, new_n6741_1_, new_n6742_,
    new_n6743_, new_n6745_, new_n6746_1_, new_n6747_, new_n6748_,
    new_n6751_1_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_1_, new_n6757_, new_n6758_, new_n6760_, new_n6761_1_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_1_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_1_, new_n6772_,
    new_n6773_, new_n6774_, new_n6776_1_, new_n6777_, new_n6778_,
    new_n6779_, new_n6780_, new_n6781_1_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_1_, new_n6787_, new_n6788_,
    new_n6790_, new_n6791_1_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_1_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_1_, new_n6807_, new_n6808_, new_n6809_, new_n6810_1_,
    new_n6811_, new_n6812_, new_n6813_, new_n6814_1_, new_n6815_,
    new_n6816_, new_n6817_, new_n6819_1_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_1_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_1_, new_n6830_, new_n6831_, new_n6832_,
    new_n6833_, new_n6834_1_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_1_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_1_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_1_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_1_, new_n6855_, new_n6856_, new_n6857_, new_n6859_1_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_1_, new_n6864_,
    new_n6865_, new_n6867_, new_n6868_1_, new_n6869_, new_n6870_,
    new_n6871_, new_n6873_1_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_1_, new_n6879_, new_n6881_, new_n6882_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_1_,
    new_n6889_, new_n6890_, new_n6891_, new_n6893_1_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_1_, new_n6899_,
    new_n6900_, new_n6901_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_1_, new_n6908_, new_n6909_, new_n6911_, new_n6912_1_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_1_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_1_, new_n6922_,
    new_n6923_, new_n6924_, new_n6925_, new_n6926_1_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_1_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_1_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_1_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_1_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_1_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_1_, new_n6957_,
    new_n6958_, new_n6959_, new_n6960_, new_n6961_1_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_1_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_1_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_1_, new_n6977_,
    new_n6978_, new_n6979_, new_n6980_, new_n6981_1_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_1_, new_n6987_,
    new_n6988_, new_n6989_, new_n6990_, new_n6991_1_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_1_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_1_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_1_, new_n7007_,
    new_n7009_, new_n7010_, new_n7011_1_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7017_, new_n7018_, new_n7019_1_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_1_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_1_, new_n7028_, new_n7029_,
    new_n7030_, new_n7031_1_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_1_, new_n7042_, new_n7043_, new_n7044_, new_n7046_1_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_1_, new_n7051_,
    new_n7052_, new_n7053_, new_n7055_1_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_1_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_1_, new_n7072_, new_n7073_, new_n7074_, new_n7075_1_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_1_,
    new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_1_, new_n7090_, new_n7091_, new_n7092_,
    new_n7093_1_, new_n7095_, new_n7096_, new_n7097_, new_n7098_1_,
    new_n7099_, new_n7100_, new_n7101_, new_n7103_1_, new_n7104_,
    new_n7105_, new_n7106_, new_n7107_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_1_, new_n7114_, new_n7115_, new_n7117_,
    new_n7118_1_, new_n7119_, new_n7120_, new_n7121_, new_n7123_1_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_1_,
    new_n7129_, new_n7130_, new_n7132_, new_n7133_1_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_1_, new_n7144_, new_n7146_, new_n7147_,
    new_n7148_1_, new_n7150_, new_n7151_, new_n7152_, new_n7153_1_,
    new_n7154_, new_n7155_, new_n7156_, new_n7158_1_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_1_, new_n7164_,
    new_n7166_, new_n7167_, new_n7168_1_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_1_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_1_, new_n7179_, new_n7180_,
    new_n7181_, new_n7182_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_1_, new_n7189_, new_n7190_, new_n7191_, new_n7192_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_1_,
    new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_1_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_1_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_1_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_1_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_1_, new_n7223_, new_n7225_,
    new_n7226_, new_n7227_1_, new_n7228_, new_n7229_, new_n7230_,
    new_n7231_, new_n7232_1_, new_n7233_, new_n7234_, new_n7235_,
    new_n7237_1_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_1_, new_n7243_, new_n7244_, new_n7245_, new_n7246_,
    new_n7247_1_, new_n7248_, new_n7249_, new_n7251_, new_n7252_1_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_1_, new_n7258_,
    new_n7259_, new_n7260_, new_n7261_, new_n7262_1_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_1_, new_n7267_, new_n7268_,
    new_n7271_1_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7277_, new_n7278_, new_n7279_, new_n7280_1_, new_n7281_,
    new_n7282_, new_n7284_1_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_1_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_1_, new_n7295_, new_n7296_, new_n7298_,
    new_n7299_1_, new_n7301_, new_n7302_, new_n7303_, new_n7304_1_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_1_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_1_,
    new_n7315_, new_n7316_, new_n7318_, new_n7319_1_, new_n7320_,
    new_n7321_, new_n7322_, new_n7323_, new_n7324_1_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_1_, new_n7330_,
    new_n7332_, new_n7333_, new_n7334_1_, new_n7335_, new_n7336_,
    new_n7337_, new_n7338_, new_n7339_1_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_1_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_1_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_1_, new_n7355_, new_n7356_,
    new_n7357_, new_n7359_1_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_1_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_1_, new_n7375_, new_n7377_, new_n7378_, new_n7379_1_,
    new_n7380_, new_n7381_, new_n7382_, new_n7384_, new_n7385_, new_n7386_,
    new_n7388_1_, new_n7389_, new_n7390_, new_n7391_, new_n7392_1_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_1_, new_n7403_, new_n7404_,
    new_n7406_, new_n7407_1_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_1_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_1_, new_n7418_, new_n7419_, new_n7420_,
    new_n7421_, new_n7422_1_, new_n7424_, new_n7425_, new_n7426_1_,
    new_n7427_, new_n7428_, new_n7429_, new_n7430_1_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_1_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_1_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_1_, new_n7446_, new_n7448_,
    new_n7449_, new_n7450_1_, new_n7451_, new_n7452_, new_n7453_,
    new_n7455_1_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_1_, new_n7461_, new_n7463_, new_n7464_, new_n7466_,
    new_n7467_, new_n7468_, new_n7470_1_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_1_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_1_, new_n7481_, new_n7483_,
    new_n7484_, new_n7485_1_, new_n7487_, new_n7488_, new_n7490_1_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_1_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_1_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_1_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_1_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_1_, new_n7520_, new_n7521_, new_n7522_,
    new_n7523_, new_n7524_1_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_1_, new_n7530_, new_n7531_, new_n7533_1_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_1_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_1_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_1_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_1_, new_n7557_, new_n7558_, new_n7559_, new_n7560_,
    new_n7561_1_, new_n7562_, new_n7563_, new_n7565_, new_n7566_1_,
    new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_1_,
    new_n7573_, new_n7574_, new_n7575_, new_n7576_1_, new_n7577_,
    new_n7579_, new_n7580_1_, new_n7581_, new_n7582_, new_n7583_,
    new_n7584_1_, new_n7585_, new_n7586_, new_n7588_, new_n7589_1_,
    new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7595_, new_n7596_,
    new_n7597_, new_n7598_, new_n7599_1_, new_n7601_, new_n7602_,
    new_n7603_1_, new_n7604_, new_n7605_, new_n7606_, new_n7607_1_,
    new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_1_,
    new_n7614_, new_n7615_, new_n7616_, new_n7617_1_, new_n7618_,
    new_n7619_, new_n7621_, new_n7622_1_, new_n7623_, new_n7624_,
    new_n7625_, new_n7627_1_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_1_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7638_, new_n7639_, new_n7640_, new_n7641_1_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_1_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_1_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_1_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7696_, new_n7697_, new_n7698_,
    new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7757_, new_n7758_,
    new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_,
    new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7864_, new_n7865_, new_n7866_,
    new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8017_, new_n8018_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8066_,
    new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_,
    new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_,
    new_n8133_, new_n8134_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8182_, new_n8183_, new_n8184_,
    new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8282_,
    new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8316_,
    new_n8317_, new_n8319_, new_n8320_, new_n8321_, new_n8323_, new_n8324_,
    new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8330_, new_n8331_,
    new_n8332_, new_n8333_, new_n8334_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8379_,
    new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8427_, new_n8428_, new_n8429_, new_n8431_, new_n8432_, new_n8433_,
    new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8439_, new_n8440_,
    new_n8441_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8470_, new_n8471_, new_n8472_, new_n8473_,
    new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8479_, new_n8480_,
    new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_,
    new_n8487_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8497_, new_n8498_, new_n8499_, new_n8500_,
    new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_,
    new_n8507_, new_n8508_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8525_, new_n8526_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8532_, new_n8533_, new_n8534_,
    new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_,
    new_n8541_, new_n8542_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_,
    new_n8601_, new_n8602_, new_n8603_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8645_, new_n8646_, new_n8647_, new_n8648_,
    new_n8649_, new_n8650_, new_n8651_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8711_, new_n8712_, new_n8713_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8720_, new_n8721_, new_n8722_,
    new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_,
    new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_,
    new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8741_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8765_, new_n8766_, new_n8767_, new_n8769_,
    new_n8770_, new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_,
    new_n8777_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8803_, new_n8804_,
    new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8821_, new_n8822_, new_n8823_, new_n8824_,
    new_n8825_, new_n8826_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8845_,
    new_n8846_, new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_,
    new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_,
    new_n8859_, new_n8861_, new_n8862_, new_n8864_, new_n8865_, new_n8866_,
    new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8896_, new_n8897_, new_n8899_, new_n8900_,
    new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_,
    new_n8907_, new_n8908_, new_n8909_, new_n8911_, new_n8912_, new_n8913_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8923_, new_n8924_, new_n8926_, new_n8927_, new_n8928_,
    new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8961_, new_n8962_, new_n8964_, new_n8965_, new_n8966_,
    new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_,
    new_n8999_, new_n9000_, new_n9003_, new_n9004_, new_n9005_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9023_, new_n9024_, new_n9025_, new_n9026_,
    new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9038_, new_n9039_, new_n9040_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_,
    new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_,
    new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_,
    new_n9101_, new_n9102_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9151_, new_n9152_, new_n9153_, new_n9154_,
    new_n9155_, new_n9156_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9162_, new_n9163_, new_n9164_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9196_, new_n9197_, new_n9199_, new_n9200_, new_n9201_, new_n9202_,
    new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9209_,
    new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_,
    new_n9216_, new_n9217_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_,
    new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_,
    new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_,
    new_n9269_, new_n9270_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9286_, new_n9287_, new_n9288_, new_n9290_,
    new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_,
    new_n9311_, new_n9312_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9337_, new_n9338_,
    new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_,
    new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_,
    new_n9365_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9375_, new_n9376_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9385_, new_n9386_,
    new_n9387_, new_n9388_, new_n9389_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9427_, new_n9428_,
    new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9462_,
    new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9480_, new_n9481_, new_n9482_,
    new_n9483_, new_n9484_, new_n9485_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9529_, new_n9530_, new_n9531_, new_n9532_,
    new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_,
    new_n9539_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9563_, new_n9564_, new_n9565_, new_n9566_,
    new_n9567_, new_n9568_, new_n9569_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9580_,
    new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9603_, new_n9604_, new_n9605_, new_n9607_, new_n9608_,
    new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_,
    new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9800_,
    new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_,
    new_n9833_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9843_, new_n9844_, new_n9845_, new_n9846_,
    new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9858_, new_n9859_, new_n9860_,
    new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9873_, new_n9874_,
    new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9891_, new_n9892_, new_n9893_, new_n9894_,
    new_n9895_, new_n9896_, new_n9897_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_,
    new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_,
    new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_,
    new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_,
    new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10042_, new_n10043_, new_n10044_, new_n10045_, new_n10046_,
    new_n10047_, new_n10048_, new_n10050_, new_n10051_, new_n10052_,
    new_n10053_, new_n10054_, new_n10055_, new_n10056_, new_n10058_,
    new_n10059_, new_n10060_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10079_, new_n10080_, new_n10081_,
    new_n10082_, new_n10083_, new_n10084_, new_n10085_, new_n10086_,
    new_n10087_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10097_, new_n10098_,
    new_n10099_, new_n10100_, new_n10101_, new_n10102_, new_n10103_,
    new_n10104_, new_n10105_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10123_, new_n10124_, new_n10125_, new_n10126_,
    new_n10127_, new_n10128_, new_n10129_, new_n10130_, new_n10131_,
    new_n10133_, new_n10134_, new_n10135_, new_n10136_, new_n10137_,
    new_n10138_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10185_, new_n10186_,
    new_n10187_, new_n10188_, new_n10189_, new_n10190_, new_n10191_,
    new_n10192_, new_n10193_, new_n10194_, new_n10195_, new_n10196_,
    new_n10197_, new_n10198_, new_n10199_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10205_, new_n10207_, new_n10208_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10311_,
    new_n10312_, new_n10313_, new_n10315_, new_n10316_, new_n10317_,
    new_n10318_, new_n10319_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10338_, new_n10339_, new_n10340_, new_n10342_,
    new_n10343_, new_n10344_, new_n10345_, new_n10346_, new_n10347_,
    new_n10348_, new_n10349_, new_n10351_, new_n10352_, new_n10353_,
    new_n10354_, new_n10355_, new_n10356_, new_n10357_, new_n10358_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10378_, new_n10379_, new_n10380_, new_n10381_,
    new_n10382_, new_n10384_, new_n10385_, new_n10387_, new_n10388_,
    new_n10389_, new_n10390_, new_n10391_, new_n10392_, new_n10393_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10409_, new_n10410_, new_n10411_,
    new_n10412_, new_n10413_, new_n10414_, new_n10416_, new_n10417_,
    new_n10418_, new_n10419_, new_n10420_, new_n10422_, new_n10423_,
    new_n10424_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10446_,
    new_n10447_, new_n10448_, new_n10449_, new_n10450_, new_n10451_,
    new_n10452_, new_n10454_, new_n10455_, new_n10456_, new_n10457_,
    new_n10458_, new_n10459_, new_n10460_, new_n10461_, new_n10462_,
    new_n10464_, new_n10465_, new_n10466_, new_n10467_, new_n10468_,
    new_n10469_, new_n10470_, new_n10471_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10500_, new_n10501_,
    new_n10502_, new_n10503_, new_n10505_, new_n10506_, new_n10507_,
    new_n10508_, new_n10509_, new_n10510_, new_n10511_, new_n10512_,
    new_n10513_, new_n10514_, new_n10516_, new_n10517_, new_n10518_,
    new_n10519_, new_n10520_, new_n10521_, new_n10522_, new_n10523_,
    new_n10524_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10548_, new_n10549_, new_n10550_, new_n10551_, new_n10552_,
    new_n10553_, new_n10555_, new_n10556_, new_n10557_, new_n10558_,
    new_n10559_, new_n10560_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10580_, new_n10581_, new_n10582_,
    new_n10583_, new_n10584_, new_n10585_, new_n10587_, new_n10588_,
    new_n10589_, new_n10590_, new_n10591_, new_n10592_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10622_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10628_,
    new_n10629_, new_n10630_, new_n10631_, new_n10632_, new_n10633_,
    new_n10634_, new_n10635_, new_n10636_, new_n10637_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10666_, new_n10667_,
    new_n10668_, new_n10669_, new_n10670_, new_n10671_, new_n10673_,
    new_n10674_, new_n10675_, new_n10676_, new_n10677_, new_n10678_,
    new_n10679_, new_n10680_, new_n10681_, new_n10682_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10702_,
    new_n10703_, new_n10704_, new_n10705_, new_n10706_, new_n10707_,
    new_n10708_, new_n10709_, new_n10711_, new_n10712_, new_n10713_,
    new_n10714_, new_n10715_, new_n10716_, new_n10717_, new_n10718_,
    new_n10719_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10758_,
    new_n10759_, new_n10760_, new_n10761_, new_n10762_, new_n10764_,
    new_n10765_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10802_, new_n10803_,
    new_n10804_, new_n10805_, new_n10806_, new_n10807_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10824_, new_n10825_, new_n10826_,
    new_n10827_, new_n10828_, new_n10829_, new_n10830_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10844_, new_n10845_, new_n10846_, new_n10847_, new_n10848_,
    new_n10849_, new_n10850_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10869_, new_n10870_, new_n10871_,
    new_n10872_, new_n10873_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10881_, new_n10882_, new_n10883_,
    new_n10884_, new_n10885_, new_n10886_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10900_, new_n10901_,
    new_n10902_, new_n10903_, new_n10904_, new_n10905_, new_n10907_,
    new_n10908_, new_n10909_, new_n10910_, new_n10911_, new_n10912_,
    new_n10913_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10949_, new_n10950_, new_n10951_, new_n10952_,
    new_n10954_, new_n10955_, new_n10956_, new_n10957_, new_n10958_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10975_,
    new_n10976_, new_n10977_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10988_, new_n10989_, new_n10990_, new_n10991_, new_n10992_,
    new_n10993_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11025_, new_n11026_, new_n11027_,
    new_n11028_, new_n11029_, new_n11030_, new_n11031_, new_n11032_,
    new_n11033_, new_n11034_, new_n11035_, new_n11036_, new_n11038_,
    new_n11039_, new_n11040_, new_n11041_, new_n11042_, new_n11043_,
    new_n11044_, new_n11045_, new_n11046_, new_n11048_, new_n11049_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11093_,
    new_n11094_, new_n11095_, new_n11096_, new_n11097_, new_n11098_,
    new_n11099_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11125_, new_n11126_, new_n11127_,
    new_n11129_, new_n11130_, new_n11131_, new_n11132_, new_n11133_,
    new_n11134_, new_n11135_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11177_,
    new_n11178_, new_n11179_, new_n11180_, new_n11181_, new_n11182_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11189_, new_n11190_, new_n11191_, new_n11192_, new_n11193_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11228_,
    new_n11229_, new_n11230_, new_n11231_, new_n11232_, new_n11233_,
    new_n11234_, new_n11235_, new_n11236_, new_n11237_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11270_, new_n11272_, new_n11273_,
    new_n11274_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11309_, new_n11310_, new_n11311_, new_n11312_, new_n11313_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11349_, new_n11350_, new_n11352_, new_n11353_, new_n11354_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11384_, new_n11385_, new_n11386_, new_n11387_, new_n11388_,
    new_n11389_, new_n11390_, new_n11391_, new_n11392_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11413_, new_n11414_, new_n11415_, new_n11416_, new_n11417_,
    new_n11418_, new_n11420_, new_n11421_, new_n11422_, new_n11423_,
    new_n11424_, new_n11425_, new_n11426_, new_n11427_, new_n11428_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11455_, new_n11456_, new_n11457_,
    new_n11459_, new_n11460_, new_n11461_, new_n11462_, new_n11463_,
    new_n11464_, new_n11466_, new_n11467_, new_n11468_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11476_,
    new_n11477_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11485_, new_n11486_, new_n11487_, new_n11488_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11517_, new_n11518_,
    new_n11519_, new_n11520_, new_n11521_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11536_,
    new_n11537_, new_n11538_, new_n11539_, new_n11540_, new_n11541_,
    new_n11542_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11551_, new_n11552_, new_n11553_,
    new_n11554_, new_n11555_, new_n11556_, new_n11557_, new_n11558_,
    new_n11559_, new_n11560_, new_n11562_, new_n11563_, new_n11564_,
    new_n11565_, new_n11566_, new_n11567_, new_n11568_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11576_,
    new_n11577_, new_n11578_, new_n11579_, new_n11580_, new_n11581_,
    new_n11582_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11592_, new_n11593_,
    new_n11594_, new_n11595_, new_n11596_, new_n11597_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11623_, new_n11624_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11632_, new_n11633_, new_n11634_,
    new_n11635_, new_n11636_, new_n11637_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11658_,
    new_n11659_, new_n11660_, new_n11661_, new_n11662_, new_n11663_,
    new_n11664_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11677_, new_n11678_, new_n11679_, new_n11680_, new_n11681_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11690_, new_n11691_, new_n11692_, new_n11693_,
    new_n11694_, new_n11695_, new_n11697_, new_n11698_, new_n11699_,
    new_n11700_, new_n11701_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11728_,
    new_n11729_, new_n11730_, new_n11731_, new_n11732_, new_n11733_,
    new_n11734_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11772_, new_n11773_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11796_, new_n11797_, new_n11798_,
    new_n11799_, new_n11800_, new_n11801_, new_n11802_, new_n11803_,
    new_n11804_, new_n11805_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11822_, new_n11823_, new_n11824_, new_n11826_,
    new_n11827_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11899_, new_n11900_, new_n11901_,
    new_n11902_, new_n11903_, new_n11904_, new_n11905_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11949_, new_n11950_, new_n11951_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11976_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11997_, new_n11998_, new_n11999_,
    new_n12000_, new_n12001_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12023_, new_n12024_, new_n12025_, new_n12026_, new_n12027_,
    new_n12028_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12037_, new_n12038_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12075_, new_n12076_, new_n12077_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12127_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12149_, new_n12150_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12171_, new_n12172_, new_n12173_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12184_, new_n12185_, new_n12186_,
    new_n12187_, new_n12188_, new_n12189_, new_n12190_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12222_, new_n12224_, new_n12225_, new_n12226_,
    new_n12227_, new_n12228_, new_n12229_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12239_, new_n12240_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12248_, new_n12249_, new_n12251_,
    new_n12252_, new_n12253_, new_n12254_, new_n12255_, new_n12256_,
    new_n12257_, new_n12258_, new_n12259_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12294_, new_n12295_, new_n12296_,
    new_n12297_, new_n12298_, new_n12299_, new_n12300_, new_n12301_,
    new_n12302_, new_n12303_, new_n12304_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12384_, new_n12385_, new_n12386_,
    new_n12387_, new_n12388_, new_n12389_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12421_,
    new_n12422_, new_n12423_, new_n12424_, new_n12425_, new_n12426_,
    new_n12427_, new_n12428_, new_n12429_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12463_, new_n12464_, new_n12465_, new_n12466_,
    new_n12467_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12498_, new_n12499_, new_n12500_, new_n12501_,
    new_n12502_, new_n12503_, new_n12504_, new_n12505_, new_n12506_,
    new_n12507_, new_n12508_, new_n12509_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12523_,
    new_n12524_, new_n12525_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12539_, new_n12540_, new_n12541_,
    new_n12542_, new_n12543_, new_n12544_, new_n12546_, new_n12547_,
    new_n12548_, new_n12549_, new_n12550_, new_n12551_, new_n12552_,
    new_n12553_, new_n12554_, new_n12555_, new_n12556_, new_n12557_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12587_, new_n12588_, new_n12589_, new_n12590_, new_n12591_,
    new_n12592_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12599_, new_n12600_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12609_,
    new_n12610_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12637_, new_n12638_,
    new_n12639_, new_n12640_, new_n12641_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12664_, new_n12665_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12674_, new_n12675_, new_n12676_, new_n12677_, new_n12678_,
    new_n12679_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12693_, new_n12694_, new_n12695_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12734_, new_n12735_, new_n12736_, new_n12737_, new_n12738_,
    new_n12739_, new_n12740_, new_n12741_, new_n12742_, new_n12743_,
    new_n12744_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12769_, new_n12770_, new_n12771_,
    new_n12772_, new_n12773_, new_n12774_, new_n12775_, new_n12776_,
    new_n12777_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12786_, new_n12787_, new_n12788_,
    new_n12789_, new_n12790_, new_n12791_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12809_, new_n12810_, new_n12811_,
    new_n12812_, new_n12813_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12850_, new_n12851_,
    new_n12852_, new_n12853_, new_n12854_, new_n12855_, new_n12857_,
    new_n12858_, new_n12859_, new_n12860_, new_n12861_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12884_, new_n12885_, new_n12886_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12918_, new_n12919_, new_n12920_, new_n12922_,
    new_n12923_, new_n12924_, new_n12925_, new_n12926_, new_n12927_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12955_, new_n12956_,
    new_n12957_, new_n12958_, new_n12959_, new_n12960_, new_n12961_,
    new_n12963_, new_n12964_, new_n12965_, new_n12966_, new_n12967_,
    new_n12968_, new_n12969_, new_n12970_, new_n12971_, new_n12973_,
    new_n12974_, new_n12975_, new_n12976_, new_n12977_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13077_, new_n13078_, new_n13079_, new_n13080_, new_n13081_,
    new_n13082_, new_n13084_, new_n13085_, new_n13086_, new_n13087_,
    new_n13088_, new_n13090_, new_n13091_, new_n13092_, new_n13093_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13113_, new_n13114_, new_n13115_, new_n13116_,
    new_n13117_, new_n13119_, new_n13120_, new_n13121_, new_n13122_,
    new_n13123_, new_n13124_, new_n13125_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13134_, new_n13135_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13141_, new_n13142_,
    new_n13143_, new_n13144_, new_n13145_, new_n13146_, new_n13147_,
    new_n13148_, new_n13149_, new_n13150_, new_n13151_, new_n13152_,
    new_n13153_, new_n13154_, new_n13155_, new_n13156_, new_n13157_,
    new_n13158_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13168_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13176_, new_n13178_, new_n13179_, new_n13180_, new_n13181_,
    new_n13182_, new_n13184_, new_n13185_, new_n13186_, new_n13187_,
    new_n13188_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13213_, new_n13214_, new_n13215_, new_n13216_,
    new_n13217_, new_n13218_, new_n13219_, new_n13221_, new_n13222_,
    new_n13223_, new_n13224_, new_n13225_, new_n13226_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13234_,
    new_n13235_, new_n13236_, new_n13237_, new_n13238_, new_n13239_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13247_, new_n13248_, new_n13250_, new_n13251_, new_n13252_,
    new_n13253_, new_n13254_, new_n13255_, new_n13256_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13264_,
    new_n13265_, new_n13266_, new_n13267_, new_n13268_, new_n13269_,
    new_n13270_, new_n13271_, new_n13272_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13280_, new_n13281_,
    new_n13283_, new_n13284_, new_n13285_, new_n13286_, new_n13287_,
    new_n13288_, new_n13289_, new_n13290_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13298_, new_n13299_,
    new_n13300_, new_n13301_, new_n13302_, new_n13303_, new_n13305_,
    new_n13306_, new_n13307_, new_n13309_, new_n13310_, new_n13311_,
    new_n13312_, new_n13313_, new_n13314_, new_n13315_, new_n13316_,
    new_n13318_, new_n13319_, new_n13320_, new_n13321_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13355_, new_n13356_, new_n13357_,
    new_n13358_, new_n13359_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13385_, new_n13386_,
    new_n13387_, new_n13388_, new_n13389_, new_n13390_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13396_, new_n13397_,
    new_n13398_, new_n13399_, new_n13400_, new_n13401_, new_n13402_,
    new_n13403_, new_n13404_, new_n13405_, new_n13406_, new_n13407_,
    new_n13408_, new_n13410_, new_n13411_, new_n13412_, new_n13413_,
    new_n13414_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13431_,
    new_n13432_, new_n13433_, new_n13435_, new_n13436_, new_n13437_,
    new_n13438_, new_n13439_, new_n13440_, new_n13441_, new_n13443_,
    new_n13444_, new_n13445_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13461_,
    new_n13462_, new_n13463_, new_n13465_, new_n13466_, new_n13467_,
    new_n13468_, new_n13469_, new_n13470_, new_n13471_, new_n13473_,
    new_n13474_, new_n13475_, new_n13476_, new_n13477_, new_n13478_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13502_,
    new_n13503_, new_n13504_, new_n13505_, new_n13506_, new_n13508_,
    new_n13509_, new_n13510_, new_n13511_, new_n13512_, new_n13513_,
    new_n13514_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13541_, new_n13542_,
    new_n13543_, new_n13544_, new_n13545_, new_n13546_, new_n13547_,
    new_n13548_, new_n13549_, new_n13550_, new_n13551_, new_n13552_,
    new_n13553_, new_n13554_, new_n13555_, new_n13556_, new_n13557_,
    new_n13558_, new_n13559_, new_n13560_, new_n13562_, new_n13563_,
    new_n13564_, new_n13565_, new_n13566_, new_n13567_, new_n13568_,
    new_n13569_, new_n13570_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13606_, new_n13607_,
    new_n13608_, new_n13609_, new_n13610_, new_n13611_, new_n13612_,
    new_n13614_, new_n13615_, new_n13616_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13625_,
    new_n13626_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13647_,
    new_n13649_, new_n13650_, new_n13651_, new_n13652_, new_n13653_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13674_, new_n13675_, new_n13676_, new_n13677_,
    new_n13678_, new_n13680_, new_n13681_, new_n13682_, new_n13683_,
    new_n13684_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13715_, new_n13716_, new_n13717_,
    new_n13718_, new_n13719_, new_n13720_, new_n13722_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13745_, new_n13746_, new_n13747_,
    new_n13748_, new_n13749_, new_n13750_, new_n13752_, new_n13753_,
    new_n13754_, new_n13755_, new_n13756_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13784_, new_n13785_, new_n13786_, new_n13787_,
    new_n13788_, new_n13789_, new_n13791_, new_n13792_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13811_,
    new_n13812_, new_n13813_, new_n13815_, new_n13816_, new_n13817_,
    new_n13818_, new_n13819_, new_n13820_, new_n13821_, new_n13823_,
    new_n13824_, new_n13825_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13848_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13856_, new_n13857_, new_n13858_,
    new_n13859_, new_n13860_, new_n13861_, new_n13862_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13880_, new_n13882_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13891_, new_n13892_, new_n13893_,
    new_n13894_, new_n13895_, new_n13898_, new_n13899_, new_n13901_,
    new_n13902_, new_n13904_, new_n13905_, new_n13906_, new_n13907_,
    new_n13908_, new_n13909_, new_n13910_, new_n13912_, new_n13913_,
    new_n13914_, new_n13915_, new_n13916_, new_n13917_, new_n13918_,
    new_n13919_, new_n13920_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13940_, new_n13941_, new_n13942_,
    new_n13943_, new_n13944_, new_n13945_, new_n13947_, new_n13948_,
    new_n13949_, new_n13950_, new_n13951_, new_n13953_, new_n13954_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13989_, new_n13990_, new_n13991_, new_n13992_, new_n13993_,
    new_n13994_, new_n13995_, new_n13996_, new_n13997_, new_n13998_,
    new_n14000_, new_n14001_, new_n14002_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14032_, new_n14033_,
    new_n14034_, new_n14035_, new_n14036_, new_n14038_, new_n14039_,
    new_n14040_, new_n14041_, new_n14042_, new_n14043_, new_n14044_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14067_, new_n14068_,
    new_n14069_, new_n14070_, new_n14071_, new_n14073_, new_n14074_,
    new_n14075_, new_n14076_, new_n14077_, new_n14078_, new_n14079_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14098_,
    new_n14099_, new_n14100_, new_n14101_, new_n14102_, new_n14103_,
    new_n14105_, new_n14106_, new_n14107_, new_n14108_, new_n14109_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14133_,
    new_n14134_, new_n14135_, new_n14136_, new_n14137_, new_n14139_,
    new_n14140_, new_n14141_, new_n14142_, new_n14143_, new_n14144_,
    new_n14145_, new_n14146_, new_n14148_, new_n14149_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14158_, new_n14159_, new_n14160_, new_n14161_, new_n14162_,
    new_n14163_, new_n14164_, new_n14165_, new_n14166_, new_n14167_,
    new_n14168_, new_n14169_, new_n14171_, new_n14172_, new_n14173_,
    new_n14174_, new_n14175_, new_n14176_, new_n14177_, new_n14178_,
    new_n14179_, new_n14180_, new_n14181_, new_n14182_, new_n14183_,
    new_n14184_, new_n14185_, new_n14186_, new_n14187_, new_n14188_,
    new_n14189_, new_n14190_, new_n14192_, new_n14193_, new_n14194_,
    new_n14195_, new_n14196_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14212_,
    new_n14213_, new_n14214_, new_n14215_, new_n14216_, new_n14218_,
    new_n14219_, new_n14220_, new_n14221_, new_n14222_, new_n14223_,
    new_n14224_, new_n14225_, new_n14227_, new_n14228_, new_n14229_,
    new_n14230_, new_n14231_, new_n14232_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14248_, new_n14249_, new_n14251_, new_n14252_, new_n14254_,
    new_n14255_, new_n14256_, new_n14257_, new_n14258_, new_n14259_,
    new_n14260_, new_n14261_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14285_, new_n14286_, new_n14287_, new_n14289_,
    new_n14290_, new_n14291_, new_n14292_, new_n14293_, new_n14294_,
    new_n14295_, new_n14296_, new_n14297_, new_n14298_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14307_, new_n14308_, new_n14309_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14325_, new_n14326_, new_n14327_, new_n14328_, new_n14329_,
    new_n14330_, new_n14331_, new_n14332_, new_n14333_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14363_, new_n14364_,
    new_n14365_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14395_, new_n14396_, new_n14397_, new_n14398_, new_n14399_,
    new_n14400_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14436_, new_n14437_, new_n14438_, new_n14439_,
    new_n14440_, new_n14441_, new_n14442_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14466_, new_n14467_, new_n14468_,
    new_n14469_, new_n14470_, new_n14471_, new_n14472_, new_n14474_,
    new_n14475_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14488_, new_n14489_, new_n14490_, new_n14491_, new_n14492_,
    new_n14493_, new_n14494_, new_n14495_, new_n14498_, new_n14499_,
    new_n14500_, new_n14501_, new_n14502_, new_n14503_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14520_, new_n14521_, new_n14522_, new_n14523_,
    new_n14524_, new_n14525_, new_n14527_, new_n14528_, new_n14529_,
    new_n14530_, new_n14531_, new_n14532_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14541_,
    new_n14542_, new_n14543_, new_n14545_, new_n14546_, new_n14548_,
    new_n14549_, new_n14550_, new_n14551_, new_n14552_, new_n14553_,
    new_n14554_, new_n14556_, new_n14557_, new_n14558_, new_n14559_,
    new_n14560_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14576_, new_n14577_,
    new_n14578_, new_n14579_, new_n14580_, new_n14581_, new_n14583_,
    new_n14584_, new_n14585_, new_n14586_, new_n14587_, new_n14588_,
    new_n14590_, new_n14591_, new_n14592_, new_n14593_, new_n14594_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14628_,
    new_n14629_, new_n14630_, new_n14631_, new_n14632_, new_n14634_,
    new_n14635_, new_n14636_, new_n14637_, new_n14638_, new_n14639_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14647_, new_n14648_, new_n14649_, new_n14650_, new_n14651_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14661_, new_n14662_, new_n14663_,
    new_n14664_, new_n14665_, new_n14666_, new_n14667_, new_n14669_,
    new_n14670_, new_n14671_, new_n14672_, new_n14673_, new_n14674_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14682_, new_n14683_, new_n14684_, new_n14685_, new_n14686_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14694_,
    new_n14695_, new_n14696_, new_n14697_, new_n14698_, new_n14699_,
    new_n14701_, new_n14702_, new_n14704_, new_n14705_, new_n14706_,
    new_n14707_, new_n14708_, new_n14709_, new_n14710_, new_n14711_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14720_, new_n14721_, new_n14722_, new_n14723_,
    new_n14724_, new_n14725_, new_n14726_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14733_, new_n14734_,
    new_n14735_, new_n14736_, new_n14737_, new_n14738_, new_n14739_,
    new_n14740_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14764_, new_n14765_, new_n14766_, new_n14767_, new_n14768_,
    new_n14769_, new_n14770_, new_n14771_, new_n14773_, new_n14774_,
    new_n14775_, new_n14776_, new_n14777_, new_n14778_, new_n14779_,
    new_n14780_, new_n14781_, new_n14782_, new_n14783_, new_n14784_,
    new_n14785_, new_n14786_, new_n14787_, new_n14788_, new_n14789_,
    new_n14790_, new_n14791_, new_n14792_, new_n14793_, new_n14794_,
    new_n14795_, new_n14796_, new_n14797_, new_n14798_, new_n14799_,
    new_n14800_, new_n14801_, new_n14802_, new_n14803_, new_n14804_,
    new_n14805_, new_n14806_, new_n14807_, new_n14808_, new_n14809_,
    new_n14810_, new_n14811_, new_n14812_, new_n14813_, new_n14814_,
    new_n14815_, new_n14816_, new_n14817_, new_n14818_, new_n14819_,
    new_n14820_, new_n14821_, new_n14822_, new_n14823_, new_n14824_,
    new_n14825_, new_n14826_, new_n14827_, new_n14828_, new_n14829_,
    new_n14830_, new_n14831_, new_n14832_, new_n14833_, new_n14834_,
    new_n14835_, new_n14836_, new_n14837_, new_n14838_, new_n14839_,
    new_n14840_, new_n14841_, new_n14842_, new_n14843_, new_n14844_,
    new_n14845_, new_n14846_, new_n14847_, new_n14848_, new_n14849_,
    new_n14850_, new_n14851_, new_n14852_, new_n14853_, new_n14854_,
    new_n14855_, new_n14856_, new_n14857_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14872_,
    new_n14873_, new_n14874_, new_n14875_, new_n14876_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14886_, new_n14887_, new_n14888_, new_n14889_,
    new_n14890_, new_n14891_, new_n14892_, new_n14893_, new_n14894_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14910_, new_n14911_, new_n14912_,
    new_n14913_, new_n14914_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14923_, new_n14924_,
    new_n14925_, new_n14926_, new_n14927_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14942_,
    new_n14943_, new_n14944_, new_n14945_, new_n14946_, new_n14947_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14974_, new_n14975_, new_n14976_,
    new_n14978_, new_n14979_, new_n14980_, new_n14981_, new_n14982_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14992_, new_n14993_, new_n14994_,
    new_n14995_, new_n14996_, new_n14997_, new_n14998_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15014_, new_n15015_, new_n15016_, new_n15017_,
    new_n15018_, new_n15019_, new_n15020_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15029_,
    new_n15030_, new_n15031_, new_n15032_, new_n15033_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15066_, new_n15068_, new_n15069_,
    new_n15070_, new_n15071_, new_n15072_, new_n15073_, new_n15074_,
    new_n15075_, new_n15076_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15093_, new_n15094_, new_n15095_, new_n15096_, new_n15097_,
    new_n15098_, new_n15099_, new_n15101_, new_n15102_, new_n15104_,
    new_n15105_, new_n15106_, new_n15107_, new_n15108_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15132_, new_n15133_, new_n15134_,
    new_n15135_, new_n15136_, new_n15137_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15145_, new_n15146_,
    new_n15148_, new_n15149_, new_n15150_, new_n15151_, new_n15152_,
    new_n15154_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15160_, new_n15161_, new_n15162_, new_n15164_, new_n15165_,
    new_n15166_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15175_, new_n15176_, new_n15177_,
    new_n15178_, new_n15179_, new_n15180_, new_n15181_, new_n15182_,
    new_n15183_, new_n15184_, new_n15185_, new_n15186_, new_n15187_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15196_, new_n15197_, new_n15198_, new_n15199_,
    new_n15200_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15213_, new_n15214_, new_n15216_, new_n15217_,
    new_n15218_, new_n15219_, new_n15220_, new_n15221_, new_n15222_,
    new_n15223_, new_n15224_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15233_, new_n15234_,
    new_n15235_, new_n15236_, new_n15237_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15245_, new_n15246_,
    new_n15247_, new_n15248_, new_n15249_, new_n15251_, new_n15252_,
    new_n15253_, new_n15254_, new_n15255_, new_n15257_, new_n15258_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15281_, new_n15282_,
    new_n15283_, new_n15284_, new_n15285_, new_n15286_, new_n15288_,
    new_n15289_, new_n15290_, new_n15291_, new_n15292_, new_n15293_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15309_, new_n15310_, new_n15311_,
    new_n15312_, new_n15313_, new_n15314_, new_n15315_, new_n15317_,
    new_n15318_, new_n15319_, new_n15320_, new_n15321_, new_n15322_,
    new_n15324_, new_n15325_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15358_, new_n15359_, new_n15360_, new_n15361_, new_n15362_,
    new_n15364_, new_n15365_, new_n15366_, new_n15367_, new_n15368_,
    new_n15369_, new_n15370_, new_n15371_, new_n15372_, new_n15373_,
    new_n15374_, new_n15375_, new_n15377_, new_n15378_, new_n15379_,
    new_n15380_, new_n15381_, new_n15382_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15399_, new_n15400_, new_n15401_, new_n15402_,
    new_n15403_, new_n15404_, new_n15405_, new_n15407_, new_n15408_,
    new_n15409_, new_n15410_, new_n15411_, new_n15413_, new_n15414_,
    new_n15415_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15434_, new_n15436_, new_n15437_, new_n15438_,
    new_n15439_, new_n15440_, new_n15441_, new_n15442_, new_n15444_,
    new_n15445_, new_n15446_, new_n15447_, new_n15448_, new_n15449_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15465_, new_n15466_, new_n15467_,
    new_n15468_, new_n15469_, new_n15470_, new_n15471_, new_n15472_,
    new_n15473_, new_n15475_, new_n15476_, new_n15477_, new_n15478_,
    new_n15479_, new_n15481_, new_n15482_, new_n15483_, new_n15484_,
    new_n15485_, new_n15486_, new_n15487_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15503_, new_n15504_, new_n15505_, new_n15506_, new_n15507_,
    new_n15508_, new_n15510_, new_n15511_, new_n15512_, new_n15513_,
    new_n15514_, new_n15515_, new_n15516_, new_n15517_, new_n15518_,
    new_n15519_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15543_, new_n15544_, new_n15545_, new_n15547_, new_n15548_,
    new_n15549_, new_n15550_, new_n15551_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15573_, new_n15574_, new_n15575_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15581_, new_n15582_,
    new_n15583_, new_n15584_, new_n15585_, new_n15586_, new_n15587_,
    new_n15588_, new_n15589_, new_n15591_, new_n15592_, new_n15593_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15602_, new_n15603_, new_n15604_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15612_,
    new_n15613_, new_n15614_, new_n15615_, new_n15616_, new_n15618_,
    new_n15619_, new_n15620_, new_n15621_, new_n15622_, new_n15624_,
    new_n15625_, new_n15626_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15635_, new_n15636_,
    new_n15637_, new_n15638_, new_n15639_, new_n15641_, new_n15642_,
    new_n15643_, new_n15644_, new_n15645_, new_n15646_, new_n15647_,
    new_n15648_, new_n15649_, new_n15650_, new_n15652_, new_n15653_,
    new_n15654_, new_n15655_, new_n15656_, new_n15657_, new_n15658_,
    new_n15659_, new_n15660_, new_n15661_, new_n15662_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15682_, new_n15683_, new_n15684_, new_n15685_, new_n15686_,
    new_n15687_, new_n15688_, new_n15690_, new_n15691_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15698_,
    new_n15699_, new_n15700_, new_n15701_, new_n15702_, new_n15703_,
    new_n15704_, new_n15705_, new_n15706_, new_n15707_, new_n15708_,
    new_n15709_, new_n15710_, new_n15712_, new_n15713_, new_n15714_,
    new_n15715_, new_n15716_, new_n15717_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15725_, new_n15726_,
    new_n15728_, new_n15729_, new_n15730_, new_n15731_, new_n15732_,
    new_n15733_, new_n15735_, new_n15736_, new_n15737_, new_n15738_,
    new_n15739_, new_n15740_, new_n15741_, new_n15743_, new_n15744_,
    new_n15745_, new_n15746_, new_n15747_, new_n15748_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15757_, new_n15758_, new_n15759_, new_n15760_, new_n15761_,
    new_n15762_, new_n15764_, new_n15765_, new_n15766_, new_n15767_,
    new_n15768_, new_n15769_, new_n15770_, new_n15772_, new_n15773_,
    new_n15774_, new_n15775_, new_n15776_, new_n15777_, new_n15778_,
    new_n15780_, new_n15781_, new_n15782_, new_n15783_, new_n15784_,
    new_n15785_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15798_, new_n15799_, new_n15800_, new_n15801_,
    new_n15802_, new_n15804_, new_n15805_, new_n15806_, new_n15807_,
    new_n15808_, new_n15809_, new_n15811_, new_n15812_, new_n15813_,
    new_n15814_, new_n15815_, new_n15816_, new_n15817_, new_n15818_,
    new_n15819_, new_n15821_, new_n15822_, new_n15823_, new_n15824_,
    new_n15825_, new_n15826_, new_n15827_, new_n15828_, new_n15829_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15851_, new_n15852_,
    new_n15853_, new_n15854_, new_n15855_, new_n15856_, new_n15857_,
    new_n15859_, new_n15860_, new_n15861_, new_n15862_, new_n15863_,
    new_n15865_, new_n15866_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15887_,
    new_n15888_, new_n15889_, new_n15890_, new_n15891_, new_n15892_,
    new_n15894_, new_n15895_, new_n15896_, new_n15897_, new_n15898_,
    new_n15899_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15924_, new_n15925_, new_n15926_, new_n15927_,
    new_n15928_, new_n15929_, new_n15930_, new_n15932_, new_n15933_,
    new_n15934_, new_n15935_, new_n15936_, new_n15937_, new_n15938_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15954_, new_n15955_, new_n15956_, new_n15957_,
    new_n15958_, new_n15959_, new_n15960_, new_n15961_, new_n15962_,
    new_n15963_, new_n15964_, new_n15965_, new_n15966_, new_n15967_,
    new_n15968_, new_n15969_, new_n15970_, new_n15971_, new_n15972_,
    new_n15974_, new_n15975_, new_n15976_, new_n15977_, new_n15978_,
    new_n15979_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16002_,
    new_n16003_, new_n16004_, new_n16005_, new_n16006_, new_n16008_,
    new_n16009_, new_n16010_, new_n16011_, new_n16012_, new_n16014_,
    new_n16015_, new_n16016_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16048_,
    new_n16049_, new_n16050_, new_n16051_, new_n16052_, new_n16053_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16083_, new_n16084_, new_n16086_, new_n16087_, new_n16088_,
    new_n16089_, new_n16090_, new_n16091_, new_n16092_, new_n16093_,
    new_n16094_, new_n16095_, new_n16097_, new_n16098_, new_n16099_,
    new_n16100_, new_n16101_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16134_, new_n16135_, new_n16136_, new_n16138_,
    new_n16139_, new_n16140_, new_n16141_, new_n16142_, new_n16143_,
    new_n16145_, new_n16146_, new_n16147_, new_n16148_, new_n16149_,
    new_n16150_, new_n16151_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16162_, new_n16164_, new_n16165_, new_n16166_, new_n16167_,
    new_n16168_, new_n16169_, new_n16171_, new_n16172_, new_n16173_,
    new_n16174_, new_n16175_, new_n16177_, new_n16178_, new_n16179_,
    new_n16180_, new_n16181_, new_n16182_, new_n16183_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16199_, new_n16200_, new_n16201_, new_n16202_,
    new_n16203_, new_n16204_, new_n16206_, new_n16207_, new_n16208_,
    new_n16209_, new_n16210_, new_n16211_, new_n16212_, new_n16214_,
    new_n16215_, new_n16216_, new_n16217_, new_n16218_, new_n16219_,
    new_n16220_, new_n16221_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16240_, new_n16241_, new_n16242_,
    new_n16243_, new_n16244_, new_n16245_, new_n16246_, new_n16247_,
    new_n16249_, new_n16250_, new_n16251_, new_n16252_, new_n16253_,
    new_n16254_, new_n16256_, new_n16257_, new_n16258_, new_n16259_,
    new_n16260_, new_n16261_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16281_, new_n16282_,
    new_n16283_, new_n16284_, new_n16285_, new_n16287_, new_n16288_,
    new_n16289_, new_n16290_, new_n16292_, new_n16293_, new_n16294_,
    new_n16295_, new_n16296_, new_n16297_, new_n16298_, new_n16300_,
    new_n16301_, new_n16302_, new_n16303_, new_n16304_, new_n16306_,
    new_n16307_, new_n16308_, new_n16309_, new_n16310_, new_n16311_,
    new_n16312_, new_n16314_, new_n16315_, new_n16316_, new_n16317_,
    new_n16318_, new_n16319_, new_n16320_, new_n16321_, new_n16322_,
    new_n16323_, new_n16324_, new_n16325_, new_n16326_, new_n16327_,
    new_n16328_, new_n16329_, new_n16330_, new_n16331_, new_n16333_,
    new_n16334_, new_n16335_, new_n16336_, new_n16337_, new_n16338_,
    new_n16339_, new_n16340_, new_n16341_, new_n16342_, new_n16343_,
    new_n16344_, new_n16345_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16354_, new_n16355_,
    new_n16356_, new_n16357_, new_n16358_, new_n16359_, new_n16360_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16369_, new_n16370_, new_n16371_, new_n16372_,
    new_n16373_, new_n16374_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16384_,
    new_n16385_, new_n16386_, new_n16387_, new_n16388_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16408_, new_n16409_, new_n16410_, new_n16411_, new_n16412_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16421_, new_n16422_, new_n16423_, new_n16424_,
    new_n16425_, new_n16426_, new_n16427_, new_n16429_, new_n16430_,
    new_n16431_, new_n16432_, new_n16433_, new_n16434_, new_n16435_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16448_, new_n16449_, new_n16450_, new_n16451_, new_n16452_,
    new_n16453_, new_n16454_, new_n16455_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16461_, new_n16462_, new_n16464_,
    new_n16465_, new_n16466_, new_n16467_, new_n16468_, new_n16470_,
    new_n16471_, new_n16472_, new_n16473_, new_n16474_, new_n16475_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16491_, new_n16492_,
    new_n16493_, new_n16494_, new_n16495_, new_n16496_, new_n16498_,
    new_n16499_, new_n16500_, new_n16501_, new_n16502_, new_n16503_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16513_, new_n16514_, new_n16515_,
    new_n16516_, new_n16517_, new_n16518_, new_n16519_, new_n16520_,
    new_n16521_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16531_, new_n16532_,
    new_n16533_, new_n16534_, new_n16535_, new_n16536_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16585_, new_n16586_,
    new_n16587_, new_n16589_, new_n16590_, new_n16591_, new_n16592_,
    new_n16593_, new_n16594_, new_n16595_, new_n16596_, new_n16597_,
    new_n16599_, new_n16600_, new_n16601_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16624_, new_n16625_, new_n16626_, new_n16627_,
    new_n16628_, new_n16629_, new_n16630_, new_n16631_, new_n16632_,
    new_n16634_, new_n16635_, new_n16636_, new_n16637_, new_n16638_,
    new_n16639_, new_n16640_, new_n16641_, new_n16642_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16651_, new_n16652_, new_n16653_, new_n16654_, new_n16655_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16664_, new_n16665_, new_n16666_, new_n16667_,
    new_n16668_, new_n16669_, new_n16670_, new_n16672_, new_n16673_,
    new_n16674_, new_n16675_, new_n16676_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16684_, new_n16685_,
    new_n16686_, new_n16687_, new_n16688_, new_n16689_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16724_, new_n16725_, new_n16726_, new_n16727_, new_n16728_,
    new_n16730_, new_n16731_, new_n16732_, new_n16733_, new_n16734_,
    new_n16735_, new_n16737_, new_n16738_, new_n16739_, new_n16740_,
    new_n16741_, new_n16743_, new_n16745_, new_n16746_, new_n16747_,
    new_n16749_, new_n16750_, new_n16751_, new_n16752_, new_n16753_,
    new_n16754_, new_n16756_, new_n16757_, new_n16758_, new_n16759_,
    new_n16760_, new_n16761_, new_n16763_, new_n16764_, new_n16765_,
    new_n16766_, new_n16767_, new_n16768_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16783_,
    new_n16784_, new_n16786_, new_n16787_, new_n16788_, new_n16789_,
    new_n16790_, new_n16791_, new_n16793_, new_n16794_, new_n16795_,
    new_n16796_, new_n16797_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16818_, new_n16819_, new_n16820_, new_n16821_, new_n16822_,
    new_n16823_, new_n16824_, new_n16825_, new_n16826_, new_n16828_,
    new_n16829_, new_n16830_, new_n16831_, new_n16832_, new_n16833_,
    new_n16834_, new_n16835_, new_n16836_, new_n16837_, new_n16838_,
    new_n16839_, new_n16840_, new_n16842_, new_n16843_, new_n16844_,
    new_n16845_, new_n16846_, new_n16847_, new_n16849_, new_n16850_,
    new_n16851_, new_n16852_, new_n16853_, new_n16854_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16863_, new_n16864_, new_n16865_, new_n16866_, new_n16867_,
    new_n16868_, new_n16869_, new_n16871_, new_n16872_, new_n16873_,
    new_n16874_, new_n16875_, new_n16876_, new_n16878_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16887_, new_n16888_, new_n16889_, new_n16891_, new_n16892_,
    new_n16893_, new_n16894_, new_n16895_, new_n16896_, new_n16898_,
    new_n16899_, new_n16900_, new_n16901_, new_n16902_, new_n16903_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16922_, new_n16923_, new_n16924_, new_n16926_, new_n16927_,
    new_n16929_, new_n16930_, new_n16931_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16939_, new_n16940_,
    new_n16941_, new_n16942_, new_n16943_, new_n16944_, new_n16946_,
    new_n16947_, new_n16948_, new_n16949_, new_n16950_, new_n16951_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16960_, new_n16961_, new_n16963_, new_n16964_,
    new_n16965_, new_n16966_, new_n16967_, new_n16968_, new_n16969_,
    new_n16970_, new_n16971_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, n688, n693, n698,
    n703, n708, n713, n718, n723, n728, n733, n738, n743, n748, n753, n758,
    n763, n768, n773, n778, n783, n788, n793, n798, n803, n808, n813, n818,
    n823, n828, n833, n838, n843, n848, n853, n858, n863, n868, n873, n878,
    n883, n888, n893, n898, n903, n908, n913, n918, n923, n928, n933, n938,
    n943, n948, n953, n958, n963, n968, n973, n978, n983, n988, n993, n998,
    n1003, n1008, n1013, n1018, n1023, n1028, n1033, n1038, n1043, n1048,
    n1053, n1058, n1063, n1068, n1073, n1078, n1083, n1088, n1093, n1098,
    n1103, n1108, n1113, n1118, n1123, n1128, n1133, n1138, n1143, n1148,
    n1153, n1158, n1163, n1168, n1173, n1178, n1183, n1188, n1193, n1198,
    n1203, n1208, n1213, n1218, n1223, n1228, n1233, n1238, n1243, n1248,
    n1253, n1258, n1263, n1268, n1273, n1278, n1283, n1288, n1293, n1298,
    n1303, n1308, n1313, n1318, n1323, n1328, n1333, n1338, n1343, n1348,
    n1353, n1358, n1363, n1368, n1373, n1378, n1382, n1387, n1392, n1397,
    n1402, n1407, n1412, n1417, n1422, n1427, n1432, n1437, n1442, n1447,
    n1452, n1457, n1462, n1467, n1472, n1477, n1482, n1486, n1491, n1496,
    n1501, n1506, n1511, n1516, n1521, n1526, n1531, n1536, n1541, n1546,
    n1551, n1556, n1560, n1565, n1570, n1575, n1580, n1585, n1590, n1595,
    n1600, n1605, n1610, n1615, n1620, n1625, n1630, n1635, n1640, n1645,
    n1650, n1655, n1660, n1665, n1670, n1675, n1680, n1685, n1690, n1695,
    n1700, n1705, n1710, n1715, n1720, n1725, n1730, n1735, n1740, n1745,
    n1750, n1754, n1759, n1764, n1769, n1774, n1779, n1784, n1789, n1794,
    n1799, n1804, n1809, n1814, n1819, n1824, n1829, n1834, n1839, n1844,
    n1849, n1854, n1859, n1864, n1869, n1873, n1878, n1883, n1888, n1893,
    n1897, n1902, n1907, n1912, n1917, n1922, n1926, n1931, n1936, n1941,
    n1946, n1951, n1956, n1960, n1965, n1970, n1975, n1980, n1985, n1990,
    n1995, n2000, n2005, n2010, n2015, n2020, n2025, n2030, n2035, n2040,
    n2045, n2050, n2055, n2060, n2065, n2070, n2075, n2080, n2085, n2090,
    n2095, n2100, n2105, n2110, n2115, n2119, n2124, n2129, n2134, n2139,
    n2144, n2149, n2153, n2158, n2163, n2168, n2173, n2178, n2183, n2187,
    n2192, n2197, n2202, n2207, n2212, n2217, n2222, n2227, n2232, n2237,
    n2242, n2247, n2252, n2257, n2262, n2267, n2272, n2277, n2282, n2287,
    n2292, n2297, n2302, n2307, n2312, n2317, n2322, n2327, n2332, n2337,
    n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2381, n2386,
    n2391, n2396, n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436,
    n2441, n2446, n2451, n2456, n2461, n2466, n2471, n2476, n2481, n2486,
    n2490, n2495, n2500, n2505, n2510, n2515, n2520, n2525, n2530, n2535,
    n2540, n2545, n2550, n2555, n2560, n2565, n2570, n2575, n2580, n2585,
    n2590, n2595, n2600, n2605, n2609, n2614, n2619, n2624, n2629, n2634,
    n2639, n2644, n2649, n2654, n2659, n2664, n2669, n2673, n2678, n2683,
    n2688, n2693, n2698, n2703, n2708, n2713, n2718, n2723, n2728, n2733,
    n2738, n2743, n2748, n2753, n2758, n2762, n2767, n2772, n2777, n2782,
    n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832,
    n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882,
    n2887, n2892, n2896, n2901, n2906, n2911, n2916, n2921, n2926, n2931,
    n2936, n2941, n2944, n2948, n2953, n2958, n2963, n2968, n2973, n2978,
    n2983, n2988, n2993, n2998, n3003, n3008, n3013, n3018, n3023, n3028,
    n3033, n3038, n3043, n3048, n3053, n3058, n3063, n3068, n3073, n3078,
    n3083, n3088, n3093, n3097, n3101, n3106, n3111, n3116, n3121, n3126,
    n3131, n3136, n3141, n3146, n3151, n3156, n3161, n3166, n3171, n3176,
    n3181, n3186, n3191, n3196, n3201, n3206, n3211, n3216, n3221, n3226,
    n3231, n3236, n3241, n3246, n3251, n3256, n3261, n3265, n3270, n3275,
    n3280, n3285, n3290, n3295, n3300, n3305, n3310, n3315, n3320, n3325,
    n3330, n3335, n3340, n3345, n3350, n3355, n3360, n3365, n3370, n3375,
    n3380, n3385, n3390, n3395, n3400, n3404, n3409, n3414, n3419, n3424,
    n3429, n3434, n3439, n3444, n3449, n3454, n3459, n3464, n3469, n3474,
    n3479, n3484, n3489, n3494, n3499, n3504, n3509, n3514, n3519, n3524,
    n3529, n3534, n3538, n3543, n3548, n3553, n3558, n3563, n3568, n3573,
    n3578, n3583, n3588, n3593, n3598, n3603, n3608, n3613, n3618, n3623,
    n3628, n3633, n3638, n3643, n3648, n3652, n3657, n3662, n3667, n3672,
    n3676, n3681, n3686, n3691, n3696, n3700, n3705, n3710, n3715, n3720,
    n3725, n3730, n3735, n3738, n3742, n3747, n3752, n3757, n3762, n3767,
    n3772, n3776, n3781, n3786, n3791, n3796, n3801, n3806, n3811, n3816,
    n3821, n3825, n3829, n3834, n3839, n3844, n3849, n3854, n3859, n3864,
    n3869, n3874, n3879, n3884, n3889, n3894, n3899, n3904, n3909, n3914,
    n3919, n3924, n3929, n3934, n3939, n3944, n3949, n3954, n3959, n3964,
    n3969, n3974, n3979, n3984, n3989, n3994, n3999, n4004, n4009, n4014,
    n4018, n4023, n4028, n4033, n4037, n4042, n4047, n4052, n4057, n4062,
    n4067, n4072, n4077, n4082, n4087, n4092, n4097, n4102, n4106, n4111,
    n4116, n4121, n4126, n4131, n4136, n4141, n4146, n4151, n4156, n4161,
    n4166, n4171, n4176, n4180, n4185, n4190, n4195, n4200, n4205, n4210,
    n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4259,
    n4264, n4269, n4274, n4279, n4284, n4289, n4294, n4299, n4304, n4309,
    n4314, n4319, n4324, n4329, n4334, n4338, n4343, n4348, n4353, n4358,
    n4363, n4368, n4373, n4378, n4383, n4388, n4393, n4397, n4402, n4407,
    n4412, n4416, n4420, n4424, n4429, n4434, n4439, n4443, n4447, n4451,
    n4456, n4460, n4465, n4470, n4475, n4480, n4485, n4490, n4494, n4499,
    n4504, n4509, n4514, n4519, n4524, n4529, n4534, n4539, n4544, n4549,
    n4554, n4559, n4564, n4569, n4574, n4579, n4584, n4589, n4594, n4599,
    n4604, n4608, n4613, n4618, n4623, n4628, n4633, n4638, n4643, n4648,
    n4653, n4658, n4663, n4668, n4673, n4678, n4682, n4687, n4691, n4696,
    n4701, n4706, n4710, n4714, n4718, n4722, n4727, n4732, n4737, n4742,
    n4747, n4752, n4757, n4762, n4767, n4771, n4776, n4781, n4786, n4791,
    n4796, n4800, n4805, n4810, n4815, n4820, n4825, n4830, n4835, n4839,
    n4844, n4848, n4852, n4857, n4862, n4867, n4872, n4877, n4882, n4887,
    n4891, n4896, n4901, n4906, n4911, n4916, n4921, n4926, n4931, n4936,
    n4940, n4945, n4950, n4955, n4960, n4965, n4970, n4975, n4980, n4985,
    n4990, n4995, n5000, n5005, n5010, n5015, n5020, n5025, n5030, n5035,
    n5040, n5045, n5050, n5054, n5058, n5063, n5068, n5073, n5077, n5082,
    n5087, n5092, n5097, n5102, n5107, n5112, n5117, n5122, n5127, n5131,
    n5136, n5141, n5146, n5151, n5156, n5161, n5166, n5171, n5176, n5181,
    n5186, n5191, n5196, n5201, n5206, n5211, n5216, n5221, n5226, n5231,
    n5235, n5240, n5245, n5249, n5254, n5258, n5263, n5268, n5273, n5278,
    n5283, n5288, n5293, n5298, n5303, n5308, n5312, n5316, n5321, n5326,
    n5330, n5334, n5339, n5344, n5349, n5353, n5358, n5363, n5368, n5373,
    n5378, n5383, n5387, n5392, n5397, n5402, n5407, n5412, n5417, n5422,
    n5427, n5432, n5437, n5442, n5447, n5452, n5457, n5462, n5467, n5472,
    n5477, n5480, n5485, n5490, n5495, n5500, n5505, n5509, n5514, n5519,
    n5524, n5529, n5533, n5537, n5542, n5547, n5552, n5557, n5562, n5566,
    n5570, n5575, n5580, n5585, n5590, n5594, n5598, n5603, n5608, n5613,
    n5618, n5623, n5628, n5633, n5638, n5643, n5648, n5653, n5658, n5663,
    n5668, n5672, n5677, n5682, n5687, n5692, n5697, n5702, n5707, n5712,
    n5717, n5722, n5727, n5732, n5737, n5742, n5747, n5752, n5757, n5762,
    n5766, n5771, n5776, n5781, n5785, n5789, n5794, n5799, n5804, n5809,
    n5814, n5819, n5824, n5829, n5834, n5838, n5843, n5848, n5853, n5858,
    n5863, n5868, n5873, n5878, n5883, n5888, n5893, n5898, n5902, n5907,
    n5912, n5917, n5921, n5925, n5930, n5935, n5940, n5945, n5950, n5955,
    n5960, n5965, n5969, n5974, n5979, n5983, n5988, n5993, n5998, n6003,
    n6008, n6013, n6018, n6023, n6028, n6033, n6037, n6041, n6045, n6050,
    n6055, n6060, n6065, n6069, n6074, n6079, n6084, n6088, n6092, n6096,
    n6101, n6105, n6109, n6114, n6119, n6124, n6129, n6134, n6139, n6144,
    n6149, n6154, n6159, n6164, n6169, n6174, n6179, n6184, n6188, n6192,
    n6197, n6202, n6207, n6212, n6216, n6220, n6225, n6230, n6235, n6240,
    n6245, n6250, n6255, n6260, n6265, n6270, n6275, n6280, n6285, n6290,
    n6295, n6300, n6304, n6308, n6313, n6318, n6323, n6328, n6333, n6338,
    n6342, n6347, n6352, n6357, n6362, n6367, n6372, n6377, n6382, n6387,
    n6392, n6397, n6402, n6407, n6411, n6416, n6420, n6425, n6430, n6435,
    n6440, n6445, n6450, n6455, n6460, n6465, n6470, n6475, n6480, n6485,
    n6489, n6493, n6498, n6503, n6508, n6513, n6518, n6523, n6527, n6532,
    n6537, n6542, n6547, n6552, n6557, n6562, n6566, n6571, n6576, n6581,
    n6586, n6591, n6596, n6600, n6604, n6609, n6614, n6619, n6624, n6628,
    n6632, n6637, n6642, n6647, n6652, n6657, n6662, n6667, n6672, n6677,
    n6682, n6687, n6691, n6696, n6701, n6706, n6711, n6716, n6721, n6726,
    n6731, n6736, n6741, n6746, n6751, n6756, n6761, n6766, n6771, n6776,
    n6781, n6786, n6791, n6796, n6801, n6806, n6810, n6814, n6819, n6824,
    n6829, n6834, n6839, n6844, n6849, n6854, n6859, n6863, n6868, n6873,
    n6878, n6883, n6888, n6893, n6898, n6902, n6907, n6912, n6916, n6921,
    n6926, n6931, n6936, n6941, n6946, n6951, n6956, n6961, n6966, n6971,
    n6976, n6981, n6986, n6991, n6996, n7001, n7006, n7011, n7016, n7019,
    n7023, n7027, n7031, n7036, n7041, n7046, n7050, n7055, n7060, n7065,
    n7070, n7075, n7080, n7085, n7089, n7093, n7098, n7103, n7108, n7113,
    n7118, n7123, n7128, n7133, n7138, n7143, n7148, n7153, n7158, n7163,
    n7168, n7173, n7178, n7183, n7188, n7193, n7198, n7203, n7208, n7213,
    n7218, n7222, n7227, n7232, n7237, n7242, n7247, n7252, n7257, n7262,
    n7266, n7271, n7276, n7280, n7284, n7289, n7294, n7299, n7304, n7309,
    n7314, n7319, n7324, n7329, n7334, n7339, n7344, n7349, n7354, n7359,
    n7364, n7369, n7374, n7379, n7383, n7388, n7392, n7397, n7402, n7407,
    n7412, n7417, n7422, n7426, n7430, n7435, n7440, n7445, n7450, n7455,
    n7460, n7465, n7470, n7475, n7480, n7485, n7490, n7495, n7500, n7505,
    n7509, n7514, n7519, n7524, n7529, n7533, n7537, n7542, n7547, n7551,
    n7556, n7561, n7566, n7571, n7576, n7580, n7584, n7589, n7594, n7599,
    n7603, n7607, n7612, n7617, n7622, n7627, n7632, n7637, n7641, n7646,
    n7651, n7656, n7660;
  assign new_n4623_1_ = ~ng6191 & ~ng6177;
  assign new_n4624_ = pg35 & ~new_n4623_1_;
  assign new_n4625_ = ~ng5485 & ~ng5499;
  assign new_n4626_ = pg35 & ~new_n4625_;
  assign new_n4627_ = ~ng5831 & ~ng5845;
  assign new_n4628_1_ = pg35 & ~new_n4627_;
  assign new_n4629_ = ~ng5138 & ~ng5152;
  assign new_n4630_ = pg35 & ~new_n4629_;
  assign new_n4631_ = ~new_n4624_ & ~new_n4626_;
  assign new_n4632_ = ~new_n4628_1_ & new_n4631_;
  assign new_n4633_1_ = ~new_n4630_ & new_n4632_;
  assign new_n4634_ = ~ng3845 & ~ng3831;
  assign new_n4635_ = pg35 & ~new_n4634_;
  assign new_n4636_ = ~ng3143 & ~ng3129;
  assign new_n4637_ = pg35 & ~new_n4636_;
  assign new_n4638_1_ = ~ng3480 & ~ng3494;
  assign new_n4639_ = pg35 & ~new_n4638_1_;
  assign new_n4640_ = ~ng6537 & ~ng6523;
  assign new_n4641_ = pg35 & ~new_n4640_;
  assign new_n4642_ = ~new_n4635_ & ~new_n4637_;
  assign new_n4643_1_ = ~new_n4639_ & new_n4642_;
  assign new_n4644_ = new_n4641_ & new_n4643_1_;
  assign new_n4645_ = new_n4633_1_ & new_n4644_;
  assign new_n4646_ = ~new_n4626_ & ~new_n4641_;
  assign new_n4647_ = ~new_n4624_ & new_n4646_;
  assign new_n4648_1_ = ~new_n4630_ & new_n4647_;
  assign new_n4649_ = new_n4628_1_ & new_n4643_1_;
  assign new_n4650_ = new_n4648_1_ & new_n4649_;
  assign new_n4651_ = ~new_n4628_1_ & new_n4646_;
  assign new_n4652_ = ~new_n4630_ & new_n4651_;
  assign new_n4653_1_ = new_n4624_ & new_n4643_1_;
  assign new_n4654_ = new_n4652_ & new_n4653_1_;
  assign new_n4655_ = ~new_n4628_1_ & ~new_n4641_;
  assign new_n4656_ = ~new_n4624_ & new_n4655_;
  assign new_n4657_ = ~new_n4630_ & new_n4656_;
  assign new_n4658_1_ = new_n4626_ & new_n4643_1_;
  assign new_n4659_ = new_n4657_ & new_n4658_1_;
  assign new_n4660_ = ~new_n4645_ & ~new_n4650_;
  assign new_n4661_ = ~new_n4654_ & ~new_n4659_;
  assign new_n4662_ = new_n4660_ & new_n4661_;
  assign new_n4663_1_ = ~new_n4626_ & new_n4656_;
  assign new_n4664_ = new_n4630_ & new_n4643_1_;
  assign new_n4665_ = new_n4663_1_ & new_n4664_;
  assign new_n4666_ = ~new_n4630_ & ~new_n4637_;
  assign new_n4667_ = ~new_n4635_ & new_n4666_;
  assign new_n4668_1_ = new_n4639_ & new_n4667_;
  assign new_n4669_ = new_n4663_1_ & new_n4668_1_;
  assign new_n4670_ = ~new_n4639_ & new_n4666_;
  assign new_n4671_ = new_n4635_ & new_n4670_;
  assign new_n4672_ = new_n4663_1_ & new_n4671_;
  assign new_n4673_1_ = ~new_n4630_ & ~new_n4639_;
  assign new_n4674_ = ~new_n4635_ & new_n4673_1_;
  assign new_n4675_ = new_n4637_ & new_n4674_;
  assign new_n4676_ = new_n4663_1_ & new_n4675_;
  assign new_n4677_ = ~new_n4665_ & ~new_n4669_;
  assign new_n4678_1_ = ~new_n4672_ & ~new_n4676_;
  assign new_n4679_ = new_n4677_ & new_n4678_1_;
  assign new_n4680_ = new_n4662_ & new_n4679_;
  assign new_n4681_ = new_n4631_ & new_n4655_;
  assign new_n4682_1_ = new_n4642_ & new_n4673_1_;
  assign new_n4683_ = new_n4681_ & new_n4682_1_;
  assign pg28030 = ~new_n4680_ | new_n4683_;
  assign new_n4685_ = ~ng969 & ~ng1008;
  assign new_n4686_ = ng1193 & ~new_n4685_;
  assign new_n4687_1_ = pg35 & ~new_n4686_;
  assign new_n4688_ = ~ng1312 & ~ng1351;
  assign new_n4689_ = ng1536 & ~new_n4688_;
  assign new_n4690_ = pg35 & ~new_n4689_;
  assign new_n4691_1_ = ~new_n4687_1_ & new_n4690_;
  assign new_n4692_ = new_n4687_1_ & ~new_n4690_;
  assign new_n4693_ = ~new_n4691_1_ & ~new_n4692_;
  assign new_n4694_ = ~new_n4687_1_ & ~new_n4690_;
  assign pg28041 = ~new_n4693_ | new_n4694_;
  assign new_n4696_1_ = ~ng1216 & ~ng1205;
  assign new_n4697_ = ~ng1221 & new_n4696_1_;
  assign new_n4698_ = ~ng1211 & new_n4697_;
  assign new_n4699_ = ng1171 & ~ng1183;
  assign new_n4700_ = ng1061 & new_n4698_;
  assign new_n4701_1_ = ng979 & new_n4699_;
  assign new_n4702_ = new_n4700_ & new_n4701_1_;
  assign pg33533 = ng1075 & ~new_n4702_;
  assign pg34437 = ~pg113 | ~ng2868;
  assign new_n4705_ = ~ng4064 & ~ng4057;
  assign new_n4706_1_ = ~ng4141 & ~ng4082;
  assign new_n4707_ = ~ng4087 & ~ng4093;
  assign new_n4708_ = ~ng4098 & new_n4707_;
  assign new_n4709_ = ng4076 & new_n4708_;
  assign new_n4710_1_ = ng4112 & new_n4709_;
  assign new_n4711_ = new_n4706_1_ & ~new_n4710_1_;
  assign new_n4712_ = new_n4705_ & ~new_n4711_;
  assign pg31521 = ~ng4125 & new_n4712_;
  assign new_n4714_1_ = ng2724 & ~ng2787;
  assign new_n4715_ = ~ng2724 & ~ng2783;
  assign new_n4716_ = ~new_n4714_1_ & ~new_n4715_;
  assign new_n4717_ = ng2729 & new_n4716_;
  assign new_n4718_1_ = ~ng2775 & ng2724;
  assign new_n4719_ = ~ng2724 & ~ng2771;
  assign new_n4720_ = ~new_n4718_1_ & ~new_n4719_;
  assign new_n4721_ = ~ng2729 & new_n4720_;
  assign pg33435 = ~new_n4717_ & ~new_n4721_;
  assign new_n4723_ = pg99 & ng37;
  assign new_n4724_ = ~pg134 & ~new_n4723_;
  assign new_n4725_ = pg72 & ng4322;
  assign new_n4726_ = ng4322 & ~new_n4725_;
  assign new_n4727_1_ = pg72 & ~new_n4725_;
  assign new_n4728_ = ~new_n4726_ & ~new_n4727_1_;
  assign new_n4729_ = pg73 & ng4332;
  assign new_n4730_ = ng4332 & ~new_n4729_;
  assign new_n4731_ = pg73 & ~new_n4729_;
  assign new_n4732_1_ = ~new_n4730_ & ~new_n4731_;
  assign new_n4733_ = new_n4728_ & new_n4732_1_;
  assign new_n4734_ = ~ng4311 & new_n4733_;
  assign new_n4735_ = ng4311 & new_n4733_;
  assign new_n4736_ = ~new_n4734_ & ~new_n4735_;
  assign new_n4737_1_ = pg113 & ~new_n4724_;
  assign new_n4738_ = ~new_n4736_ & new_n4737_1_;
  assign new_n4739_ = ~ng4349 & ~ng4358;
  assign new_n4740_ = new_n4734_ & new_n4739_;
  assign pg25114 = ng5297 & ng5357;
  assign new_n4742_1_ = new_n4740_ & pg25114;
  assign new_n4743_ = ~ng4349 & ng4358;
  assign new_n4744_ = new_n4734_ & new_n4743_;
  assign new_n4745_ = ng5990 & ng6049;
  assign new_n4746_ = new_n4744_ & new_n4745_;
  assign new_n4747_1_ = ng4349 & ~ng4358;
  assign new_n4748_ = new_n4734_ & new_n4747_1_;
  assign new_n4749_ = ng5703 & ng5644;
  assign new_n4750_ = new_n4748_ & new_n4749_;
  assign new_n4751_ = ng4349 & ng4358;
  assign new_n4752_1_ = new_n4734_ & new_n4751_;
  assign new_n4753_ = ng6336 & ng6395;
  assign new_n4754_ = new_n4752_1_ & new_n4753_;
  assign new_n4755_ = ~new_n4742_1_ & ~new_n4746_;
  assign new_n4756_ = ~new_n4750_ & ~new_n4754_;
  assign new_n4757_1_ = new_n4755_ & new_n4756_;
  assign new_n4758_ = new_n4735_ & new_n4739_;
  assign new_n4759_ = ng6741 & ng6682;
  assign new_n4760_ = new_n4758_ & new_n4759_;
  assign new_n4761_ = new_n4735_ & new_n4743_;
  assign new_n4762_1_ = ng3703 & ng3639;
  assign new_n4763_ = new_n4761_ & new_n4762_1_;
  assign new_n4764_ = new_n4735_ & new_n4747_1_;
  assign new_n4765_ = ng3352 & ng3288;
  assign new_n4766_ = new_n4764_ & new_n4765_;
  assign new_n4767_1_ = new_n4735_ & new_n4751_;
  assign new_n4768_ = ng4054 & ng3990;
  assign new_n4769_ = new_n4767_1_ & new_n4768_;
  assign new_n4770_ = ~new_n4760_ & ~new_n4763_;
  assign new_n4771_1_ = ~new_n4766_ & ~new_n4769_;
  assign new_n4772_ = new_n4770_ & new_n4771_1_;
  assign new_n4773_ = new_n4757_1_ & new_n4772_;
  assign new_n4774_ = new_n4738_ & ~new_n4773_;
  assign pg34425 = ~new_n4738_ | new_n4774_;
  assign new_n4776_1_ = pg35 & ng3817;
  assign new_n4777_ = pg35 & ng3115;
  assign new_n4778_ = pg35 & ng3466;
  assign new_n4779_ = pg35 & ng4420;
  assign new_n4780_ = pg35 & ng4427;
  assign new_n4781_1_ = ~new_n4779_ & ~new_n4780_;
  assign new_n4782_ = ~new_n4776_1_ & ~new_n4777_;
  assign new_n4783_ = ~new_n4778_ & new_n4782_;
  assign new_n4784_ = ~new_n4781_1_ & new_n4783_;
  assign new_n4785_ = pg35 & ng6163;
  assign new_n4786_1_ = pg35 & ng5471;
  assign new_n4787_ = pg35 & ng5817;
  assign new_n4788_ = pg35 & ng5124;
  assign new_n4789_ = ~new_n4785_ & ~new_n4786_1_;
  assign new_n4790_ = ~new_n4787_ & new_n4789_;
  assign new_n4791_1_ = ~new_n4788_ & new_n4790_;
  assign new_n4792_ = pg35 & ng6509;
  assign new_n4793_ = new_n4784_ & new_n4791_1_;
  assign new_n4794_ = ~new_n4792_ & new_n4793_;
  assign new_n4795_ = ~new_n4777_ & new_n4781_1_;
  assign new_n4796_1_ = ~new_n4776_1_ & new_n4795_;
  assign new_n4797_ = new_n4778_ & new_n4796_1_;
  assign new_n4798_ = new_n4791_1_ & new_n4797_;
  assign new_n4799_ = ~new_n4792_ & new_n4798_;
  assign new_n4800_1_ = ~new_n4778_ & new_n4795_;
  assign new_n4801_ = new_n4776_1_ & new_n4800_1_;
  assign new_n4802_ = new_n4791_1_ & new_n4801_;
  assign new_n4803_ = ~new_n4792_ & new_n4802_;
  assign new_n4804_ = ~new_n4778_ & new_n4781_1_;
  assign new_n4805_1_ = ~new_n4776_1_ & new_n4804_;
  assign new_n4806_ = new_n4777_ & new_n4805_1_;
  assign new_n4807_ = new_n4791_1_ & new_n4806_;
  assign new_n4808_ = ~new_n4792_ & new_n4807_;
  assign new_n4809_ = ~new_n4794_ & ~new_n4799_;
  assign new_n4810_1_ = ~new_n4803_ & ~new_n4808_;
  assign new_n4811_ = new_n4809_ & new_n4810_1_;
  assign new_n4812_ = new_n4783_ & new_n4785_;
  assign new_n4813_ = ~new_n4787_ & ~new_n4788_;
  assign new_n4814_ = ~new_n4786_1_ & new_n4813_;
  assign new_n4815_1_ = new_n4781_1_ & new_n4814_;
  assign new_n4816_ = new_n4812_ & new_n4815_1_;
  assign new_n4817_ = ~new_n4792_ & new_n4816_;
  assign new_n4818_ = new_n4783_ & new_n4786_1_;
  assign new_n4819_ = ~new_n4785_ & ~new_n4788_;
  assign new_n4820_1_ = ~new_n4787_ & new_n4819_;
  assign new_n4821_ = new_n4781_1_ & new_n4820_1_;
  assign new_n4822_ = new_n4818_ & new_n4821_;
  assign new_n4823_ = ~new_n4792_ & new_n4822_;
  assign new_n4824_ = new_n4783_ & new_n4787_;
  assign new_n4825_1_ = ~new_n4786_1_ & new_n4819_;
  assign new_n4826_ = new_n4781_1_ & new_n4825_1_;
  assign new_n4827_ = new_n4824_ & new_n4826_;
  assign new_n4828_ = ~new_n4792_ & new_n4827_;
  assign new_n4829_ = new_n4783_ & new_n4788_;
  assign new_n4830_1_ = new_n4781_1_ & new_n4790_;
  assign new_n4831_ = new_n4829_ & new_n4830_1_;
  assign new_n4832_ = ~new_n4792_ & new_n4831_;
  assign new_n4833_ = ~new_n4817_ & ~new_n4823_;
  assign new_n4834_ = ~new_n4828_ & ~new_n4832_;
  assign new_n4835_1_ = new_n4833_ & new_n4834_;
  assign new_n4836_ = new_n4783_ & new_n4792_;
  assign new_n4837_ = new_n4815_1_ & new_n4836_;
  assign new_n4838_ = ~new_n4785_ & new_n4837_;
  assign new_n4839_1_ = new_n4811_ & new_n4835_1_;
  assign new_n4840_ = ~new_n4838_ & new_n4839_1_;
  assign new_n4841_ = new_n4782_ & new_n4804_;
  assign new_n4842_ = new_n4789_ & new_n4813_;
  assign new_n4843_ = new_n4841_ & new_n4842_;
  assign new_n4844_1_ = ~new_n4792_ & new_n4843_;
  assign pg31793 = ~new_n4840_ | new_n4844_1_;
  assign pg34436 = ~pg113 | ~ng2873;
  assign pg21727 = ~pg35 & ng3003;
  assign new_n4848_1_ = ~ng1710 & ~ng1724;
  assign new_n4849_ = ~ng1992 & ~ng1978;
  assign new_n4850_ = ~ng1858 & ~ng1844;
  assign new_n4851_ = ~ng2112 & ~ng2126;
  assign new_n4852_1_ = new_n4848_1_ & new_n4849_;
  assign new_n4853_ = new_n4850_ & new_n4852_1_;
  assign new_n4854_ = new_n4851_ & new_n4853_;
  assign new_n4855_ = pg35 & ~new_n4854_;
  assign new_n4856_ = ~ng2269 & ~ng2283;
  assign new_n4857_1_ = ~ng2537 & ~ng2551;
  assign new_n4858_ = ~ng2417 & ~ng2403;
  assign new_n4859_ = ~ng2671 & ~ng2685;
  assign new_n4860_ = new_n4856_ & new_n4857_1_;
  assign new_n4861_ = new_n4858_ & new_n4860_;
  assign new_n4862_1_ = new_n4859_ & new_n4861_;
  assign new_n4863_ = pg35 & ~new_n4862_1_;
  assign new_n4864_ = ~new_n4855_ & new_n4863_;
  assign new_n4865_ = new_n4855_ & ~new_n4863_;
  assign new_n4866_ = ~new_n4864_ & ~new_n4865_;
  assign new_n4867_1_ = ~new_n4855_ & ~new_n4863_;
  assign pg26876 = ~new_n4866_ | new_n4867_1_;
  assign new_n4869_ = ~pg73 & ng490;
  assign new_n4870_ = ~pg73 & ~new_n4869_;
  assign new_n4871_ = ng490 & ~new_n4869_;
  assign new_n4872_1_ = ~new_n4870_ & ~new_n4871_;
  assign new_n4873_ = ~pg72 & ng482;
  assign new_n4874_ = ~pg72 & ~new_n4873_;
  assign new_n4875_ = ng482 & ~new_n4873_;
  assign new_n4876_ = ~new_n4874_ & ~new_n4875_;
  assign new_n4877_1_ = ng479 & ~new_n4872_1_;
  assign new_n4878_ = ~ng528 & ~new_n4876_;
  assign new_n4879_ = new_n4877_1_ & new_n4878_;
  assign pg33894 = ng890 & ~new_n4879_;
  assign new_n4881_ = ~ng7 & ~ng6;
  assign new_n4882_1_ = ~ng8 & new_n4881_;
  assign new_n4883_ = ~ng31 & ng28;
  assign new_n4884_ = new_n4882_1_ & new_n4883_;
  assign new_n4885_ = ~ng16 & new_n4884_;
  assign new_n4886_ = ~ng9 & new_n4885_;
  assign new_n4887_1_ = ng19 & new_n4886_;
  assign new_n4888_ = pg54 & ~ng34;
  assign new_n4889_ = ~pg53 & new_n4888_;
  assign new_n4890_ = ~pg57 & new_n4889_;
  assign new_n4891_1_ = ~pg56 & new_n4890_;
  assign n3414 = pg54 & new_n4891_1_;
  assign new_n4893_ = new_n4887_1_ & n3414;
  assign new_n4894_ = ~pg53 & ~n3414;
  assign new_n4895_ = ng31 & ~ng28;
  assign new_n4896_1_ = new_n4882_1_ & new_n4895_;
  assign new_n4897_ = ~ng16 & new_n4896_1_;
  assign new_n4898_ = ~ng9 & new_n4897_;
  assign new_n4899_ = ng19 & new_n4898_;
  assign new_n4900_ = ~ng19 & new_n4886_;
  assign new_n4901_1_ = ng31 & ng28;
  assign new_n4902_ = new_n4882_1_ & new_n4901_1_;
  assign new_n4903_ = ~ng16 & new_n4902_;
  assign new_n4904_ = ~ng9 & new_n4903_;
  assign new_n4905_ = ~ng19 & new_n4904_;
  assign new_n4906_1_ = ~ng31 & ~ng28;
  assign new_n4907_ = new_n4882_1_ & new_n4906_1_;
  assign new_n4908_ = ~ng16 & new_n4907_;
  assign new_n4909_ = ~ng9 & new_n4908_;
  assign new_n4910_ = ~ng19 & new_n4909_;
  assign new_n4911_1_ = ~new_n4900_ & ~new_n4905_;
  assign new_n4912_ = ~new_n4910_ & new_n4911_1_;
  assign new_n4913_ = ng19 & new_n4909_;
  assign new_n4914_ = ~new_n4899_ & new_n4912_;
  assign new_n4915_ = ~new_n4913_ & new_n4914_;
  assign new_n4916_1_ = n3414 & ~new_n4915_;
  assign new_n4917_ = ng16 & new_n4907_;
  assign new_n4918_ = ~ng9 & new_n4917_;
  assign new_n4919_ = ~ng19 & new_n4918_;
  assign new_n4920_ = n3414 & new_n4919_;
  assign new_n4921_1_ = ~new_n4893_ & ~new_n4894_;
  assign new_n4922_ = ~new_n4916_1_ & new_n4921_1_;
  assign new_n4923_ = new_n4920_ & new_n4922_;
  assign new_n4924_ = ng19 & new_n4918_;
  assign new_n4925_ = n3414 & new_n4924_;
  assign new_n4926_1_ = ng9 & new_n4908_;
  assign new_n4927_ = ~ng19 & new_n4926_1_;
  assign new_n4928_ = n3414 & new_n4927_;
  assign new_n4929_ = ng9 & new_n4885_;
  assign new_n4930_ = ng19 & new_n4929_;
  assign new_n4931_1_ = n3414 & new_n4930_;
  assign new_n4932_ = ng7 & ng6;
  assign new_n4933_ = ng8 & new_n4932_;
  assign new_n4934_ = new_n4906_1_ & new_n4933_;
  assign new_n4935_ = ~ng16 & new_n4934_;
  assign new_n4936_1_ = ng9 & new_n4935_;
  assign new_n4937_ = ~ng19 & new_n4936_1_;
  assign new_n4938_ = new_n4883_ & new_n4933_;
  assign new_n4939_ = ~ng16 & new_n4938_;
  assign new_n4940_1_ = ng9 & new_n4939_;
  assign new_n4941_ = ng19 & new_n4940_1_;
  assign new_n4942_ = ~ng19 & new_n4940_1_;
  assign new_n4943_ = ng16 & new_n4934_;
  assign new_n4944_ = ng9 & new_n4943_;
  assign new_n4945_1_ = ~ng19 & new_n4944_;
  assign new_n4946_ = ~new_n4937_ & ~new_n4941_;
  assign new_n4947_ = ~new_n4942_ & new_n4946_;
  assign new_n4948_ = ~new_n4945_1_ & new_n4947_;
  assign new_n4949_ = ng16 & new_n4902_;
  assign new_n4950_1_ = ~ng9 & new_n4949_;
  assign new_n4951_ = ~ng19 & new_n4950_1_;
  assign new_n4952_ = ng16 & new_n4884_;
  assign new_n4953_ = ~ng9 & new_n4952_;
  assign new_n4954_ = ~ng19 & new_n4953_;
  assign new_n4955_1_ = ~ng19 & new_n4929_;
  assign new_n4956_ = ~new_n4951_ & ~new_n4954_;
  assign new_n4957_ = ~new_n4955_1_ & new_n4956_;
  assign new_n4958_ = new_n4948_ & new_n4957_;
  assign new_n4959_ = n3414 & ~new_n4958_;
  assign new_n4960_1_ = ~new_n4925_ & ~new_n4928_;
  assign new_n4961_ = ~new_n4931_1_ & new_n4960_1_;
  assign new_n4962_ = ~new_n4959_ & new_n4961_;
  assign new_n4963_ = ng19 & new_n4953_;
  assign new_n4964_ = n3414 & new_n4963_;
  assign new_n4965_1_ = new_n4923_ & new_n4962_;
  assign new_n4966_ = ~new_n4964_ & new_n4965_1_;
  assign new_n4967_ = ~new_n4894_ & ~new_n4920_;
  assign new_n4968_ = ~new_n4893_ & new_n4967_;
  assign new_n4969_ = new_n4916_1_ & new_n4968_;
  assign new_n4970_1_ = new_n4962_ & new_n4969_;
  assign new_n4971_ = ~new_n4964_ & new_n4970_1_;
  assign new_n4972_ = ~new_n4916_1_ & new_n4967_;
  assign new_n4973_ = new_n4893_ & new_n4972_;
  assign new_n4974_ = new_n4962_ & new_n4973_;
  assign new_n4975_1_ = ~new_n4964_ & new_n4974_;
  assign new_n4976_ = ~new_n4916_1_ & ~new_n4920_;
  assign new_n4977_ = ~new_n4893_ & new_n4976_;
  assign new_n4978_ = new_n4894_ & new_n4977_;
  assign new_n4979_ = new_n4962_ & new_n4978_;
  assign new_n4980_1_ = ~new_n4964_ & new_n4979_;
  assign new_n4981_ = ~new_n4966_ & ~new_n4971_;
  assign new_n4982_ = ~new_n4975_1_ & ~new_n4980_1_;
  assign new_n4983_ = new_n4981_ & new_n4982_;
  assign new_n4984_ = new_n4922_ & new_n4925_;
  assign new_n4985_1_ = ~new_n4931_1_ & ~new_n4959_;
  assign new_n4986_ = ~new_n4928_ & new_n4985_1_;
  assign new_n4987_ = ~new_n4920_ & new_n4986_;
  assign new_n4988_ = new_n4984_ & new_n4987_;
  assign new_n4989_ = ~new_n4964_ & new_n4988_;
  assign new_n4990_1_ = new_n4922_ & new_n4928_;
  assign new_n4991_ = ~new_n4925_ & ~new_n4959_;
  assign new_n4992_ = ~new_n4931_1_ & new_n4991_;
  assign new_n4993_ = ~new_n4920_ & new_n4992_;
  assign new_n4994_ = new_n4990_1_ & new_n4993_;
  assign new_n4995_1_ = ~new_n4964_ & new_n4994_;
  assign new_n4996_ = new_n4922_ & new_n4931_1_;
  assign new_n4997_ = ~new_n4928_ & new_n4991_;
  assign new_n4998_ = ~new_n4920_ & new_n4997_;
  assign new_n4999_ = new_n4996_ & new_n4998_;
  assign new_n5000_1_ = ~new_n4964_ & new_n4999_;
  assign new_n5001_ = new_n4922_ & new_n4959_;
  assign new_n5002_ = ~new_n4920_ & new_n4961_;
  assign new_n5003_ = new_n5001_ & new_n5002_;
  assign new_n5004_ = ~new_n4964_ & new_n5003_;
  assign new_n5005_1_ = ~new_n4989_ & ~new_n4995_1_;
  assign new_n5006_ = ~new_n5000_1_ & ~new_n5004_;
  assign new_n5007_ = new_n5005_1_ & new_n5006_;
  assign new_n5008_ = new_n4922_ & new_n4964_;
  assign new_n5009_ = new_n4987_ & new_n5008_;
  assign new_n5010_1_ = ~new_n4925_ & new_n5009_;
  assign new_n5011_ = new_n4983_ & new_n5007_;
  assign new_n5012_ = ~new_n5010_1_ & new_n5011_;
  assign new_n5013_ = new_n4921_1_ & new_n4976_;
  assign new_n5014_ = new_n4960_1_ & new_n4985_1_;
  assign new_n5015_1_ = new_n5013_ & new_n5014_;
  assign new_n5016_ = ~new_n4964_ & new_n5015_1_;
  assign pg34239 = ~new_n5012_ | new_n5016_;
  assign new_n5018_ = ~ng1664 & ~ng1644;
  assign new_n5019_ = ~ng1913 & ~ng1932;
  assign new_n5020_1_ = ~ng1779 & ~ng1798;
  assign new_n5021_ = ~ng2047 & ~ng2066;
  assign new_n5022_ = new_n5018_ & new_n5019_;
  assign new_n5023_ = new_n5020_1_ & new_n5022_;
  assign new_n5024_ = new_n5021_ & new_n5023_;
  assign new_n5025_1_ = pg35 & ~new_n5024_;
  assign new_n5026_ = ~ng2204 & ~ng2223;
  assign new_n5027_ = ~ng2472 & ~ng2491;
  assign new_n5028_ = ~ng2338 & ~ng2357;
  assign new_n5029_ = ~ng2606 & ~ng2625;
  assign new_n5030_1_ = new_n5026_ & new_n5027_;
  assign new_n5031_ = new_n5028_ & new_n5030_1_;
  assign new_n5032_ = new_n5029_ & new_n5031_;
  assign new_n5033_ = pg35 & ~new_n5032_;
  assign new_n5034_ = ~new_n5025_1_ & new_n5033_;
  assign new_n5035_1_ = new_n5025_1_ & ~new_n5033_;
  assign new_n5036_ = ~new_n5034_ & ~new_n5035_1_;
  assign new_n5037_ = ~new_n5025_1_ & ~new_n5033_;
  assign pg26877 = ~new_n5036_ | new_n5037_;
  assign new_n5039_ = ng2902 & ng2907;
  assign new_n5040_1_ = ng2912 & ng2917;
  assign new_n5041_ = ~new_n5039_ & ~new_n5040_1_;
  assign new_n5042_ = ng2927 & ng2922;
  assign new_n5043_ = new_n5041_ & ~new_n5042_;
  assign new_n5044_ = ng2941 & ng2936;
  assign new_n5045_1_ = new_n5043_ & ~new_n5044_;
  assign new_n5046_ = ng2950 & ng2955;
  assign new_n5047_ = new_n5045_1_ & ~new_n5046_;
  assign new_n5048_ = ng2960 & ng2965;
  assign new_n5049_ = new_n5047_ & ~new_n5048_;
  assign new_n5050_1_ = ng2975 & ng2970;
  assign pg32185 = new_n5049_ & ~new_n5050_1_;
  assign pg23190 = ~ng22 & ~ng25;
  assign new_n5053_ = ng5188 & ng5180;
  assign pg26801 = ng5176 & new_n5053_;
  assign new_n5055_ = ng4507 & ~new_n4724_;
  assign new_n5056_ = ng66 & new_n5055_;
  assign pg33874 = ~new_n5055_ | new_n5056_;
  assign new_n5058_1_ = ng9 & new_n4897_;
  assign new_n5059_ = ng19 & new_n5058_1_;
  assign new_n5060_ = n3414 & new_n5059_;
  assign new_n5061_ = ng19 & new_n4926_1_;
  assign new_n5062_ = n3414 & new_n5061_;
  assign new_n5063_1_ = ~new_n4928_ & ~new_n5060_;
  assign new_n5064_ = ~new_n4959_ & new_n5063_1_;
  assign new_n5065_ = ~new_n5062_ & new_n5064_;
  assign new_n5066_ = new_n4923_ & new_n5065_;
  assign new_n5067_ = ~new_n4931_1_ & new_n5066_;
  assign new_n5068_1_ = new_n4969_ & new_n5065_;
  assign new_n5069_ = ~new_n4931_1_ & new_n5068_1_;
  assign new_n5070_ = new_n4973_ & new_n5065_;
  assign new_n5071_ = ~new_n4931_1_ & new_n5070_;
  assign new_n5072_ = new_n4978_ & new_n5065_;
  assign new_n5073_1_ = ~new_n4931_1_ & new_n5072_;
  assign new_n5074_ = ~new_n5067_ & ~new_n5069_;
  assign new_n5075_ = ~new_n5071_ & ~new_n5073_1_;
  assign new_n5076_ = new_n5074_ & new_n5075_;
  assign new_n5077_1_ = ~new_n4959_ & ~new_n5062_;
  assign new_n5078_ = ~new_n5060_ & new_n5077_1_;
  assign new_n5079_ = ~new_n4920_ & new_n5078_;
  assign new_n5080_ = new_n4990_1_ & new_n5079_;
  assign new_n5081_ = ~new_n4931_1_ & new_n5080_;
  assign new_n5082_1_ = new_n4922_ & new_n5060_;
  assign new_n5083_ = ~new_n4928_ & ~new_n5062_;
  assign new_n5084_ = ~new_n4959_ & new_n5083_;
  assign new_n5085_ = ~new_n4920_ & new_n5084_;
  assign new_n5086_ = new_n5082_1_ & new_n5085_;
  assign new_n5087_1_ = ~new_n4931_1_ & new_n5086_;
  assign new_n5088_ = ~new_n5060_ & new_n5083_;
  assign new_n5089_ = ~new_n4920_ & new_n5088_;
  assign new_n5090_ = new_n5001_ & new_n5089_;
  assign new_n5091_ = ~new_n4931_1_ & new_n5090_;
  assign new_n5092_1_ = new_n4922_ & new_n5062_;
  assign new_n5093_ = ~new_n4920_ & new_n5064_;
  assign new_n5094_ = new_n5092_1_ & new_n5093_;
  assign new_n5095_ = ~new_n4931_1_ & new_n5094_;
  assign new_n5096_ = ~new_n5081_ & ~new_n5087_1_;
  assign new_n5097_1_ = ~new_n5091_ & ~new_n5095_;
  assign new_n5098_ = new_n5096_ & new_n5097_1_;
  assign new_n5099_ = new_n4996_ & new_n5079_;
  assign new_n5100_ = ~new_n4928_ & new_n5099_;
  assign new_n5101_ = new_n5076_ & new_n5098_;
  assign new_n5102_1_ = ~new_n5100_ & new_n5101_;
  assign new_n5103_ = new_n5063_1_ & new_n5077_1_;
  assign new_n5104_ = new_n5013_ & new_n5103_;
  assign new_n5105_ = ~new_n4931_1_ & new_n5104_;
  assign pg34237 = ~new_n5102_1_ | new_n5105_;
  assign new_n5107_1_ = pg35 & ~ng962;
  assign new_n5108_ = pg35 & ~ng1306;
  assign new_n5109_ = ~new_n5107_1_ & new_n5108_;
  assign new_n5110_ = new_n5107_1_ & ~new_n5108_;
  assign new_n5111_ = ~new_n5109_ & ~new_n5110_;
  assign new_n5112_1_ = ~new_n5107_1_ & ~new_n5108_;
  assign pg28042 = ~new_n5111_ | new_n5112_1_;
  assign new_n5114_ = ~new_n4927_ & ~new_n4954_;
  assign new_n5115_ = ~new_n4951_ & new_n5114_;
  assign new_n5116_ = ~new_n4955_1_ & new_n5115_;
  assign new_n5117_1_ = new_n4948_ & new_n5116_;
  assign new_n5118_ = n3414 & ~new_n5117_1_;
  assign new_n5119_ = ~new_n4964_ & ~new_n5060_;
  assign new_n5120_ = ~new_n4925_ & new_n5119_;
  assign new_n5121_ = ~new_n5118_ & new_n5120_;
  assign new_n5122_1_ = new_n4923_ & new_n5121_;
  assign new_n5123_ = ~new_n5062_ & new_n5122_1_;
  assign new_n5124_ = new_n4969_ & new_n5121_;
  assign new_n5125_ = ~new_n5062_ & new_n5124_;
  assign new_n5126_ = new_n4973_ & new_n5121_;
  assign new_n5127_1_ = ~new_n5062_ & new_n5126_;
  assign new_n5128_ = new_n4978_ & new_n5121_;
  assign new_n5129_ = ~new_n5062_ & new_n5128_;
  assign new_n5130_ = ~new_n5123_ & ~new_n5125_;
  assign new_n5131_1_ = ~new_n5127_1_ & ~new_n5129_;
  assign new_n5132_ = new_n5130_ & new_n5131_1_;
  assign new_n5133_ = ~new_n4925_ & ~new_n5118_;
  assign new_n5134_ = ~new_n5060_ & new_n5133_;
  assign new_n5135_ = ~new_n4920_ & new_n5134_;
  assign new_n5136_1_ = new_n5008_ & new_n5135_;
  assign new_n5137_ = ~new_n5062_ & new_n5136_1_;
  assign new_n5138_ = ~new_n4964_ & ~new_n5118_;
  assign new_n5139_ = ~new_n4925_ & new_n5138_;
  assign new_n5140_ = ~new_n4920_ & new_n5139_;
  assign new_n5141_1_ = new_n5082_1_ & new_n5140_;
  assign new_n5142_ = ~new_n5062_ & new_n5141_1_;
  assign new_n5143_ = ~new_n5060_ & new_n5138_;
  assign new_n5144_ = ~new_n4920_ & new_n5143_;
  assign new_n5145_ = new_n4984_ & new_n5144_;
  assign new_n5146_1_ = ~new_n5062_ & new_n5145_;
  assign new_n5147_ = new_n4922_ & new_n5118_;
  assign new_n5148_ = ~new_n4920_ & new_n5120_;
  assign new_n5149_ = new_n5147_ & new_n5148_;
  assign new_n5150_ = ~new_n5062_ & new_n5149_;
  assign new_n5151_1_ = ~new_n5137_ & ~new_n5142_;
  assign new_n5152_ = ~new_n5146_1_ & ~new_n5150_;
  assign new_n5153_ = new_n5151_1_ & new_n5152_;
  assign new_n5154_ = new_n5092_1_ & new_n5135_;
  assign new_n5155_ = ~new_n4964_ & new_n5154_;
  assign new_n5156_1_ = new_n5132_ & new_n5153_;
  assign new_n5157_ = ~new_n5155_ & new_n5156_1_;
  assign new_n5158_ = new_n5119_ & new_n5133_;
  assign new_n5159_ = new_n5013_ & new_n5158_;
  assign new_n5160_ = ~new_n5062_ & new_n5159_;
  assign pg34235 = ~new_n5157_ | new_n5160_;
  assign new_n5162_ = pg72 & ~ng2759;
  assign new_n5163_ = pg72 & ~new_n5162_;
  assign new_n5164_ = ~ng2759 & ~new_n5162_;
  assign new_n5165_ = ~new_n5163_ & ~new_n5164_;
  assign new_n5166_1_ = pg73 & ~ng2763;
  assign new_n5167_ = pg73 & ~new_n5166_1_;
  assign new_n5168_ = ~ng2763 & ~new_n5166_1_;
  assign new_n5169_ = ~new_n5167_ & ~new_n5168_;
  assign new_n5170_ = ~new_n5165_ & ~new_n5169_;
  assign new_n5171_1_ = ~ng2756 & ~ng2741;
  assign new_n5172_ = ~ng2748 & new_n5171_1_;
  assign new_n5173_ = new_n5170_ & new_n5172_;
  assign new_n5174_ = ng2748 & new_n5171_1_;
  assign new_n5175_ = new_n5170_ & new_n5174_;
  assign new_n5176_1_ = ~ng2756 & ng2741;
  assign new_n5177_ = ~ng2748 & new_n5176_1_;
  assign new_n5178_ = new_n5170_ & new_n5177_;
  assign new_n5179_ = ng2748 & new_n5176_1_;
  assign new_n5180_ = new_n5170_ & new_n5179_;
  assign new_n5181_1_ = ~new_n5173_ & ~new_n5175_;
  assign new_n5182_ = ~new_n5178_ & ~new_n5180_;
  assign new_n5183_ = new_n5181_1_ & new_n5182_;
  assign new_n5184_ = pg113 & ~new_n5183_;
  assign new_n5185_ = ~new_n4724_ & new_n5184_;
  assign new_n5186_1_ = ng2756 & ~ng2741;
  assign new_n5187_ = ~ng2748 & new_n5186_1_;
  assign new_n5188_ = new_n5170_ & new_n5187_;
  assign new_n5189_ = ng2748 & new_n5186_1_;
  assign new_n5190_ = new_n5170_ & new_n5189_;
  assign new_n5191_1_ = ng2756 & ng2741;
  assign new_n5192_ = ~ng2748 & new_n5191_1_;
  assign new_n5193_ = new_n5170_ & new_n5192_;
  assign new_n5194_ = ng2748 & new_n5191_1_;
  assign new_n5195_ = new_n5170_ & new_n5194_;
  assign new_n5196_1_ = ~new_n5188_ & ~new_n5190_;
  assign new_n5197_ = ~new_n5193_ & ~new_n5195_;
  assign new_n5198_ = new_n5196_1_ & new_n5197_;
  assign new_n5199_ = pg113 & ~new_n5198_;
  assign new_n5200_ = ~new_n4724_ & new_n5199_;
  assign new_n5201_1_ = ~new_n5185_ & ~new_n5200_;
  assign pg25167 = ~ng1657 & ng1648;
  assign new_n5203_ = new_n5173_ & pg25167;
  assign new_n5204_ = ~ng1926 & ng1917;
  assign new_n5205_ = new_n5175_ & new_n5204_;
  assign new_n5206_1_ = ng1783 & ~ng1792;
  assign new_n5207_ = new_n5178_ & new_n5206_1_;
  assign new_n5208_ = ng2051 & ~ng2060;
  assign new_n5209_ = new_n5180_ & new_n5208_;
  assign new_n5210_ = ~new_n5203_ & ~new_n5205_;
  assign new_n5211_1_ = ~new_n5207_ & ~new_n5209_;
  assign new_n5212_ = new_n5210_ & new_n5211_1_;
  assign new_n5213_ = ~ng2217 & ng2208;
  assign new_n5214_ = new_n5188_ & new_n5213_;
  assign new_n5215_ = ~ng2485 & ng2476;
  assign new_n5216_1_ = new_n5190_ & new_n5215_;
  assign new_n5217_ = ng2342 & ~ng2351;
  assign new_n5218_ = new_n5193_ & new_n5217_;
  assign new_n5219_ = ng2610 & ~ng2619;
  assign new_n5220_ = new_n5195_ & new_n5219_;
  assign new_n5221_1_ = ~new_n5214_ & ~new_n5216_1_;
  assign new_n5222_ = ~new_n5218_ & ~new_n5220_;
  assign new_n5223_ = new_n5221_1_ & new_n5222_;
  assign new_n5224_ = new_n5212_ & new_n5223_;
  assign new_n5225_ = ~new_n5201_1_ & ~new_n5224_;
  assign pg34201 = new_n5201_1_ | new_n5225_;
  assign new_n5227_ = ~new_n4925_ & ~new_n5062_;
  assign new_n5228_ = ~new_n4964_ & new_n5227_;
  assign new_n5229_ = ~new_n5118_ & new_n5228_;
  assign new_n5230_ = new_n4923_ & new_n5229_;
  assign new_n5231_1_ = ~new_n5060_ & new_n5230_;
  assign new_n5232_ = new_n4969_ & new_n5229_;
  assign new_n5233_ = ~new_n5060_ & new_n5232_;
  assign new_n5234_ = new_n4973_ & new_n5229_;
  assign new_n5235_1_ = ~new_n5060_ & new_n5234_;
  assign new_n5236_ = new_n4978_ & new_n5229_;
  assign new_n5237_ = ~new_n5060_ & new_n5236_;
  assign new_n5238_ = ~new_n5231_1_ & ~new_n5233_;
  assign new_n5239_ = ~new_n5235_1_ & ~new_n5237_;
  assign new_n5240_1_ = new_n5238_ & new_n5239_;
  assign new_n5241_ = new_n5092_1_ & new_n5140_;
  assign new_n5242_ = ~new_n5060_ & new_n5241_;
  assign new_n5243_ = ~new_n5062_ & ~new_n5118_;
  assign new_n5244_ = ~new_n4964_ & new_n5243_;
  assign new_n5245_1_ = ~new_n4920_ & new_n5244_;
  assign new_n5246_ = new_n4984_ & new_n5245_1_;
  assign new_n5247_ = ~new_n5060_ & new_n5246_;
  assign new_n5248_ = ~new_n4925_ & new_n5243_;
  assign new_n5249_1_ = ~new_n4920_ & new_n5248_;
  assign new_n5250_ = new_n5008_ & new_n5249_1_;
  assign new_n5251_ = ~new_n5060_ & new_n5250_;
  assign new_n5252_ = ~new_n4920_ & new_n5228_;
  assign new_n5253_ = new_n5147_ & new_n5252_;
  assign new_n5254_1_ = ~new_n5060_ & new_n5253_;
  assign new_n5255_ = ~new_n5242_ & ~new_n5247_;
  assign new_n5256_ = ~new_n5251_ & ~new_n5254_1_;
  assign new_n5257_ = new_n5255_ & new_n5256_;
  assign new_n5258_1_ = new_n5240_1_ & new_n5257_;
  assign new_n5259_ = ~new_n5142_ & new_n5258_1_;
  assign new_n5260_ = new_n5138_ & new_n5227_;
  assign new_n5261_ = new_n5013_ & new_n5260_;
  assign new_n5262_ = ~new_n5060_ & new_n5261_;
  assign pg34236 = ~new_n5259_ | new_n5262_;
  assign new_n5264_ = ~pg56 & pg54;
  assign new_n5265_ = ng55 & ~new_n5264_;
  assign new_n5266_ = ng1300 & ~ng1291;
  assign new_n5267_ = new_n4920_ & new_n5266_;
  assign new_n5268_1_ = ng538 & new_n4910_;
  assign new_n5269_ = pg35 & ~ng595;
  assign new_n5270_ = new_n4899_ & ~new_n5269_;
  assign new_n5271_ = pg35 & ~ng632;
  assign new_n5272_ = new_n4913_ & ~new_n5271_;
  assign new_n5273_1_ = ~new_n5270_ & ~new_n5272_;
  assign new_n5274_ = pg35 & ~ng776;
  assign new_n5275_ = new_n4905_ & ~new_n5274_;
  assign new_n5276_ = ~new_n5268_1_ & new_n5273_1_;
  assign new_n5277_ = ~new_n5275_ & new_n5276_;
  assign new_n5278_1_ = new_n4916_1_ & ~new_n5277_;
  assign new_n5279_ = ~ng947 & ng956;
  assign new_n5280_ = new_n4893_ & new_n5279_;
  assign new_n5281_ = ng45 & new_n4894_;
  assign new_n5282_ = ~new_n5267_ & ~new_n5278_1_;
  assign new_n5283_1_ = ~new_n5280_ & ~new_n5281_;
  assign new_n5284_ = new_n5282_ & new_n5283_1_;
  assign new_n5285_ = ng4917 & new_n4964_;
  assign new_n5286_ = ng3853 & new_n5060_;
  assign new_n5287_ = ng4727 & new_n4925_;
  assign new_n5288_1_ = ng2907 & new_n4942_;
  assign new_n5289_ = ng2902 & new_n4937_;
  assign new_n5290_ = ~new_n5288_1_ & ~new_n5289_;
  assign new_n5291_ = ng2844 & new_n4927_;
  assign new_n5292_ = ng2848 & new_n4955_1_;
  assign new_n5293_1_ = ~new_n5291_ & ~new_n5292_;
  assign new_n5294_ = new_n5290_ & new_n5293_1_;
  assign new_n5295_ = new_n5118_ & ~new_n5294_;
  assign new_n5296_ = ~new_n5285_ & ~new_n5286_;
  assign new_n5297_ = ~new_n5287_ & ~new_n5295_;
  assign new_n5298_1_ = new_n5296_ & new_n5297_;
  assign new_n5299_ = ng6199 & new_n5062_;
  assign new_n5300_ = new_n5284_ & new_n5298_1_;
  assign n4955 = new_n5299_ | ~new_n5300_;
  assign new_n5302_ = ng1472 & ~ng1291;
  assign new_n5303_1_ = new_n4920_ & new_n5302_;
  assign new_n5304_ = pg35 & ~ng590;
  assign new_n5305_ = new_n4899_ & ~new_n5304_;
  assign new_n5306_ = pg35 & ~ng626;
  assign new_n5307_ = new_n4913_ & ~new_n5306_;
  assign new_n5308_1_ = ~new_n5305_ & ~new_n5307_;
  assign new_n5309_ = pg35 & ~ng772;
  assign new_n5310_ = new_n4905_ & ~new_n5309_;
  assign new_n5311_ = new_n5308_1_ & ~new_n5310_;
  assign new_n5312_1_ = new_n4916_1_ & ~new_n5311_;
  assign new_n5313_ = ~ng947 & ng1129;
  assign new_n5314_ = new_n4893_ & new_n5313_;
  assign new_n5315_ = ng46 & new_n4894_;
  assign new_n5316_1_ = ~new_n5303_1_ & ~new_n5312_1_;
  assign new_n5317_ = ~new_n5314_ & ~new_n5315_;
  assign new_n5318_ = new_n5316_1_ & new_n5317_;
  assign new_n5319_ = ng4922 & new_n4964_;
  assign new_n5320_ = ng3502 & new_n5060_;
  assign new_n5321_1_ = ng4732 & new_n4925_;
  assign new_n5322_ = ng2912 & new_n4942_;
  assign new_n5323_ = ng2917 & new_n4937_;
  assign new_n5324_ = ~new_n5322_ & ~new_n5323_;
  assign new_n5325_ = ng2852 & new_n4927_;
  assign new_n5326_1_ = ng2999 & new_n4954_;
  assign new_n5327_ = ng2856 & new_n4955_1_;
  assign new_n5328_ = ~new_n5325_ & ~new_n5326_1_;
  assign new_n5329_ = ~new_n5327_ & new_n5328_;
  assign new_n5330_1_ = new_n5324_ & new_n5329_;
  assign new_n5331_ = new_n5118_ & ~new_n5330_1_;
  assign new_n5332_ = ~new_n5319_ & ~new_n5320_;
  assign new_n5333_ = ~new_n5321_1_ & ~new_n5331_;
  assign new_n5334_1_ = new_n5332_ & new_n5333_;
  assign new_n5335_ = ng5853 & new_n5062_;
  assign new_n5336_ = new_n5318_ & new_n5334_1_;
  assign n3583 = new_n5335_ | ~new_n5336_;
  assign new_n5338_ = n4955 & n3583;
  assign new_n5339_1_ = n4955 & ~new_n5338_;
  assign new_n5340_ = n3583 & ~new_n5338_;
  assign new_n5341_ = ~new_n5339_1_ & ~new_n5340_;
  assign new_n5342_ = ng1448 & ~ng1291;
  assign new_n5343_ = new_n4920_ & new_n5342_;
  assign new_n5344_1_ = pg35 & ~ng582;
  assign new_n5345_ = new_n4899_ & ~new_n5344_1_;
  assign new_n5346_ = pg35 & ~ng622;
  assign new_n5347_ = new_n4913_ & ~new_n5346_;
  assign new_n5348_ = ~new_n5345_ & ~new_n5347_;
  assign new_n5349_1_ = pg35 & ~ng554;
  assign new_n5350_ = new_n4900_ & ~new_n5349_1_;
  assign new_n5351_ = ng546 & new_n4910_;
  assign new_n5352_ = pg35 & ~ng767;
  assign new_n5353_1_ = new_n4905_ & ~new_n5352_;
  assign new_n5354_ = new_n5348_ & ~new_n5350_;
  assign new_n5355_ = ~new_n5351_ & ~new_n5353_1_;
  assign new_n5356_ = new_n5354_ & new_n5355_;
  assign new_n5357_ = new_n4916_1_ & ~new_n5356_;
  assign new_n5358_1_ = ~ng947 & ng1105;
  assign new_n5359_ = new_n4893_ & new_n5358_1_;
  assign new_n5360_ = ng47 & new_n4894_;
  assign new_n5361_ = ~new_n5343_ & ~new_n5357_;
  assign new_n5362_ = ~new_n5359_ & ~new_n5360_;
  assign new_n5363_1_ = new_n5361_ & new_n5362_;
  assign new_n5364_ = ng4907 & new_n4964_;
  assign new_n5365_ = ng3151 & new_n5060_;
  assign new_n5366_ = ng4717 & new_n4925_;
  assign new_n5367_ = ng2922 & new_n4942_;
  assign new_n5368_1_ = ng2927 & new_n4937_;
  assign new_n5369_ = ~new_n5367_ & ~new_n5368_1_;
  assign new_n5370_ = ng2860 & new_n4927_;
  assign new_n5371_ = ~ng2994 & new_n4954_;
  assign new_n5372_ = ng2864 & new_n4955_1_;
  assign new_n5373_1_ = ~new_n5370_ & ~new_n5371_;
  assign new_n5374_ = ~new_n5372_ & new_n5373_1_;
  assign new_n5375_ = new_n5369_ & new_n5374_;
  assign new_n5376_ = new_n5118_ & ~new_n5375_;
  assign new_n5377_ = ~new_n5364_ & ~new_n5365_;
  assign new_n5378_1_ = ~new_n5366_ & ~new_n5376_;
  assign new_n5379_ = new_n5377_ & new_n5378_1_;
  assign new_n5380_ = ng5507 & new_n5062_;
  assign new_n5381_ = new_n5363_1_ & new_n5379_;
  assign n5814 = new_n5380_ | ~new_n5381_;
  assign new_n5383_1_ = ng1478 & ~ng1291;
  assign new_n5384_ = new_n4920_ & new_n5383_1_;
  assign new_n5385_ = pg35 & ~ng577;
  assign new_n5386_ = new_n4899_ & ~new_n5385_;
  assign new_n5387_1_ = pg35 & ~ng617;
  assign new_n5388_ = new_n4913_ & ~new_n5387_1_;
  assign new_n5389_ = ~new_n5386_ & ~new_n5388_;
  assign new_n5390_ = pg35 & ~ng807;
  assign new_n5391_ = new_n4900_ & ~new_n5390_;
  assign new_n5392_1_ = ng542 & new_n4910_;
  assign new_n5393_ = pg35 & ~ng763;
  assign new_n5394_ = new_n4905_ & ~new_n5393_;
  assign new_n5395_ = new_n5389_ & ~new_n5391_;
  assign new_n5396_ = ~new_n5392_1_ & ~new_n5394_;
  assign new_n5397_1_ = new_n5395_ & new_n5396_;
  assign new_n5398_ = new_n4916_1_ & ~new_n5397_1_;
  assign new_n5399_ = ng1135 & ~ng947;
  assign new_n5400_ = new_n4893_ & new_n5399_;
  assign new_n5401_ = ng48 & new_n4894_;
  assign new_n5402_1_ = ~new_n5384_ & ~new_n5398_;
  assign new_n5403_ = ~new_n5400_ & ~new_n5401_;
  assign new_n5404_ = new_n5402_1_ & new_n5403_;
  assign new_n5405_ = ng5160 & new_n5062_;
  assign new_n5406_ = ng4722 & new_n4925_;
  assign new_n5407_1_ = ng4912 & new_n4964_;
  assign new_n5408_ = ng2941 & new_n4937_;
  assign new_n5409_ = ng2936 & new_n4942_;
  assign new_n5410_ = ~new_n5408_ & ~new_n5409_;
  assign new_n5411_ = ~new_n4941_ & new_n5410_;
  assign new_n5412_1_ = ng2894 & new_n4927_;
  assign new_n5413_ = ng2988 & new_n4954_;
  assign new_n5414_ = ng2898 & new_n4955_1_;
  assign new_n5415_ = ~new_n5412_1_ & ~new_n5413_;
  assign new_n5416_ = ~new_n5414_ & new_n5415_;
  assign new_n5417_1_ = new_n5411_ & new_n5416_;
  assign new_n5418_ = new_n5118_ & ~new_n5417_1_;
  assign new_n5419_ = ~new_n5405_ & ~new_n5406_;
  assign new_n5420_ = ~new_n5407_1_ & ~new_n5418_;
  assign new_n5421_ = new_n5419_ & new_n5420_;
  assign new_n5422_1_ = ng6545 & new_n5060_;
  assign new_n5423_ = new_n5404_ & new_n5421_;
  assign n2287 = new_n5422_1_ | ~new_n5423_;
  assign new_n5425_ = n5814 & n2287;
  assign new_n5426_ = n5814 & ~new_n5425_;
  assign new_n5427_1_ = n2287 & ~new_n5425_;
  assign new_n5428_ = ~new_n5426_ & ~new_n5427_1_;
  assign new_n5429_ = ~new_n5341_ & ~new_n5428_;
  assign new_n5430_ = ~new_n5341_ & ~new_n5429_;
  assign new_n5431_ = ~new_n5428_ & ~new_n5429_;
  assign new_n5432_1_ = ~new_n5430_ & ~new_n5431_;
  assign new_n5433_ = ng1291 & new_n4920_;
  assign new_n5434_ = pg35 & ~ng586;
  assign new_n5435_ = new_n4899_ & ~new_n5434_;
  assign new_n5436_ = pg35 & ~ng613;
  assign new_n5437_1_ = new_n4913_ & ~new_n5436_;
  assign new_n5438_ = ~new_n5435_ & ~new_n5437_1_;
  assign new_n5439_ = pg35 & ~ng794;
  assign new_n5440_ = new_n4900_ & ~new_n5439_;
  assign new_n5441_ = ng534 & new_n4910_;
  assign new_n5442_1_ = pg35 & ~ng758;
  assign new_n5443_ = new_n4905_ & ~new_n5442_1_;
  assign new_n5444_ = new_n5438_ & ~new_n5440_;
  assign new_n5445_ = ~new_n5441_ & ~new_n5443_;
  assign new_n5446_ = new_n5444_ & new_n5445_;
  assign new_n5447_1_ = new_n4916_1_ & ~new_n5446_;
  assign new_n5448_ = ng947 & new_n4893_;
  assign new_n5449_ = ng49 & new_n4894_;
  assign new_n5450_ = ~new_n5433_ & ~new_n5447_1_;
  assign new_n5451_ = ~new_n5448_ & ~new_n5449_;
  assign new_n5452_1_ = new_n5450_ & new_n5451_;
  assign new_n5453_ = ~ng4737 & new_n4925_;
  assign new_n5454_ = ng4172 & new_n4928_;
  assign new_n5455_ = ng4300 & new_n4931_1_;
  assign new_n5456_ = ng2955 & new_n4937_;
  assign new_n5457_1_ = ng2950 & new_n4942_;
  assign new_n5458_ = ~new_n5456_ & ~new_n5457_1_;
  assign new_n5459_ = ~new_n4941_ & new_n5458_;
  assign new_n5460_ = ng37 & new_n4951_;
  assign new_n5461_ = ng2868 & new_n4954_;
  assign new_n5462_1_ = ng2882 & new_n4955_1_;
  assign new_n5463_ = ~new_n5460_ & ~new_n5461_;
  assign new_n5464_ = ~new_n5462_1_ & new_n5463_;
  assign new_n5465_ = new_n5459_ & new_n5464_;
  assign new_n5466_ = new_n4959_ & ~new_n5465_;
  assign new_n5467_1_ = ~new_n5453_ & ~new_n5454_;
  assign new_n5468_ = ~new_n5455_ & ~new_n5466_;
  assign new_n5469_ = new_n5467_1_ & new_n5468_;
  assign new_n5470_ = ~ng4927 & new_n4964_;
  assign new_n5471_ = new_n5452_1_ & new_n5469_;
  assign n6079 = new_n5470_ | ~new_n5471_;
  assign new_n5473_ = ~ng1296 & new_n4920_;
  assign new_n5474_ = pg35 & ~ng572;
  assign new_n5475_ = new_n4899_ & ~new_n5474_;
  assign new_n5476_ = pg35 & ~ng608;
  assign new_n5477_1_ = new_n4913_ & ~new_n5476_;
  assign new_n5478_ = ~new_n5475_ & ~new_n5477_1_;
  assign new_n5479_ = pg35 & ~ng790;
  assign new_n5480_1_ = new_n4900_ & ~new_n5479_;
  assign new_n5481_ = ~ng550 & new_n4910_;
  assign new_n5482_ = pg35 & ~ng749;
  assign new_n5483_ = new_n4905_ & ~new_n5482_;
  assign new_n5484_ = new_n5478_ & ~new_n5480_1_;
  assign new_n5485_1_ = ~new_n5481_ & ~new_n5483_;
  assign new_n5486_ = new_n5484_ & new_n5485_1_;
  assign new_n5487_ = new_n4916_1_ & ~new_n5486_;
  assign new_n5488_ = ~ng952 & new_n4893_;
  assign new_n5489_ = ng50 & new_n4894_;
  assign new_n5490_1_ = ~new_n5473_ & ~new_n5487_;
  assign new_n5491_ = ~new_n5488_ & ~new_n5489_;
  assign new_n5492_ = new_n5490_1_ & new_n5491_;
  assign new_n5493_ = ng4176 & new_n4928_;
  assign new_n5494_ = ng2689 & new_n5060_;
  assign new_n5495_1_ = ng2960 & new_n4942_;
  assign new_n5496_ = ng2965 & new_n4937_;
  assign new_n5497_ = ~new_n5495_1_ & ~new_n5496_;
  assign new_n5498_ = ng94 & new_n4951_;
  assign new_n5499_ = ng2873 & new_n4954_;
  assign new_n5500_1_ = ng2878 & new_n4955_1_;
  assign new_n5501_ = ~new_n5498_ & ~new_n5499_;
  assign new_n5502_ = ~new_n5500_1_ & new_n5501_;
  assign new_n5503_ = new_n5497_ & new_n5502_;
  assign new_n5504_ = new_n4959_ & ~new_n5503_;
  assign new_n5505_1_ = ng2130 & new_n5062_;
  assign new_n5506_ = ~new_n5493_ & ~new_n5494_;
  assign new_n5507_ = ~new_n5504_ & ~new_n5505_1_;
  assign new_n5508_ = new_n5506_ & new_n5507_;
  assign new_n5509_1_ = ng4253 & new_n4931_1_;
  assign new_n5510_ = new_n5492_ & new_n5508_;
  assign n4465 = new_n5509_1_ | ~new_n5510_;
  assign new_n5512_ = n6079 & n4465;
  assign new_n5513_ = n6079 & ~new_n5512_;
  assign new_n5514_1_ = n4465 & ~new_n5512_;
  assign new_n5515_ = ~new_n5513_ & ~new_n5514_1_;
  assign new_n5516_ = ng1283 & new_n4920_;
  assign new_n5517_ = pg35 & ~ng568;
  assign new_n5518_ = new_n4899_ & ~new_n5517_;
  assign new_n5519_1_ = pg35 & ~ng604;
  assign new_n5520_ = new_n4913_ & ~new_n5519_1_;
  assign new_n5521_ = ~new_n5518_ & ~new_n5520_;
  assign new_n5522_ = pg35 & ~ng785;
  assign new_n5523_ = new_n4900_ & ~new_n5522_;
  assign new_n5524_1_ = ng136 & new_n4910_;
  assign new_n5525_ = pg35 & ~ng744;
  assign new_n5526_ = new_n4905_ & ~new_n5525_;
  assign new_n5527_ = new_n5521_ & ~new_n5523_;
  assign new_n5528_ = ~new_n5524_1_ & ~new_n5526_;
  assign new_n5529_1_ = new_n5527_ & new_n5528_;
  assign new_n5530_ = new_n4916_1_ & ~new_n5529_1_;
  assign new_n5531_ = ng939 & new_n4893_;
  assign new_n5532_ = ng51 & new_n4894_;
  assign new_n5533_1_ = ~new_n5516_ & ~new_n5530_;
  assign new_n5534_ = ~new_n5531_ & ~new_n5532_;
  assign new_n5535_ = new_n5533_1_ & new_n5534_;
  assign new_n5536_ = ng4146 & new_n4928_;
  assign new_n5537_1_ = ng2697 & new_n5060_;
  assign new_n5538_ = ng2975 & new_n4937_;
  assign new_n5539_ = ng2970 & new_n4942_;
  assign new_n5540_ = ng2980 & new_n4945_1_;
  assign new_n5541_ = ~new_n5538_ & ~new_n5539_;
  assign new_n5542_1_ = ~new_n5540_ & new_n5541_;
  assign new_n5543_ = pg92 & new_n4951_;
  assign new_n5544_ = pg127 & new_n4954_;
  assign new_n5545_ = ng2886 & new_n4955_1_;
  assign new_n5546_ = ~new_n5543_ & ~new_n5544_;
  assign new_n5547_1_ = ~new_n5545_ & new_n5546_;
  assign new_n5548_ = new_n5542_1_ & new_n5547_1_;
  assign new_n5549_ = new_n4959_ & ~new_n5548_;
  assign new_n5550_ = ng2138 & new_n5062_;
  assign new_n5551_ = ~new_n5536_ & ~new_n5537_1_;
  assign new_n5552_1_ = ~new_n5549_ & ~new_n5550_;
  assign new_n5553_ = new_n5551_ & new_n5552_1_;
  assign new_n5554_ = ng4249 & new_n4931_1_;
  assign new_n5555_ = new_n5535_ & new_n5553_;
  assign n5005 = new_n5554_ | ~new_n5555_;
  assign new_n5557_1_ = ng1287 & new_n4920_;
  assign new_n5558_ = pg35 & ~ng562;
  assign new_n5559_ = new_n4899_ & ~new_n5558_;
  assign new_n5560_ = pg35 & ~ng599;
  assign new_n5561_ = new_n4913_ & ~new_n5560_;
  assign new_n5562_1_ = ~new_n5559_ & ~new_n5561_;
  assign new_n5563_ = pg35 & ~ng739;
  assign new_n5564_ = new_n4905_ & ~new_n5563_;
  assign new_n5565_ = pg35 & ~ng781;
  assign new_n5566_1_ = new_n4900_ & ~new_n5565_;
  assign new_n5567_ = ng199 & new_n4910_;
  assign new_n5568_ = new_n5562_1_ & ~new_n5564_;
  assign new_n5569_ = ~new_n5566_1_ & ~new_n5567_;
  assign new_n5570_1_ = new_n5568_ & new_n5569_;
  assign new_n5571_ = new_n4916_1_ & ~new_n5570_1_;
  assign new_n5572_ = ng943 & new_n4893_;
  assign new_n5573_ = ng52 & new_n4894_;
  assign new_n5574_ = ~new_n5557_1_ & ~new_n5571_;
  assign new_n5575_1_ = ~new_n5572_ & ~new_n5573_;
  assign new_n5576_ = new_n5574_ & new_n5575_1_;
  assign new_n5577_ = ng4157 & new_n4928_;
  assign new_n5578_ = ng2704 & new_n5060_;
  assign new_n5579_ = ng2984 & new_n4945_1_;
  assign new_n5580_1_ = ~new_n4941_ & ~new_n5579_;
  assign new_n5581_ = ng2890 & new_n4954_;
  assign new_n5582_ = pg100 & new_n4951_;
  assign new_n5583_ = ~new_n5581_ & ~new_n5582_;
  assign new_n5584_ = new_n5580_1_ & new_n5583_;
  assign new_n5585_1_ = new_n4959_ & ~new_n5584_;
  assign new_n5586_ = ng2145 & new_n5062_;
  assign new_n5587_ = ~new_n5577_ & ~new_n5578_;
  assign new_n5588_ = ~new_n5585_1_ & ~new_n5586_;
  assign new_n5589_ = new_n5587_ & new_n5588_;
  assign new_n5590_1_ = ng4245 & new_n4931_1_;
  assign new_n5591_ = new_n5576_ & new_n5589_;
  assign n2272 = new_n5590_1_ | ~new_n5591_;
  assign new_n5593_ = n5005 & n2272;
  assign new_n5594_1_ = n5005 & ~new_n5593_;
  assign new_n5595_ = n2272 & ~new_n5593_;
  assign new_n5596_ = ~new_n5594_1_ & ~new_n5595_;
  assign new_n5597_ = ~new_n5515_ & ~new_n5596_;
  assign new_n5598_1_ = ~new_n5515_ & ~new_n5597_;
  assign new_n5599_ = ~new_n5596_ & ~new_n5597_;
  assign new_n5600_ = ~new_n5598_1_ & ~new_n5599_;
  assign new_n5601_ = ~new_n5432_1_ & ~new_n5600_;
  assign new_n5602_ = ~new_n5432_1_ & ~new_n5601_;
  assign new_n5603_1_ = ~new_n5600_ & ~new_n5601_;
  assign new_n5604_ = ~new_n5602_ & ~new_n5603_1_;
  assign new_n5605_ = ~new_n5265_ & ~new_n5604_;
  assign new_n5606_ = ~new_n5265_ & ~new_n5605_;
  assign new_n5607_ = ~new_n5604_ & ~new_n5605_;
  assign n3854 = new_n5606_ | new_n5607_;
  assign new_n5609_ = ng22 & n3854;
  assign pg34972 = ~ng22 | new_n5609_;
  assign new_n5611_ = ng4322 & ~ng4311;
  assign new_n5612_ = ng4332 & new_n5611_;
  assign new_n5613_1_ = pg72 & ~new_n5612_;
  assign new_n5614_ = ~ng4322 & ~ng4311;
  assign new_n5615_ = ng4332 & new_n5614_;
  assign new_n5616_ = ~pg72 & ~new_n5615_;
  assign new_n5617_ = ~new_n5613_1_ & ~new_n5616_;
  assign new_n5618_1_ = pg73 & new_n5617_;
  assign new_n5619_ = ~ng4332 & new_n5611_;
  assign new_n5620_ = pg72 & ~new_n5619_;
  assign new_n5621_ = ~ng4332 & new_n5614_;
  assign new_n5622_ = ~pg72 & ~new_n5621_;
  assign new_n5623_1_ = ~new_n5620_ & ~new_n5622_;
  assign new_n5624_ = ~pg73 & new_n5623_1_;
  assign new_n5625_ = ~new_n5618_1_ & ~new_n5624_;
  assign new_n5626_ = ~ng4366 & ~new_n5625_;
  assign pg34956 = ng4369 & ~new_n5626_;
  assign new_n5628_1_ = pg73 & ng490;
  assign new_n5629_ = ng490 & ~new_n5628_1_;
  assign new_n5630_ = pg73 & ~new_n5628_1_;
  assign new_n5631_ = ~new_n5629_ & ~new_n5630_;
  assign new_n5632_ = pg72 & ng482;
  assign new_n5633_1_ = ng482 & ~new_n5632_;
  assign new_n5634_ = pg72 & ~new_n5632_;
  assign new_n5635_ = ~new_n5633_1_ & ~new_n5634_;
  assign new_n5636_ = new_n5631_ & new_n5635_;
  assign new_n5637_ = ~ng504 & new_n5636_;
  assign new_n5638_1_ = ~ng518 & new_n5637_;
  assign new_n5639_ = ~ng528 & new_n5638_1_;
  assign new_n5640_ = ng504 & new_n5636_;
  assign new_n5641_ = ng518 & new_n5640_;
  assign new_n5642_ = ~ng528 & new_n5641_;
  assign new_n5643_1_ = ~ng518 & new_n5640_;
  assign new_n5644_ = ~ng528 & new_n5643_1_;
  assign new_n5645_ = ng518 & new_n5637_;
  assign new_n5646_ = ~ng528 & new_n5645_;
  assign new_n5647_ = ~new_n5639_ & ~new_n5642_;
  assign new_n5648_1_ = ~new_n5644_ & ~new_n5646_;
  assign new_n5649_ = new_n5647_ & new_n5648_1_;
  assign new_n5650_ = pg113 & ~new_n5649_;
  assign new_n5651_ = ~new_n4724_ & new_n5650_;
  assign new_n5652_ = ng528 & new_n5638_1_;
  assign new_n5653_1_ = ng528 & new_n5641_;
  assign new_n5654_ = ng528 & new_n5643_1_;
  assign new_n5655_ = ng528 & new_n5645_;
  assign new_n5656_ = ~new_n5652_ & ~new_n5653_1_;
  assign new_n5657_ = ~new_n5654_ & ~new_n5655_;
  assign new_n5658_1_ = new_n5656_ & new_n5657_;
  assign new_n5659_ = pg113 & ~new_n5658_1_;
  assign new_n5660_ = ~new_n4724_ & new_n5659_;
  assign new_n5661_ = ~new_n5651_ & ~new_n5660_;
  assign new_n5662_ = new_n4734_ & new_n4737_1_;
  assign new_n5663_1_ = new_n4735_ & new_n4737_1_;
  assign new_n5664_ = ~new_n5662_ & ~new_n5663_1_;
  assign new_n5665_ = ng4785 & ng4709;
  assign new_n5666_ = ~ng4801 & ng4793;
  assign new_n5667_ = ng4776 & new_n5666_;
  assign new_n5668_1_ = ng4653 & ng4659;
  assign new_n5669_ = ng4669 & new_n5668_1_;
  assign new_n5670_ = ng4688 & new_n5669_;
  assign new_n5671_ = new_n4734_ & new_n5665_;
  assign new_n5672_1_ = new_n5667_ & new_n5671_;
  assign new_n5673_ = new_n5670_ & new_n5672_1_;
  assign new_n5674_ = ng4975 & ng4899;
  assign new_n5675_ = ~ng4991 & ng4983;
  assign new_n5676_ = ng4966 & new_n5675_;
  assign new_n5677_1_ = ng4849 & ng4843;
  assign new_n5678_ = ng4859 & new_n5677_1_;
  assign new_n5679_ = ng4878 & new_n5678_;
  assign new_n5680_ = new_n4735_ & new_n5674_;
  assign new_n5681_ = new_n5676_ & new_n5680_;
  assign new_n5682_1_ = new_n5679_ & new_n5681_;
  assign new_n5683_ = ~new_n5673_ & ~new_n5682_1_;
  assign new_n5684_ = ~new_n5664_ & ~new_n5683_;
  assign pg34221 = new_n5664_ | new_n5684_;
  assign pg25259 = ng1668 & ~ng1636;
  assign new_n5687_1_ = ng5002 & ng5005;
  assign new_n5688_ = ~new_n4724_ & new_n5687_1_;
  assign new_n5689_ = ~ng4801 & ~ng4793;
  assign new_n5690_ = ng4776 & new_n5689_;
  assign new_n5691_ = ~ng4785 & new_n5690_;
  assign new_n5692_1_ = ~ng4709 & new_n5691_;
  assign new_n5693_ = new_n5669_ & new_n5692_1_;
  assign new_n5694_ = ng4698 & new_n5693_;
  assign pg33959 = ng4646 & ~new_n5694_;
  assign new_n5696_ = ng22 & n5005;
  assign pg34927 = ~ng22 | new_n5696_;
  assign new_n5698_ = ng22 & n3583;
  assign pg34917 = ~ng22 | new_n5698_;
  assign new_n5700_ = ng4812 & ng4815;
  assign new_n5701_ = ~new_n4724_ & new_n5700_;
  assign new_n5702_1_ = ng22 & n5814;
  assign pg34919 = ~ng22 | new_n5702_1_;
  assign new_n5704_ = ng1668 & new_n5639_;
  assign new_n5705_ = ~ng1636 & new_n5704_;
  assign new_n5706_ = ng1936 & new_n5642_;
  assign new_n5707_1_ = ~ng1906 & new_n5706_;
  assign new_n5708_ = ng1802 & new_n5644_;
  assign new_n5709_ = ~ng1772 & new_n5708_;
  assign new_n5710_ = ng2070 & new_n5646_;
  assign new_n5711_ = ~ng2040 & new_n5710_;
  assign new_n5712_1_ = ~new_n5705_ & ~new_n5707_1_;
  assign new_n5713_ = ~new_n5709_ & ~new_n5711_;
  assign new_n5714_ = new_n5712_1_ & new_n5713_;
  assign new_n5715_ = ng2227 & new_n5652_;
  assign new_n5716_ = ~ng2197 & new_n5715_;
  assign new_n5717_1_ = ng2495 & new_n5653_1_;
  assign new_n5718_ = ~ng2465 & new_n5717_1_;
  assign new_n5719_ = ng2361 & new_n5654_;
  assign new_n5720_ = ~ng2331 & new_n5719_;
  assign new_n5721_ = ng2629 & new_n5655_;
  assign new_n5722_1_ = ~ng2599 & new_n5721_;
  assign new_n5723_ = ~new_n5716_ & ~new_n5718_;
  assign new_n5724_ = ~new_n5720_ & ~new_n5722_1_;
  assign new_n5725_ = new_n5723_ & new_n5724_;
  assign new_n5726_ = new_n5714_ & new_n5725_;
  assign new_n5727_1_ = ~new_n5661_ & ~new_n5726_;
  assign pg34383 = new_n5661_ | new_n5727_1_;
  assign new_n5729_ = ng22 & n6079;
  assign pg34923 = ~ng22 | new_n5729_;
  assign new_n5731_ = ~ng2819 & ng2724;
  assign new_n5732_1_ = ~ng2815 & ~ng2724;
  assign new_n5733_ = ~new_n5731_ & ~new_n5732_1_;
  assign new_n5734_ = ng2729 & new_n5733_;
  assign new_n5735_ = ng2724 & ~ng2807;
  assign new_n5736_ = ~ng2803 & ~ng2724;
  assign new_n5737_1_ = ~new_n5735_ & ~new_n5736_;
  assign new_n5738_ = ~ng2729 & new_n5737_1_;
  assign pg33079 = ~new_n5734_ & ~new_n5738_;
  assign new_n5740_ = ng22 & n4955;
  assign pg34913 = ~ng22 | new_n5740_;
  assign new_n5742_1_ = ~ng4975 & ~ng4899;
  assign new_n5743_ = ng4888 & new_n5742_1_;
  assign new_n5744_ = ~ng4975 & ng4899;
  assign new_n5745_ = ng4944 & new_n5744_;
  assign new_n5746_ = ng4975 & ~ng4899;
  assign new_n5747_1_ = ng4933 & new_n5746_;
  assign new_n5748_ = ng4955 & new_n5674_;
  assign new_n5749_ = ~new_n5743_ & ~new_n5745_;
  assign new_n5750_ = ~new_n5747_1_ & ~new_n5748_;
  assign new_n5751_ = new_n5749_ & new_n5750_;
  assign new_n5752_1_ = new_n5688_ & ~new_n5751_;
  assign pg33935 = ~new_n5688_ | new_n5752_1_;
  assign new_n5754_ = ng22 & n4465;
  assign pg34925 = ~ng22 | new_n5754_;
  assign new_n5756_ = ng22 & n2272;
  assign pg34915 = ~ng22 | new_n5756_;
  assign new_n5758_ = pg72 & ~ng4108;
  assign new_n5759_ = pg72 & ~new_n5758_;
  assign new_n5760_ = ~ng4108 & ~new_n5758_;
  assign new_n5761_ = ~new_n5759_ & ~new_n5760_;
  assign new_n5762_1_ = pg73 & ~ng4104;
  assign new_n5763_ = pg73 & ~new_n5762_1_;
  assign new_n5764_ = ~ng4104 & ~new_n5762_1_;
  assign new_n5765_ = ~new_n5763_ & ~new_n5764_;
  assign new_n5766_1_ = ~new_n5761_ & ~new_n5765_;
  assign new_n5767_ = new_n4737_1_ & new_n5766_1_;
  assign new_n5768_ = ~ng4087 & ~ng4098;
  assign new_n5769_ = ~ng4093 & new_n5768_;
  assign new_n5770_ = new_n5766_1_ & new_n5769_;
  assign new_n5771_1_ = ng5180 & new_n5770_;
  assign new_n5772_ = ng5188 & new_n5771_1_;
  assign new_n5773_ = ng5176 & new_n5772_;
  assign new_n5774_ = ng4093 & new_n5768_;
  assign new_n5775_ = new_n5766_1_ & new_n5774_;
  assign new_n5776_1_ = ng5873 & new_n5775_;
  assign new_n5777_ = ng5881 & new_n5776_1_;
  assign new_n5778_ = ng5869 & new_n5777_;
  assign new_n5779_ = ng4087 & ~ng4098;
  assign new_n5780_ = ~ng4093 & new_n5779_;
  assign new_n5781_1_ = new_n5766_1_ & new_n5780_;
  assign new_n5782_ = ng5527 & new_n5781_1_;
  assign new_n5783_ = ng5535 & new_n5782_;
  assign new_n5784_ = ng5523 & new_n5783_;
  assign new_n5785_1_ = ng4093 & new_n5779_;
  assign new_n5786_ = new_n5766_1_ & new_n5785_1_;
  assign new_n5787_ = ng6219 & new_n5786_;
  assign new_n5788_ = ng6227 & new_n5787_;
  assign new_n5789_1_ = ng6215 & new_n5788_;
  assign new_n5790_ = ~new_n5773_ & ~new_n5778_;
  assign new_n5791_ = ~new_n5784_ & ~new_n5789_1_;
  assign new_n5792_ = new_n5790_ & new_n5791_;
  assign new_n5793_ = ~ng4087 & ng4098;
  assign new_n5794_1_ = ~ng4093 & new_n5793_;
  assign new_n5795_ = new_n5766_1_ & new_n5794_1_;
  assign new_n5796_ = ng6565 & new_n5795_;
  assign new_n5797_ = ng6573 & new_n5796_;
  assign new_n5798_ = ng6561 & new_n5797_;
  assign new_n5799_1_ = ng4093 & new_n5793_;
  assign new_n5800_ = new_n5766_1_ & new_n5799_1_;
  assign new_n5801_ = ng3522 & new_n5800_;
  assign new_n5802_ = ng3530 & new_n5801_;
  assign new_n5803_ = ng3518 & new_n5802_;
  assign new_n5804_1_ = ng4087 & ng4098;
  assign new_n5805_ = ~ng4093 & new_n5804_1_;
  assign new_n5806_ = new_n5766_1_ & new_n5805_;
  assign new_n5807_ = ng3171 & new_n5806_;
  assign new_n5808_ = ng3179 & new_n5807_;
  assign new_n5809_1_ = ng3167 & new_n5808_;
  assign new_n5810_ = ng4093 & new_n5804_1_;
  assign new_n5811_ = new_n5766_1_ & new_n5810_;
  assign new_n5812_ = ng3873 & new_n5811_;
  assign new_n5813_ = ng3881 & new_n5812_;
  assign new_n5814_1_ = ng3869 & new_n5813_;
  assign new_n5815_ = ~new_n5798_ & ~new_n5803_;
  assign new_n5816_ = ~new_n5809_1_ & ~new_n5814_1_;
  assign new_n5817_ = new_n5815_ & new_n5816_;
  assign new_n5818_ = new_n5792_ & new_n5817_;
  assign new_n5819_1_ = new_n5767_ & ~new_n5818_;
  assign pg33659 = ~new_n5767_ | new_n5819_1_;
  assign new_n5821_ = ng22 & n2287;
  assign pg34921 = ~ng22 | new_n5821_;
  assign new_n5823_ = ~ng1964 & ~ng1696;
  assign new_n5824_1_ = ~ng1830 & new_n5823_;
  assign new_n5825_ = ~ng2098 & new_n5824_1_;
  assign new_n5826_ = pg35 & ~new_n5825_;
  assign new_n5827_ = ~ng2255 & ~ng2523;
  assign new_n5828_ = ~ng2389 & new_n5827_;
  assign new_n5829_1_ = ~ng2657 & new_n5828_;
  assign new_n5830_ = pg35 & ~new_n5829_1_;
  assign new_n5831_ = ~new_n5826_ & new_n5830_;
  assign new_n5832_ = new_n5826_ & ~new_n5830_;
  assign new_n5833_ = ~new_n5831_ & ~new_n5832_;
  assign new_n5834_1_ = ~new_n5826_ & ~new_n5830_;
  assign pg26875 = ~new_n5833_ | new_n5834_1_;
  assign new_n5836_ = ~ng4785 & ~ng4709;
  assign new_n5837_ = ng4698 & new_n5836_;
  assign new_n5838_1_ = ~ng4785 & ng4709;
  assign new_n5839_ = ng4754 & new_n5838_1_;
  assign new_n5840_ = ng4785 & ~ng4709;
  assign new_n5841_ = ng4743 & new_n5840_;
  assign new_n5842_ = ng4765 & new_n5665_;
  assign new_n5843_1_ = ~new_n5837_ & ~new_n5839_;
  assign new_n5844_ = ~new_n5841_ & ~new_n5842_;
  assign new_n5845_ = new_n5843_1_ & new_n5844_;
  assign new_n5846_ = new_n5701_ & ~new_n5845_;
  assign pg33636 = ~new_n5701_ | new_n5846_;
  assign new_n5848_1_ = ~pg35 & ng6209;
  assign new_n5849_ = ng6209 & ng6203;
  assign new_n5850_ = ~pg113 & new_n5786_;
  assign new_n5851_ = ~new_n4724_ & new_n5850_;
  assign new_n5852_ = ng43 & new_n5851_;
  assign new_n5853_1_ = ~ng6215 & ~new_n5852_;
  assign new_n5854_ = new_n5849_ & new_n5853_1_;
  assign new_n5855_ = ng6215 & new_n5853_1_;
  assign new_n5856_ = ~new_n5849_ & new_n5855_;
  assign new_n5857_ = ~new_n5854_ & ~new_n5856_;
  assign new_n5858_1_ = pg35 & ~new_n5857_;
  assign n688 = new_n5848_1_ | new_n5858_1_;
  assign new_n5860_ = ~pg35 & ng4322;
  assign new_n5861_ = ~ng4639 & ng4621;
  assign new_n5862_ = ng4628 & new_n5861_;
  assign new_n5863_1_ = ng4340 & ng4349;
  assign new_n5864_ = ng4358 & new_n5863_1_;
  assign new_n5865_ = new_n5862_ & new_n5864_;
  assign new_n5866_ = ng4311 & new_n5865_;
  assign new_n5867_ = ng4322 & new_n5866_;
  assign new_n5868_1_ = ng4322 & new_n5865_;
  assign new_n5869_ = ng4332 & new_n5868_1_;
  assign new_n5870_ = ~pg113 & ~new_n4724_;
  assign new_n5871_ = ~pg73 & ~pg72;
  assign new_n5872_ = ~new_n5870_ & new_n5871_;
  assign new_n5873_1_ = ng65 & ~new_n5872_;
  assign new_n5874_ = ~new_n5869_ & ~new_n5873_1_;
  assign new_n5875_ = ~ng4332 & new_n5874_;
  assign new_n5876_ = new_n5867_ & new_n5875_;
  assign new_n5877_ = ng4332 & new_n5874_;
  assign new_n5878_1_ = ~new_n5867_ & new_n5877_;
  assign new_n5879_ = ~new_n5876_ & ~new_n5878_1_;
  assign new_n5880_ = pg35 & ~new_n5879_;
  assign n693 = new_n5860_ | new_n5880_;
  assign new_n5882_ = pg35 & ng2711;
  assign new_n5883_1_ = ~pg35 & new_n5882_;
  assign new_n5884_ = pg125 & pg35;
  assign n698 = new_n5883_1_ | new_n5884_;
  assign new_n5886_ = ~pg35 & ng1094;
  assign new_n5887_ = ng1116 & new_n4699_;
  assign new_n5888_1_ = ~ng1152 & ng1099;
  assign new_n5889_ = new_n5887_ & new_n5888_1_;
  assign new_n5890_ = ng1135 & ng1094;
  assign new_n5891_ = ng1135 & ~new_n5890_;
  assign new_n5892_ = ng1094 & ~new_n5890_;
  assign new_n5893_1_ = ~new_n5891_ & ~new_n5892_;
  assign new_n5894_ = new_n5889_ & ~new_n5893_1_;
  assign new_n5895_ = ng1135 & ~new_n5889_;
  assign new_n5896_ = ~new_n5894_ & ~new_n5895_;
  assign new_n5897_ = pg35 & ~new_n5896_;
  assign n703 = new_n5886_ | new_n5897_;
  assign new_n5899_ = ~pg35 & ng2491;
  assign new_n5900_ = ~ng2741 & ~ng2748;
  assign new_n5901_ = ~ng2756 & new_n5900_;
  assign new_n5902_1_ = ng2735 & new_n5901_;
  assign new_n5903_ = ~ng2815 & new_n5902_1_;
  assign new_n5904_ = ~ng2724 & ~ng2729;
  assign new_n5905_ = ~new_n5903_ & new_n5904_;
  assign new_n5906_ = ~ng2715 & ~new_n5905_;
  assign new_n5907_1_ = ng2719 & new_n5906_;
  assign new_n5908_ = ~pg113 & new_n5190_;
  assign new_n5909_ = ng110 & ~new_n4724_;
  assign new_n5910_ = new_n5908_ & new_n5909_;
  assign new_n5911_ = ~ng2476 & ~new_n5910_;
  assign new_n5912_1_ = new_n5907_1_ & ~new_n5911_;
  assign new_n5913_ = ng2485 & ~new_n5907_1_;
  assign new_n5914_ = ~new_n5912_1_ & ~new_n5913_;
  assign new_n5915_ = pg35 & ~new_n5914_;
  assign n708 = new_n5899_ | new_n5915_;
  assign new_n5917_1_ = ~pg35 & ng4427;
  assign new_n5918_ = pg35 & ng4423;
  assign n713 = new_n5917_1_ | new_n5918_;
  assign new_n5920_ = pg35 & ng1;
  assign new_n5921_1_ = ~pg35 & new_n5920_;
  assign new_n5922_ = ng4304 & ng4308;
  assign new_n5923_ = ng4304 & ~new_n5922_;
  assign new_n5924_ = ng4308 & ~new_n5922_;
  assign new_n5925_1_ = ~new_n5923_ & ~new_n5924_;
  assign new_n5926_ = ~ng4304 & ~new_n5925_1_;
  assign new_n5927_ = ~new_n5925_1_ & ~new_n5926_;
  assign new_n5928_ = ~ng4304 & ~new_n5926_;
  assign new_n5929_ = ~new_n5927_ & ~new_n5928_;
  assign new_n5930_1_ = pg35 & ~new_n5929_;
  assign n718 = new_n5921_1_ | new_n5930_1_;
  assign new_n5932_ = pg35 & ng979;
  assign new_n5933_ = ~pg35 & new_n5932_;
  assign new_n5934_ = ng1178 & ng996;
  assign new_n5935_1_ = ~ng1189 & new_n5934_;
  assign new_n5936_ = ng979 & ng996;
  assign new_n5937_ = ng979 & ~new_n5936_;
  assign new_n5938_ = ng996 & ~new_n5936_;
  assign new_n5939_ = ~new_n5937_ & ~new_n5938_;
  assign new_n5940_1_ = ~ng990 & ~ng979;
  assign new_n5941_ = ng1036 & ng1024;
  assign new_n5942_ = ng1002 & new_n5941_;
  assign new_n5943_ = new_n5939_ & ~new_n5940_1_;
  assign new_n5944_ = new_n5942_ & new_n5943_;
  assign new_n5945_1_ = ~ng1008 & ~new_n5944_;
  assign new_n5946_ = ~ng969 & new_n5945_1_;
  assign new_n5947_ = ng1157 & new_n5935_1_;
  assign new_n5948_ = ~new_n5946_ & new_n5947_;
  assign new_n5949_ = ~ng1193 & new_n5948_;
  assign new_n5950_1_ = ~ng1171 & ng1183;
  assign new_n5951_ = new_n5948_ & new_n5950_1_;
  assign new_n5952_ = ng1193 & new_n5951_;
  assign new_n5953_ = ~new_n5949_ & ~new_n5952_;
  assign new_n5954_ = ng1171 & new_n5953_;
  assign new_n5955_1_ = ng1157 & ~new_n5954_;
  assign new_n5956_ = ~ng1171 & new_n5953_;
  assign new_n5957_ = ~ng1157 & ~new_n5956_;
  assign new_n5958_ = ~new_n5955_1_ & ~new_n5957_;
  assign new_n5959_ = pg35 & ~new_n5958_;
  assign n723 = new_n5933_ | new_n5959_;
  assign new_n5961_ = ~pg35 & ng3219;
  assign new_n5962_ = ng3171 & ~ng3179;
  assign new_n5963_ = ng3161 & ~ng3155;
  assign new_n5964_ = new_n5962_ & new_n5963_;
  assign new_n5965_1_ = ng3235 & ~new_n5964_;
  assign new_n5966_ = ~ng4284 & ng4180;
  assign new_n5967_ = new_n5964_ & ~new_n5966_;
  assign new_n5968_ = ~new_n5965_1_ & ~new_n5967_;
  assign new_n5969_1_ = pg35 & ~new_n5968_;
  assign n728 = new_n5961_ | new_n5969_1_;
  assign new_n5971_ = ~pg35 & ng2844;
  assign new_n5972_ = ng12 & new_n4927_;
  assign new_n5973_ = n3583 & new_n5972_;
  assign new_n5974_1_ = ng2852 & ~new_n5972_;
  assign new_n5975_ = ~new_n5973_ & ~new_n5974_1_;
  assign new_n5976_ = pg35 & ~new_n5975_;
  assign n733 = new_n5971_ | new_n5976_;
  assign new_n5978_ = ~pg35 & ng4132;
  assign new_n5979_1_ = ~ng4064 & ng4057;
  assign new_n5980_ = ~ng4076 & new_n4708_;
  assign new_n5981_ = new_n4706_1_ & new_n5979_1_;
  assign new_n5982_ = new_n5980_ & new_n5981_;
  assign new_n5983_1_ = ng4135 & ~new_n5982_;
  assign new_n5984_ = ng4164 & new_n5982_;
  assign new_n5985_ = ~new_n5983_1_ & ~new_n5984_;
  assign new_n5986_ = pg35 & ~new_n5985_;
  assign n738 = new_n5978_ | new_n5986_;
  assign new_n5988_1_ = ~pg35 & ng301;
  assign new_n5989_ = ~ng499 & ~ng518;
  assign new_n5990_ = ~ng482 & ~ng528;
  assign new_n5991_ = ~ng490 & new_n5990_;
  assign new_n5992_ = ng385 & ~ng370;
  assign new_n5993_1_ = ng358 & ng376;
  assign new_n5994_ = new_n5992_ & new_n5993_1_;
  assign new_n5995_ = new_n5989_ & new_n5991_;
  assign new_n5996_ = new_n5994_ & new_n5995_;
  assign new_n5997_ = ~ng718 & ~ng753;
  assign new_n5998_1_ = ~ng655 & new_n5997_;
  assign new_n5999_ = ng718 & ng753;
  assign new_n6000_ = ng655 & new_n5999_;
  assign new_n6001_ = ng554 & ng807;
  assign new_n6002_ = new_n5996_ & ~new_n5998_1_;
  assign new_n6003_1_ = ~new_n6000_ & new_n6002_;
  assign new_n6004_ = ~new_n6001_ & new_n6003_1_;
  assign new_n6005_ = ~ng262 & ~ng255;
  assign new_n6006_ = ng232 & new_n6005_;
  assign new_n6007_ = ng225 & new_n6006_;
  assign new_n6008_1_ = ~ng269 & new_n6007_;
  assign new_n6009_ = ng246 & new_n6008_1_;
  assign new_n6010_ = ng239 & new_n6009_;
  assign new_n6011_ = ng278 & new_n6010_;
  assign new_n6012_ = ng262 & ng255;
  assign new_n6013_1_ = ~ng232 & new_n6012_;
  assign new_n6014_ = ~ng225 & new_n6013_1_;
  assign new_n6015_ = ng269 & new_n6014_;
  assign new_n6016_ = ~ng246 & new_n6015_;
  assign new_n6017_ = ~ng239 & new_n6016_;
  assign new_n6018_1_ = ~ng278 & new_n6017_;
  assign new_n6019_ = ~new_n6011_ & ~new_n6018_1_;
  assign new_n6020_ = ~new_n6004_ & ~new_n6019_;
  assign new_n6021_ = ng691 & new_n6020_;
  assign new_n6022_ = ng283 & new_n6021_;
  assign new_n6023_1_ = new_n6021_ & new_n6022_;
  assign new_n6024_ = ng287 & new_n6023_1_;
  assign new_n6025_ = new_n6021_ & new_n6024_;
  assign new_n6026_ = ng291 & new_n6025_;
  assign new_n6027_ = new_n6021_ & new_n6026_;
  assign new_n6028_1_ = ng294 & new_n6027_;
  assign new_n6029_ = new_n6021_ & new_n6028_1_;
  assign new_n6030_ = ng298 & new_n6029_;
  assign new_n6031_ = ng142 & new_n6030_;
  assign new_n6032_ = pg35 & new_n6031_;
  assign n743 = new_n5988_1_ | new_n6032_;
  assign new_n6034_ = pg35 & ng391;
  assign new_n6035_ = ~pg35 & new_n6034_;
  assign new_n6036_ = ~ng365 & ~ng358;
  assign new_n6037_1_ = pg35 & new_n6036_;
  assign n748 = new_n6035_ | new_n6037_1_;
  assign new_n6039_ = ~pg35 & ng2819;
  assign new_n6040_ = ng2735 & ng2748;
  assign new_n6041_1_ = new_n5191_1_ & new_n6040_;
  assign new_n6042_ = ~ng2724 & ng2729;
  assign new_n6043_ = new_n6041_1_ & new_n6042_;
  assign new_n6044_ = ng2815 & ~new_n6043_;
  assign new_n6045_1_ = ng111 & new_n5870_;
  assign new_n6046_ = ng2823 & ~new_n5870_;
  assign new_n6047_ = ~new_n6045_1_ & ~new_n6046_;
  assign new_n6048_ = new_n6043_ & new_n6047_;
  assign new_n6049_ = ~new_n6044_ & ~new_n6048_;
  assign new_n6050_1_ = pg35 & ~new_n6049_;
  assign n753 = new_n6039_ | new_n6050_1_;
  assign new_n6052_ = ~pg35 & ng4894;
  assign new_n6053_ = new_n5674_ & new_n5676_;
  assign new_n6054_ = ~ng5008 & ~ng4999;
  assign new_n6055_1_ = ~new_n4724_ & new_n6054_;
  assign new_n6056_ = ~new_n6053_ & ~new_n6055_1_;
  assign new_n6057_ = ng4894 & ~new_n6055_1_;
  assign new_n6058_ = ng71 & new_n6055_1_;
  assign new_n6059_ = ~new_n6057_ & ~new_n6058_;
  assign new_n6060_1_ = ~new_n6056_ & ~new_n6059_;
  assign new_n6061_ = ng4888 & new_n6056_;
  assign new_n6062_ = ~new_n6060_1_ & ~new_n6061_;
  assign new_n6063_ = pg35 & ~new_n6062_;
  assign n758 = new_n6052_ | new_n6063_;
  assign new_n6065_1_ = ~pg35 & ng437;
  assign new_n6066_ = ng385 & ng370;
  assign new_n6067_ = new_n5993_1_ & new_n6066_;
  assign new_n6068_ = ng433 & ~new_n6067_;
  assign new_n6069_1_ = ng269 & new_n6067_;
  assign new_n6070_ = ~new_n6068_ & ~new_n6069_1_;
  assign new_n6071_ = pg35 & ~new_n6070_;
  assign n763 = new_n6065_1_ | new_n6071_;
  assign new_n6073_ = ~pg35 & ng3731;
  assign new_n6074_1_ = ng3712 & ~ng3706;
  assign new_n6075_ = ~ng3719 & new_n6074_1_;
  assign new_n6076_ = ~ng3723 & new_n6075_;
  assign new_n6077_ = ~ng3727 & new_n6076_;
  assign new_n6078_ = ~ng3731 & new_n6077_;
  assign new_n6079_1_ = ng3752 & ng3706;
  assign new_n6080_ = ng3719 & new_n6079_1_;
  assign new_n6081_ = ng3723 & new_n6080_;
  assign new_n6082_ = ng3727 & new_n6081_;
  assign new_n6083_ = ng3731 & new_n6082_;
  assign new_n6084_1_ = ~new_n6078_ & ~new_n6083_;
  assign new_n6085_ = ~ng3736 & ~new_n6084_1_;
  assign new_n6086_ = ~ng3736 & ng3747;
  assign new_n6087_ = ~ng3731 & new_n6086_;
  assign new_n6088_1_ = pg84 & new_n6087_;
  assign new_n6089_ = ng3712 & new_n6088_1_;
  assign new_n6090_ = ng3736 & ~ng3747;
  assign new_n6091_ = ng3731 & new_n6090_;
  assign new_n6092_1_ = pg84 & new_n6091_;
  assign new_n6093_ = ng3752 & new_n6092_1_;
  assign new_n6094_ = ng3747 & ~ng3742;
  assign new_n6095_ = ~ng3736 & new_n6094_;
  assign new_n6096_1_ = ~pg84 & new_n6095_;
  assign new_n6097_ = ng3712 & new_n6096_1_;
  assign new_n6098_ = ~ng3747 & ng3742;
  assign new_n6099_ = ng3736 & new_n6098_;
  assign new_n6100_ = ~pg84 & new_n6099_;
  assign new_n6101_1_ = ng3752 & new_n6100_;
  assign new_n6102_ = ~new_n6089_ & ~new_n6093_;
  assign new_n6103_ = ~new_n6097_ & ~new_n6101_1_;
  assign new_n6104_ = new_n6102_ & new_n6103_;
  assign new_n6105_1_ = ng3736 & new_n6104_;
  assign new_n6106_ = new_n6084_1_ & new_n6105_1_;
  assign new_n6107_ = ~new_n6085_ & ~new_n6106_;
  assign new_n6108_ = pg35 & ~new_n6107_;
  assign n768 = new_n6073_ | new_n6108_;
  assign new_n6110_ = ~pg35 & ng269;
  assign new_n6111_ = ~ng862 & ng890;
  assign new_n6112_ = ~ng896 & new_n6111_;
  assign new_n6113_ = ng887 & new_n6112_;
  assign new_n6114_1_ = ng246 & ~new_n6112_;
  assign new_n6115_ = ~new_n6113_ & ~new_n6114_1_;
  assign new_n6116_ = pg35 & ~new_n6115_;
  assign n773 = new_n6110_ | new_n6116_;
  assign new_n6118_ = ~pg35 & ng479;
  assign new_n6119_1_ = pg72 & ng225;
  assign new_n6120_ = ~pg72 & ng232;
  assign new_n6121_ = ~new_n6119_1_ & ~new_n6120_;
  assign new_n6122_ = pg73 & new_n6121_;
  assign new_n6123_ = pg72 & ng239;
  assign new_n6124_1_ = ~pg72 & ng246;
  assign new_n6125_ = ~new_n6123_ & ~new_n6124_1_;
  assign new_n6126_ = ~pg73 & new_n6125_;
  assign new_n6127_ = ~new_n6122_ & ~new_n6126_;
  assign new_n6128_ = pg35 & new_n6127_;
  assign n778 = new_n6118_ | new_n6128_;
  assign new_n6130_ = ~pg35 & ng1024;
  assign new_n6131_ = ~ng1008 & ~new_n5939_;
  assign new_n6132_ = ng1030 & ng1018;
  assign new_n6133_ = new_n5939_ & new_n6132_;
  assign new_n6134_1_ = ng1008 & new_n6133_;
  assign new_n6135_ = ng1046 & ~new_n5939_;
  assign new_n6136_ = ~new_n6131_ & ~new_n6134_1_;
  assign new_n6137_ = ~ng969 & ~new_n6135_;
  assign new_n6138_ = new_n6136_ & new_n6137_;
  assign new_n6139_1_ = ~ng1002 & new_n6138_;
  assign new_n6140_ = ~new_n5940_1_ & ~new_n6139_1_;
  assign new_n6141_ = ~ng1018 & new_n6138_;
  assign new_n6142_ = new_n6140_ & ~new_n6141_;
  assign new_n6143_ = ~ng1024 & new_n6138_;
  assign new_n6144_1_ = new_n6142_ & ~new_n6143_;
  assign new_n6145_ = ng1030 & ~new_n6144_1_;
  assign new_n6146_ = ~ng1030 & new_n6138_;
  assign new_n6147_ = new_n6144_1_ & new_n6146_;
  assign new_n6148_ = ~new_n6145_ & ~new_n6147_;
  assign new_n6149_1_ = pg35 & ~new_n6148_;
  assign n783 = new_n6130_ | new_n6149_1_;
  assign new_n6151_ = ~new_n5201_1_ & pg34201;
  assign new_n6152_ = new_n5201_1_ & ~new_n5224_;
  assign n788 = new_n6151_ | new_n6152_;
  assign new_n6154_1_ = ~pg35 & ng4793;
  assign new_n6155_ = ng4793 & new_n5670_;
  assign new_n6156_ = ng4793 & ng4776;
  assign new_n6157_ = new_n5670_ & new_n6156_;
  assign new_n6158_ = ~pg113 & ng63;
  assign new_n6159_1_ = ~new_n4724_ & new_n4734_;
  assign new_n6160_ = new_n6158_ & new_n6159_1_;
  assign new_n6161_ = ~new_n6157_ & ~new_n6160_;
  assign new_n6162_ = ng4801 & new_n6161_;
  assign new_n6163_ = ~new_n6155_ & new_n6162_;
  assign new_n6164_1_ = ~ng4801 & new_n6161_;
  assign new_n6165_ = new_n6155_ & new_n6164_1_;
  assign new_n6166_ = ~new_n6163_ & ~new_n6165_;
  assign new_n6167_ = pg35 & ~new_n6166_;
  assign n798 = new_n6154_1_ | new_n6167_;
  assign new_n6169_1_ = ~pg35 & ng4040;
  assign new_n6170_ = ng4012 & ng4005;
  assign new_n6171_ = ng3983 & ng3969;
  assign new_n6172_ = new_n6170_ & new_n6171_;
  assign new_n6173_ = ng4040 & new_n6172_;
  assign new_n6174_1_ = ~ng4049 & ~new_n6173_;
  assign new_n6175_ = pg35 & new_n6174_1_;
  assign n803 = new_n6169_1_ | new_n6175_;
  assign new_n6177_ = ~pg35 & ng4165;
  assign new_n6178_ = pg35 & ng4165;
  assign n808 = new_n6177_ | new_n6178_;
  assign new_n6180_ = ~pg35 & ng2138;
  assign new_n6181_ = ng12 & new_n5061_;
  assign new_n6182_ = n2272 & new_n6181_;
  assign new_n6183_ = ng2145 & ~new_n6181_;
  assign new_n6184_1_ = ~new_n6182_ & ~new_n6183_;
  assign new_n6185_ = pg35 & ~new_n6184_1_;
  assign n813 = new_n6180_ | new_n6185_;
  assign new_n6187_ = ~pg35 & ng5134;
  assign new_n6188_1_ = ng5357 & ng5343;
  assign new_n6189_ = ng5283 & new_n6188_1_;
  assign new_n6190_ = ng5297 & new_n6189_;
  assign new_n6191_ = pg33959 & new_n6190_;
  assign new_n6192_1_ = ng5138 & ~new_n6191_;
  assign new_n6193_ = ng5128 & ~ng5134;
  assign new_n6194_ = ng5128 & ~new_n6193_;
  assign new_n6195_ = ~ng5134 & ~new_n6193_;
  assign new_n6196_ = ~new_n6194_ & ~new_n6195_;
  assign new_n6197_1_ = new_n6191_ & ~new_n6196_;
  assign new_n6198_ = ~new_n6192_1_ & ~new_n6197_1_;
  assign new_n6199_ = pg35 & ~new_n6198_;
  assign n818 = new_n6187_ | new_n6199_;
  assign new_n6201_ = ~pg35 & ng3869;
  assign new_n6202_1_ = ~pg113 & new_n5811_;
  assign new_n6203_ = ~new_n4724_ & new_n6202_1_;
  assign new_n6204_ = ng43 & new_n6203_;
  assign new_n6205_ = ng3873 & ~new_n6204_;
  assign new_n6206_ = ~ng3869 & new_n6205_;
  assign new_n6207_1_ = ~ng3873 & ~new_n6204_;
  assign new_n6208_ = ng3869 & new_n6207_1_;
  assign new_n6209_ = ~new_n6206_ & ~new_n6208_;
  assign new_n6210_ = pg35 & ~new_n6209_;
  assign n823 = new_n6201_ | new_n6210_;
  assign new_n6212_1_ = ~pg35 & ng3802;
  assign new_n6213_ = ~ng3802 & ng3794;
  assign new_n6214_ = ~ng3752 & ~new_n6213_;
  assign new_n6215_ = ~ng3798 & ~new_n6214_;
  assign new_n6216_1_ = pg35 & new_n6215_;
  assign n828 = new_n6212_1_ | new_n6216_1_;
  assign new_n6218_ = ~pg35 & ng550;
  assign new_n6219_ = ng12 & new_n4910_;
  assign new_n6220_1_ = n5005 & new_n6219_;
  assign new_n6221_ = ng136 & ~new_n6219_;
  assign new_n6222_ = ~new_n6220_1_ & ~new_n6221_;
  assign new_n6223_ = pg35 & ~new_n6222_;
  assign n833 = new_n6218_ | new_n6223_;
  assign new_n6225_1_ = ~pg35 & ng1779;
  assign new_n6226_ = ~ng2138 & ng2130;
  assign new_n6227_ = ng2145 & new_n6226_;
  assign new_n6228_ = ~ng209 & ng691;
  assign new_n6229_ = new_n4686_ & new_n6228_;
  assign new_n6230_1_ = ~pg134 & ~new_n6229_;
  assign new_n6231_ = ~new_n5358_1_ & ~new_n6230_1_;
  assign new_n6232_ = ~new_n6227_ & new_n6231_;
  assign new_n6233_ = ng979 & new_n5950_1_;
  assign new_n6234_ = new_n4700_ & new_n6233_;
  assign new_n6235_1_ = ng1079 & ~new_n6234_;
  assign new_n6236_ = new_n6232_ & ~new_n6235_1_;
  assign new_n6237_ = ~new_n4724_ & new_n5644_;
  assign new_n6238_ = ~pg113 & new_n6237_;
  assign new_n6239_ = ng112 & new_n6238_;
  assign new_n6240_1_ = ng1728 & ~new_n6239_;
  assign new_n6241_ = ~new_n6236_ & new_n6240_1_;
  assign new_n6242_ = ng1772 & new_n6236_;
  assign new_n6243_ = ~new_n6241_ & ~new_n6242_;
  assign new_n6244_ = pg35 & ~new_n6243_;
  assign n838 = new_n6225_1_ | new_n6244_;
  assign new_n6246_ = ~pg35 & ng3167;
  assign new_n6247_ = ~pg113 & new_n5806_;
  assign new_n6248_ = ~new_n4724_ & new_n6247_;
  assign new_n6249_ = ng43 & new_n6248_;
  assign new_n6250_1_ = ng3171 & ~new_n6249_;
  assign new_n6251_ = ~ng3167 & new_n6250_1_;
  assign new_n6252_ = ~ng3171 & ~new_n6249_;
  assign new_n6253_ = ng3167 & new_n6252_;
  assign new_n6254_ = ~new_n6251_ & ~new_n6253_;
  assign new_n6255_1_ = pg35 & ~new_n6254_;
  assign n848 = new_n6246_ | new_n6255_1_;
  assign new_n6257_ = ~pg35 & ng174;
  assign new_n6258_ = ng168 & ~new_n5994_;
  assign new_n6259_ = ng174 & new_n5994_;
  assign new_n6260_1_ = ~new_n6258_ & ~new_n6259_;
  assign new_n6261_ = pg35 & ~new_n6260_1_;
  assign n853 = new_n6257_ | new_n6261_;
  assign new_n6263_ = ~pg35 & ng475;
  assign new_n6264_ = ng441 & ~new_n6067_;
  assign new_n6265_1_ = ng475 & new_n6067_;
  assign new_n6266_ = ~new_n6264_ & ~new_n6265_1_;
  assign new_n6267_ = pg35 & ~new_n6266_;
  assign n858 = new_n6263_ | new_n6267_;
  assign new_n6269_ = ~pg35 & ng157;
  assign new_n6270_1_ = ~ng513 & ng518;
  assign new_n6271_ = ng203 & new_n6270_1_;
  assign new_n6272_ = ~ng182 & ~ng174;
  assign new_n6273_ = ~ng168 & new_n6272_;
  assign new_n6274_ = new_n6271_ & ~new_n6273_;
  assign new_n6275_1_ = ng691 & ~new_n6004_;
  assign new_n6276_ = ~new_n6274_ & new_n6275_1_;
  assign new_n6277_ = new_n6271_ & new_n6276_;
  assign new_n6278_ = ng146 & new_n6277_;
  assign new_n6279_ = new_n6276_ & new_n6278_;
  assign new_n6280_1_ = ng164 & new_n6279_;
  assign new_n6281_ = new_n6276_ & new_n6280_1_;
  assign new_n6282_ = ng150 & new_n6281_;
  assign new_n6283_ = new_n6276_ & new_n6282_;
  assign new_n6284_ = ng153 & new_n6283_;
  assign new_n6285_1_ = new_n6276_ & new_n6284_;
  assign new_n6286_ = ng157 & new_n6285_1_;
  assign new_n6287_ = ~ng160 & new_n6286_;
  assign new_n6288_ = ng160 & new_n6276_;
  assign new_n6289_ = ~new_n6286_ & new_n6288_;
  assign new_n6290_1_ = ~new_n6287_ & ~new_n6289_;
  assign new_n6291_ = pg35 & ~new_n6290_1_;
  assign n863 = new_n6269_ | new_n6291_;
  assign new_n6293_ = ~pg35 & ng1345;
  assign new_n6294_ = ~ng1322 & ~ng1333;
  assign new_n6295_1_ = ng1322 & ng1339;
  assign new_n6296_ = ng1322 & ~new_n6295_1_;
  assign new_n6297_ = ng1339 & ~new_n6295_1_;
  assign new_n6298_ = ~new_n6296_ & ~new_n6297_;
  assign new_n6299_ = ~ng1351 & ~new_n6298_;
  assign new_n6300_1_ = ng1361 & ng1373;
  assign new_n6301_ = new_n6298_ & new_n6300_1_;
  assign new_n6302_ = ng1351 & new_n6301_;
  assign new_n6303_ = ng1389 & ~new_n6298_;
  assign new_n6304_1_ = ~new_n6299_ & ~new_n6302_;
  assign new_n6305_ = ~ng1312 & ~new_n6303_;
  assign new_n6306_ = new_n6304_1_ & new_n6305_;
  assign new_n6307_ = ~ng1345 & new_n6306_;
  assign new_n6308_1_ = ~new_n6294_ & ~new_n6307_;
  assign new_n6309_ = ng1361 & ~new_n6308_1_;
  assign new_n6310_ = ~ng1361 & new_n6306_;
  assign new_n6311_ = new_n6308_1_ & new_n6310_;
  assign new_n6312_ = ~new_n6309_ & ~new_n6311_;
  assign new_n6313_1_ = pg35 & ~new_n6312_;
  assign n873 = new_n6293_ | new_n6313_1_;
  assign new_n6315_ = ~pg35 & ng6601;
  assign new_n6316_ = ng6573 & ng6565;
  assign new_n6317_ = ~ng6555 & ng6549;
  assign new_n6318_1_ = new_n6316_ & new_n6317_;
  assign new_n6319_ = ng6621 & ~new_n6318_1_;
  assign new_n6320_ = ~new_n5966_ & new_n6318_1_;
  assign new_n6321_ = ~new_n6319_ & ~new_n6320_;
  assign new_n6322_ = pg35 & ~new_n6321_;
  assign n878 = new_n6315_ | new_n6322_;
  assign new_n6324_ = ~pg35 & ng5685;
  assign new_n6325_ = ng5666 & ng5659;
  assign new_n6326_ = ng5637 & ng5623;
  assign new_n6327_ = new_n6325_ & new_n6326_;
  assign new_n6328_1_ = ng5689 & ~new_n6327_;
  assign new_n6329_ = ~ng5689 & new_n6327_;
  assign new_n6330_ = ~new_n6328_1_ & ~new_n6329_;
  assign new_n6331_ = pg35 & ~new_n6330_;
  assign n883 = new_n6324_ | new_n6331_;
  assign new_n6333_1_ = ~pg35 & ng6597;
  assign new_n6334_ = ng6573 & ~ng6565;
  assign new_n6335_ = ~ng6555 & ~ng6549;
  assign new_n6336_ = ~ng6561 & new_n6335_;
  assign new_n6337_ = new_n6334_ & new_n6336_;
  assign new_n6338_1_ = ng6593 & ~new_n6337_;
  assign new_n6339_ = ~new_n5966_ & new_n6337_;
  assign new_n6340_ = ~new_n6338_1_ & ~new_n6339_;
  assign new_n6341_ = pg35 & ~new_n6340_;
  assign n888 = new_n6333_1_ | new_n6341_;
  assign new_n6343_ = ng22 & pg34972;
  assign new_n6344_ = ~ng22 & n3854;
  assign n893 = new_n6343_ | new_n6344_;
  assign new_n6346_ = ~pg35 & ng5821;
  assign new_n6347_1_ = ng6035 & ng6049;
  assign new_n6348_ = ng5976 & new_n6347_1_;
  assign new_n6349_ = ng5990 & new_n6348_;
  assign new_n6350_ = ng4709 & new_n5691_;
  assign new_n6351_ = new_n5669_ & new_n6350_;
  assign new_n6352_1_ = ng4754 & new_n6351_;
  assign new_n6353_ = ng4681 & ~new_n6352_1_;
  assign new_n6354_ = new_n6349_ & new_n6353_;
  assign new_n6355_ = ng5827 & ~new_n6354_;
  assign new_n6356_ = ng5821 & new_n6354_;
  assign new_n6357_1_ = ~new_n6355_ & ~new_n6356_;
  assign new_n6358_ = pg35 & ~new_n6357_1_;
  assign n898 = new_n6346_ | new_n6358_;
  assign new_n6360_ = ~pg35 & ng355;
  assign new_n6361_ = ~ng333 & ~ng355;
  assign new_n6362_1_ = ng351 & new_n6361_;
  assign new_n6363_ = ~ng74 & ~ng351;
  assign new_n6364_ = ~new_n6362_1_ & ~new_n6363_;
  assign new_n6365_ = pg35 & new_n6364_;
  assign n908 = new_n6360_ | new_n6365_;
  assign new_n6367_1_ = ~pg35 & ng5377;
  assign new_n6368_ = ~ng5360 & ng5366;
  assign new_n6369_ = ~ng5373 & new_n6368_;
  assign new_n6370_ = ~ng5377 & new_n6369_;
  assign new_n6371_ = ng5406 & ng5360;
  assign new_n6372_1_ = ng5373 & new_n6371_;
  assign new_n6373_ = ng5377 & new_n6372_1_;
  assign new_n6374_ = ~new_n6370_ & ~new_n6373_;
  assign new_n6375_ = ~ng5381 & ~new_n6374_;
  assign new_n6376_ = ng5401 & ~ng5390;
  assign new_n6377_1_ = ~ng5385 & new_n6376_;
  assign new_n6378_ = pg84 & new_n6377_1_;
  assign new_n6379_ = ng5366 & new_n6378_;
  assign new_n6380_ = ~ng5401 & ng5390;
  assign new_n6381_ = ng5385 & new_n6380_;
  assign new_n6382_1_ = pg84 & new_n6381_;
  assign new_n6383_ = ng5406 & new_n6382_1_;
  assign new_n6384_ = ~ng5396 & ng5401;
  assign new_n6385_ = ~ng5390 & new_n6384_;
  assign new_n6386_ = ~pg84 & new_n6385_;
  assign new_n6387_1_ = ng5366 & new_n6386_;
  assign new_n6388_ = ng5396 & ~ng5401;
  assign new_n6389_ = ng5390 & new_n6388_;
  assign new_n6390_ = ~pg84 & new_n6389_;
  assign new_n6391_ = ng5406 & new_n6390_;
  assign new_n6392_1_ = ~new_n6379_ & ~new_n6383_;
  assign new_n6393_ = ~new_n6387_1_ & ~new_n6391_;
  assign new_n6394_ = new_n6392_1_ & new_n6393_;
  assign new_n6395_ = ng5381 & new_n6394_;
  assign new_n6396_ = new_n6374_ & new_n6395_;
  assign new_n6397_1_ = ~new_n6375_ & ~new_n6396_;
  assign new_n6398_ = pg35 & ~new_n6397_1_;
  assign n913 = new_n6367_1_ | new_n6398_;
  assign new_n6400_ = ~pg35 & ng5719;
  assign new_n6401_ = ng5712 & ~ng5706;
  assign new_n6402_1_ = ~ng5719 & new_n6401_;
  assign new_n6403_ = ng5752 & ng5706;
  assign new_n6404_ = ng5719 & new_n6403_;
  assign new_n6405_ = ~new_n6402_1_ & ~new_n6404_;
  assign new_n6406_ = ng5747 & ~ng5736;
  assign new_n6407_1_ = ~ng5731 & new_n6406_;
  assign new_n6408_ = pg84 & new_n6407_1_;
  assign new_n6409_ = ng5712 & new_n6408_;
  assign new_n6410_ = ~ng5747 & ng5736;
  assign new_n6411_1_ = ng5731 & new_n6410_;
  assign new_n6412_ = pg84 & new_n6411_1_;
  assign new_n6413_ = ng5752 & new_n6412_;
  assign new_n6414_ = ng5747 & ~ng5742;
  assign new_n6415_ = ~ng5736 & new_n6414_;
  assign new_n6416_1_ = ~pg84 & new_n6415_;
  assign new_n6417_ = ng5712 & new_n6416_1_;
  assign new_n6418_ = ~ng5747 & ng5742;
  assign new_n6419_ = ng5736 & new_n6418_;
  assign new_n6420_1_ = ~pg84 & new_n6419_;
  assign new_n6421_ = ng5752 & new_n6420_1_;
  assign new_n6422_ = ~new_n6409_ & ~new_n6413_;
  assign new_n6423_ = ~new_n6417_ & ~new_n6421_;
  assign new_n6424_ = new_n6422_ & new_n6423_;
  assign new_n6425_1_ = ng5723 & new_n6424_;
  assign new_n6426_ = new_n6405_ & new_n6425_1_;
  assign new_n6427_ = ~ng5723 & ~new_n6405_;
  assign new_n6428_ = ~new_n6426_ & ~new_n6427_;
  assign new_n6429_ = pg35 & ~new_n6428_;
  assign n918 = new_n6400_ | new_n6429_;
  assign new_n6431_ = ~pg35 & ng1472;
  assign new_n6432_ = ~ng1514 & ~ng1526;
  assign new_n6433_ = ng1459 & new_n6432_;
  assign new_n6434_ = ng1484 & ~new_n6433_;
  assign new_n6435_1_ = ~ng1442 & ~ng1489;
  assign new_n6436_ = ~ng1319 & new_n4689_;
  assign new_n6437_ = ng1300 & new_n6436_;
  assign new_n6438_ = ng1300 & ~new_n6437_;
  assign new_n6439_ = new_n6436_ & ~new_n6437_;
  assign new_n6440_1_ = ~new_n6438_ & ~new_n6439_;
  assign new_n6441_ = ng1484 & ~new_n6440_1_;
  assign new_n6442_ = ~new_n6435_1_ & new_n6441_;
  assign new_n6443_ = new_n6435_1_ & ~new_n6440_1_;
  assign new_n6444_ = ~new_n6442_ & ~new_n6443_;
  assign new_n6445_1_ = new_n6433_ & ~new_n6444_;
  assign new_n6446_ = ~new_n6434_ & ~new_n6445_1_;
  assign new_n6447_ = pg35 & ~new_n6446_;
  assign n933 = new_n6431_ | new_n6447_;
  assign new_n6449_ = ~pg35 & ng6040;
  assign new_n6450_1_ = ng6012 & ng6005;
  assign new_n6451_ = ng5969 & ng5983;
  assign new_n6452_ = new_n6450_1_ & new_n6451_;
  assign new_n6453_ = ng6035 & new_n6452_;
  assign new_n6454_ = ng6040 & ~new_n6453_;
  assign new_n6455_1_ = pg35 & new_n6454_;
  assign n938 = new_n6449_ | new_n6455_1_;
  assign new_n6457_ = ~pg35 & ng3808;
  assign new_n6458_ = ng4040 & ng4054;
  assign new_n6459_ = ng3976 & new_n6458_;
  assign new_n6460_1_ = ng3990 & new_n6459_;
  assign new_n6461_ = ~ng4991 & ~ng4983;
  assign new_n6462_ = ng4966 & new_n6461_;
  assign new_n6463_ = ng4975 & new_n6462_;
  assign new_n6464_ = ng4899 & new_n6463_;
  assign new_n6465_1_ = new_n5678_ & new_n6464_;
  assign new_n6466_ = ng4955 & new_n6465_1_;
  assign new_n6467_ = ng4878 & ~new_n6466_;
  assign new_n6468_ = new_n6460_1_ & new_n6467_;
  assign new_n6469_ = ng3817 & ~new_n6468_;
  assign new_n6470_1_ = ng3808 & ng3813;
  assign new_n6471_ = ng3813 & ~new_n6470_1_;
  assign new_n6472_ = ng3808 & ~new_n6470_1_;
  assign new_n6473_ = ~new_n6471_ & ~new_n6472_;
  assign new_n6474_ = new_n6468_ & ~new_n6473_;
  assign new_n6475_1_ = ~new_n6469_ & ~new_n6474_;
  assign new_n6476_ = pg35 & ~new_n6475_1_;
  assign n943 = new_n6457_ | new_n6476_;
  assign new_n6478_ = ~pg35 & ng324;
  assign new_n6479_ = ng305 & ng324;
  assign new_n6480_1_ = ~ng324 & ng311;
  assign new_n6481_ = ~new_n6479_ & ~new_n6480_1_;
  assign new_n6482_ = pg35 & ~new_n6481_;
  assign n948 = new_n6478_ | new_n6482_;
  assign new_n6484_ = ~pg35 & ng3072;
  assign new_n6485_1_ = ~ng3080 & ng3072;
  assign new_n6486_ = ng3080 & ~ng3072;
  assign new_n6487_ = ~new_n6485_1_ & ~new_n6486_;
  assign new_n6488_ = pg35 & ~new_n6487_;
  assign n958 = new_n6484_ | new_n6488_;
  assign new_n6490_ = pg35 & ng714;
  assign new_n6491_ = ~pg35 & new_n6490_;
  assign new_n6492_ = ng385 & ~ng376;
  assign new_n6493_1_ = ng358 & new_n6492_;
  assign new_n6494_ = ng667 & ~ng686;
  assign new_n6495_ = ng499 & ~ng513;
  assign new_n6496_ = ng518 & ~new_n6494_;
  assign new_n6497_ = ~new_n6495_ & new_n6496_;
  assign new_n6498_1_ = new_n6493_1_ & ~new_n6497_;
  assign new_n6499_ = ng499 & ~new_n6493_1_;
  assign new_n6500_ = ~new_n6498_1_ & ~new_n6499_;
  assign new_n6501_ = pg35 & ~new_n6500_;
  assign n963 = new_n6491_ | new_n6501_;
  assign new_n6503_1_ = pg35 & ng3639;
  assign new_n6504_ = ~pg35 & new_n6503_1_;
  assign new_n6505_ = pg35 & ng3530;
  assign n973 = new_n6504_ | new_n6505_;
  assign new_n6507_ = ~pg35 & ng2265;
  assign new_n6508_1_ = ng2689 & ~ng2697;
  assign new_n6509_ = ~ng2704 & new_n6508_1_;
  assign new_n6510_ = new_n4689_ & new_n6228_;
  assign new_n6511_ = ~pg134 & ~new_n6510_;
  assign new_n6512_ = ~new_n5383_1_ & ~new_n6511_;
  assign new_n6513_1_ = ~new_n6509_ & new_n6512_;
  assign new_n6514_ = ~ng1548 & ~ng1559;
  assign new_n6515_ = ~ng1564 & new_n6514_;
  assign new_n6516_ = ~ng1554 & new_n6515_;
  assign new_n6517_ = ng1514 & ~ng1526;
  assign new_n6518_1_ = ng1404 & new_n6516_;
  assign new_n6519_ = ng1322 & new_n6517_;
  assign new_n6520_ = new_n6518_1_ & new_n6519_;
  assign new_n6521_ = ng1418 & ~new_n6520_;
  assign new_n6522_ = new_n6513_1_ & ~new_n6521_;
  assign new_n6523_1_ = ~ng2153 & ~ng2227;
  assign new_n6524_ = ~new_n6522_ & new_n6523_1_;
  assign new_n6525_ = ng2269 & ~new_n6524_;
  assign new_n6526_ = ng2259 & ~ng2265;
  assign new_n6527_1_ = ng2259 & ~new_n6526_;
  assign new_n6528_ = ~ng2265 & ~new_n6526_;
  assign new_n6529_ = ~new_n6527_1_ & ~new_n6528_;
  assign new_n6530_ = new_n6524_ & ~new_n6529_;
  assign new_n6531_ = ~new_n6525_ & ~new_n6530_;
  assign new_n6532_1_ = pg35 & ~new_n6531_;
  assign n978 = new_n6507_ | new_n6532_1_;
  assign new_n6534_ = ~pg35 & ng2917;
  assign new_n6535_ = ng12 & n5814;
  assign new_n6536_ = new_n4937_ & new_n6535_;
  assign new_n6537_1_ = pg44 & ~ng2932;
  assign new_n6538_ = ~ng2927 & new_n6537_1_;
  assign new_n6539_ = ~new_n6536_ & ~new_n6538_;
  assign new_n6540_ = pg35 & new_n6539_;
  assign n983 = new_n6534_ | new_n6540_;
  assign new_n6542_1_ = ~pg35 & ng586;
  assign new_n6543_ = ng637 & ~ng640;
  assign new_n6544_ = ng74 & ~new_n6543_;
  assign new_n6545_ = ~ng559 & ng640;
  assign new_n6546_ = new_n6544_ & ~new_n6545_;
  assign new_n6547_1_ = ng562 & new_n6546_;
  assign new_n6548_ = ~new_n6545_ & new_n6547_1_;
  assign new_n6549_ = ng568 & new_n6548_;
  assign new_n6550_ = ~new_n6545_ & new_n6549_;
  assign new_n6551_ = ng572 & new_n6550_;
  assign new_n6552_1_ = ~new_n6545_ & new_n6551_;
  assign new_n6553_ = ng586 & new_n6552_1_;
  assign new_n6554_ = ~ng577 & new_n6553_;
  assign new_n6555_ = ng577 & ~new_n6545_;
  assign new_n6556_ = ~new_n6553_ & new_n6555_;
  assign new_n6557_1_ = ~new_n6554_ & ~new_n6556_;
  assign new_n6558_ = pg35 & ~new_n6557_1_;
  assign n988 = new_n6542_1_ | new_n6558_;
  assign new_n6560_ = ~pg35 & ng595;
  assign new_n6561_ = ~new_n6545_ & new_n6553_;
  assign new_n6562_1_ = ng577 & new_n6561_;
  assign new_n6563_ = ~new_n6545_ & new_n6562_1_;
  assign new_n6564_ = ng582 & new_n6563_;
  assign new_n6565_ = ~new_n6545_ & new_n6564_;
  assign new_n6566_1_ = ng590 & new_n6565_;
  assign new_n6567_ = ~new_n6545_ & new_n6566_1_;
  assign new_n6568_ = ng595 & new_n6567_;
  assign new_n6569_ = ~ng599 & new_n6568_;
  assign new_n6570_ = ng599 & ~new_n6545_;
  assign new_n6571_1_ = ~new_n6568_ & new_n6570_;
  assign new_n6572_ = ~new_n6569_ & ~new_n6571_1_;
  assign new_n6573_ = pg35 & ~new_n6572_;
  assign n993 = new_n6560_ | new_n6573_;
  assign new_n6575_ = ~pg35 & ng776;
  assign new_n6576_1_ = ng799 & ~ng802;
  assign new_n6577_ = new_n6004_ & ~new_n6576_1_;
  assign new_n6578_ = ~ng736 & ng802;
  assign new_n6579_ = new_n6577_ & ~new_n6578_;
  assign new_n6580_ = ng739 & new_n6579_;
  assign new_n6581_1_ = ~new_n6578_ & new_n6580_;
  assign new_n6582_ = ng744 & new_n6581_1_;
  assign new_n6583_ = ~new_n6578_ & new_n6582_;
  assign new_n6584_ = ng749 & new_n6583_;
  assign new_n6585_ = ~new_n6578_ & new_n6584_;
  assign new_n6586_1_ = ng758 & new_n6585_;
  assign new_n6587_ = ~new_n6578_ & new_n6586_1_;
  assign new_n6588_ = ng763 & new_n6587_;
  assign new_n6589_ = ~new_n6578_ & new_n6588_;
  assign new_n6590_ = ng767 & new_n6589_;
  assign new_n6591_1_ = ~new_n6578_ & new_n6590_;
  assign new_n6592_ = ng772 & new_n6591_1_;
  assign new_n6593_ = ~new_n6578_ & new_n6592_;
  assign new_n6594_ = ng776 & new_n6593_;
  assign new_n6595_ = ng781 & ~new_n6578_;
  assign new_n6596_1_ = ~new_n6594_ & new_n6595_;
  assign new_n6597_ = ~ng781 & new_n6594_;
  assign new_n6598_ = ~new_n6596_1_ & ~new_n6597_;
  assign new_n6599_ = pg35 & ~new_n6598_;
  assign n1003 = new_n6575_ | new_n6599_;
  assign new_n6601_ = ~pg35 & ng6423;
  assign new_n6602_ = ~ng6398 & ng6404;
  assign new_n6603_ = ~ng6411 & new_n6602_;
  assign new_n6604_1_ = ~ng6415 & new_n6603_;
  assign new_n6605_ = ~ng6419 & new_n6604_1_;
  assign new_n6606_ = ~ng6423 & new_n6605_;
  assign new_n6607_ = ng6398 & ng6444;
  assign new_n6608_ = ng6411 & new_n6607_;
  assign new_n6609_1_ = ng6415 & new_n6608_;
  assign new_n6610_ = ng6419 & new_n6609_1_;
  assign new_n6611_ = ng6423 & new_n6610_;
  assign new_n6612_ = ~new_n6606_ & ~new_n6611_;
  assign new_n6613_ = ~ng6428 & ~new_n6612_;
  assign new_n6614_1_ = ~ng6428 & ng6439;
  assign new_n6615_ = ~ng6423 & new_n6614_1_;
  assign new_n6616_ = pg84 & new_n6615_;
  assign new_n6617_ = ng6404 & new_n6616_;
  assign new_n6618_ = ng6428 & ~ng6439;
  assign new_n6619_1_ = ng6423 & new_n6618_;
  assign new_n6620_ = pg84 & new_n6619_1_;
  assign new_n6621_ = ng6444 & new_n6620_;
  assign new_n6622_ = ~ng6434 & ng6439;
  assign new_n6623_ = ~ng6428 & new_n6622_;
  assign new_n6624_1_ = ~pg84 & new_n6623_;
  assign new_n6625_ = ng6404 & new_n6624_1_;
  assign new_n6626_ = ng6434 & ~ng6439;
  assign new_n6627_ = ng6428 & new_n6626_;
  assign new_n6628_1_ = ~pg84 & new_n6627_;
  assign new_n6629_ = ng6444 & new_n6628_1_;
  assign new_n6630_ = ~new_n6617_ & ~new_n6621_;
  assign new_n6631_ = ~new_n6625_ & ~new_n6629_;
  assign new_n6632_1_ = new_n6630_ & new_n6631_;
  assign new_n6633_ = ng6428 & new_n6632_1_;
  assign new_n6634_ = new_n6612_ & new_n6633_;
  assign new_n6635_ = ~new_n6613_ & ~new_n6634_;
  assign new_n6636_ = pg35 & ~new_n6635_;
  assign n1008 = new_n6601_ | new_n6636_;
  assign new_n6638_ = ~pg35 & ng2756;
  assign new_n6639_ = ng2715 & ng2719;
  assign new_n6640_ = ng2724 & new_n6639_;
  assign new_n6641_ = ng2729 & new_n6640_;
  assign new_n6642_1_ = ng2735 & new_n6641_;
  assign new_n6643_ = ng2741 & new_n6642_1_;
  assign new_n6644_ = ng2748 & new_n6643_;
  assign new_n6645_ = ng2756 & new_n6644_;
  assign new_n6646_ = ng2759 & ~new_n6645_;
  assign new_n6647_1_ = ~ng2759 & new_n6645_;
  assign new_n6648_ = ~new_n6646_ & ~new_n6647_1_;
  assign new_n6649_ = ng2841 & ~new_n6648_;
  assign new_n6650_ = ng2841 & ~new_n6649_;
  assign new_n6651_ = pg35 & ~new_n6650_;
  assign n1013 = new_n6638_ | new_n6651_;
  assign new_n6653_ = ~pg35 & ng2712;
  assign new_n6654_ = ~ng2715 & ng2841;
  assign new_n6655_ = ng2841 & ~new_n6654_;
  assign new_n6656_ = pg35 & ~new_n6655_;
  assign n1018 = new_n6653_ | new_n6656_;
  assign new_n6658_ = ~pg35 & ng1874;
  assign new_n6659_ = ng2138 & ng2130;
  assign new_n6660_ = ~ng2145 & new_n6659_;
  assign new_n6661_ = ~new_n5313_ & ~new_n6230_1_;
  assign new_n6662_1_ = ~new_n6660_ & new_n6661_;
  assign new_n6663_ = ng1171 & ng1183;
  assign new_n6664_ = ng979 & new_n6663_;
  assign new_n6665_ = new_n4700_ & new_n6664_;
  assign new_n6666_ = ng1083 & ~new_n6665_;
  assign new_n6667_1_ = new_n6662_1_ & ~new_n6666_;
  assign new_n6668_ = ng1862 & ~ng1906;
  assign new_n6669_ = ~new_n6667_1_ & new_n6668_;
  assign new_n6670_ = ng1870 & ~new_n6669_;
  assign new_n6671_ = ng4180 & new_n6661_;
  assign new_n6672_1_ = ~new_n6662_1_ & ~new_n6671_;
  assign new_n6673_ = ng1242 & new_n6662_1_;
  assign new_n6674_ = ~new_n6672_1_ & ~new_n6673_;
  assign new_n6675_ = new_n6669_ & ~new_n6674_;
  assign new_n6676_ = ~new_n6670_ & ~new_n6675_;
  assign new_n6677_1_ = pg35 & ~new_n6676_;
  assign n1023 = new_n6658_ | new_n6677_1_;
  assign new_n6679_ = ~pg35 & ng1748;
  assign new_n6680_ = ~ng2775 & new_n5902_1_;
  assign new_n6681_ = new_n5904_ & ~new_n6680_;
  assign new_n6682_1_ = ng2715 & ~new_n6681_;
  assign new_n6683_ = ~ng2719 & new_n6682_1_;
  assign new_n6684_ = new_n5206_1_ & new_n6683_;
  assign new_n6685_ = ng1768 & ~new_n6684_;
  assign new_n6686_ = ng1772 & ~ng1728;
  assign new_n6687_1_ = new_n6684_ & ~new_n6686_;
  assign new_n6688_ = ~new_n6685_ & ~new_n6687_1_;
  assign new_n6689_ = pg35 & ~new_n6688_;
  assign n1028 = new_n6679_ | new_n6689_;
  assign new_n6691_1_ = ~pg35 & ng6177;
  assign new_n6692_ = ng6381 & ng6395;
  assign new_n6693_ = ng6322 & new_n6692_;
  assign new_n6694_ = ng6336 & new_n6693_;
  assign new_n6695_ = ng4785 & new_n5690_;
  assign new_n6696_1_ = ng4709 & new_n6695_;
  assign new_n6697_ = new_n5669_ & new_n6696_1_;
  assign new_n6698_ = ng4765 & new_n6697_;
  assign new_n6699_ = ng4688 & ~new_n6698_;
  assign new_n6700_ = new_n6694_ & new_n6699_;
  assign new_n6701_1_ = ng6181 & ~new_n6700_;
  assign new_n6702_ = ~ng6181 & new_n6700_;
  assign new_n6703_ = ~new_n6701_1_ & ~new_n6702_;
  assign new_n6704_ = pg35 & ~new_n6703_;
  assign n1038 = new_n6691_1_ | new_n6704_;
  assign new_n6706_1_ = ~pg35 & ng5727;
  assign new_n6707_ = ~ng5723 & new_n6402_1_;
  assign new_n6708_ = ~ng5727 & new_n6707_;
  assign new_n6709_ = ng5723 & new_n6404_;
  assign new_n6710_ = ng5727 & new_n6709_;
  assign new_n6711_1_ = ~new_n6708_ & ~new_n6710_;
  assign new_n6712_ = ng5731 & new_n6424_;
  assign new_n6713_ = new_n6711_1_ & new_n6712_;
  assign new_n6714_ = ~ng5731 & ~new_n6711_1_;
  assign new_n6715_ = ~new_n6713_ & ~new_n6714_;
  assign new_n6716_1_ = pg35 & ~new_n6715_;
  assign n1043 = new_n6706_1_ | new_n6716_1_;
  assign new_n6718_ = ~pg35 & ng2177;
  assign new_n6719_ = ng2153 & ng2227;
  assign new_n6720_ = ~new_n6522_ & new_n6719_;
  assign new_n6721_1_ = ng2173 & ~new_n6720_;
  assign new_n6722_ = ng4180 & new_n6512_;
  assign new_n6723_ = ~new_n6513_1_ & ~new_n6722_;
  assign new_n6724_ = ng1585 & new_n6513_1_;
  assign new_n6725_ = ~new_n6723_ & ~new_n6724_;
  assign new_n6726_1_ = new_n6720_ & ~new_n6725_;
  assign new_n6727_ = ~new_n6721_1_ & ~new_n6726_1_;
  assign new_n6728_ = pg35 & ~new_n6727_;
  assign n1048 = new_n6718_ | new_n6728_;
  assign new_n6730_ = ~pg35 & ng1760;
  assign new_n6731_1_ = ~pg113 & new_n5178_;
  assign new_n6732_ = new_n5909_ & new_n6731_1_;
  assign new_n6733_ = ~ng1760 & ~new_n6732_;
  assign new_n6734_ = new_n6683_ & ~new_n6733_;
  assign new_n6735_ = ng1783 & ~new_n6683_;
  assign new_n6736_1_ = ~new_n6734_ & ~new_n6735_;
  assign new_n6737_ = pg35 & ~new_n6736_1_;
  assign n1053 = new_n6730_ | new_n6737_;
  assign new_n6739_ = ~pg35 & ng6151;
  assign new_n6740_ = ~ng6151 & ng6144;
  assign new_n6741_1_ = ~ng6058 & ~new_n6740_;
  assign new_n6742_ = ~ng6140 & ~new_n6741_1_;
  assign new_n6743_ = pg35 & new_n6742_;
  assign n1058 = new_n6739_ | new_n6743_;
  assign new_n6745_ = ~pg35 & ng74;
  assign new_n6746_1_ = ng329 & new_n6481_;
  assign new_n6747_ = ~ng341 & new_n6746_1_;
  assign new_n6748_ = pg35 & new_n6747_;
  assign n1063 = new_n6745_ | new_n6748_;
  assign n1068 = ~pg35 & ng2710;
  assign new_n6751_1_ = ~pg35 & ng2807;
  assign new_n6752_ = new_n5904_ & new_n6041_1_;
  assign new_n6753_ = ng2803 & ~new_n6752_;
  assign new_n6754_ = ng2799 & ~new_n5870_;
  assign new_n6755_ = ~new_n6045_1_ & ~new_n6754_;
  assign new_n6756_1_ = new_n6752_ & new_n6755_;
  assign new_n6757_ = ~new_n6753_ & ~new_n6756_1_;
  assign new_n6758_ = pg35 & ~new_n6757_;
  assign n1073 = new_n6751_1_ | new_n6758_;
  assign new_n6760_ = ~pg35 & ng6287;
  assign new_n6761_1_ = ng6227 & ~ng6219;
  assign new_n6762_ = new_n5849_ & new_n6761_1_;
  assign new_n6763_ = ng6303 & ~new_n6762_;
  assign new_n6764_ = ~new_n5966_ & new_n6762_;
  assign new_n6765_ = ~new_n6763_ & ~new_n6764_;
  assign new_n6766_1_ = pg35 & ~new_n6765_;
  assign n1078 = new_n6760_ | new_n6766_1_;
  assign new_n6768_ = ~pg35 & ng3498;
  assign new_n6769_ = ng3530 & ng3522;
  assign new_n6770_ = ng3518 & new_n6769_;
  assign new_n6771_1_ = ng3462 & ~new_n6770_;
  assign new_n6772_ = ng3498 & new_n6770_;
  assign new_n6773_ = ~new_n6771_1_ & ~new_n6772_;
  assign new_n6774_ = pg35 & ~new_n6773_;
  assign n1083 = new_n6768_ | new_n6774_;
  assign new_n6776_1_ = ~pg35 & ng528;
  assign new_n6777_ = ~ng513 & new_n6493_1_;
  assign new_n6778_ = ng518 & new_n6777_;
  assign new_n6779_ = ng482 & ng490;
  assign new_n6780_ = ~ng528 & new_n6779_;
  assign new_n6781_1_ = ~ng528 & ~new_n6780_;
  assign new_n6782_ = new_n6778_ & ~new_n6781_1_;
  assign new_n6783_ = ng482 & ~new_n6494_;
  assign new_n6784_ = new_n6782_ & ~new_n6783_;
  assign new_n6785_ = ~ng482 & ~new_n6494_;
  assign new_n6786_1_ = ~new_n6782_ & ~new_n6785_;
  assign new_n6787_ = ~new_n6784_ & ~new_n6786_1_;
  assign new_n6788_ = pg35 & ~new_n6787_;
  assign n1088 = new_n6776_1_ | new_n6788_;
  assign new_n6790_ = ~pg35 & ng3080;
  assign new_n6791_1_ = ng3080 & ng3072;
  assign new_n6792_ = ng3085 & ~new_n6791_1_;
  assign new_n6793_ = ~ng3085 & new_n6791_1_;
  assign new_n6794_ = ~new_n6792_ & ~new_n6793_;
  assign new_n6795_ = pg35 & ~new_n6794_;
  assign n1093 = new_n6790_ | new_n6795_;
  assign new_n6797_ = ~pg35 & ng1792;
  assign new_n6798_ = ~ng1783 & ng1760;
  assign new_n6799_ = ng1752 & new_n6798_;
  assign new_n6800_ = ~ng1792 & ~ng1760;
  assign new_n6801_1_ = ng1748 & new_n6800_;
  assign new_n6802_ = ng1756 & new_n5206_1_;
  assign new_n6803_ = ~new_n6799_ & ~new_n6801_1_;
  assign new_n6804_ = ~new_n6802_ & new_n6803_;
  assign new_n6805_ = ng1783 & ~ng1760;
  assign new_n6806_1_ = ng1736 & new_n6805_;
  assign new_n6807_ = ng1792 & ng1760;
  assign new_n6808_ = ng1740 & new_n6807_;
  assign new_n6809_ = ~ng1783 & ng1792;
  assign new_n6810_1_ = ng1744 & new_n6809_;
  assign new_n6811_ = new_n6804_ & ~new_n6806_1_;
  assign new_n6812_ = ~new_n6808_ & ~new_n6810_1_;
  assign new_n6813_ = new_n6811_ & new_n6812_;
  assign new_n6814_1_ = new_n6683_ & ~new_n6813_;
  assign new_n6815_ = ng1811 & ~new_n6683_;
  assign new_n6816_ = ~new_n6814_1_ & ~new_n6815_;
  assign new_n6817_ = pg35 & ~new_n6816_;
  assign n1098 = new_n6797_ | new_n6817_;
  assign new_n6819_1_ = ~pg35 & ng2873;
  assign new_n6820_ = ng12 & n2272;
  assign new_n6821_ = new_n4954_ & new_n6820_;
  assign new_n6822_ = pg44 & ~ng2890;
  assign new_n6823_ = ~new_n6821_ & ~new_n6822_;
  assign new_n6824_1_ = pg35 & new_n6823_;
  assign n1103 = new_n6819_1_ | new_n6824_1_;
  assign new_n6826_ = ~pg35 & ng1536;
  assign new_n6827_ = ~ng1514 & ng1526;
  assign new_n6828_ = ng1521 & ng1339;
  assign new_n6829_1_ = ~ng1532 & new_n6828_;
  assign new_n6830_ = ng1500 & new_n6827_;
  assign new_n6831_ = ~new_n6829_1_ & new_n6830_;
  assign new_n6832_ = ng1367 & ng1379;
  assign new_n6833_ = ng1345 & new_n6832_;
  assign new_n6834_1_ = ~new_n6294_ & new_n6298_;
  assign new_n6835_ = new_n6833_ & new_n6834_1_;
  assign new_n6836_ = ~ng1351 & ~new_n6835_;
  assign new_n6837_ = ~ng1312 & new_n6836_;
  assign new_n6838_ = ng1500 & new_n6829_1_;
  assign new_n6839_1_ = ~new_n6837_ & new_n6838_;
  assign new_n6840_ = ~ng1536 & new_n6839_1_;
  assign new_n6841_ = new_n6827_ & new_n6839_1_;
  assign new_n6842_ = ng1536 & new_n6841_;
  assign new_n6843_ = ~new_n6840_ & ~new_n6842_;
  assign new_n6844_1_ = ~ng1542 & new_n6843_;
  assign new_n6845_ = new_n6831_ & new_n6844_1_;
  assign new_n6846_ = ng1542 & new_n6843_;
  assign new_n6847_ = ~new_n6831_ & new_n6846_;
  assign new_n6848_ = ~new_n6845_ & ~new_n6847_;
  assign new_n6849_1_ = pg35 & ~new_n6848_;
  assign n1108 = new_n6826_ | new_n6849_1_;
  assign new_n6851_ = ~pg35 & ng2165;
  assign new_n6852_ = ~ng2197 & ng2153;
  assign new_n6853_ = ~new_n6522_ & new_n6852_;
  assign new_n6854_1_ = ng2161 & ~new_n6853_;
  assign new_n6855_ = ~new_n6725_ & new_n6853_;
  assign new_n6856_ = ~new_n6854_1_ & ~new_n6855_;
  assign new_n6857_ = pg35 & ~new_n6856_;
  assign n1118 = new_n6851_ | new_n6857_;
  assign new_n6859_1_ = pg35 & ng956;
  assign new_n6860_ = ~pg35 & new_n6859_1_;
  assign new_n6861_ = ng12 & new_n4887_1_;
  assign new_n6862_ = n6079 & new_n6861_;
  assign new_n6863_1_ = ng947 & ~new_n6861_;
  assign new_n6864_ = ~new_n6862_ & ~new_n6863_1_;
  assign new_n6865_ = pg35 & ~new_n6864_;
  assign n1123 = new_n6860_ | new_n6865_;
  assign new_n6867_ = ~pg35 & ng538;
  assign new_n6868_1_ = new_n4910_ & new_n6535_;
  assign new_n6869_ = ~ng546 & ng691;
  assign new_n6870_ = ~new_n6868_1_ & ~new_n6869_;
  assign new_n6871_ = pg35 & new_n6870_;
  assign n1128 = new_n6867_ | new_n6871_;
  assign new_n6873_1_ = ~pg35 & ng3957;
  assign new_n6874_ = ~ng3873 & ng3881;
  assign new_n6875_ = ng3869 & new_n6874_;
  assign new_n6876_ = ng3913 & ~new_n6875_;
  assign new_n6877_ = ~new_n5966_ & new_n6875_;
  assign new_n6878_1_ = ~new_n6876_ & ~new_n6877_;
  assign new_n6879_ = pg35 & ~new_n6878_1_;
  assign n1133 = new_n6873_1_ | new_n6879_;
  assign new_n6881_ = ~pg35 & ng1554;
  assign new_n6882_ = pg35 & ng496;
  assign n1138 = new_n6881_ | new_n6882_;
  assign new_n6884_ = ~pg35 & ng5583;
  assign new_n6885_ = ng5535 & ng5527;
  assign new_n6886_ = ~ng5511 & ng5517;
  assign new_n6887_ = new_n6885_ & new_n6886_;
  assign new_n6888_1_ = ng5599 & ~new_n6887_;
  assign new_n6889_ = ~new_n5966_ & new_n6887_;
  assign new_n6890_ = ~new_n6888_1_ & ~new_n6889_;
  assign new_n6891_ = pg35 & ~new_n6890_;
  assign n1148 = new_n6884_ | new_n6891_;
  assign new_n6893_1_ = ~pg35 & ng3897;
  assign new_n6894_ = ng3873 & ~ng3881;
  assign new_n6895_ = ~ng3857 & ~ng3863;
  assign new_n6896_ = ~ng3869 & new_n6895_;
  assign new_n6897_ = new_n6894_ & new_n6896_;
  assign new_n6898_1_ = ng3893 & ~new_n6897_;
  assign new_n6899_ = ~new_n5966_ & new_n6897_;
  assign new_n6900_ = ~new_n6898_1_ & ~new_n6899_;
  assign new_n6901_ = pg35 & ~new_n6900_;
  assign n1153 = new_n6893_1_ | new_n6901_;
  assign new_n6903_ = ~pg35 & ng4057;
  assign new_n6904_ = ng4064 & ng4057;
  assign new_n6905_ = ng4141 & ~new_n6904_;
  assign new_n6906_ = ~ng4141 & new_n6904_;
  assign new_n6907_1_ = ~new_n6905_ & ~new_n6906_;
  assign new_n6908_ = ng4169 & ~new_n6907_1_;
  assign new_n6909_ = pg35 & new_n6908_;
  assign n1158 = new_n6903_ | new_n6909_;
  assign new_n6911_ = ~pg35 & ng3111;
  assign new_n6912_1_ = ~ng4899 & new_n6463_;
  assign new_n6913_ = new_n5678_ & new_n6912_1_;
  assign new_n6914_ = ng4933 & new_n6913_;
  assign new_n6915_ = ng4864 & ~new_n6914_;
  assign new_n6916_1_ = ng3352 & ng3338;
  assign new_n6917_ = ng3274 & new_n6916_1_;
  assign new_n6918_ = ng3288 & new_n6917_;
  assign new_n6919_ = ng3106 & ~new_n6918_;
  assign new_n6920_ = ~ng3352 & ~ng3288;
  assign new_n6921_1_ = ~ng3338 & new_n6920_;
  assign new_n6922_ = ng3239 & ng3321;
  assign new_n6923_ = new_n6921_1_ & new_n6922_;
  assign new_n6924_ = ~ng3352 & ng3288;
  assign new_n6925_ = ~ng3338 & new_n6924_;
  assign new_n6926_1_ = ng3211 & ng3329;
  assign new_n6927_ = new_n6925_ & new_n6926_1_;
  assign new_n6928_ = ng3352 & ~ng3288;
  assign new_n6929_ = ~ng3338 & new_n6928_;
  assign new_n6930_ = ng3255 & ng3325;
  assign new_n6931_1_ = new_n6929_ & new_n6930_;
  assign new_n6932_ = ~ng3338 & new_n4765_;
  assign new_n6933_ = ng3207 & ng3303;
  assign new_n6934_ = new_n6932_ & new_n6933_;
  assign new_n6935_ = ~new_n6923_ & ~new_n6927_;
  assign new_n6936_1_ = ~new_n6931_1_ & ~new_n6934_;
  assign new_n6937_ = new_n6935_ & new_n6936_1_;
  assign new_n6938_ = ng3338 & new_n6920_;
  assign new_n6939_ = ng3195 & ng3329;
  assign new_n6940_ = new_n6938_ & new_n6939_;
  assign new_n6941_1_ = ng3338 & ng3303;
  assign new_n6942_ = ng3303 & ~new_n6941_1_;
  assign new_n6943_ = ng3338 & ~new_n6941_1_;
  assign new_n6944_ = ~new_n6942_ & ~new_n6943_;
  assign new_n6945_ = new_n6924_ & new_n6944_;
  assign new_n6946_1_ = ng3219 & ng3281;
  assign new_n6947_ = new_n6945_ & new_n6946_1_;
  assign new_n6948_ = ng3338 & new_n6928_;
  assign new_n6949_ = ng3191 & ng3303;
  assign new_n6950_ = new_n6948_ & new_n6949_;
  assign new_n6951_1_ = new_n4765_ & new_n6944_;
  assign new_n6952_ = ng3235 & ng3310;
  assign new_n6953_ = new_n6951_1_ & new_n6952_;
  assign new_n6954_ = ~new_n6940_ & ~new_n6947_;
  assign new_n6955_ = ~new_n6950_ & ~new_n6953_;
  assign new_n6956_1_ = new_n6954_ & new_n6955_;
  assign new_n6957_ = ng3298 & ng3187;
  assign new_n6958_ = new_n6938_ & new_n6957_;
  assign new_n6959_ = ng3338 & new_n6924_;
  assign new_n6960_ = ng3231 & ng3321;
  assign new_n6961_1_ = new_n6959_ & new_n6960_;
  assign new_n6962_ = ng3317 & ng3215;
  assign new_n6963_ = new_n6948_ & new_n6962_;
  assign new_n6964_ = ng3338 & new_n4765_;
  assign new_n6965_ = ng3325 & ng3247;
  assign new_n6966_1_ = new_n6964_ & new_n6965_;
  assign new_n6967_ = ~new_n6958_ & ~new_n6961_1_;
  assign new_n6968_ = ~new_n6963_ & ~new_n6966_1_;
  assign new_n6969_ = new_n6967_ & new_n6968_;
  assign new_n6970_ = new_n6920_ & new_n6944_;
  assign new_n6971_1_ = ng3251 & ng3267;
  assign new_n6972_ = new_n6970_ & new_n6971_1_;
  assign new_n6973_ = ng3298 & ng3199;
  assign new_n6974_ = new_n6925_ & new_n6973_;
  assign new_n6975_ = ng3203 & ng3274;
  assign new_n6976_1_ = new_n6929_ & new_n6975_;
  assign new_n6977_ = ng3317 & ng3223;
  assign new_n6978_ = new_n6932_ & new_n6977_;
  assign new_n6979_ = ~new_n6972_ & ~new_n6974_;
  assign new_n6980_ = ~new_n6976_1_ & ~new_n6978_;
  assign new_n6981_1_ = new_n6979_ & new_n6980_;
  assign new_n6982_ = new_n6956_1_ & new_n6969_;
  assign new_n6983_ = new_n6981_1_ & new_n6982_;
  assign new_n6984_ = new_n6920_ & ~new_n6944_;
  assign new_n6985_ = ng3281 & ng3227;
  assign new_n6986_1_ = new_n6984_ & new_n6985_;
  assign new_n6987_ = new_n6924_ & ~new_n6944_;
  assign new_n6988_ = ng3259 & ng3267;
  assign new_n6989_ = new_n6987_ & new_n6988_;
  assign new_n6990_ = new_n6928_ & ~new_n6944_;
  assign new_n6991_1_ = ng3243 & ng3310;
  assign new_n6992_ = new_n6990_ & new_n6991_1_;
  assign new_n6993_ = ng3263 & ng3274;
  assign new_n6994_ = new_n6964_ & new_n6993_;
  assign new_n6995_ = ~new_n6986_1_ & ~new_n6989_;
  assign new_n6996_1_ = ~new_n6992_ & ~new_n6994_;
  assign new_n6997_ = new_n6995_ & new_n6996_1_;
  assign new_n6998_ = new_n6937_ & new_n6983_;
  assign new_n6999_ = new_n6997_ & new_n6998_;
  assign new_n7000_ = new_n6919_ & ~new_n6999_;
  assign new_n7001_1_ = new_n6919_ & ~new_n7000_;
  assign new_n7002_ = ~new_n6999_ & ~new_n7000_;
  assign new_n7003_ = ~new_n7001_1_ & ~new_n7002_;
  assign new_n7004_ = new_n6915_ & ~new_n7003_;
  assign new_n7005_ = ng3106 & ~new_n6915_;
  assign new_n7006_1_ = ~new_n7004_ & ~new_n7005_;
  assign new_n7007_ = pg35 & ~new_n7006_1_;
  assign n1163 = new_n6911_ | new_n7007_;
  assign new_n7009_ = ~pg35 & ng3835;
  assign new_n7010_ = ng3873 & ng3881;
  assign new_n7011_1_ = ng3869 & new_n7010_;
  assign new_n7012_ = ng3841 & ~new_n7011_1_;
  assign new_n7013_ = ng3835 & new_n7011_1_;
  assign new_n7014_ = ~new_n7012_ & ~new_n7013_;
  assign new_n7015_ = pg35 & ~new_n7014_;
  assign n1168 = new_n7009_ | new_n7015_;
  assign new_n7017_ = ~pg35 & ng2008;
  assign new_n7018_ = ng2145 & new_n6659_;
  assign new_n7019_1_ = ~new_n5279_ & ~new_n6230_1_;
  assign new_n7020_ = ~new_n7018_ & new_n7019_1_;
  assign new_n7021_ = ~ng1171 & ~ng1183;
  assign new_n7022_ = ng979 & new_n7021_;
  assign new_n7023_1_ = new_n4700_ & new_n7022_;
  assign new_n7024_ = ng1087 & ~new_n7023_1_;
  assign new_n7025_ = new_n7020_ & ~new_n7024_;
  assign new_n7026_ = ng1996 & ~ng2040;
  assign new_n7027_1_ = ~new_n7025_ & new_n7026_;
  assign new_n7028_ = ng2004 & ~new_n7027_1_;
  assign new_n7029_ = ng4180 & new_n7019_1_;
  assign new_n7030_ = ~new_n7020_ & ~new_n7029_;
  assign new_n7031_1_ = ~ng1242 & new_n7020_;
  assign new_n7032_ = ~new_n7030_ & ~new_n7031_1_;
  assign new_n7033_ = new_n7027_1_ & ~new_n7032_;
  assign new_n7034_ = ~new_n7028_ & ~new_n7033_;
  assign new_n7035_ = pg35 & ~new_n7034_;
  assign n1173 = new_n7017_ | new_n7035_;
  assign new_n7037_ = ~pg35 & ng3570;
  assign new_n7038_ = ~ng3530 & ng3522;
  assign new_n7039_ = ~ng3506 & ng3512;
  assign new_n7040_ = new_n7038_ & new_n7039_;
  assign new_n7041_1_ = ng3586 & ~new_n7040_;
  assign new_n7042_ = ~new_n5966_ & new_n7040_;
  assign new_n7043_ = ~new_n7041_1_ & ~new_n7042_;
  assign new_n7044_ = pg35 & ~new_n7043_;
  assign n1178 = new_n7037_ | new_n7044_;
  assign new_n7046_1_ = ~pg35 & ng4129;
  assign new_n7047_ = ng4064 & ~ng4057;
  assign new_n7048_ = new_n4706_1_ & new_n7047_;
  assign new_n7049_ = new_n5980_ & new_n7048_;
  assign new_n7050_1_ = ng4132 & ~new_n7049_;
  assign new_n7051_ = ng4164 & new_n7049_;
  assign new_n7052_ = ~new_n7050_1_ & ~new_n7051_;
  assign new_n7053_ = pg35 & ~new_n7052_;
  assign n1183 = new_n7046_1_ | new_n7053_;
  assign new_n7055_1_ = ~pg35 & ng952;
  assign new_n7056_ = n5005 & new_n6861_;
  assign new_n7057_ = ~ng939 & ~ng933;
  assign new_n7058_ = ~new_n7056_ & ~new_n7057_;
  assign new_n7059_ = pg35 & new_n7058_;
  assign n1188 = new_n7055_1_ | new_n7059_;
  assign new_n7061_ = pg35 & ng4826;
  assign new_n7062_ = ~pg35 & new_n7061_;
  assign new_n7063_ = ng6227 & ng6219;
  assign new_n7064_ = ng6215 & new_n7063_;
  assign new_n7065_1_ = ng6195 & ~new_n7064_;
  assign new_n7066_ = ~new_n5966_ & new_n7065_1_;
  assign new_n7067_ = new_n7065_1_ & ~new_n7066_;
  assign new_n7068_ = ~new_n5966_ & ~new_n7066_;
  assign new_n7069_ = ~new_n7067_ & ~new_n7068_;
  assign new_n7070_1_ = pg35 & ~new_n7069_;
  assign n1193 = new_n7062_ | new_n7070_1_;
  assign new_n7072_ = ~pg35 & ng918;
  assign new_n7073_ = ng904 & ng1227;
  assign new_n7074_ = ng921 & new_n7073_;
  assign new_n7075_1_ = ng936 & new_n7074_;
  assign new_n7076_ = ng907 & new_n7075_1_;
  assign new_n7077_ = ng911 & new_n7076_;
  assign new_n7078_ = ng914 & new_n7077_;
  assign new_n7079_ = ng918 & new_n7078_;
  assign new_n7080_1_ = ~ng925 & new_n7079_;
  assign new_n7081_ = ng925 & ng1227;
  assign new_n7082_ = ~new_n7079_ & new_n7081_;
  assign new_n7083_ = ~new_n7080_1_ & ~new_n7082_;
  assign new_n7084_ = pg35 & ~new_n7083_;
  assign n1198 = new_n7072_ | new_n7084_;
  assign new_n7086_ = ~pg35 & ng6259;
  assign new_n7087_ = ~ng6209 & ~ng6203;
  assign new_n7088_ = ~ng6215 & new_n7087_;
  assign new_n7089_1_ = new_n7063_ & new_n7088_;
  assign new_n7090_ = ng6255 & ~new_n7089_1_;
  assign new_n7091_ = ~new_n5966_ & new_n7089_1_;
  assign new_n7092_ = ~new_n7090_ & ~new_n7091_;
  assign new_n7093_1_ = pg35 & ~new_n7092_;
  assign n1203 = new_n7086_ | new_n7093_1_;
  assign new_n7095_ = ~pg35 & ng2181;
  assign new_n7096_ = ng2197 & ~ng2153;
  assign new_n7097_ = ~new_n6522_ & new_n7096_;
  assign new_n7098_1_ = ng2177 & ~new_n7097_;
  assign new_n7099_ = ~new_n6725_ & new_n7097_;
  assign new_n7100_ = ~new_n7098_1_ & ~new_n7099_;
  assign new_n7101_ = pg35 & ~new_n7100_;
  assign n1208 = new_n7095_ | new_n7101_;
  assign new_n7103_1_ = ~pg35 & ng5831;
  assign new_n7104_ = ng5835 & ~new_n6354_;
  assign new_n7105_ = ~ng5835 & new_n6354_;
  assign new_n7106_ = ~new_n7104_ & ~new_n7105_;
  assign new_n7107_ = pg35 & ~new_n7106_;
  assign n1213 = new_n7103_1_ | new_n7107_;
  assign new_n7109_ = ~pg35 & ng4540;
  assign new_n7110_ = pg73 & ~pg72;
  assign new_n7111_ = ~ng4578 & new_n7110_;
  assign new_n7112_ = ng4581 & ~new_n7111_;
  assign new_n7113_1_ = ~ng4581 & ng4540;
  assign new_n7114_ = ~new_n7112_ & ~new_n7113_1_;
  assign new_n7115_ = pg35 & ~new_n7114_;
  assign n1218 = new_n7109_ | new_n7115_;
  assign new_n7117_ = ~pg35 & ng5084;
  assign new_n7118_1_ = ~ng5092 & ng5084;
  assign new_n7119_ = ng5092 & ~ng5084;
  assign new_n7120_ = ~new_n7118_1_ & ~new_n7119_;
  assign new_n7121_ = pg35 & ~new_n7120_;
  assign n1228 = new_n7117_ | new_n7121_;
  assign new_n7123_1_ = ~pg35 & ng3917;
  assign new_n7124_ = ~ng3873 & ~ng3881;
  assign new_n7125_ = ~ng3857 & ng3863;
  assign new_n7126_ = new_n7124_ & new_n7125_;
  assign new_n7127_ = ng3933 & ~new_n7126_;
  assign new_n7128_1_ = ~new_n5966_ & new_n7126_;
  assign new_n7129_ = ~new_n7127_ & ~new_n7128_1_;
  assign new_n7130_ = pg35 & ~new_n7129_;
  assign n1233 = new_n7123_1_ | new_n7130_;
  assign new_n7132_ = ~pg35 & ng907;
  assign new_n7133_1_ = ng911 & ng1227;
  assign new_n7134_ = ~new_n7076_ & new_n7133_1_;
  assign new_n7135_ = ~ng911 & new_n7076_;
  assign new_n7136_ = ~new_n7134_ & ~new_n7135_;
  assign new_n7137_ = pg35 & ~new_n7136_;
  assign n1243 = new_n7132_ | new_n7137_;
  assign new_n7139_ = ~pg35 & ng3905;
  assign new_n7140_ = new_n6874_ & new_n6896_;
  assign new_n7141_ = ng3901 & ~new_n7140_;
  assign new_n7142_ = ~new_n5966_ & new_n7140_;
  assign new_n7143_1_ = ~new_n7141_ & ~new_n7142_;
  assign new_n7144_ = pg35 & ~new_n7143_1_;
  assign n1248 = new_n7139_ | new_n7144_;
  assign new_n7146_ = ~pg35 & ng4045;
  assign new_n7147_ = ng4045 & ~new_n6173_;
  assign new_n7148_1_ = pg35 & new_n7147_;
  assign n1263 = new_n7146_ | new_n7148_1_;
  assign new_n7150_ = ~pg35 & ng3133;
  assign new_n7151_ = ng3171 & ng3179;
  assign new_n7152_ = ng3167 & new_n7151_;
  assign new_n7153_1_ = ng3139 & ~new_n7152_;
  assign new_n7154_ = ng3133 & new_n7152_;
  assign new_n7155_ = ~new_n7153_1_ & ~new_n7154_;
  assign new_n7156_ = pg35 & ~new_n7155_;
  assign n1268 = new_n7150_ | new_n7156_;
  assign new_n7158_1_ = ~pg35 & ng6633;
  assign new_n7159_ = ng6555 & ng6549;
  assign new_n7160_ = new_n6334_ & new_n7159_;
  assign new_n7161_ = ng6649 & ~new_n7160_;
  assign new_n7162_ = ~new_n5966_ & new_n7160_;
  assign new_n7163_1_ = ~new_n7161_ & ~new_n7162_;
  assign new_n7164_ = pg35 & ~new_n7163_1_;
  assign n1278 = new_n7158_1_ | new_n7164_;
  assign new_n7166_ = ~pg35 & ng2606;
  assign new_n7167_ = ng2689 & ng2697;
  assign new_n7168_1_ = ng2704 & new_n7167_;
  assign new_n7169_ = ~new_n5266_ & ~new_n6511_;
  assign new_n7170_ = ~new_n7168_1_ & new_n7169_;
  assign new_n7171_ = ng1322 & new_n6432_;
  assign new_n7172_ = new_n6518_1_ & new_n7171_;
  assign new_n7173_1_ = ng1430 & ~new_n7172_;
  assign new_n7174_ = new_n7170_ & ~new_n7173_1_;
  assign new_n7175_ = ~new_n4724_ & new_n5655_;
  assign new_n7176_ = ~pg113 & new_n7175_;
  assign new_n7177_ = ng112 & new_n7176_;
  assign new_n7178_1_ = ng2555 & ~new_n7177_;
  assign new_n7179_ = ~new_n7174_ & new_n7178_1_;
  assign new_n7180_ = ng2599 & new_n7174_;
  assign new_n7181_ = ~new_n7179_ & ~new_n7180_;
  assign new_n7182_ = pg35 & ~new_n7181_;
  assign n1283 = new_n7166_ | new_n7182_;
  assign new_n7184_ = ~pg35 & ng4076;
  assign new_n7185_ = ng4141 & new_n6904_;
  assign new_n7186_ = ng4082 & new_n7185_;
  assign new_n7187_ = ng4076 & new_n7186_;
  assign new_n7188_1_ = ~ng4087 & new_n7187_;
  assign new_n7189_ = ng4087 & ~new_n7187_;
  assign new_n7190_ = ~new_n7188_1_ & ~new_n7189_;
  assign new_n7191_ = ng4169 & ~new_n7190_;
  assign new_n7192_ = pg35 & new_n7191_;
  assign n1288 = new_n7184_ | new_n7192_;
  assign new_n7194_ = ~pg35 & ng1448;
  assign new_n7195_ = ng1514 & ng1526;
  assign new_n7196_ = ng1459 & new_n7195_;
  assign new_n7197_ = ng1467 & ~new_n7196_;
  assign new_n7198_1_ = ng1472 & new_n6436_;
  assign new_n7199_ = ng1472 & ~new_n7198_1_;
  assign new_n7200_ = new_n6436_ & ~new_n7198_1_;
  assign new_n7201_ = ~new_n7199_ & ~new_n7200_;
  assign new_n7202_ = ng1467 & ~new_n7201_;
  assign new_n7203_1_ = ~new_n6435_1_ & new_n7202_;
  assign new_n7204_ = new_n6435_1_ & ~new_n7201_;
  assign new_n7205_ = ~new_n7203_1_ & ~new_n7204_;
  assign new_n7206_ = new_n7196_ & ~new_n7205_;
  assign new_n7207_ = ~new_n7197_ & ~new_n7206_;
  assign new_n7208_1_ = pg35 & ~new_n7207_;
  assign n1293 = new_n7194_ | new_n7208_1_;
  assign new_n7210_ = ~pg35 & ng6513;
  assign new_n7211_ = ng6741 & ng6727;
  assign new_n7212_ = ng6668 & new_n7211_;
  assign new_n7213_1_ = ng6682 & new_n7212_;
  assign new_n7214_ = ~ng4975 & new_n6462_;
  assign new_n7215_ = ~ng4899 & new_n7214_;
  assign new_n7216_ = new_n5678_ & new_n7215_;
  assign new_n7217_ = ng4888 & new_n7216_;
  assign new_n7218_1_ = ng4836 & ~new_n7217_;
  assign new_n7219_ = new_n7213_1_ & new_n7218_1_;
  assign new_n7220_ = ng6519 & ~new_n7219_;
  assign new_n7221_ = ng6513 & new_n7219_;
  assign new_n7222_1_ = ~new_n7220_ & ~new_n7221_;
  assign new_n7223_ = pg35 & ~new_n7222_1_;
  assign n1298 = new_n7210_ | new_n7223_;
  assign new_n7225_ = ~pg35 & ng1696;
  assign new_n7226_ = ng1624 & ng1657;
  assign new_n7227_1_ = ~ng2771 & new_n5902_1_;
  assign new_n7228_ = new_n5904_ & ~new_n7227_1_;
  assign new_n7229_ = ~ng2715 & ~new_n7228_;
  assign new_n7230_ = ~ng2719 & new_n7229_;
  assign new_n7231_ = new_n7226_ & new_n7230_;
  assign new_n7232_1_ = ng1700 & ~new_n7231_;
  assign new_n7233_ = ~ng1700 & new_n7231_;
  assign new_n7234_ = ~new_n7232_1_ & ~new_n7233_;
  assign new_n7235_ = pg35 & ~new_n7234_;
  assign n1303 = new_n7225_ | new_n7235_;
  assign new_n7237_1_ = ~pg35 & ng1936;
  assign new_n7238_ = ~ng1936 & ~ng1862;
  assign new_n7239_ = ng1950 & ~new_n7238_;
  assign new_n7240_ = ng1246 & new_n6662_1_;
  assign new_n7241_ = ~new_n6672_1_ & ~new_n7240_;
  assign new_n7242_1_ = new_n7239_ & ~new_n7241_;
  assign new_n7243_ = new_n7239_ & ~new_n7242_1_;
  assign new_n7244_ = ~new_n7241_ & ~new_n7242_1_;
  assign new_n7245_ = ~new_n7243_ & ~new_n7244_;
  assign new_n7246_ = ~new_n6667_1_ & ~new_n7245_;
  assign new_n7247_1_ = ng1950 & new_n6667_1_;
  assign new_n7248_ = ~new_n7246_ & ~new_n7247_1_;
  assign new_n7249_ = pg35 & ~new_n7248_;
  assign n1308 = new_n7237_1_ | new_n7249_;
  assign new_n7251_ = ng22 & pg34917;
  assign new_n7252_1_ = ~ng22 & n3583;
  assign n1318 = new_n7251_ | new_n7252_1_;
  assign new_n7254_ = ~pg35 & ng2413;
  assign new_n7255_ = ng2319 & ng2351;
  assign new_n7256_ = ~ng2807 & new_n5902_1_;
  assign new_n7257_1_ = new_n5904_ & ~new_n7256_;
  assign new_n7258_ = ng2715 & ~new_n7257_1_;
  assign new_n7259_ = ~ng2719 & new_n7258_;
  assign new_n7260_ = new_n7255_ & new_n7259_;
  assign new_n7261_ = ng2417 & ~new_n7260_;
  assign new_n7262_1_ = ng2407 & ~ng2413;
  assign new_n7263_ = ng2407 & ~new_n7262_1_;
  assign new_n7264_ = ~ng2413 & ~new_n7262_1_;
  assign new_n7265_ = ~new_n7263_ & ~new_n7264_;
  assign new_n7266_1_ = new_n7260_ & ~new_n7265_;
  assign new_n7267_ = ~new_n7261_ & ~new_n7266_1_;
  assign new_n7268_ = pg35 & ~new_n7267_;
  assign n1323 = new_n7254_ | new_n7268_;
  assign n1328 = ~pg35 & ng4737;
  assign new_n7271_1_ = ~pg35 & ng424;
  assign new_n7272_ = ng475 & ~new_n6067_;
  assign new_n7273_ = ng246 & new_n6067_;
  assign new_n7274_ = ~new_n7272_ & ~new_n7273_;
  assign new_n7275_ = pg35 & ~new_n7274_;
  assign n1333 = new_n7271_1_ | new_n7275_;
  assign new_n7277_ = ~pg35 & ng3782;
  assign new_n7278_ = ng3774 & ng3782;
  assign new_n7279_ = ng3787 & ~new_n7278_;
  assign new_n7280_1_ = ~ng3787 & new_n7278_;
  assign new_n7281_ = ~new_n7279_ & ~new_n7280_1_;
  assign new_n7282_ = pg35 & ~new_n7281_;
  assign n1338 = new_n7277_ | new_n7282_;
  assign new_n7284_1_ = ~pg35 & ng329;
  assign new_n7285_ = ng319 & ~new_n6481_;
  assign new_n7286_ = ng305 & ~new_n6481_;
  assign new_n7287_ = ng336 & new_n7286_;
  assign new_n7288_ = ~ng305 & ~ng311;
  assign new_n7289_1_ = ~ng319 & new_n7288_;
  assign new_n7290_ = ~ng329 & new_n7289_1_;
  assign new_n7291_ = ng311 & ~new_n6481_;
  assign new_n7292_ = ~ng336 & new_n7291_;
  assign new_n7293_ = ~new_n7285_ & ~new_n7287_;
  assign new_n7294_1_ = ~new_n7290_ & ~new_n7292_;
  assign new_n7295_ = new_n7293_ & new_n7294_1_;
  assign new_n7296_ = pg35 & ~new_n7295_;
  assign n1343 = new_n7284_1_ | new_n7296_;
  assign new_n7298_ = ~pg35 & ng5062;
  assign new_n7299_1_ = pg35 & ng5343;
  assign n1348 = new_n7298_ | new_n7299_1_;
  assign new_n7301_ = pg35 & ng5853;
  assign new_n7302_ = ~pg35 & new_n7301_;
  assign new_n7303_ = ~ng6322 & ng6346;
  assign new_n7304_1_ = ~ng6315 & ng6322;
  assign new_n7305_ = ng6351 & ng6358;
  assign new_n7306_ = ng6315 & ng6329;
  assign new_n7307_ = new_n7305_ & new_n7306_;
  assign new_n7308_ = ~new_n7303_ & ~new_n7304_1_;
  assign new_n7309_1_ = ~new_n7307_ & new_n7308_;
  assign new_n7310_ = ~ng6329 & ng6358;
  assign new_n7311_ = ~ng6351 & ng6329;
  assign new_n7312_ = ng6315 & ~ng6358;
  assign new_n7313_ = new_n7309_1_ & ~new_n7310_;
  assign new_n7314_1_ = ~new_n7311_ & new_n7313_;
  assign new_n7315_ = ~new_n7312_ & new_n7314_1_;
  assign new_n7316_ = pg35 & new_n7315_;
  assign n1353 = new_n7302_ | new_n7316_;
  assign new_n7318_ = ~pg35 & ng1728;
  assign new_n7319_1_ = ~pg113 & new_n5644_;
  assign new_n7320_ = ~new_n4724_ & new_n7319_1_;
  assign new_n7321_ = new_n6235_1_ & new_n7320_;
  assign new_n7322_ = ~ng1772 & ng1802;
  assign new_n7323_ = ng112 & new_n7322_;
  assign new_n7324_1_ = ng112 & ~new_n7323_;
  assign new_n7325_ = new_n7322_ & ~new_n7323_;
  assign new_n7326_ = ~new_n7324_1_ & ~new_n7325_;
  assign new_n7327_ = new_n7321_ & ~new_n7326_;
  assign new_n7328_ = ng1779 & ~new_n7321_;
  assign new_n7329_1_ = ~new_n7327_ & ~new_n7328_;
  assign new_n7330_ = pg35 & ~new_n7329_1_;
  assign n1358 = new_n7318_ | new_n7330_;
  assign new_n7332_ = ~pg35 & ng2803;
  assign new_n7333_ = ~ng2735 & new_n5901_;
  assign new_n7334_1_ = ~ng2724 & new_n7333_;
  assign new_n7335_ = ~ng2729 & new_n7334_1_;
  assign new_n7336_ = ng2715 & ~ng2819;
  assign new_n7337_ = ~ng2815 & ~ng2715;
  assign new_n7338_ = ~new_n7336_ & ~new_n7337_;
  assign new_n7339_1_ = ng2719 & new_n7338_;
  assign new_n7340_ = ng2715 & ~ng2807;
  assign new_n7341_ = ~ng2715 & ~ng2803;
  assign new_n7342_ = ~new_n7340_ & ~new_n7341_;
  assign new_n7343_ = ~ng2719 & new_n7342_;
  assign new_n7344_1_ = ~new_n7339_1_ & ~new_n7343_;
  assign new_n7345_ = new_n7335_ & new_n7344_1_;
  assign new_n7346_ = ng2715 & ng2638;
  assign new_n7347_ = ~ng2715 & ng2504;
  assign new_n7348_ = ~new_n7346_ & ~new_n7347_;
  assign new_n7349_1_ = ng2719 & new_n7348_;
  assign new_n7350_ = ng2715 & ng2370;
  assign new_n7351_ = ~ng2715 & ng2236;
  assign new_n7352_ = ~new_n7350_ & ~new_n7351_;
  assign new_n7353_ = ~ng2719 & new_n7352_;
  assign new_n7354_1_ = ~new_n7349_1_ & ~new_n7353_;
  assign new_n7355_ = ~new_n7335_ & new_n7354_1_;
  assign new_n7356_ = ~new_n7345_ & ~new_n7355_;
  assign new_n7357_ = pg35 & ~new_n7356_;
  assign n1363 = new_n7332_ | new_n7357_;
  assign new_n7359_1_ = ~pg35 & ng3466;
  assign new_n7360_ = ng3470 & ~new_n6770_;
  assign new_n7361_ = ~ng3470 & new_n6770_;
  assign new_n7362_ = ~new_n7360_ & ~new_n7361_;
  assign new_n7363_ = pg35 & ~new_n7362_;
  assign n1368 = new_n7359_1_ | new_n7363_;
  assign new_n7365_ = ~pg35 & ng5180;
  assign new_n7366_ = ng5176 & ng5180;
  assign new_n7367_ = ~pg113 & new_n5770_;
  assign new_n7368_ = ~new_n4724_ & new_n7367_;
  assign new_n7369_1_ = ng43 & new_n7368_;
  assign new_n7370_ = ~ng5188 & ~new_n7369_1_;
  assign new_n7371_ = new_n7366_ & new_n7370_;
  assign new_n7372_ = ng5188 & ~new_n7369_1_;
  assign new_n7373_ = ~new_n7366_ & new_n7372_;
  assign new_n7374_1_ = ~new_n7371_ & ~new_n7373_;
  assign new_n7375_ = pg35 & ~new_n7374_1_;
  assign n1373 = new_n7365_ | new_n7375_;
  assign new_n7377_ = ~pg35 & ng499;
  assign new_n7378_ = ~ng499 & ~new_n6494_;
  assign new_n7379_1_ = new_n6493_1_ & ~new_n7378_;
  assign new_n7380_ = ng504 & ~new_n6493_1_;
  assign new_n7381_ = ~new_n7379_1_ & ~new_n7380_;
  assign new_n7382_ = pg35 & ~new_n7381_;
  assign n1382 = new_n7377_ | new_n7382_;
  assign new_n7384_ = ~pg35 & ng3763;
  assign new_n7385_ = ng3763 & ng3759;
  assign new_n7386_ = pg35 & new_n7385_;
  assign n1387 = new_n7384_ | new_n7386_;
  assign new_n7388_1_ = pg35 & ng5011;
  assign new_n7389_ = ~pg35 & new_n7388_1_;
  assign new_n7390_ = ng6561 & new_n6316_;
  assign new_n7391_ = ng6541 & ~new_n7390_;
  assign new_n7392_1_ = ~new_n5966_ & new_n7391_;
  assign new_n7393_ = new_n7391_ & ~new_n7392_1_;
  assign new_n7394_ = ~new_n5966_ & ~new_n7392_1_;
  assign new_n7395_ = ~new_n7393_ & ~new_n7394_;
  assign new_n7396_ = pg35 & ~new_n7395_;
  assign n1392 = new_n7389_ | new_n7396_;
  assign new_n7398_ = ~pg35 & ng6203;
  assign new_n7399_ = ng6209 & ~new_n5852_;
  assign new_n7400_ = ~ng6203 & new_n7399_;
  assign new_n7401_ = ~ng6209 & ~new_n5852_;
  assign new_n7402_1_ = ng6203 & new_n7401_;
  assign new_n7403_ = ~new_n7400_ & ~new_n7402_1_;
  assign new_n7404_ = pg35 & ~new_n7403_;
  assign n1397 = new_n7398_ | new_n7404_;
  assign new_n7406_ = ~pg35 & ng996;
  assign new_n7407_1_ = ~ng990 & ~ng1239;
  assign new_n7408_ = ~ng1157 & new_n7407_1_;
  assign new_n7409_ = ~ng1116 & new_n7408_;
  assign new_n7410_ = ~ng1056 & new_n7409_;
  assign new_n7411_ = ng979 & ~ng1236;
  assign new_n7412_1_ = ~ng1236 & ~new_n7411_;
  assign new_n7413_ = ng979 & ~new_n7411_;
  assign new_n7414_ = ~new_n7412_1_ & ~new_n7413_;
  assign new_n7415_ = ~ng969 & ~new_n5940_1_;
  assign new_n7416_ = new_n6131_ & new_n7415_;
  assign new_n7417_1_ = new_n7414_ & new_n7416_;
  assign new_n7418_ = new_n7410_ & new_n7417_1_;
  assign new_n7419_ = new_n7410_ & ~new_n7418_;
  assign new_n7420_ = new_n7417_1_ & ~new_n7418_;
  assign new_n7421_ = ~new_n7419_ & ~new_n7420_;
  assign new_n7422_1_ = pg35 & ~new_n7421_;
  assign n1407 = new_n7406_ | new_n7422_1_;
  assign new_n7424_ = ~pg35 & ng3457;
  assign new_n7425_ = ng3689 & ng3703;
  assign new_n7426_1_ = ng3625 & new_n7425_;
  assign new_n7427_ = ng3639 & new_n7426_1_;
  assign new_n7428_ = ng4899 & new_n7214_;
  assign new_n7429_ = new_n5678_ & new_n7428_;
  assign new_n7430_1_ = ng4944 & new_n7429_;
  assign new_n7431_ = ng4871 & ~new_n7430_1_;
  assign new_n7432_ = new_n7427_ & new_n7431_;
  assign new_n7433_ = ng3466 & ~new_n7432_;
  assign new_n7434_ = ng3462 & ng3457;
  assign new_n7435_1_ = ng3462 & ~new_n7434_;
  assign new_n7436_ = ng3457 & ~new_n7434_;
  assign new_n7437_ = ~new_n7435_1_ & ~new_n7436_;
  assign new_n7438_ = new_n7432_ & ~new_n7437_;
  assign new_n7439_ = ~new_n7433_ & ~new_n7438_;
  assign new_n7440_1_ = pg35 & ~new_n7439_;
  assign n1412 = new_n7424_ | new_n7440_1_;
  assign new_n7442_ = ~pg35 & ng3263;
  assign new_n7443_ = new_n6915_ & ~new_n6999_;
  assign new_n7444_ = ng3333 & ~new_n6915_;
  assign new_n7445_1_ = ~new_n7443_ & ~new_n7444_;
  assign new_n7446_ = pg35 & ~new_n7445_1_;
  assign n1417 = new_n7442_ | new_n7446_;
  assign new_n7448_ = ~pg35 & ng4917;
  assign new_n7449_ = ng12 & new_n4963_;
  assign new_n7450_1_ = ng4922 & ~new_n7449_;
  assign new_n7451_ = n3583 & new_n7449_;
  assign new_n7452_ = ~new_n7450_1_ & ~new_n7451_;
  assign new_n7453_ = pg35 & ~new_n7452_;
  assign n1422 = new_n7448_ | new_n7453_;
  assign new_n7455_1_ = ~pg35 & ng6585;
  assign new_n7456_ = ~ng6573 & ng6565;
  assign new_n7457_ = new_n6317_ & new_n7456_;
  assign new_n7458_ = ng6613 & ~new_n7457_;
  assign new_n7459_ = ~new_n5966_ & new_n7457_;
  assign new_n7460_1_ = ~new_n7458_ & ~new_n7459_;
  assign new_n7461_ = pg35 & ~new_n7460_1_;
  assign n1427 = new_n7455_1_ | new_n7461_;
  assign new_n7463_ = new_n4738_ & pg34425;
  assign new_n7464_ = ~new_n4738_ & ~new_n4773_;
  assign n1432 = new_n7463_ | new_n7464_;
  assign new_n7466_ = pg35 & ng341;
  assign new_n7467_ = ~pg35 & new_n7466_;
  assign new_n7468_ = pg64 & pg35;
  assign n1437 = new_n7467_ | new_n7468_;
  assign new_n7470_1_ = ~pg35 & ng1437;
  assign new_n7471_ = ng1459 & new_n6517_;
  assign new_n7472_ = ~ng1495 & ng1442;
  assign new_n7473_ = new_n7471_ & new_n7472_;
  assign new_n7474_ = ng1478 & ng1437;
  assign new_n7475_1_ = ng1478 & ~new_n7474_;
  assign new_n7476_ = ng1437 & ~new_n7474_;
  assign new_n7477_ = ~new_n7475_1_ & ~new_n7476_;
  assign new_n7478_ = new_n7473_ & ~new_n7477_;
  assign new_n7479_ = ng1478 & ~new_n7473_;
  assign new_n7480_1_ = ~new_n7478_ & ~new_n7479_;
  assign new_n7481_ = pg35 & ~new_n7480_1_;
  assign n1447 = new_n7470_1_ | new_n7481_;
  assign new_n7483_ = ~pg35 & ng5401;
  assign new_n7484_ = ~new_n6379_ & ~new_n6387_1_;
  assign new_n7485_1_ = pg35 & new_n7484_;
  assign n1452 = new_n7483_ | new_n7485_1_;
  assign new_n7487_ = ~new_n5664_ & pg34221;
  assign new_n7488_ = new_n5664_ & ~new_n5683_;
  assign n1457 = new_n7487_ | new_n7488_;
  assign new_n7490_1_ = ~pg35 & ng2629;
  assign new_n7491_ = ~ng2555 & ~ng2629;
  assign new_n7492_ = ng2643 & ~new_n7491_;
  assign new_n7493_ = ng4180 & new_n7169_;
  assign new_n7494_ = ~new_n7170_ & ~new_n7493_;
  assign new_n7495_1_ = ~ng1589 & new_n7170_;
  assign new_n7496_ = ~new_n7494_ & ~new_n7495_1_;
  assign new_n7497_ = new_n7492_ & ~new_n7496_;
  assign new_n7498_ = new_n7492_ & ~new_n7497_;
  assign new_n7499_ = ~new_n7496_ & ~new_n7497_;
  assign new_n7500_1_ = ~new_n7498_ & ~new_n7499_;
  assign new_n7501_ = ~new_n7174_ & ~new_n7500_1_;
  assign new_n7502_ = ng2643 & new_n7174_;
  assign new_n7503_ = ~new_n7501_ & ~new_n7502_;
  assign new_n7504_ = pg35 & ~new_n7503_;
  assign n1462 = new_n7490_1_ | new_n7504_;
  assign new_n7506_ = ~pg35 & ng6058;
  assign new_n7507_ = ~ng6058 & ~ng6098;
  assign new_n7508_ = ng6052 & new_n7507_;
  assign new_n7509_1_ = ~ng6082 & ng6093;
  assign new_n7510_ = ~ng6077 & new_n7509_1_;
  assign new_n7511_ = pg84 & new_n7510_;
  assign new_n7512_ = ng6058 & new_n7511_;
  assign new_n7513_ = ng6082 & ~ng6093;
  assign new_n7514_1_ = ng6077 & new_n7513_;
  assign new_n7515_ = pg84 & new_n7514_1_;
  assign new_n7516_ = ng6098 & new_n7515_;
  assign new_n7517_ = ~ng6088 & ng6093;
  assign new_n7518_ = ~ng6082 & new_n7517_;
  assign new_n7519_1_ = ~pg84 & new_n7518_;
  assign new_n7520_ = ng6058 & new_n7519_1_;
  assign new_n7521_ = ng6088 & ~ng6093;
  assign new_n7522_ = ng6082 & new_n7521_;
  assign new_n7523_ = ~pg84 & new_n7522_;
  assign new_n7524_1_ = ng6098 & new_n7523_;
  assign new_n7525_ = ~new_n7512_ & ~new_n7516_;
  assign new_n7526_ = ~new_n7520_ & ~new_n7524_1_;
  assign new_n7527_ = new_n7525_ & new_n7526_;
  assign new_n7528_ = ~ng6052 & new_n7527_;
  assign new_n7529_1_ = ~new_n7507_ & new_n7528_;
  assign new_n7530_ = ~new_n7508_ & ~new_n7529_1_;
  assign new_n7531_ = pg35 & ~new_n7530_;
  assign n1472 = new_n7506_ | new_n7531_;
  assign new_n7533_1_ = ~pg35 & ng1608;
  assign new_n7534_ = ~ng2145 & new_n6226_;
  assign new_n7535_ = ~new_n5399_ & ~new_n6230_1_;
  assign new_n7536_ = ~new_n7534_ & new_n7535_;
  assign new_n7537_1_ = ~pg33533 & new_n7536_;
  assign new_n7538_ = pg25259 & ~new_n7537_1_;
  assign new_n7539_ = ng1620 & ~new_n7538_;
  assign new_n7540_ = ng4180 & new_n7535_;
  assign new_n7541_ = ~new_n7536_ & ~new_n7540_;
  assign new_n7542_1_ = ng1242 & new_n7536_;
  assign new_n7543_ = ~new_n7541_ & ~new_n7542_1_;
  assign new_n7544_ = new_n7538_ & ~new_n7543_;
  assign new_n7545_ = ~new_n7539_ & ~new_n7544_;
  assign new_n7546_ = pg35 & ~new_n7545_;
  assign n1477 = new_n7533_1_ | new_n7546_;
  assign new_n7548_ = ~pg35 & ng2465;
  assign new_n7549_ = ~ng2704 & new_n7167_;
  assign new_n7550_ = ~new_n5302_ & ~new_n6511_;
  assign new_n7551_1_ = ~new_n7549_ & new_n7550_;
  assign new_n7552_ = ng1322 & new_n7195_;
  assign new_n7553_ = new_n6518_1_ & new_n7552_;
  assign new_n7554_ = ng1426 & ~new_n7553_;
  assign new_n7555_ = new_n7551_1_ & ~new_n7554_;
  assign new_n7556_1_ = ~new_n4724_ & new_n5653_1_;
  assign new_n7557_ = ~pg113 & new_n7556_1_;
  assign new_n7558_ = ng112 & new_n7557_;
  assign new_n7559_ = ng2465 & ~new_n7558_;
  assign new_n7560_ = ~new_n7555_ & new_n7559_;
  assign new_n7561_1_ = ng2495 & new_n7555_;
  assign new_n7562_ = ~new_n7560_ & ~new_n7561_1_;
  assign new_n7563_ = pg35 & ~new_n7562_;
  assign n1486 = new_n7548_ | new_n7563_;
  assign new_n7565_ = ~pg35 & ng5563;
  assign new_n7566_1_ = ng5511 & ~ng5517;
  assign new_n7567_ = new_n6885_ & new_n7566_1_;
  assign new_n7568_ = ng5583 & ~new_n7567_;
  assign new_n7569_ = ~new_n5966_ & new_n7567_;
  assign new_n7570_ = ~new_n7568_ & ~new_n7569_;
  assign new_n7571_1_ = pg35 & ~new_n7570_;
  assign n1491 = new_n7565_ | new_n7571_1_;
  assign new_n7573_ = ~pg35 & ng2130;
  assign new_n7574_ = n5005 & new_n6181_;
  assign new_n7575_ = ng2138 & ~new_n6181_;
  assign new_n7576_1_ = ~new_n7574_ & ~new_n7575_;
  assign new_n7577_ = pg35 & ~new_n7576_1_;
  assign n1496 = new_n7573_ | new_n7577_;
  assign new_n7579_ = ~pg35 & ng5228;
  assign new_n7580_1_ = ~ng5188 & ng5180;
  assign new_n7581_ = ng5170 & ~ng5164;
  assign new_n7582_ = new_n7580_1_ & new_n7581_;
  assign new_n7583_ = ng5244 & ~new_n7582_;
  assign new_n7584_1_ = ~new_n5966_ & new_n7582_;
  assign new_n7585_ = ~new_n7583_ & ~new_n7584_1_;
  assign new_n7586_ = pg35 & ~new_n7585_;
  assign n1501 = new_n7579_ | new_n7586_;
  assign new_n7588_ = ~pg35 & ng921;
  assign new_n7589_1_ = ng936 & ng1227;
  assign new_n7590_ = ~new_n7074_ & new_n7589_1_;
  assign new_n7591_ = ~ng936 & new_n7074_;
  assign new_n7592_ = ~new_n7590_ & ~new_n7591_;
  assign new_n7593_ = pg35 & ~new_n7592_;
  assign n1506 = new_n7588_ | new_n7593_;
  assign new_n7595_ = ~pg35 & ng433;
  assign new_n7596_ = ng429 & ~new_n6067_;
  assign new_n7597_ = ng433 & new_n6067_;
  assign new_n7598_ = ~new_n7596_ & ~new_n7597_;
  assign new_n7599_1_ = pg35 & ~new_n7598_;
  assign n1511 = new_n7595_ | new_n7599_1_;
  assign new_n7601_ = ~pg35 & ng4849;
  assign new_n7602_ = ng4843 & ng4878;
  assign new_n7603_1_ = ng4849 & new_n7602_;
  assign new_n7604_ = ng63 & new_n5870_;
  assign new_n7605_ = new_n4735_ & new_n7604_;
  assign new_n7606_ = ~new_n5679_ & ~new_n7605_;
  assign new_n7607_1_ = ~ng4854 & new_n7606_;
  assign new_n7608_ = new_n7603_1_ & new_n7607_1_;
  assign new_n7609_ = ng4854 & new_n7606_;
  assign new_n7610_ = ~new_n7603_1_ & new_n7609_;
  assign new_n7611_ = ~new_n7608_ & ~new_n7610_;
  assign new_n7612_1_ = pg35 & ~new_n7611_;
  assign n1516 = new_n7601_ | new_n7612_1_;
  assign new_n7614_ = ~pg35 & ng2894;
  assign new_n7615_ = ng12 & new_n4951_;
  assign new_n7616_ = n6079 & new_n7615_;
  assign new_n7617_1_ = ng37 & ~new_n7615_;
  assign new_n7618_ = ~new_n7616_ & ~new_n7617_1_;
  assign new_n7619_ = pg35 & ~new_n7618_;
  assign n1521 = new_n7614_ | new_n7619_;
  assign new_n7621_ = ~pg35 & ng6377;
  assign new_n7622_1_ = ng6381 & ~new_n7307_;
  assign new_n7623_ = ~ng6381 & new_n7307_;
  assign new_n7624_ = ~new_n7622_1_ & ~new_n7623_;
  assign new_n7625_ = pg35 & ~new_n7624_;
  assign n1526 = new_n7621_ | new_n7625_;
  assign new_n7627_1_ = ~pg35 & ng4284;
  assign new_n7628_ = ng4287 & ng4291;
  assign new_n7629_ = ng4287 & ~new_n7628_;
  assign new_n7630_ = ng4291 & ~new_n7628_;
  assign new_n7631_ = ~new_n7629_ & ~new_n7630_;
  assign new_n7632_1_ = ~ng4287 & ~new_n7631_;
  assign new_n7633_ = ~new_n7631_ & ~new_n7632_1_;
  assign new_n7634_ = ~ng4287 & ~new_n7632_1_;
  assign new_n7635_ = ~new_n7633_ & ~new_n7634_;
  assign new_n7636_ = pg35 & ~new_n7635_;
  assign n1536 = new_n7627_1_ | new_n7636_;
  assign new_n7638_ = ~pg35 & ng2763;
  assign new_n7639_ = ng2741 & ~ng2748;
  assign new_n7640_ = ~ng2756 & new_n7639_;
  assign new_n7641_1_ = ~ng2756 & ~ng2748;
  assign new_n7642_ = ~new_n6041_1_ & ~new_n7641_1_;
  assign new_n7643_ = ~ng1632 & new_n7642_;
  assign new_n7644_ = ~ng2767 & ~new_n7643_;
  assign new_n7645_ = ~new_n7640_ & ~new_n7644_;
  assign new_n7646_1_ = pg35 & new_n7645_;
  assign n1541 = new_n7638_ | new_n7646_1_;
  assign new_n7648_ = ~pg35 & ng5893;
  assign new_n7649_ = ~ng5881 & ng5873;
  assign new_n7650_ = ng5857 & ~ng5863;
  assign new_n7651_1_ = new_n7649_ & new_n7650_;
  assign new_n7652_ = ng5921 & ~new_n7651_1_;
  assign new_n7653_ = ~new_n5966_ & new_n7651_1_;
  assign new_n7654_ = ~new_n7652_ & ~new_n7653_;
  assign new_n7655_ = pg35 & ~new_n7654_;
  assign n1551 = new_n7648_ | new_n7655_;
  assign new_n7657_ = ~pg35 & ng5057;
  assign new_n7658_ = ~ng5046 & ng5057;
  assign new_n7659_ = ~ng5041 & new_n7658_;
  assign new_n7660_1_ = pg84 & new_n7659_;
  assign new_n7661_ = ng5022 & new_n7660_1_;
  assign new_n7662_ = ~ng5052 & ng5057;
  assign new_n7663_ = ~ng5046 & new_n7662_;
  assign new_n7664_ = ~pg84 & new_n7663_;
  assign new_n7665_ = ng5022 & new_n7664_;
  assign new_n7666_ = ~new_n7661_ & ~new_n7665_;
  assign new_n7667_ = pg35 & new_n7666_;
  assign n1565 = new_n7657_ | new_n7667_;
  assign new_n7669_ = ~pg35 & ng1052;
  assign new_n7670_ = ~ng990 & ~ng1056;
  assign new_n7671_ = ~ng1157 & new_n7670_;
  assign new_n7672_ = ng1227 & ~new_n7671_;
  assign new_n7673_ = ng1052 & new_n7672_;
  assign new_n7674_ = ng1061 & new_n7673_;
  assign new_n7675_ = ~ng1061 & ~new_n7673_;
  assign new_n7676_ = ~new_n7674_ & ~new_n7675_;
  assign new_n7677_ = ~ng979 & new_n7676_;
  assign new_n7678_ = pg35 & new_n7677_;
  assign n1570 = new_n7669_ | new_n7678_;
  assign new_n7680_ = ~pg35 & ng4405;
  assign new_n7681_ = ~ng4414 & ~ng4405;
  assign new_n7682_ = ~ng4411 & new_n7681_;
  assign new_n7683_ = ~ng4375 & new_n7682_;
  assign new_n7684_ = ~ng4408 & new_n7683_;
  assign new_n7685_ = ~ng4392 & new_n7684_;
  assign new_n7686_ = ng4388 & new_n7685_;
  assign new_n7687_ = ~ng4405 & ~new_n7686_;
  assign new_n7688_ = pg35 & ~new_n7687_;
  assign n1575 = new_n7680_ | new_n7688_;
  assign new_n7690_ = ~pg35 & ng3423;
  assign new_n7691_ = ~ng3431 & ng3423;
  assign new_n7692_ = ng3431 & ~ng3423;
  assign new_n7693_ = ~new_n7691_ & ~new_n7692_;
  assign new_n7694_ = pg35 & ~new_n7693_;
  assign n1585 = new_n7690_ | new_n7694_;
  assign new_n7696_ = ~pg35 & ng3594;
  assign new_n7697_ = ng3506 & ng3512;
  assign new_n7698_ = new_n6769_ & new_n7697_;
  assign new_n7699_ = ng3610 & ~new_n7698_;
  assign new_n7700_ = ~new_n5966_ & new_n7698_;
  assign new_n7701_ = ~new_n7699_ & ~new_n7700_;
  assign new_n7702_ = pg35 & ~new_n7701_;
  assign n1590 = new_n7696_ | new_n7702_;
  assign new_n7704_ = ~pg35 & ng4966;
  assign new_n7705_ = ng4966 & ng4983;
  assign new_n7706_ = new_n5679_ & new_n7705_;
  assign new_n7707_ = ~new_n4724_ & new_n4735_;
  assign new_n7708_ = new_n6158_ & new_n7707_;
  assign new_n7709_ = ng4975 & ~new_n7708_;
  assign new_n7710_ = ~new_n7706_ & new_n7709_;
  assign new_n7711_ = ~ng4975 & ~new_n7708_;
  assign new_n7712_ = new_n7706_ & new_n7711_;
  assign new_n7713_ = ~new_n7710_ & ~new_n7712_;
  assign new_n7714_ = pg35 & ~new_n7713_;
  assign n1595 = new_n7704_ | new_n7714_;
  assign new_n7716_ = ~pg35 & ng4430;
  assign new_n7717_ = ng4401 & ng4434;
  assign new_n7718_ = ng4401 & ~new_n7717_;
  assign new_n7719_ = ng4434 & ~new_n7717_;
  assign new_n7720_ = ~new_n7718_ & ~new_n7719_;
  assign new_n7721_ = ng4388 & ng4430;
  assign new_n7722_ = ng4430 & ~new_n7721_;
  assign new_n7723_ = ng4388 & ~new_n7721_;
  assign new_n7724_ = ~new_n7722_ & ~new_n7723_;
  assign new_n7725_ = new_n7720_ & new_n7724_;
  assign new_n7726_ = pg35 & ~new_n7725_;
  assign n1600 = new_n7716_ | new_n7726_;
  assign new_n7728_ = ~pg35 & ng4104;
  assign new_n7729_ = pg124 & ng4146;
  assign new_n7730_ = pg120 & ~ng4146;
  assign new_n7731_ = ~new_n7729_ & ~new_n7730_;
  assign new_n7732_ = pg35 & ~new_n7731_;
  assign n1605 = new_n7728_ | new_n7732_;
  assign new_n7734_ = ~pg35 & ng1830;
  assign new_n7735_ = new_n6683_ & new_n6807_;
  assign new_n7736_ = ng1834 & ~new_n7735_;
  assign new_n7737_ = ~ng1834 & new_n7735_;
  assign new_n7738_ = ~new_n7736_ & ~new_n7737_;
  assign new_n7739_ = pg35 & ~new_n7738_;
  assign n1610 = new_n7734_ | new_n7739_;
  assign new_n7741_ = ~pg35 & ng5698;
  assign new_n7742_ = ~ng4709 & new_n6695_;
  assign new_n7743_ = new_n5669_ & new_n7742_;
  assign new_n7744_ = ng4743 & new_n7743_;
  assign new_n7745_ = ng4674 & ~new_n7744_;
  assign new_n7746_ = ng93 & ~new_n4724_;
  assign new_n7747_ = ~pg113 & new_n7746_;
  assign new_n7748_ = new_n4747_1_ & new_n7747_;
  assign new_n7749_ = new_n7745_ & new_n7748_;
  assign new_n7750_ = new_n4734_ & new_n7749_;
  assign new_n7751_ = ~ng5703 & ~new_n7750_;
  assign new_n7752_ = new_n7745_ & new_n7751_;
  assign new_n7753_ = ng5703 & ~new_n7745_;
  assign new_n7754_ = ~new_n7752_ & ~new_n7753_;
  assign new_n7755_ = pg35 & ~new_n7754_;
  assign n1615 = new_n7741_ | new_n7755_;
  assign new_n7757_ = ~pg35 & ng4492;
  assign new_n7758_ = ~ng59 & new_n5871_;
  assign new_n7759_ = ng4581 & ~new_n7758_;
  assign new_n7760_ = ng4512 & ~ng4581;
  assign new_n7761_ = ~new_n7759_ & ~new_n7760_;
  assign new_n7762_ = ~new_n5871_ & new_n7761_;
  assign new_n7763_ = ng4483 & ng4489;
  assign new_n7764_ = ng4486 & new_n7763_;
  assign new_n7765_ = ng4492 & new_n7764_;
  assign new_n7766_ = ~ng2988 & ~new_n7765_;
  assign new_n7767_ = new_n5871_ & new_n7766_;
  assign new_n7768_ = ~new_n7762_ & ~new_n7767_;
  assign new_n7769_ = pg35 & new_n7768_;
  assign n1620 = new_n7757_ | new_n7769_;
  assign new_n7771_ = ~pg35 & ng1129;
  assign new_n7772_ = ng1116 & new_n7021_;
  assign new_n7773_ = ng1141 & ~new_n7772_;
  assign new_n7774_ = ~ng1146 & ~ng1099;
  assign new_n7775_ = ~ng976 & new_n4686_;
  assign new_n7776_ = ng956 & new_n7775_;
  assign new_n7777_ = ng956 & ~new_n7776_;
  assign new_n7778_ = new_n7775_ & ~new_n7776_;
  assign new_n7779_ = ~new_n7777_ & ~new_n7778_;
  assign new_n7780_ = ng1141 & ~new_n7779_;
  assign new_n7781_ = ~new_n7774_ & new_n7780_;
  assign new_n7782_ = new_n7774_ & ~new_n7779_;
  assign new_n7783_ = ~new_n7781_ & ~new_n7782_;
  assign new_n7784_ = new_n7772_ & ~new_n7783_;
  assign new_n7785_ = ~new_n7773_ & ~new_n7784_;
  assign new_n7786_ = pg35 & ~new_n7785_;
  assign n1625 = new_n7771_ | new_n7786_;
  assign new_n7788_ = ~pg35 & ng6116;
  assign new_n7789_ = ng6113 & ~ng6105;
  assign new_n7790_ = ~ng6116 & ~new_n7789_;
  assign new_n7791_ = ~ng6120 & new_n7790_;
  assign new_n7792_ = ng6120 & ng6116;
  assign new_n7793_ = ng6113 & ~ng6109;
  assign new_n7794_ = ~new_n7791_ & ~new_n7792_;
  assign new_n7795_ = ~new_n7793_ & new_n7794_;
  assign new_n7796_ = pg35 & ~new_n7795_;
  assign n1630 = new_n7788_ | new_n7796_;
  assign new_n7798_ = ~pg35 & ng4504;
  assign new_n7799_ = ~ng4572 & new_n5871_;
  assign new_n7800_ = ng4581 & ~new_n7799_;
  assign new_n7801_ = ng4504 & ~ng4581;
  assign new_n7802_ = ~new_n7800_ & ~new_n7801_;
  assign new_n7803_ = pg35 & ~new_n7802_;
  assign n1635 = new_n7798_ | new_n7803_;
  assign new_n7805_ = ~pg35 & ng4300;
  assign new_n7806_ = ng12 & new_n4930_;
  assign new_n7807_ = n4465 & new_n7806_;
  assign new_n7808_ = ng4253 & ~new_n7806_;
  assign new_n7809_ = ~new_n7807_ & ~new_n7808_;
  assign new_n7810_ = pg35 & ~new_n7809_;
  assign n1640 = new_n7805_ | new_n7810_;
  assign new_n7812_ = ~pg35 & ng4552;
  assign new_n7813_ = ~ng4575 & new_n5871_;
  assign new_n7814_ = ng4581 & ~new_n7813_;
  assign new_n7815_ = ng4552 & ~ng4581;
  assign new_n7816_ = ~new_n7814_ & ~new_n7815_;
  assign new_n7817_ = pg35 & ~new_n7816_;
  assign n1645 = new_n7812_ | new_n7817_;
  assign new_n7819_ = ~pg35 & ng1430;
  assign new_n7820_ = ~ng1548 & ng1430;
  assign new_n7821_ = ng1548 & ~ng1430;
  assign new_n7822_ = ~new_n7820_ & ~new_n7821_;
  assign new_n7823_ = pg35 & ~new_n7822_;
  assign n1650 = new_n7819_ | new_n7823_;
  assign new_n7825_ = ~pg35 & ng4281;
  assign new_n7826_ = ng4281 & ng4277;
  assign new_n7827_ = ng4277 & ~new_n7826_;
  assign new_n7828_ = ng4281 & ~new_n7826_;
  assign new_n7829_ = ~new_n7827_ & ~new_n7828_;
  assign new_n7830_ = pg35 & ~new_n7829_;
  assign n1655 = new_n7825_ | new_n7830_;
  assign new_n7832_ = ~pg35 & ng376;
  assign new_n7833_ = ~ng385 & ~new_n5993_1_;
  assign new_n7834_ = ~new_n5993_1_ & ~new_n7833_;
  assign new_n7835_ = ~ng385 & ~new_n7833_;
  assign new_n7836_ = ~new_n7834_ & ~new_n7835_;
  assign new_n7837_ = pg35 & ~new_n7836_;
  assign n1660 = new_n7832_ | new_n7837_;
  assign new_n7839_ = ~pg35 & ng287;
  assign new_n7840_ = ng291 & new_n6021_;
  assign new_n7841_ = ~new_n6024_ & new_n7840_;
  assign new_n7842_ = ~ng291 & new_n6024_;
  assign new_n7843_ = ~new_n7841_ & ~new_n7842_;
  assign new_n7844_ = pg35 & ~new_n7843_;
  assign n1665 = new_n7839_ | new_n7844_;
  assign new_n7846_ = ~pg35 & ng3147;
  assign new_n7847_ = ng3111 & ~new_n7152_;
  assign new_n7848_ = ng3147 & new_n7152_;
  assign new_n7849_ = ~new_n7847_ & ~new_n7848_;
  assign new_n7850_ = pg35 & ~new_n7849_;
  assign n1675 = new_n7846_ | new_n7850_;
  assign new_n7852_ = ~pg35 & ng655;
  assign new_n7853_ = ng691 & ~new_n5989_;
  assign new_n7854_ = ~ng411 & ng417;
  assign new_n7855_ = ~ng424 & new_n7854_;
  assign new_n7856_ = ~ng691 & ~new_n7855_;
  assign new_n7857_ = ~new_n7853_ & ~new_n7856_;
  assign new_n7858_ = new_n5994_ & new_n7857_;
  assign new_n7859_ = ng718 & ~new_n7858_;
  assign new_n7860_ = ng655 & new_n7858_;
  assign new_n7861_ = ~new_n7859_ & ~new_n7860_;
  assign new_n7862_ = pg35 & ~new_n7861_;
  assign n1680 = new_n7852_ | new_n7862_;
  assign new_n7864_ = ~pg35 & ng6239;
  assign new_n7865_ = ~ng6227 & ng6219;
  assign new_n7866_ = ~ng6209 & ng6203;
  assign new_n7867_ = new_n7865_ & new_n7866_;
  assign new_n7868_ = ng6267 & ~new_n7867_;
  assign new_n7869_ = ~new_n5966_ & new_n7867_;
  assign new_n7870_ = ~new_n7868_ & ~new_n7869_;
  assign new_n7871_ = pg35 & ~new_n7870_;
  assign n1690 = new_n7864_ | new_n7871_;
  assign new_n7873_ = ~pg35 & ng3103;
  assign new_n7874_ = ~ng3103 & ng3096;
  assign new_n7875_ = ~ng3010 & ~new_n7874_;
  assign new_n7876_ = ~ng3092 & ~new_n7875_;
  assign new_n7877_ = pg35 & new_n7876_;
  assign n1695 = new_n7873_ | new_n7877_;
  assign new_n7879_ = ~pg35 & ng2393;
  assign new_n7880_ = ng2704 & new_n6508_1_;
  assign new_n7881_ = ~new_n5342_ & ~new_n6511_;
  assign new_n7882_ = ~new_n7880_ & new_n7881_;
  assign new_n7883_ = ng1322 & new_n6827_;
  assign new_n7884_ = new_n6518_1_ & new_n7883_;
  assign new_n7885_ = ng1422 & ~new_n7884_;
  assign new_n7886_ = new_n7882_ & ~new_n7885_;
  assign new_n7887_ = ~ng2361 & ~ng2287;
  assign new_n7888_ = ~new_n7886_ & new_n7887_;
  assign new_n7889_ = ng2399 & ~new_n7888_;
  assign new_n7890_ = ng2393 & new_n7888_;
  assign new_n7891_ = ~new_n7889_ & ~new_n7890_;
  assign new_n7892_ = pg35 & ~new_n7891_;
  assign n1700 = new_n7879_ | new_n7892_;
  assign new_n7894_ = ~pg35 & ng2864;
  assign new_n7895_ = ng12 & new_n4955_1_;
  assign new_n7896_ = n2287 & new_n7895_;
  assign new_n7897_ = ~ng2898 & new_n4683_;
  assign new_n7898_ = ~new_n7896_ & ~new_n7897_;
  assign new_n7899_ = pg35 & new_n7898_;
  assign n1705 = new_n7894_ | new_n7899_;
  assign new_n7901_ = ~pg35 & ng4375;
  assign new_n7902_ = ng4392 & new_n7684_;
  assign new_n7903_ = ng4375 & ng4382;
  assign new_n7904_ = ~new_n7684_ & new_n7903_;
  assign new_n7905_ = ~new_n7902_ & ~new_n7904_;
  assign new_n7906_ = pg35 & ~new_n7905_;
  assign n1710 = new_n7901_ | new_n7906_;
  assign new_n7908_ = ~pg35 & ng5965;
  assign new_n7909_ = ~ng5990 & ~ng6049;
  assign new_n7910_ = ~ng6035 & new_n7909_;
  assign new_n7911_ = ng6023 & ng5941;
  assign new_n7912_ = new_n7910_ & new_n7911_;
  assign new_n7913_ = ng5990 & ~ng6049;
  assign new_n7914_ = ~ng6035 & new_n7913_;
  assign new_n7915_ = ng5913 & ng6031;
  assign new_n7916_ = new_n7914_ & new_n7915_;
  assign new_n7917_ = ~ng5990 & ng6049;
  assign new_n7918_ = ~ng6035 & new_n7917_;
  assign new_n7919_ = ng6027 & ng5957;
  assign new_n7920_ = new_n7918_ & new_n7919_;
  assign new_n7921_ = ~ng6035 & new_n4745_;
  assign new_n7922_ = ng6005 & ng5909;
  assign new_n7923_ = new_n7921_ & new_n7922_;
  assign new_n7924_ = ~new_n7912_ & ~new_n7916_;
  assign new_n7925_ = ~new_n7920_ & ~new_n7923_;
  assign new_n7926_ = new_n7924_ & new_n7925_;
  assign new_n7927_ = ng6035 & new_n7909_;
  assign new_n7928_ = ng5897 & ng6031;
  assign new_n7929_ = new_n7927_ & new_n7928_;
  assign new_n7930_ = ng6035 & ng6005;
  assign new_n7931_ = ng6005 & ~new_n7930_;
  assign new_n7932_ = ng6035 & ~new_n7930_;
  assign new_n7933_ = ~new_n7931_ & ~new_n7932_;
  assign new_n7934_ = new_n7913_ & new_n7933_;
  assign new_n7935_ = ng5921 & ng5983;
  assign new_n7936_ = new_n7934_ & new_n7935_;
  assign new_n7937_ = ng6035 & new_n7917_;
  assign new_n7938_ = ng5893 & ng6005;
  assign new_n7939_ = new_n7937_ & new_n7938_;
  assign new_n7940_ = new_n4745_ & new_n7933_;
  assign new_n7941_ = ng6012 & ng5937;
  assign new_n7942_ = new_n7940_ & new_n7941_;
  assign new_n7943_ = ~new_n7929_ & ~new_n7936_;
  assign new_n7944_ = ~new_n7939_ & ~new_n7942_;
  assign new_n7945_ = new_n7943_ & new_n7944_;
  assign new_n7946_ = ng5889 & ng6000;
  assign new_n7947_ = new_n7927_ & new_n7946_;
  assign new_n7948_ = ng6035 & new_n7913_;
  assign new_n7949_ = ng6023 & ng5933;
  assign new_n7950_ = new_n7948_ & new_n7949_;
  assign new_n7951_ = ng5917 & ng6019;
  assign new_n7952_ = new_n7937_ & new_n7951_;
  assign new_n7953_ = ng6035 & new_n4745_;
  assign new_n7954_ = ng6027 & ng5949;
  assign new_n7955_ = new_n7953_ & new_n7954_;
  assign new_n7956_ = ~new_n7947_ & ~new_n7950_;
  assign new_n7957_ = ~new_n7952_ & ~new_n7955_;
  assign new_n7958_ = new_n7956_ & new_n7957_;
  assign new_n7959_ = new_n7909_ & new_n7933_;
  assign new_n7960_ = ng5953 & ng5969;
  assign new_n7961_ = new_n7959_ & new_n7960_;
  assign new_n7962_ = ng5901 & ng6000;
  assign new_n7963_ = new_n7914_ & new_n7962_;
  assign new_n7964_ = ng5976 & ng5905;
  assign new_n7965_ = new_n7918_ & new_n7964_;
  assign new_n7966_ = ng6019 & ng5925;
  assign new_n7967_ = new_n7921_ & new_n7966_;
  assign new_n7968_ = ~new_n7961_ & ~new_n7963_;
  assign new_n7969_ = ~new_n7965_ & ~new_n7967_;
  assign new_n7970_ = new_n7968_ & new_n7969_;
  assign new_n7971_ = new_n7945_ & new_n7958_;
  assign new_n7972_ = new_n7970_ & new_n7971_;
  assign new_n7973_ = new_n7909_ & ~new_n7933_;
  assign new_n7974_ = ng5929 & ng5983;
  assign new_n7975_ = new_n7973_ & new_n7974_;
  assign new_n7976_ = new_n7913_ & ~new_n7933_;
  assign new_n7977_ = ng5969 & ng5961;
  assign new_n7978_ = new_n7976_ & new_n7977_;
  assign new_n7979_ = new_n7917_ & ~new_n7933_;
  assign new_n7980_ = ng6012 & ng5945;
  assign new_n7981_ = new_n7979_ & new_n7980_;
  assign new_n7982_ = ng5976 & ng5965;
  assign new_n7983_ = new_n7953_ & new_n7982_;
  assign new_n7984_ = ~new_n7975_ & ~new_n7978_;
  assign new_n7985_ = ~new_n7981_ & ~new_n7983_;
  assign new_n7986_ = new_n7984_ & new_n7985_;
  assign new_n7987_ = new_n7926_ & new_n7972_;
  assign new_n7988_ = new_n7986_ & new_n7987_;
  assign new_n7989_ = new_n6353_ & ~new_n7988_;
  assign new_n7990_ = ng4831 & ~new_n6353_;
  assign new_n7991_ = ~new_n7989_ & ~new_n7990_;
  assign new_n7992_ = pg35 & ~new_n7991_;
  assign n1715 = new_n7908_ | new_n7992_;
  assign new_n7994_ = ~pg35 & ng5881;
  assign new_n7995_ = ~ng5881 & ~ng5873;
  assign new_n7996_ = ~ng5857 & ~ng5863;
  assign new_n7997_ = ~ng5869 & new_n7996_;
  assign new_n7998_ = new_n7995_ & new_n7997_;
  assign new_n7999_ = ng5889 & ~new_n7998_;
  assign new_n8000_ = ~new_n5966_ & new_n7998_;
  assign new_n8001_ = ~new_n7999_ & ~new_n8000_;
  assign new_n8002_ = pg35 & ~new_n8001_;
  assign n1720 = new_n7994_ | new_n8002_;
  assign new_n8004_ = ~pg35 & ng832;
  assign new_n8005_ = ng817 & new_n6067_;
  assign new_n8006_ = ng832 & new_n8005_;
  assign new_n8007_ = ng812 & ng847;
  assign new_n8008_ = ~ng837 & ng847;
  assign new_n8009_ = ~new_n8007_ & ~new_n8008_;
  assign new_n8010_ = ng822 & new_n8009_;
  assign new_n8011_ = ~new_n8006_ & new_n8010_;
  assign new_n8012_ = ~ng822 & new_n8009_;
  assign new_n8013_ = new_n8006_ & new_n8012_;
  assign new_n8014_ = ~new_n8011_ & ~new_n8013_;
  assign new_n8015_ = pg35 & ~new_n8014_;
  assign n1725 = new_n8004_ | new_n8015_;
  assign new_n8017_ = new_n5767_ & pg33659;
  assign new_n8018_ = ~new_n5767_ & ~new_n5818_;
  assign n1730 = new_n8017_ | new_n8018_;
  assign new_n8020_ = ~pg35 & ng2108;
  assign new_n8021_ = ~ng2070 & ~ng1996;
  assign new_n8022_ = ~new_n7025_ & new_n8021_;
  assign new_n8023_ = ng2112 & ~new_n8022_;
  assign new_n8024_ = ng2102 & ~ng2108;
  assign new_n8025_ = ng2102 & ~new_n8024_;
  assign new_n8026_ = ~ng2108 & ~new_n8024_;
  assign new_n8027_ = ~new_n8025_ & ~new_n8026_;
  assign new_n8028_ = new_n8022_ & ~new_n8027_;
  assign new_n8029_ = ~new_n8023_ & ~new_n8028_;
  assign new_n8030_ = pg35 & ~new_n8029_;
  assign n1740 = new_n8020_ | new_n8030_;
  assign new_n8032_ = ~pg35 & ng5535;
  assign new_n8033_ = ~ng5535 & ~ng5527;
  assign new_n8034_ = ~ng5511 & ~ng5517;
  assign new_n8035_ = ~ng5523 & new_n8034_;
  assign new_n8036_ = new_n8033_ & new_n8035_;
  assign new_n8037_ = ng5543 & ~new_n8036_;
  assign new_n8038_ = ~new_n5966_ & new_n8036_;
  assign new_n8039_ = ~new_n8037_ & ~new_n8038_;
  assign new_n8040_ = pg35 & ~new_n8039_;
  assign n1745 = new_n8032_ | new_n8040_;
  assign new_n8042_ = ~pg35 & ng4438;
  assign new_n8043_ = ~ng4449 & ~ng4452;
  assign new_n8044_ = ~ng4443 & new_n8043_;
  assign new_n8045_ = ~ng4438 & new_n8044_;
  assign new_n8046_ = ~ng4446 & new_n8045_;
  assign new_n8047_ = ng4392 & new_n8046_;
  assign new_n8048_ = ng4382 & ng4438;
  assign new_n8049_ = ~new_n8046_ & new_n8048_;
  assign new_n8050_ = ~new_n8047_ & ~new_n8049_;
  assign new_n8051_ = pg35 & ~new_n8050_;
  assign n1750 = new_n8042_ | new_n8051_;
  assign new_n8053_ = ~pg35 & ng298;
  assign new_n8054_ = ~ng142 & new_n6030_;
  assign new_n8055_ = ng142 & new_n6021_;
  assign new_n8056_ = ~new_n6030_ & new_n8055_;
  assign new_n8057_ = ~new_n8054_ & ~new_n8056_;
  assign new_n8058_ = pg35 & ~new_n8057_;
  assign n1754 = new_n8053_ | new_n8058_;
  assign new_n8060_ = ~pg35 & ng5112;
  assign new_n8061_ = ng5105 & ~ng5112;
  assign new_n8062_ = ~ng5022 & ~new_n8061_;
  assign new_n8063_ = ~ng5101 & ~new_n8062_;
  assign new_n8064_ = pg35 & new_n8063_;
  assign n1759 = new_n8060_ | new_n8064_;
  assign new_n8066_ = ~pg35 & ng1454;
  assign new_n8067_ = ng1459 & new_n6827_;
  assign new_n8068_ = new_n7472_ & new_n8067_;
  assign new_n8069_ = ng1448 & ng1454;
  assign new_n8070_ = ng1448 & ~new_n8069_;
  assign new_n8071_ = ng1454 & ~new_n8069_;
  assign new_n8072_ = ~new_n8070_ & ~new_n8071_;
  assign new_n8073_ = new_n8068_ & ~new_n8072_;
  assign new_n8074_ = ng1448 & ~new_n8068_;
  assign new_n8075_ = ~new_n8073_ & ~new_n8074_;
  assign new_n8076_ = pg35 & ~new_n8075_;
  assign n1769 = new_n8066_ | new_n8076_;
  assign new_n8078_ = ~pg35 & ng3945;
  assign new_n8079_ = ng3857 & ng3863;
  assign new_n8080_ = new_n7010_ & new_n8079_;
  assign new_n8081_ = ng3961 & ~new_n8080_;
  assign new_n8082_ = ~new_n5966_ & new_n8080_;
  assign new_n8083_ = ~new_n8081_ & ~new_n8082_;
  assign new_n8084_ = pg35 & ~new_n8083_;
  assign n1774 = new_n8078_ | new_n8084_;
  assign new_n8086_ = ~pg35 & ng1002;
  assign new_n8087_ = ng1018 & ~new_n6140_;
  assign new_n8088_ = new_n6140_ & new_n6141_;
  assign new_n8089_ = ~new_n8087_ & ~new_n8088_;
  assign new_n8090_ = pg35 & ~new_n8089_;
  assign n1779 = new_n8086_ | new_n8090_;
  assign new_n8092_ = ~pg35 & ng5016;
  assign new_n8093_ = ng5022 & ~ng5016;
  assign new_n8094_ = ng5016 & ng5062;
  assign new_n8095_ = ~new_n8093_ & ~new_n8094_;
  assign new_n8096_ = ~ng5029 & ~new_n8095_;
  assign new_n8097_ = ng5046 & ~ng5057;
  assign new_n8098_ = ng5041 & new_n8097_;
  assign new_n8099_ = pg84 & new_n8098_;
  assign new_n8100_ = ng5062 & new_n8099_;
  assign new_n8101_ = ng5052 & ~ng5057;
  assign new_n8102_ = ng5046 & new_n8101_;
  assign new_n8103_ = ~pg84 & new_n8102_;
  assign new_n8104_ = ng5062 & new_n8103_;
  assign new_n8105_ = ~new_n7661_ & ~new_n8100_;
  assign new_n8106_ = ~new_n7665_ & ~new_n8104_;
  assign new_n8107_ = new_n8105_ & new_n8106_;
  assign new_n8108_ = ng5029 & new_n8107_;
  assign new_n8109_ = new_n8095_ & new_n8108_;
  assign new_n8110_ = ~new_n8096_ & ~new_n8109_;
  assign new_n8111_ = pg35 & ~new_n8110_;
  assign n1784 = new_n8092_ | new_n8111_;
  assign new_n8113_ = ~pg35 & ng504;
  assign new_n8114_ = ng504 & ~new_n6494_;
  assign new_n8115_ = new_n6493_1_ & new_n8114_;
  assign new_n8116_ = ng513 & ~new_n6493_1_;
  assign new_n8117_ = ~new_n8115_ & ~new_n8116_;
  assign new_n8118_ = pg35 & ~new_n8117_;
  assign n1789 = new_n8113_ | new_n8118_;
  assign new_n8120_ = ~pg35 & ng2020;
  assign new_n8121_ = ng2070 & ng1996;
  assign new_n8122_ = ~new_n7025_ & new_n8121_;
  assign new_n8123_ = ng2016 & ~new_n8122_;
  assign new_n8124_ = ~new_n7032_ & new_n8122_;
  assign new_n8125_ = ~new_n8123_ & ~new_n8124_;
  assign new_n8126_ = pg35 & ~new_n8125_;
  assign n1799 = new_n8120_ | new_n8126_;
  assign new_n8128_ = ~pg35 & ng5547;
  assign new_n8129_ = ~ng5535 & ng5527;
  assign new_n8130_ = new_n7566_1_ & new_n8129_;
  assign new_n8131_ = ng5575 & ~new_n8130_;
  assign new_n8132_ = ~new_n5966_ & new_n8130_;
  assign new_n8133_ = ~new_n8131_ & ~new_n8132_;
  assign new_n8134_ = pg35 & ~new_n8133_;
  assign n1804 = new_n8128_ | new_n8134_;
  assign new_n8136_ = ~pg35 & ng5046;
  assign new_n8137_ = ~ng5029 & new_n8093_;
  assign new_n8138_ = ~ng5033 & new_n8137_;
  assign new_n8139_ = ~ng5037 & new_n8138_;
  assign new_n8140_ = ~ng5041 & new_n8139_;
  assign new_n8141_ = ~ng5046 & new_n8140_;
  assign new_n8142_ = ng5029 & new_n8094_;
  assign new_n8143_ = ng5033 & new_n8142_;
  assign new_n8144_ = ng5037 & new_n8143_;
  assign new_n8145_ = ng5041 & new_n8144_;
  assign new_n8146_ = ng5046 & new_n8145_;
  assign new_n8147_ = ~new_n8141_ & ~new_n8146_;
  assign new_n8148_ = ng5052 & new_n8107_;
  assign new_n8149_ = new_n8147_ & new_n8148_;
  assign new_n8150_ = ~ng5052 & ~new_n8147_;
  assign new_n8151_ = ~new_n8149_ & ~new_n8150_;
  assign new_n8152_ = pg35 & ~new_n8151_;
  assign n1809 = new_n8136_ | new_n8152_;
  assign new_n8154_ = ~pg35 & ng3408;
  assign new_n8155_ = ng3385 & ~ng3396;
  assign new_n8156_ = ng3380 & new_n8155_;
  assign new_n8157_ = pg84 & new_n8156_;
  assign new_n8158_ = ng3401 & new_n8157_;
  assign new_n8159_ = ng3391 & ~ng3396;
  assign new_n8160_ = ng3385 & new_n8159_;
  assign new_n8161_ = ~pg84 & new_n8160_;
  assign new_n8162_ = ng3401 & new_n8161_;
  assign new_n8163_ = ~new_n8158_ & ~new_n8162_;
  assign new_n8164_ = pg35 & new_n8163_;
  assign n1814 = new_n8154_ | new_n8164_;
  assign new_n8166_ = ~pg35 & ng1988;
  assign new_n8167_ = ng1926 & ng1894;
  assign new_n8168_ = ~ng2783 & new_n5902_1_;
  assign new_n8169_ = new_n5904_ & ~new_n8168_;
  assign new_n8170_ = ~ng2715 & ~new_n8169_;
  assign new_n8171_ = ng2719 & new_n8170_;
  assign new_n8172_ = new_n8167_ & new_n8171_;
  assign new_n8173_ = ng1992 & ~new_n8172_;
  assign new_n8174_ = ~ng1988 & ng1982;
  assign new_n8175_ = ng1982 & ~new_n8174_;
  assign new_n8176_ = ~ng1988 & ~new_n8174_;
  assign new_n8177_ = ~new_n8175_ & ~new_n8176_;
  assign new_n8178_ = new_n8172_ & ~new_n8177_;
  assign new_n8179_ = ~new_n8173_ & ~new_n8178_;
  assign new_n8180_ = pg35 & ~new_n8179_;
  assign n1819 = new_n8166_ | new_n8180_;
  assign new_n8182_ = ~pg35 & ng2970;
  assign new_n8183_ = ng12 & n4955;
  assign new_n8184_ = new_n4937_ & new_n8183_;
  assign new_n8185_ = ~ng301 & ng691;
  assign new_n8186_ = ~ng209 & new_n8185_;
  assign new_n8187_ = ~ng2902 & new_n8186_;
  assign new_n8188_ = ~new_n8184_ & ~new_n8187_;
  assign new_n8189_ = pg35 & new_n8188_;
  assign n1824 = new_n8182_ | new_n8189_;
  assign new_n8191_ = ~pg35 & ng3813;
  assign new_n8192_ = ng3808 & ~new_n6460_1_;
  assign new_n8193_ = ~ng4054 & ~ng3990;
  assign new_n8194_ = ~ng4040 & new_n8193_;
  assign new_n8195_ = ng4023 & ng3941;
  assign new_n8196_ = new_n8194_ & new_n8195_;
  assign new_n8197_ = ~ng4054 & ng3990;
  assign new_n8198_ = ~ng4040 & new_n8197_;
  assign new_n8199_ = ng4031 & ng3913;
  assign new_n8200_ = new_n8198_ & new_n8199_;
  assign new_n8201_ = ng4054 & ~ng3990;
  assign new_n8202_ = ~ng4040 & new_n8201_;
  assign new_n8203_ = ng4027 & ng3957;
  assign new_n8204_ = new_n8202_ & new_n8203_;
  assign new_n8205_ = ~ng4040 & new_n4768_;
  assign new_n8206_ = ng3909 & ng4005;
  assign new_n8207_ = new_n8205_ & new_n8206_;
  assign new_n8208_ = ~new_n8196_ & ~new_n8200_;
  assign new_n8209_ = ~new_n8204_ & ~new_n8207_;
  assign new_n8210_ = new_n8208_ & new_n8209_;
  assign new_n8211_ = ng4040 & new_n8193_;
  assign new_n8212_ = ng4031 & ng3897;
  assign new_n8213_ = new_n8211_ & new_n8212_;
  assign new_n8214_ = ng4040 & ng4005;
  assign new_n8215_ = ng4005 & ~new_n8214_;
  assign new_n8216_ = ng4040 & ~new_n8214_;
  assign new_n8217_ = ~new_n8215_ & ~new_n8216_;
  assign new_n8218_ = new_n8197_ & new_n8217_;
  assign new_n8219_ = ng3983 & ng3921;
  assign new_n8220_ = new_n8218_ & new_n8219_;
  assign new_n8221_ = ng4040 & new_n8201_;
  assign new_n8222_ = ng3893 & ng4005;
  assign new_n8223_ = new_n8221_ & new_n8222_;
  assign new_n8224_ = new_n4768_ & new_n8217_;
  assign new_n8225_ = ng4012 & ng3937;
  assign new_n8226_ = new_n8224_ & new_n8225_;
  assign new_n8227_ = ~new_n8213_ & ~new_n8220_;
  assign new_n8228_ = ~new_n8223_ & ~new_n8226_;
  assign new_n8229_ = new_n8227_ & new_n8228_;
  assign new_n8230_ = ng3889 & ng4000;
  assign new_n8231_ = new_n8211_ & new_n8230_;
  assign new_n8232_ = ng4040 & new_n8197_;
  assign new_n8233_ = ng3933 & ng4023;
  assign new_n8234_ = new_n8232_ & new_n8233_;
  assign new_n8235_ = ng4019 & ng3917;
  assign new_n8236_ = new_n8221_ & new_n8235_;
  assign new_n8237_ = ng4040 & new_n4768_;
  assign new_n8238_ = ng3949 & ng4027;
  assign new_n8239_ = new_n8237_ & new_n8238_;
  assign new_n8240_ = ~new_n8231_ & ~new_n8234_;
  assign new_n8241_ = ~new_n8236_ & ~new_n8239_;
  assign new_n8242_ = new_n8240_ & new_n8241_;
  assign new_n8243_ = new_n8193_ & new_n8217_;
  assign new_n8244_ = ng3969 & ng3953;
  assign new_n8245_ = new_n8243_ & new_n8244_;
  assign new_n8246_ = ng3901 & ng4000;
  assign new_n8247_ = new_n8198_ & new_n8246_;
  assign new_n8248_ = ng3976 & ng3905;
  assign new_n8249_ = new_n8202_ & new_n8248_;
  assign new_n8250_ = ng3925 & ng4019;
  assign new_n8251_ = new_n8205_ & new_n8250_;
  assign new_n8252_ = ~new_n8245_ & ~new_n8247_;
  assign new_n8253_ = ~new_n8249_ & ~new_n8251_;
  assign new_n8254_ = new_n8252_ & new_n8253_;
  assign new_n8255_ = new_n8229_ & new_n8242_;
  assign new_n8256_ = new_n8254_ & new_n8255_;
  assign new_n8257_ = new_n8193_ & ~new_n8217_;
  assign new_n8258_ = ng3983 & ng3929;
  assign new_n8259_ = new_n8257_ & new_n8258_;
  assign new_n8260_ = new_n8197_ & ~new_n8217_;
  assign new_n8261_ = ng3961 & ng3969;
  assign new_n8262_ = new_n8260_ & new_n8261_;
  assign new_n8263_ = new_n8201_ & ~new_n8217_;
  assign new_n8264_ = ng4012 & ng3945;
  assign new_n8265_ = new_n8263_ & new_n8264_;
  assign new_n8266_ = ng3976 & ng3965;
  assign new_n8267_ = new_n8237_ & new_n8266_;
  assign new_n8268_ = ~new_n8259_ & ~new_n8262_;
  assign new_n8269_ = ~new_n8265_ & ~new_n8267_;
  assign new_n8270_ = new_n8268_ & new_n8269_;
  assign new_n8271_ = new_n8210_ & new_n8256_;
  assign new_n8272_ = new_n8270_ & new_n8271_;
  assign new_n8273_ = new_n8192_ & ~new_n8272_;
  assign new_n8274_ = new_n8192_ & ~new_n8273_;
  assign new_n8275_ = ~new_n8272_ & ~new_n8273_;
  assign new_n8276_ = ~new_n8274_ & ~new_n8275_;
  assign new_n8277_ = new_n6467_ & ~new_n8276_;
  assign new_n8278_ = ng3808 & ~new_n6467_;
  assign new_n8279_ = ~new_n8277_ & ~new_n8278_;
  assign new_n8280_ = pg35 & ~new_n8279_;
  assign n1829 = new_n8191_ | new_n8280_;
  assign new_n8282_ = ~pg35 & ng5360;
  assign new_n8283_ = ~new_n6368_ & ~new_n6371_;
  assign new_n8284_ = ~ng5373 & ~new_n8283_;
  assign new_n8285_ = ng5373 & new_n6394_;
  assign new_n8286_ = new_n8283_ & new_n8285_;
  assign new_n8287_ = ~new_n8284_ & ~new_n8286_;
  assign new_n8288_ = pg35 & ~new_n8287_;
  assign n1834 = new_n8282_ | new_n8288_;
  assign new_n8290_ = ~pg35 & ng1600;
  assign new_n8291_ = ~ng1668 & ng1636;
  assign new_n8292_ = ~new_n7537_1_ & new_n8291_;
  assign new_n8293_ = ng1608 & ~new_n8292_;
  assign new_n8294_ = ~new_n7543_ & new_n8292_;
  assign new_n8295_ = ~new_n8293_ & ~new_n8294_;
  assign new_n8296_ = pg35 & ~new_n8295_;
  assign n1839 = new_n8290_ | new_n8296_;
  assign new_n8298_ = ~pg35 & ng5527;
  assign new_n8299_ = ng5523 & ng5527;
  assign new_n8300_ = ~pg113 & new_n5781_1_;
  assign new_n8301_ = ~new_n4724_ & new_n8300_;
  assign new_n8302_ = ng43 & new_n8301_;
  assign new_n8303_ = ~ng5535 & ~new_n8302_;
  assign new_n8304_ = new_n8299_ & new_n8303_;
  assign new_n8305_ = ng5535 & ~new_n8302_;
  assign new_n8306_ = ~new_n8299_ & new_n8305_;
  assign new_n8307_ = ~new_n8304_ & ~new_n8306_;
  assign new_n8308_ = pg35 & ~new_n8307_;
  assign n1844 = new_n8298_ | new_n8308_;
  assign new_n8310_ = ~pg35 & ng392;
  assign new_n8311_ = ng405 & ~new_n6067_;
  assign new_n8312_ = ng392 & new_n6067_;
  assign new_n8313_ = ~new_n8311_ & ~new_n8312_;
  assign new_n8314_ = pg35 & ~new_n8313_;
  assign n1849 = new_n8310_ | new_n8314_;
  assign new_n8316_ = ~pg35 & ng209;
  assign new_n8317_ = pg35 & ~ng218;
  assign n1854 = new_n8316_ | new_n8317_;
  assign new_n8319_ = pg35 & ng5644;
  assign new_n8320_ = ~pg35 & new_n8319_;
  assign new_n8321_ = pg35 & ng5535;
  assign n1859 = new_n8320_ | new_n8321_;
  assign new_n8323_ = ~pg35 & ng3251;
  assign new_n8324_ = ng3167 & new_n5962_;
  assign new_n8325_ = ng3203 & ~new_n8324_;
  assign new_n8326_ = ~new_n5966_ & new_n8324_;
  assign new_n8327_ = ~new_n8325_ & ~new_n8326_;
  assign new_n8328_ = pg35 & ~new_n8327_;
  assign n1864 = new_n8323_ | new_n8328_;
  assign new_n8330_ = ~pg35 & ng650;
  assign new_n8331_ = ng655 & ~new_n7858_;
  assign new_n8332_ = ng650 & new_n7858_;
  assign new_n8333_ = ~new_n8331_ & ~new_n8332_;
  assign new_n8334_ = pg35 & ~new_n8333_;
  assign n1869 = new_n8330_ | new_n8334_;
  assign new_n8336_ = ~pg35 & ng4628;
  assign new_n8337_ = ng4639 & ng4621;
  assign new_n8338_ = ng4628 & new_n8337_;
  assign new_n8339_ = ~ng4643 & ~new_n5873_1_;
  assign new_n8340_ = ng4633 & new_n8339_;
  assign new_n8341_ = ~new_n8338_ & new_n8340_;
  assign new_n8342_ = ~ng4633 & new_n8339_;
  assign new_n8343_ = new_n8338_ & new_n8342_;
  assign new_n8344_ = ~new_n8341_ & ~new_n8343_;
  assign new_n8345_ = pg35 & ~new_n8344_;
  assign n1878 = new_n8336_ | new_n8345_;
  assign new_n8347_ = ~pg35 & ng4112;
  assign new_n8348_ = ng4116 & ~new_n7049_;
  assign new_n8349_ = ng4145 & new_n7049_;
  assign new_n8350_ = ~new_n8348_ & ~new_n8349_;
  assign new_n8351_ = pg35 & ~new_n8350_;
  assign n1883 = new_n8347_ | new_n8351_;
  assign new_n8353_ = ~pg35 & ng294;
  assign new_n8354_ = ng298 & new_n6021_;
  assign new_n8355_ = ~new_n6028_1_ & new_n8354_;
  assign new_n8356_ = ~ng298 & new_n6028_1_;
  assign new_n8357_ = ~new_n8355_ & ~new_n8356_;
  assign new_n8358_ = pg35 & ~new_n8357_;
  assign n1888 = new_n8353_ | new_n8358_;
  assign new_n8360_ = pg35 & ng933;
  assign new_n8361_ = ~pg35 & new_n8360_;
  assign new_n8362_ = ng1221 & ng1087;
  assign new_n8363_ = ng1205 & new_n8362_;
  assign new_n8364_ = ng1211 & new_n8363_;
  assign new_n8365_ = ~new_n7416_ & new_n8364_;
  assign new_n8366_ = ~ng1075 & ~ng1083;
  assign new_n8367_ = ~ng1079 & new_n8366_;
  assign new_n8368_ = ~new_n8365_ & new_n8367_;
  assign new_n8369_ = pg35 & new_n8368_;
  assign n1893 = new_n8361_ | new_n8369_;
  assign new_n8371_ = ~pg35 & ng4498;
  assign new_n8372_ = ~pg73 & pg72;
  assign new_n8373_ = ~ng4572 & new_n8372_;
  assign new_n8374_ = ng4581 & ~new_n8373_;
  assign new_n8375_ = ~ng4581 & ng4498;
  assign new_n8376_ = ~new_n8374_ & ~new_n8375_;
  assign new_n8377_ = pg35 & ~new_n8376_;
  assign n1897 = new_n8371_ | new_n8377_;
  assign new_n8379_ = ~pg35 & ng6509;
  assign new_n8380_ = ng6513 & ~new_n7390_;
  assign new_n8381_ = ~ng6513 & new_n7390_;
  assign new_n8382_ = ~new_n8380_ & ~new_n8381_;
  assign new_n8383_ = pg35 & ~new_n8382_;
  assign n1902 = new_n8379_ | new_n8383_;
  assign new_n8385_ = ~pg35 & ng3355;
  assign new_n8386_ = ng3361 & ~ng3355;
  assign new_n8387_ = ng3401 & ng3355;
  assign new_n8388_ = ~new_n8386_ & ~new_n8387_;
  assign new_n8389_ = ~ng3368 & ~new_n8388_;
  assign new_n8390_ = ~ng3385 & ng3396;
  assign new_n8391_ = ~ng3380 & new_n8390_;
  assign new_n8392_ = pg84 & new_n8391_;
  assign new_n8393_ = ng3361 & new_n8392_;
  assign new_n8394_ = ~ng3391 & ng3396;
  assign new_n8395_ = ~ng3385 & new_n8394_;
  assign new_n8396_ = ~pg84 & new_n8395_;
  assign new_n8397_ = ng3361 & new_n8396_;
  assign new_n8398_ = ~new_n8158_ & ~new_n8393_;
  assign new_n8399_ = ~new_n8162_ & ~new_n8397_;
  assign new_n8400_ = new_n8398_ & new_n8399_;
  assign new_n8401_ = ng3368 & new_n8400_;
  assign new_n8402_ = new_n8388_ & new_n8401_;
  assign new_n8403_ = ~new_n8389_ & ~new_n8402_;
  assign new_n8404_ = pg35 & ~new_n8403_;
  assign n1907 = new_n8385_ | new_n8404_;
  assign new_n8406_ = ~pg35 & ng5224;
  assign new_n8407_ = ~ng5188 & ~ng5180;
  assign new_n8408_ = new_n7581_ & new_n8407_;
  assign new_n8409_ = ng5240 & ~new_n8408_;
  assign new_n8410_ = ~new_n5966_ & new_n8408_;
  assign new_n8411_ = ~new_n8409_ & ~new_n8410_;
  assign new_n8412_ = pg35 & ~new_n8411_;
  assign n1912 = new_n8406_ | new_n8412_;
  assign new_n8414_ = ~pg35 & ng1008;
  assign new_n8415_ = ng1002 & new_n5940_1_;
  assign new_n8416_ = ~new_n5940_1_ & new_n6139_1_;
  assign new_n8417_ = ~new_n8415_ & ~new_n8416_;
  assign new_n8418_ = pg35 & ~new_n8417_;
  assign n1917 = new_n8414_ | new_n8418_;
  assign new_n8420_ = ~pg35 & ng862;
  assign new_n8421_ = ng862 & ~ng890;
  assign new_n8422_ = ~ng890 & ~new_n8421_;
  assign new_n8423_ = ng862 & ~new_n8421_;
  assign new_n8424_ = ~new_n8422_ & ~new_n8423_;
  assign new_n8425_ = pg35 & ~new_n8424_;
  assign n1922 = new_n8420_ | new_n8425_;
  assign new_n8427_ = ~pg35 & ng2841;
  assign new_n8428_ = ng2837 & ~ng2712;
  assign new_n8429_ = pg35 & new_n8428_;
  assign n1931 = new_n8427_ | new_n8429_;
  assign new_n8431_ = ~pg35 & ng5909;
  assign new_n8432_ = ng5881 & ng5873;
  assign new_n8433_ = new_n7650_ & new_n8432_;
  assign new_n8434_ = ng5929 & ~new_n8433_;
  assign new_n8435_ = ~new_n5966_ & new_n8433_;
  assign new_n8436_ = ~new_n8434_ & ~new_n8435_;
  assign new_n8437_ = pg35 & ~new_n8436_;
  assign n1936 = new_n8431_ | new_n8437_;
  assign new_n8439_ = pg35 & ng6682;
  assign new_n8440_ = ~pg35 & new_n8439_;
  assign new_n8441_ = pg35 & ng6573;
  assign n1941 = new_n8440_ | new_n8441_;
  assign new_n8443_ = ~pg35 & ng703;
  assign new_n8444_ = ng837 & ~new_n6067_;
  assign new_n8445_ = ng827 & ng832;
  assign new_n8446_ = ~ng812 & ~new_n8445_;
  assign new_n8447_ = ng837 & new_n8446_;
  assign new_n8448_ = ng703 & ng847;
  assign new_n8449_ = ~ng837 & new_n8448_;
  assign new_n8450_ = ~ng847 & ~new_n8445_;
  assign new_n8451_ = ng837 & new_n8450_;
  assign new_n8452_ = ~new_n8447_ & ~new_n8449_;
  assign new_n8453_ = ~new_n8451_ & new_n8452_;
  assign new_n8454_ = new_n6067_ & ~new_n8453_;
  assign new_n8455_ = ~new_n8444_ & ~new_n8454_;
  assign new_n8456_ = pg35 & ~new_n8455_;
  assign n1946 = new_n8443_ | new_n8456_;
  assign new_n8458_ = ~pg35 & ng2429;
  assign new_n8459_ = ~ng2495 & ng2465;
  assign new_n8460_ = ~new_n7555_ & new_n8459_;
  assign new_n8461_ = ng2437 & ~new_n8460_;
  assign new_n8462_ = ng4180 & new_n7550_;
  assign new_n8463_ = ~new_n7551_1_ & ~new_n8462_;
  assign new_n8464_ = ng1585 & new_n7551_1_;
  assign new_n8465_ = ~new_n8463_ & ~new_n8464_;
  assign new_n8466_ = new_n8460_ & ~new_n8465_;
  assign new_n8467_ = ~new_n8461_ & ~new_n8466_;
  assign new_n8468_ = pg35 & ~new_n8467_;
  assign n1951 = new_n8458_ | new_n8468_;
  assign new_n8470_ = ~pg35 & ng781;
  assign new_n8471_ = ~new_n6578_ & new_n6594_;
  assign new_n8472_ = ng781 & new_n8471_;
  assign new_n8473_ = ~ng785 & new_n8472_;
  assign new_n8474_ = ng785 & ~new_n6578_;
  assign new_n8475_ = ~new_n8472_ & new_n8474_;
  assign new_n8476_ = ~new_n8473_ & ~new_n8475_;
  assign new_n8477_ = pg35 & ~new_n8476_;
  assign n1965 = new_n8470_ | new_n8477_;
  assign new_n8479_ = ~pg35 & ng2579;
  assign new_n8480_ = ng2555 & ng2629;
  assign new_n8481_ = ~new_n7174_ & new_n8480_;
  assign new_n8482_ = ng2575 & ~new_n8481_;
  assign new_n8483_ = ~ng1585 & new_n7170_;
  assign new_n8484_ = ~new_n7494_ & ~new_n8483_;
  assign new_n8485_ = new_n8481_ & ~new_n8484_;
  assign new_n8486_ = ~new_n8482_ & ~new_n8485_;
  assign new_n8487_ = pg35 & ~new_n8486_;
  assign n1970 = new_n8479_ | new_n8487_;
  assign new_n8489_ = ~pg35 & ng3901;
  assign new_n8490_ = ng3857 & ~ng3863;
  assign new_n8491_ = new_n6874_ & new_n8490_;
  assign new_n8492_ = ng3925 & ~new_n8491_;
  assign new_n8493_ = ~new_n5966_ & new_n8491_;
  assign new_n8494_ = ~new_n8492_ & ~new_n8493_;
  assign new_n8495_ = pg35 & ~new_n8494_;
  assign n1980 = new_n8489_ | new_n8495_;
  assign new_n8497_ = ~pg35 & ng4771;
  assign new_n8498_ = new_n5667_ & new_n5838_1_;
  assign new_n8499_ = ~ng4809 & ~ng4818;
  assign new_n8500_ = ~new_n4724_ & new_n8499_;
  assign new_n8501_ = ~new_n8498_ & ~new_n8500_;
  assign new_n8502_ = ng4771 & ~new_n8500_;
  assign new_n8503_ = ng101 & new_n8500_;
  assign new_n8504_ = ~new_n8502_ & ~new_n8503_;
  assign new_n8505_ = ~new_n8501_ & ~new_n8504_;
  assign new_n8506_ = ng4765 & new_n8501_;
  assign new_n8507_ = ~new_n8505_ & ~new_n8506_;
  assign new_n8508_ = pg35 & ~new_n8507_;
  assign n1990 = new_n8497_ | new_n8508_;
  assign new_n8510_ = ~pg35 & ng1249;
  assign new_n8511_ = ng1570 & ng1249;
  assign new_n8512_ = ~ng1266 & new_n8511_;
  assign new_n8513_ = ng1570 & ng1266;
  assign new_n8514_ = ~new_n8511_ & new_n8513_;
  assign new_n8515_ = ~new_n8512_ & ~new_n8514_;
  assign new_n8516_ = pg35 & ~new_n8515_;
  assign n1995 = new_n8510_ | new_n8516_;
  assign new_n8518_ = ~pg35 & ng6649;
  assign new_n8519_ = ng6561 & new_n6334_;
  assign new_n8520_ = ng6605 & ~new_n8519_;
  assign new_n8521_ = ~new_n5966_ & new_n8519_;
  assign new_n8522_ = ~new_n8520_ & ~new_n8521_;
  assign new_n8523_ = pg35 & ~new_n8522_;
  assign n2000 = new_n8518_ | new_n8523_;
  assign new_n8525_ = ~pg35 & ng2988;
  assign new_n8526_ = ng12 & new_n4954_;
  assign new_n8527_ = n6079 & new_n8526_;
  assign new_n8528_ = ng2868 & ~new_n8526_;
  assign new_n8529_ = ~new_n8527_ & ~new_n8528_;
  assign new_n8530_ = pg35 & ~new_n8529_;
  assign n2005 = new_n8525_ | new_n8530_;
  assign new_n8532_ = ~pg35 & ng6565;
  assign new_n8533_ = ng6561 & ng6565;
  assign new_n8534_ = ~pg113 & new_n5795_;
  assign new_n8535_ = ~new_n4724_ & new_n8534_;
  assign new_n8536_ = ng43 & new_n8535_;
  assign new_n8537_ = ~ng6573 & ~new_n8536_;
  assign new_n8538_ = new_n8533_ & new_n8537_;
  assign new_n8539_ = ng6573 & ~new_n8536_;
  assign new_n8540_ = ~new_n8533_ & new_n8539_;
  assign new_n8541_ = ~new_n8538_ & ~new_n8540_;
  assign new_n8542_ = pg35 & ~new_n8541_;
  assign n2010 = new_n8532_ | new_n8542_;
  assign new_n8544_ = ~pg35 & ng5481;
  assign new_n8545_ = ng5689 & ng5703;
  assign new_n8546_ = ng5630 & new_n8545_;
  assign new_n8547_ = ng5644 & new_n8546_;
  assign new_n8548_ = new_n7745_ & new_n8547_;
  assign new_n8549_ = ng5485 & ~new_n8548_;
  assign new_n8550_ = ~ng5481 & ng5475;
  assign new_n8551_ = ng5475 & ~new_n8550_;
  assign new_n8552_ = ~ng5481 & ~new_n8550_;
  assign new_n8553_ = ~new_n8551_ & ~new_n8552_;
  assign new_n8554_ = new_n8548_ & ~new_n8553_;
  assign new_n8555_ = ~new_n8549_ & ~new_n8554_;
  assign new_n8556_ = pg35 & ~new_n8555_;
  assign n2015 = new_n8544_ | new_n8556_;
  assign new_n8558_ = ~pg35 & ng1216;
  assign new_n8559_ = ng1087 & ng1205;
  assign new_n8560_ = ng1221 & new_n8559_;
  assign new_n8561_ = ng1216 & new_n8560_;
  assign new_n8562_ = ng1211 & ~new_n8364_;
  assign new_n8563_ = ~new_n8561_ & new_n8562_;
  assign new_n8564_ = ~ng1211 & ~new_n8364_;
  assign new_n8565_ = new_n8561_ & new_n8564_;
  assign new_n8566_ = ~new_n8563_ & ~new_n8565_;
  assign new_n8567_ = pg35 & ~new_n8566_;
  assign n2020 = new_n8558_ | new_n8567_;
  assign new_n8569_ = ~pg35 & ng1816;
  assign new_n8570_ = ~ng1728 & ~ng1802;
  assign new_n8571_ = ~new_n6236_ & new_n8570_;
  assign new_n8572_ = ng1821 & ~new_n8571_;
  assign new_n8573_ = ng1816 & new_n8571_;
  assign new_n8574_ = ~new_n8572_ & ~new_n8573_;
  assign new_n8575_ = pg35 & ~new_n8574_;
  assign n2025 = new_n8569_ | new_n8575_;
  assign new_n8577_ = ~pg35 & ng5115;
  assign new_n8578_ = ng5124 & ~new_n6191_;
  assign new_n8579_ = ng5120 & ng5115;
  assign new_n8580_ = ng5120 & ~new_n8579_;
  assign new_n8581_ = ng5115 & ~new_n8579_;
  assign new_n8582_ = ~new_n8580_ & ~new_n8581_;
  assign new_n8583_ = new_n6191_ & ~new_n8582_;
  assign new_n8584_ = ~new_n8578_ & ~new_n8583_;
  assign new_n8585_ = pg35 & ~new_n8584_;
  assign n2030 = new_n8577_ | new_n8585_;
  assign new_n8587_ = ~pg35 & ng5373;
  assign new_n8588_ = ~new_n6369_ & ~new_n6372_1_;
  assign new_n8589_ = ng5377 & new_n6394_;
  assign new_n8590_ = new_n8588_ & new_n8589_;
  assign new_n8591_ = ~ng5377 & ~new_n8588_;
  assign new_n8592_ = ~new_n8590_ & ~new_n8591_;
  assign new_n8593_ = pg35 & ~new_n8592_;
  assign n2035 = new_n8587_ | new_n8593_;
  assign new_n8595_ = ~pg35 & ng6428;
  assign new_n8596_ = ~ng6428 & new_n6606_;
  assign new_n8597_ = ng6428 & new_n6611_;
  assign new_n8598_ = ~new_n8596_ & ~new_n8597_;
  assign new_n8599_ = ng6434 & new_n6632_1_;
  assign new_n8600_ = new_n8598_ & new_n8599_;
  assign new_n8601_ = ~ng6434 & ~new_n8598_;
  assign new_n8602_ = ~new_n8600_ & ~new_n8601_;
  assign new_n8603_ = pg35 & ~new_n8602_;
  assign n2040 = new_n8595_ | new_n8603_;
  assign new_n8605_ = pg35 & ng6199;
  assign new_n8606_ = ~pg35 & new_n8605_;
  assign new_n8607_ = ng6692 & ~ng6668;
  assign new_n8608_ = ng6668 & ~ng6661;
  assign new_n8609_ = ng6697 & ng6704;
  assign new_n8610_ = ng6675 & ng6661;
  assign new_n8611_ = new_n8609_ & new_n8610_;
  assign new_n8612_ = ~new_n8607_ & ~new_n8608_;
  assign new_n8613_ = ~new_n8611_ & new_n8612_;
  assign new_n8614_ = ~ng6675 & ng6704;
  assign new_n8615_ = ~ng6697 & ng6675;
  assign new_n8616_ = ~ng6704 & ng6661;
  assign new_n8617_ = new_n8613_ & ~new_n8614_;
  assign new_n8618_ = ~new_n8615_ & new_n8617_;
  assign new_n8619_ = ~new_n8616_ & new_n8618_;
  assign new_n8620_ = pg35 & new_n8619_;
  assign n2045 = new_n8606_ | new_n8620_;
  assign n2050 = ~pg35 & ng4931;
  assign new_n8623_ = ~pg35 & ng785;
  assign new_n8624_ = ~new_n6578_ & new_n8472_;
  assign new_n8625_ = ng785 & new_n8624_;
  assign new_n8626_ = ng790 & ~new_n6578_;
  assign new_n8627_ = ~new_n8625_ & new_n8626_;
  assign new_n8628_ = ~ng790 & new_n8625_;
  assign new_n8629_ = ~new_n8627_ & ~new_n8628_;
  assign new_n8630_ = pg35 & ~new_n8629_;
  assign n2060 = new_n8623_ | new_n8630_;
  assign new_n8632_ = ~pg35 & ng5138;
  assign new_n8633_ = ng5142 & ~new_n6191_;
  assign new_n8634_ = ~ng5142 & new_n6191_;
  assign new_n8635_ = ~new_n8633_ & ~new_n8634_;
  assign new_n8636_ = pg35 & ~new_n8635_;
  assign n2065 = new_n8632_ | new_n8636_;
  assign new_n8638_ = ~pg35 & ng3578;
  assign new_n8639_ = new_n6769_ & new_n7039_;
  assign new_n8640_ = ng3594 & ~new_n8639_;
  assign new_n8641_ = ~new_n5966_ & new_n8639_;
  assign new_n8642_ = ~new_n8640_ & ~new_n8641_;
  assign new_n8643_ = pg35 & ~new_n8642_;
  assign n2070 = new_n8638_ | new_n8643_;
  assign new_n8645_ = ~pg35 & ng5937;
  assign new_n8646_ = ng5857 & ng5863;
  assign new_n8647_ = new_n7649_ & new_n8646_;
  assign new_n8648_ = ng5953 & ~new_n8647_;
  assign new_n8649_ = ~new_n5966_ & new_n8647_;
  assign new_n8650_ = ~new_n8648_ & ~new_n8649_;
  assign new_n8651_ = pg35 & ~new_n8650_;
  assign n2075 = new_n8645_ | new_n8651_;
  assign new_n8653_ = ~pg35 & ng6555;
  assign new_n8654_ = ~ng6561 & ~new_n8536_;
  assign new_n8655_ = new_n7159_ & new_n8654_;
  assign new_n8656_ = ng6561 & new_n8654_;
  assign new_n8657_ = ~new_n7159_ & new_n8656_;
  assign new_n8658_ = ~new_n8655_ & ~new_n8657_;
  assign new_n8659_ = pg35 & ~new_n8658_;
  assign n2085 = new_n8653_ | new_n8659_;
  assign new_n8661_ = ~pg35 & ng2783;
  assign new_n8662_ = ng2724 & ~ng2729;
  assign new_n8663_ = new_n6041_1_ & new_n8662_;
  assign new_n8664_ = ng2775 & ~new_n8663_;
  assign new_n8665_ = ng85 & new_n5870_;
  assign new_n8666_ = ng2779 & ~new_n5870_;
  assign new_n8667_ = ~new_n8665_ & ~new_n8666_;
  assign new_n8668_ = new_n8663_ & new_n8667_;
  assign new_n8669_ = ~new_n8664_ & ~new_n8668_;
  assign new_n8670_ = pg35 & ~new_n8669_;
  assign n2090 = new_n8661_ | new_n8670_;
  assign new_n8672_ = pg35 & ng4616;
  assign new_n8673_ = ~pg35 & new_n8672_;
  assign new_n8674_ = ~ng4584 & ~ng4593;
  assign new_n8675_ = ng4608 & new_n8674_;
  assign new_n8676_ = ng4601 & ng4593;
  assign new_n8677_ = ng4601 & ~new_n8676_;
  assign new_n8678_ = ng4593 & ~new_n8676_;
  assign new_n8679_ = ~new_n8677_ & ~new_n8678_;
  assign new_n8680_ = ng4584 & ng4608;
  assign new_n8681_ = ng4584 & ~new_n8680_;
  assign new_n8682_ = ng4608 & ~new_n8680_;
  assign new_n8683_ = ~new_n8681_ & ~new_n8682_;
  assign new_n8684_ = new_n8679_ & new_n8683_;
  assign new_n8685_ = ~ng4616 & new_n8684_;
  assign new_n8686_ = ng4584 & ng4593;
  assign new_n8687_ = ~ng4601 & ~ng4608;
  assign new_n8688_ = new_n8686_ & new_n8687_;
  assign new_n8689_ = ~new_n8675_ & ~new_n8685_;
  assign new_n8690_ = ~new_n8688_ & new_n8689_;
  assign new_n8691_ = ~pg135 & ~new_n8690_;
  assign new_n8692_ = ng4633 & new_n5861_;
  assign new_n8693_ = new_n5864_ & new_n8692_;
  assign new_n8694_ = new_n8691_ & new_n8693_;
  assign new_n8695_ = pg35 & ~new_n8694_;
  assign n2095 = new_n8673_ | new_n8695_;
  assign new_n8697_ = ~pg35 & ng5022;
  assign new_n8698_ = ~ng5022 & ~ng5062;
  assign new_n8699_ = ng5016 & new_n8698_;
  assign new_n8700_ = ~ng5016 & new_n8107_;
  assign new_n8701_ = ~new_n8698_ & new_n8700_;
  assign new_n8702_ = ~new_n8699_ & ~new_n8701_;
  assign new_n8703_ = pg35 & ~new_n8702_;
  assign n2100 = new_n8697_ | new_n8703_;
  assign new_n8705_ = ~pg35 & ng5124;
  assign new_n8706_ = ng5128 & ~pg26801;
  assign new_n8707_ = ~ng5128 & pg26801;
  assign new_n8708_ = ~new_n8706_ & ~new_n8707_;
  assign new_n8709_ = pg35 & ~new_n8708_;
  assign n2110 = new_n8705_ | new_n8709_;
  assign new_n8711_ = ~pg35 & ng3759;
  assign new_n8712_ = ~new_n6093_ & ~new_n6101_1_;
  assign new_n8713_ = pg35 & new_n8712_;
  assign n2115 = new_n8711_ | new_n8713_;
  assign new_n8715_ = ~pg35 & ng4646;
  assign new_n8716_ = new_n4734_ & new_n7604_;
  assign new_n8717_ = ng4646 & ~new_n8716_;
  assign new_n8718_ = pg35 & new_n8717_;
  assign n2124 = new_n8715_ | new_n8718_;
  assign new_n8720_ = ~pg35 & ng4122;
  assign new_n8721_ = ~pg124 & ng4146;
  assign new_n8722_ = pg126 & ~ng4146;
  assign new_n8723_ = ~new_n8721_ & ~new_n8722_;
  assign new_n8724_ = ~new_n7731_ & new_n8723_;
  assign new_n8725_ = ~new_n7731_ & ~new_n8724_;
  assign new_n8726_ = new_n8723_ & ~new_n8724_;
  assign new_n8727_ = ~new_n8725_ & ~new_n8726_;
  assign new_n8728_ = pg116 & ng4157;
  assign new_n8729_ = pg114 & ~ng4157;
  assign new_n8730_ = ~new_n8728_ & ~new_n8729_;
  assign new_n8731_ = ~pg116 & ng4157;
  assign new_n8732_ = pg115 & ~ng4157;
  assign new_n8733_ = ~new_n8731_ & ~new_n8732_;
  assign new_n8734_ = ~new_n8730_ & new_n8733_;
  assign new_n8735_ = ~new_n8730_ & ~new_n8734_;
  assign new_n8736_ = new_n8733_ & ~new_n8734_;
  assign new_n8737_ = ~new_n8735_ & ~new_n8736_;
  assign new_n8738_ = new_n8727_ & new_n8737_;
  assign new_n8739_ = pg35 & ~new_n8738_;
  assign n2129 = new_n8720_ | new_n8739_;
  assign new_n8741_ = ~pg35 & ng2834;
  assign n2134 = new_n7357_ | new_n8741_;
  assign new_n8743_ = ~pg35 & ng3223;
  assign new_n8744_ = ~ng3171 & ng3179;
  assign new_n8745_ = new_n5963_ & new_n8744_;
  assign new_n8746_ = ng3239 & ~new_n8745_;
  assign new_n8747_ = ~new_n5966_ & new_n8745_;
  assign new_n8748_ = ~new_n8746_ & ~new_n8747_;
  assign new_n8749_ = pg35 & ~new_n8748_;
  assign n2139 = new_n8743_ | new_n8749_;
  assign new_n8751_ = ~pg35 & ng1442;
  assign new_n8752_ = ng1437 & ~new_n7471_;
  assign new_n8753_ = ng1478 & new_n6436_;
  assign new_n8754_ = ng1478 & ~new_n8753_;
  assign new_n8755_ = new_n6436_ & ~new_n8753_;
  assign new_n8756_ = ~new_n8754_ & ~new_n8755_;
  assign new_n8757_ = ng1437 & ~new_n8756_;
  assign new_n8758_ = ~new_n6435_1_ & new_n8757_;
  assign new_n8759_ = new_n6435_1_ & ~new_n8756_;
  assign new_n8760_ = ~new_n8758_ & ~new_n8759_;
  assign new_n8761_ = new_n7471_ & ~new_n8760_;
  assign new_n8762_ = ~new_n8752_ & ~new_n8761_;
  assign new_n8763_ = pg35 & ~new_n8762_;
  assign n2144 = new_n8751_ | new_n8763_;
  assign new_n8765_ = pg35 & ng4575;
  assign new_n8766_ = ~pg35 & new_n8765_;
  assign new_n8767_ = pg113 & pg35;
  assign n2149 = new_n8766_ | new_n8767_;
  assign new_n8769_ = ng22 & pg34915;
  assign new_n8770_ = ~ng22 & n2272;
  assign n2153 = new_n8769_ | new_n8770_;
  assign new_n8772_ = ~pg35 & ng4264;
  assign new_n8773_ = ng4264 & ng4258;
  assign new_n8774_ = ng4269 & ~new_n8773_;
  assign new_n8775_ = ~ng4269 & new_n8773_;
  assign new_n8776_ = ~new_n8774_ & ~new_n8775_;
  assign new_n8777_ = pg35 & ~new_n8776_;
  assign n2158 = new_n8772_ | new_n8777_;
  assign new_n8779_ = ~pg35 & ng3338;
  assign new_n8780_ = ng3310 & ng3303;
  assign new_n8781_ = ng3281 & ng3267;
  assign new_n8782_ = new_n8780_ & new_n8781_;
  assign new_n8783_ = ng3338 & new_n8782_;
  assign new_n8784_ = ~ng3347 & ~new_n8783_;
  assign new_n8785_ = pg35 & new_n8784_;
  assign n2163 = new_n8779_ | new_n8785_;
  assign new_n8787_ = ~pg35 & ng2827;
  assign new_n8788_ = ng2724 & ng2729;
  assign new_n8789_ = new_n6041_1_ & new_n8788_;
  assign new_n8790_ = ng2819 & ~new_n8789_;
  assign new_n8791_ = ng2827 & ~new_n5870_;
  assign new_n8792_ = ~new_n6045_1_ & ~new_n8791_;
  assign new_n8793_ = new_n8789_ & new_n8792_;
  assign new_n8794_ = ~new_n8790_ & ~new_n8793_;
  assign new_n8795_ = pg35 & ~new_n8794_;
  assign n2168 = new_n8787_ | new_n8795_;
  assign new_n8797_ = ~pg35 & ng3100;
  assign new_n8798_ = ~ng3100 & ng3092;
  assign new_n8799_ = ~ng3050 & ~new_n8798_;
  assign new_n8800_ = ~ng3096 & ~new_n8799_;
  assign new_n8801_ = pg35 & new_n8800_;
  assign n2173 = new_n8797_ | new_n8801_;
  assign new_n8803_ = ~pg35 & ng4480;
  assign new_n8804_ = ~ng4572 & new_n7110_;
  assign new_n8805_ = ng4581 & ~new_n8804_;
  assign new_n8806_ = ~ng4581 & ng4480;
  assign new_n8807_ = ~new_n8805_ & ~new_n8806_;
  assign new_n8808_ = pg35 & ~new_n8807_;
  assign n2178 = new_n8803_ | new_n8808_;
  assign new_n8810_ = ~pg35 & ng1199;
  assign new_n8811_ = ng1157 & new_n5950_1_;
  assign new_n8812_ = ~new_n5935_1_ & new_n8811_;
  assign new_n8813_ = ng1199 & new_n8812_;
  assign new_n8814_ = ng1070 & new_n5953_;
  assign new_n8815_ = ~new_n8813_ & new_n8814_;
  assign new_n8816_ = ~ng1070 & new_n5953_;
  assign new_n8817_ = new_n8813_ & new_n8816_;
  assign new_n8818_ = ~new_n8815_ & ~new_n8817_;
  assign new_n8819_ = pg35 & ~new_n8818_;
  assign n2183 = new_n8810_ | new_n8819_;
  assign new_n8821_ = ~pg35 & ng6299;
  assign new_n8822_ = ng6215 & new_n7865_;
  assign new_n8823_ = ng6251 & ~new_n8822_;
  assign new_n8824_ = ~new_n5966_ & new_n8822_;
  assign new_n8825_ = ~new_n8823_ & ~new_n8824_;
  assign new_n8826_ = pg35 & ~new_n8825_;
  assign n2192 = new_n8821_ | new_n8826_;
  assign new_n8828_ = ~pg35 & ng1296;
  assign new_n8829_ = ng12 & new_n4919_;
  assign new_n8830_ = n5005 & new_n8829_;
  assign new_n8831_ = ~ng1283 & ~ng1277;
  assign new_n8832_ = ~new_n8830_ & ~new_n8831_;
  assign new_n8833_ = pg35 & new_n8832_;
  assign n2197 = new_n8828_ | new_n8833_;
  assign new_n8835_ = ~pg35 & ng6533;
  assign new_n8836_ = ng6537 & ~new_n7390_;
  assign new_n8837_ = ~ng6533 & ng6527;
  assign new_n8838_ = ng6527 & ~new_n8837_;
  assign new_n8839_ = ~ng6533 & ~new_n8837_;
  assign new_n8840_ = ~new_n8838_ & ~new_n8839_;
  assign new_n8841_ = new_n7390_ & ~new_n8840_;
  assign new_n8842_ = ~new_n8836_ & ~new_n8841_;
  assign new_n8843_ = pg35 & ~new_n8842_;
  assign n2202 = new_n8835_ | new_n8843_;
  assign new_n8845_ = ~pg35 & ng4308;
  assign new_n8846_ = pg35 & ~new_n5925_1_;
  assign n2207 = new_n8845_ | new_n8846_;
  assign new_n8848_ = ~pg35 & ng4332;
  assign new_n8849_ = new_n5865_ & new_n5869_;
  assign new_n8850_ = ng4616 & new_n5869_;
  assign new_n8851_ = ng4584 & new_n5865_;
  assign new_n8852_ = new_n8850_ & new_n8851_;
  assign new_n8853_ = ~new_n5873_1_ & ~new_n8852_;
  assign new_n8854_ = ~ng4584 & new_n8853_;
  assign new_n8855_ = new_n8849_ & new_n8854_;
  assign new_n8856_ = ng4584 & new_n8853_;
  assign new_n8857_ = ~new_n8849_ & new_n8856_;
  assign new_n8858_ = ~new_n8855_ & ~new_n8857_;
  assign new_n8859_ = pg35 & ~new_n8858_;
  assign n2212 = new_n8848_ | new_n8859_;
  assign new_n8861_ = ~pg35 & ng5752;
  assign new_n8862_ = pg35 & ng6035;
  assign n2222 = new_n8861_ | new_n8862_;
  assign new_n8864_ = ~pg35 & ng2980;
  assign new_n8865_ = new_n4945_1_ & new_n6820_;
  assign new_n8866_ = ~pg56 & ~pg54;
  assign new_n8867_ = ~pg53 & new_n8866_;
  assign new_n8868_ = n3854 & new_n8867_;
  assign new_n8869_ = ~ng2984 & ~new_n8868_;
  assign new_n8870_ = ~new_n8865_ & ~new_n8869_;
  assign new_n8871_ = pg35 & new_n8870_;
  assign n2232 = new_n8864_ | new_n8871_;
  assign new_n8873_ = pg35 & ng1277;
  assign new_n8874_ = ~pg35 & new_n8873_;
  assign new_n8875_ = ng1564 & ng1430;
  assign new_n8876_ = ng1548 & new_n8875_;
  assign new_n8877_ = ng1554 & new_n8876_;
  assign new_n8878_ = ~ng1312 & ~new_n6294_;
  assign new_n8879_ = new_n6299_ & new_n8878_;
  assign new_n8880_ = new_n8877_ & ~new_n8879_;
  assign new_n8881_ = ~ng1418 & ~ng1426;
  assign new_n8882_ = ~ng1422 & new_n8881_;
  assign new_n8883_ = ~new_n8880_ & new_n8882_;
  assign new_n8884_ = pg35 & new_n8883_;
  assign n2237 = new_n8874_ | new_n8884_;
  assign new_n8886_ = ~pg35 & ng1252;
  assign new_n8887_ = ng1266 & new_n8511_;
  assign new_n8888_ = ng1280 & new_n8887_;
  assign new_n8889_ = ng1252 & new_n8888_;
  assign new_n8890_ = ng1570 & ng1256;
  assign new_n8891_ = ~new_n8889_ & new_n8890_;
  assign new_n8892_ = ~ng1256 & new_n8889_;
  assign new_n8893_ = ~new_n8891_ & ~new_n8892_;
  assign new_n8894_ = pg35 & ~new_n8893_;
  assign n2242 = new_n8886_ | new_n8894_;
  assign new_n8896_ = ~pg35 & ng2837;
  assign new_n8897_ = pg35 & ng2837;
  assign n2247 = new_n8896_ | new_n8897_;
  assign new_n8899_ = ~pg35 & ng2311;
  assign new_n8900_ = ng2361 & ng2287;
  assign new_n8901_ = ~new_n7886_ & new_n8900_;
  assign new_n8902_ = ng2307 & ~new_n8901_;
  assign new_n8903_ = ng4180 & new_n7881_;
  assign new_n8904_ = ~new_n7882_ & ~new_n8903_;
  assign new_n8905_ = ~ng1585 & new_n7882_;
  assign new_n8906_ = ~new_n8904_ & ~new_n8905_;
  assign new_n8907_ = new_n8901_ & ~new_n8906_;
  assign new_n8908_ = ~new_n8902_ & ~new_n8907_;
  assign new_n8909_ = pg35 & ~new_n8908_;
  assign n2252 = new_n8899_ | new_n8909_;
  assign new_n8911_ = ~pg35 & ng5747;
  assign new_n8912_ = ~new_n6409_ & ~new_n6417_;
  assign new_n8913_ = pg35 & new_n8912_;
  assign n2257 = new_n8911_ | new_n8913_;
  assign new_n8915_ = ~pg35 & ng3706;
  assign new_n8916_ = ~new_n6074_1_ & ~new_n6079_1_;
  assign new_n8917_ = ~ng3719 & ~new_n8916_;
  assign new_n8918_ = ng3719 & new_n6104_;
  assign new_n8919_ = new_n8916_ & new_n8918_;
  assign new_n8920_ = ~new_n8917_ & ~new_n8919_;
  assign new_n8921_ = pg35 & ~new_n8920_;
  assign n2262 = new_n8915_ | new_n8921_;
  assign new_n8923_ = ~pg35 & ng5406;
  assign new_n8924_ = pg35 & ng5689;
  assign n2267 = new_n8923_ | new_n8924_;
  assign new_n8926_ = ~pg35 & ng3025;
  assign new_n8927_ = ng3010 & ~ng3004;
  assign new_n8928_ = ~ng3017 & new_n8927_;
  assign new_n8929_ = ~ng3021 & new_n8928_;
  assign new_n8930_ = ~ng3025 & new_n8929_;
  assign new_n8931_ = ng3050 & ng3004;
  assign new_n8932_ = ng3017 & new_n8931_;
  assign new_n8933_ = ng3021 & new_n8932_;
  assign new_n8934_ = ng3025 & new_n8933_;
  assign new_n8935_ = ~new_n8930_ & ~new_n8934_;
  assign new_n8936_ = ng3045 & ~ng3034;
  assign new_n8937_ = ~ng3029 & new_n8936_;
  assign new_n8938_ = pg84 & new_n8937_;
  assign new_n8939_ = ng3010 & new_n8938_;
  assign new_n8940_ = ~ng3045 & ng3034;
  assign new_n8941_ = ng3029 & new_n8940_;
  assign new_n8942_ = pg84 & new_n8941_;
  assign new_n8943_ = ng3050 & new_n8942_;
  assign new_n8944_ = ng3045 & ~ng3040;
  assign new_n8945_ = ~ng3034 & new_n8944_;
  assign new_n8946_ = ~pg84 & new_n8945_;
  assign new_n8947_ = ng3010 & new_n8946_;
  assign new_n8948_ = ~ng3045 & ng3040;
  assign new_n8949_ = ng3034 & new_n8948_;
  assign new_n8950_ = ~pg84 & new_n8949_;
  assign new_n8951_ = ng3050 & new_n8950_;
  assign new_n8952_ = ~new_n8939_ & ~new_n8943_;
  assign new_n8953_ = ~new_n8947_ & ~new_n8951_;
  assign new_n8954_ = new_n8952_ & new_n8953_;
  assign new_n8955_ = ng3029 & new_n8954_;
  assign new_n8956_ = new_n8935_ & new_n8955_;
  assign new_n8957_ = ~ng3029 & ~new_n8935_;
  assign new_n8958_ = ~new_n8956_ & ~new_n8957_;
  assign new_n8959_ = pg35 & ~new_n8958_;
  assign n2277 = new_n8926_ | new_n8959_;
  assign new_n8961_ = ~pg35 & ng4456;
  assign new_n8962_ = pg35 & ng4456;
  assign n2282 = new_n8961_ | new_n8962_;
  assign new_n8964_ = ~pg35 & ng5441;
  assign new_n8965_ = ng5428 & ng5436;
  assign new_n8966_ = ng5441 & new_n8965_;
  assign new_n8967_ = ~ng5445 & new_n8966_;
  assign new_n8968_ = ng5445 & ~new_n8966_;
  assign new_n8969_ = ~new_n8967_ & ~new_n8968_;
  assign new_n8970_ = pg35 & ~new_n8969_;
  assign n2292 = new_n8964_ | new_n8970_;
  assign new_n8972_ = pg35 & ng4933;
  assign new_n8973_ = ~pg35 & new_n8972_;
  assign new_n8974_ = new_n5676_ & new_n5746_;
  assign new_n8975_ = ~ng3694 & ~ng3639;
  assign new_n8976_ = ~ng3703 & new_n8975_;
  assign new_n8977_ = ng3694 & ng3639;
  assign new_n8978_ = ~ng3703 & new_n8977_;
  assign new_n8979_ = ~ng3639 & ~ng3698;
  assign new_n8980_ = ng3703 & new_n8979_;
  assign new_n8981_ = ng3639 & ng3698;
  assign new_n8982_ = ng3703 & new_n8981_;
  assign new_n8983_ = ~new_n8976_ & ~new_n8978_;
  assign new_n8984_ = ~new_n8980_ & ~new_n8982_;
  assign new_n8985_ = new_n8983_ & new_n8984_;
  assign new_n8986_ = ~ng4950 & new_n8985_;
  assign new_n8987_ = new_n8974_ & ~new_n8986_;
  assign new_n8988_ = new_n7431_ & new_n8987_;
  assign new_n8989_ = ng4950 & ~new_n7431_;
  assign new_n8990_ = ~new_n8988_ & ~new_n8989_;
  assign new_n8991_ = pg35 & ~new_n8990_;
  assign n2302 = new_n8973_ | new_n8991_;
  assign new_n8993_ = ~pg35 & ng5220;
  assign new_n8994_ = ~ng5170 & ~ng5164;
  assign new_n8995_ = ~ng5176 & new_n8994_;
  assign new_n8996_ = new_n5053_ & new_n8995_;
  assign new_n8997_ = ng5216 & ~new_n8996_;
  assign new_n8998_ = ~new_n5966_ & new_n8996_;
  assign new_n8999_ = ~new_n8997_ & ~new_n8998_;
  assign new_n9000_ = pg35 & ~new_n8999_;
  assign n2307 = new_n8993_ | new_n9000_;
  assign n2312 = ~pg35 & ng2704;
  assign new_n9003_ = ~pg35 & ng1906;
  assign new_n9004_ = ~new_n4724_ & new_n5642_;
  assign new_n9005_ = ~pg113 & new_n9004_;
  assign new_n9006_ = ng112 & new_n9005_;
  assign new_n9007_ = ng1906 & ~new_n9006_;
  assign new_n9008_ = ~new_n6667_1_ & new_n9007_;
  assign new_n9009_ = ng1936 & new_n6667_1_;
  assign new_n9010_ = ~new_n9008_ & ~new_n9009_;
  assign new_n9011_ = pg35 & ~new_n9010_;
  assign n2317 = new_n9003_ | new_n9011_;
  assign new_n9013_ = ~pg35 & ng1636;
  assign new_n9014_ = ~new_n4724_ & new_n5639_;
  assign new_n9015_ = ~pg113 & new_n9014_;
  assign new_n9016_ = ng112 & new_n9015_;
  assign new_n9017_ = ng1636 & ~new_n9016_;
  assign new_n9018_ = ~new_n7537_1_ & new_n9017_;
  assign new_n9019_ = ng1668 & new_n7537_1_;
  assign new_n9020_ = ~new_n9018_ & ~new_n9019_;
  assign new_n9021_ = pg35 & ~new_n9020_;
  assign n2322 = new_n9013_ | new_n9021_;
  assign new_n9023_ = ~pg35 & ng3680;
  assign new_n9024_ = ng3661 & ng3654;
  assign new_n9025_ = ng3632 & ng3618;
  assign new_n9026_ = new_n9024_ & new_n9025_;
  assign new_n9027_ = ng3689 & ~new_n9026_;
  assign new_n9028_ = ~ng3689 & new_n9026_;
  assign new_n9029_ = ~new_n9027_ & ~new_n9028_;
  assign new_n9030_ = pg35 & ~new_n9029_;
  assign n2332 = new_n9023_ | new_n9030_;
  assign new_n9032_ = ~pg35 & ng4176;
  assign new_n9033_ = n5005 & new_n5972_;
  assign new_n9034_ = ng4146 & ~new_n5972_;
  assign new_n9035_ = ~new_n9033_ & ~new_n9034_;
  assign new_n9036_ = pg35 & ~new_n9035_;
  assign n2337 = new_n9032_ | new_n9036_;
  assign new_n9038_ = ~pg35 & ng4674;
  assign new_n9039_ = ng4674 & ~new_n8716_;
  assign new_n9040_ = pg35 & new_n9039_;
  assign n2342 = new_n9038_ | new_n9040_;
  assign new_n9042_ = ~pg35 & ng3770;
  assign new_n9043_ = ng3767 & ~ng3759;
  assign new_n9044_ = ~ng3770 & ~new_n9043_;
  assign new_n9045_ = ~ng3774 & new_n9044_;
  assign new_n9046_ = ng3774 & ng3770;
  assign new_n9047_ = ng3767 & ~ng3763;
  assign new_n9048_ = ~new_n9045_ & ~new_n9046_;
  assign new_n9049_ = ~new_n9047_ & new_n9048_;
  assign new_n9050_ = pg35 & ~new_n9049_;
  assign n2347 = new_n9042_ | new_n9050_;
  assign new_n9052_ = ~pg35 & ng822;
  assign new_n9053_ = ng822 & new_n8006_;
  assign new_n9054_ = ng827 & new_n8009_;
  assign new_n9055_ = ~new_n9053_ & new_n9054_;
  assign new_n9056_ = ~ng827 & new_n8009_;
  assign new_n9057_ = new_n9053_ & new_n9056_;
  assign new_n9058_ = ~new_n9055_ & ~new_n9057_;
  assign new_n9059_ = pg35 & ~new_n9058_;
  assign n2352 = new_n9052_ | new_n9059_;
  assign new_n9061_ = ~pg35 & ng283;
  assign new_n9062_ = ~ng287 & new_n6022_;
  assign new_n9063_ = ng287 & new_n6021_;
  assign new_n9064_ = ~new_n6022_ & new_n9063_;
  assign new_n9065_ = ~new_n9062_ & ~new_n9064_;
  assign new_n9066_ = pg35 & ~new_n9065_;
  assign n2357 = new_n9061_ | new_n9066_;
  assign new_n9068_ = ~pg35 & ng1274;
  assign new_n9069_ = ng1256 & new_n8889_;
  assign new_n9070_ = ng1259 & new_n9069_;
  assign new_n9071_ = ng1263 & new_n9070_;
  assign new_n9072_ = ng1270 & new_n9071_;
  assign new_n9073_ = ng1274 & new_n9072_;
  assign new_n9074_ = ~new_n4689_ & new_n9073_;
  assign new_n9075_ = pg35 & new_n9074_;
  assign n2362 = new_n9068_ | new_n9075_;
  assign new_n9077_ = ~pg35 & ng121;
  assign new_n9078_ = ~ng2193 & new_n7642_;
  assign new_n9079_ = ~ng2799 & ~new_n9078_;
  assign new_n9080_ = ~new_n7640_ & ~new_n9079_;
  assign new_n9081_ = pg35 & new_n9080_;
  assign n2367 = new_n9077_ | new_n9081_;
  assign new_n9083_ = ~pg35 & ng1926;
  assign new_n9084_ = ~ng1917 & ng1894;
  assign new_n9085_ = ng1886 & new_n9084_;
  assign new_n9086_ = ~ng1926 & ~ng1894;
  assign new_n9087_ = ng1882 & new_n9086_;
  assign new_n9088_ = ng1890 & new_n5204_;
  assign new_n9089_ = ~new_n9085_ & ~new_n9087_;
  assign new_n9090_ = ~new_n9088_ & new_n9089_;
  assign new_n9091_ = ng1917 & ~ng1894;
  assign new_n9092_ = ng1870 & new_n9091_;
  assign new_n9093_ = ng1874 & new_n8167_;
  assign new_n9094_ = ng1926 & ~ng1917;
  assign new_n9095_ = ng1878 & new_n9094_;
  assign new_n9096_ = new_n9090_ & ~new_n9092_;
  assign new_n9097_ = ~new_n9093_ & ~new_n9095_;
  assign new_n9098_ = new_n9096_ & new_n9097_;
  assign new_n9099_ = new_n8171_ & ~new_n9098_;
  assign new_n9100_ = ng1945 & ~new_n8171_;
  assign new_n9101_ = ~new_n9099_ & ~new_n9100_;
  assign new_n9102_ = pg35 & ~new_n9101_;
  assign n2372 = new_n9083_ | new_n9102_;
  assign new_n9104_ = ~pg35 & ng772;
  assign new_n9105_ = ~ng776 & new_n6592_;
  assign new_n9106_ = ng776 & ~new_n6578_;
  assign new_n9107_ = ~new_n6592_ & new_n9106_;
  assign new_n9108_ = ~new_n9105_ & ~new_n9107_;
  assign new_n9109_ = pg35 & ~new_n9108_;
  assign n2377 = new_n9104_ | new_n9109_;
  assign n2386 = ~pg35 & ng943;
  assign new_n9112_ = ~pg35 & ng622;
  assign new_n9113_ = ~new_n6545_ & new_n6568_;
  assign new_n9114_ = ng599 & new_n9113_;
  assign new_n9115_ = ~new_n6545_ & new_n9114_;
  assign new_n9116_ = ng604 & new_n9115_;
  assign new_n9117_ = ~new_n6545_ & new_n9116_;
  assign new_n9118_ = ng608 & new_n9117_;
  assign new_n9119_ = ~new_n6545_ & new_n9118_;
  assign new_n9120_ = ng613 & new_n9119_;
  assign new_n9121_ = ~new_n6545_ & new_n9120_;
  assign new_n9122_ = ng617 & new_n9121_;
  assign new_n9123_ = ~new_n6545_ & new_n9122_;
  assign new_n9124_ = ng622 & new_n9123_;
  assign new_n9125_ = ~ng626 & new_n9124_;
  assign new_n9126_ = ng626 & ~new_n6545_;
  assign new_n9127_ = ~new_n9124_ & new_n9126_;
  assign new_n9128_ = ~new_n9125_ & ~new_n9127_;
  assign new_n9129_ = pg35 & ~new_n9128_;
  assign n2391 = new_n9112_ | new_n9129_;
  assign new_n9131_ = ~pg35 & ng4643;
  assign new_n9132_ = ~new_n5862_ & ~new_n5873_1_;
  assign new_n9133_ = ng4340 & ~new_n5873_1_;
  assign new_n9134_ = ~new_n9132_ & ~new_n9133_;
  assign new_n9135_ = ng4340 & new_n9132_;
  assign new_n9136_ = ~new_n9134_ & ~new_n9135_;
  assign new_n9137_ = pg35 & ~new_n9136_;
  assign n2396 = new_n9131_ | new_n9137_;
  assign new_n9139_ = ~pg35 & ng2016;
  assign new_n9140_ = ~ng2787 & new_n5902_1_;
  assign new_n9141_ = new_n5904_ & ~new_n9140_;
  assign new_n9142_ = ng2715 & ~new_n9141_;
  assign new_n9143_ = ng2719 & new_n9142_;
  assign new_n9144_ = new_n5208_ & new_n9143_;
  assign new_n9145_ = ng2036 & ~new_n9144_;
  assign new_n9146_ = ~ng1996 & ng2040;
  assign new_n9147_ = new_n9144_ & ~new_n9146_;
  assign new_n9148_ = ~new_n9145_ & ~new_n9147_;
  assign new_n9149_ = pg35 & ~new_n9148_;
  assign n2401 = new_n9139_ | new_n9149_;
  assign new_n9151_ = pg35 & ng218;
  assign new_n9152_ = ~pg35 & new_n9151_;
  assign new_n9153_ = ~ng1570 & new_n8511_;
  assign new_n9154_ = ng1570 & ~ng1249;
  assign new_n9155_ = ~new_n9153_ & ~new_n9154_;
  assign new_n9156_ = pg35 & ~new_n9155_;
  assign n2406 = new_n9152_ | new_n9156_;
  assign new_n9158_ = ~pg35 & ng2098;
  assign new_n9159_ = ng2060 & ng2028;
  assign new_n9160_ = new_n9143_ & new_n9159_;
  assign new_n9161_ = ng2102 & ~new_n9160_;
  assign new_n9162_ = ~ng2102 & new_n9160_;
  assign new_n9163_ = ~new_n9161_ & ~new_n9162_;
  assign new_n9164_ = pg35 & ~new_n9163_;
  assign n2411 = new_n9158_ | new_n9164_;
  assign new_n9166_ = ~pg35 & ng6167;
  assign new_n9167_ = ng6173 & ~new_n6700_;
  assign new_n9168_ = ng6167 & new_n6700_;
  assign new_n9169_ = ~new_n9167_ & ~new_n9168_;
  assign new_n9170_ = pg35 & ~new_n9169_;
  assign n2416 = new_n9166_ | new_n9170_;
  assign new_n9172_ = ~pg35 & ng2287;
  assign new_n9173_ = ~pg113 & new_n5654_;
  assign new_n9174_ = ~new_n4724_ & new_n9173_;
  assign new_n9175_ = new_n7885_ & new_n9174_;
  assign new_n9176_ = ng2361 & ~ng2331;
  assign new_n9177_ = ng112 & new_n9176_;
  assign new_n9178_ = ng112 & ~new_n9177_;
  assign new_n9179_ = new_n9176_ & ~new_n9177_;
  assign new_n9180_ = ~new_n9178_ & ~new_n9179_;
  assign new_n9181_ = new_n9175_ & ~new_n9180_;
  assign new_n9182_ = ng2338 & ~new_n9175_;
  assign new_n9183_ = ~new_n9181_ & ~new_n9182_;
  assign new_n9184_ = pg35 & ~new_n9183_;
  assign n2421 = new_n9172_ | new_n9184_;
  assign new_n9186_ = ~pg35 & ng6736;
  assign new_n9187_ = new_n4739_ & new_n7747_;
  assign new_n9188_ = new_n7218_1_ & new_n9187_;
  assign new_n9189_ = new_n4735_ & new_n9188_;
  assign new_n9190_ = ~ng6741 & ~new_n9189_;
  assign new_n9191_ = new_n7218_1_ & new_n9190_;
  assign new_n9192_ = ng6741 & ~new_n7218_1_;
  assign new_n9193_ = ~new_n9191_ & ~new_n9192_;
  assign new_n9194_ = pg35 & ~new_n9193_;
  assign n2426 = new_n9186_ | new_n9194_;
  assign new_n9196_ = new_n5055_ & pg33874;
  assign new_n9197_ = ng66 & ~new_n5055_;
  assign n2431 = new_n9196_ | new_n9197_;
  assign new_n9199_ = ~pg35 & ng6500;
  assign new_n9200_ = ng6509 & ~new_n7219_;
  assign new_n9201_ = ng6500 & ng6505;
  assign new_n9202_ = ng6505 & ~new_n9201_;
  assign new_n9203_ = ng6500 & ~new_n9201_;
  assign new_n9204_ = ~new_n9202_ & ~new_n9203_;
  assign new_n9205_ = new_n7219_ & ~new_n9204_;
  assign new_n9206_ = ~new_n9200_ & ~new_n9205_;
  assign new_n9207_ = pg35 & ~new_n9206_;
  assign n2441 = new_n9199_ | new_n9207_;
  assign new_n9209_ = ~pg35 & ng2040;
  assign new_n9210_ = ~new_n4724_ & new_n5646_;
  assign new_n9211_ = ~pg113 & new_n9210_;
  assign new_n9212_ = ng112 & new_n9211_;
  assign new_n9213_ = ng2040 & ~new_n9212_;
  assign new_n9214_ = ~new_n7025_ & new_n9213_;
  assign new_n9215_ = ng2070 & new_n7025_;
  assign new_n9216_ = ~new_n9214_ & ~new_n9215_;
  assign new_n9217_ = pg35 & ~new_n9216_;
  assign n2446 = new_n9209_ | new_n9217_;
  assign new_n9219_ = ~pg35 & ng5567;
  assign new_n9220_ = new_n6885_ & new_n8035_;
  assign new_n9221_ = ng5563 & ~new_n9220_;
  assign new_n9222_ = ~new_n5966_ & new_n9220_;
  assign new_n9223_ = ~new_n9221_ & ~new_n9222_;
  assign new_n9224_ = pg35 & ~new_n9223_;
  assign n2451 = new_n9219_ | new_n9224_;
  assign new_n9226_ = ~pg35 & ng4369;
  assign new_n9227_ = ng4473 & ~ng4462;
  assign new_n9228_ = ~ng4507 & ~new_n4724_;
  assign new_n9229_ = ~pg73 & ~new_n9228_;
  assign new_n9230_ = ~pg72 & new_n9229_;
  assign new_n9231_ = ng4474 & ~new_n9230_;
  assign new_n9232_ = ~ng4477 & new_n9231_;
  assign new_n9233_ = ~ng4459 & ~new_n9227_;
  assign new_n9234_ = ~new_n9232_ & new_n9233_;
  assign new_n9235_ = pg35 & ~new_n9234_;
  assign n2456 = new_n9226_ | new_n9235_;
  assign new_n9237_ = ~pg35 & ng2449;
  assign new_n9238_ = ~ng2421 & ng2465;
  assign new_n9239_ = ~new_n7555_ & new_n9238_;
  assign new_n9240_ = ng2445 & ~new_n9239_;
  assign new_n9241_ = ~new_n8465_ & new_n9239_;
  assign new_n9242_ = ~new_n9240_ & ~new_n9241_;
  assign new_n9243_ = pg35 & ~new_n9242_;
  assign n2461 = new_n9237_ | new_n9243_;
  assign new_n9245_ = ~pg35 & ng2403;
  assign new_n9246_ = ng2407 & ~new_n7888_;
  assign new_n9247_ = ~ng2407 & new_n7888_;
  assign new_n9248_ = ~new_n9246_ & ~new_n9247_;
  assign new_n9249_ = pg35 & ~new_n9248_;
  assign n2466 = new_n9245_ | new_n9249_;
  assign new_n9251_ = ~pg35 & ng1657;
  assign new_n9252_ = ng1624 & ~ng1648;
  assign new_n9253_ = ng1616 & new_n9252_;
  assign new_n9254_ = ~ng1624 & ~ng1657;
  assign new_n9255_ = ng1612 & new_n9254_;
  assign new_n9256_ = ng1620 & pg25167;
  assign new_n9257_ = ~new_n9253_ & ~new_n9255_;
  assign new_n9258_ = ~new_n9256_ & new_n9257_;
  assign new_n9259_ = ~ng1624 & ng1648;
  assign new_n9260_ = ng1600 & new_n9259_;
  assign new_n9261_ = ng1604 & new_n7226_;
  assign new_n9262_ = ng1657 & ~ng1648;
  assign new_n9263_ = ng1608 & new_n9262_;
  assign new_n9264_ = new_n9258_ & ~new_n9260_;
  assign new_n9265_ = ~new_n9261_ & ~new_n9263_;
  assign new_n9266_ = new_n9264_ & new_n9265_;
  assign new_n9267_ = new_n7230_ & ~new_n9266_;
  assign new_n9268_ = ng1677 & ~new_n7230_;
  assign new_n9269_ = ~new_n9267_ & ~new_n9268_;
  assign new_n9270_ = pg35 & ~new_n9269_;
  assign n2471 = new_n9251_ | new_n9270_;
  assign new_n9272_ = ~pg35 & ng5097;
  assign new_n9273_ = ng5092 & ng5084;
  assign new_n9274_ = ng5097 & new_n9273_;
  assign new_n9275_ = ~ng86 & new_n9274_;
  assign new_n9276_ = ng86 & ~new_n9274_;
  assign new_n9277_ = ~new_n9275_ & ~new_n9276_;
  assign new_n9278_ = pg35 & ~new_n9277_;
  assign n2476 = new_n9272_ | new_n9278_;
  assign new_n9280_ = ~pg35 & ng2823;
  assign new_n9281_ = ~ng2595 & new_n7642_;
  assign new_n9282_ = ~ng2827 & ~new_n9281_;
  assign new_n9283_ = ~new_n7640_ & ~new_n9282_;
  assign new_n9284_ = pg35 & new_n9283_;
  assign n2481 = new_n9280_ | new_n9284_;
  assign new_n9286_ = ~pg35 & ng6439;
  assign new_n9287_ = ~new_n6617_ & ~new_n6625_;
  assign new_n9288_ = pg35 & new_n9287_;
  assign n2486 = new_n9286_ | new_n9288_;
  assign new_n9290_ = ~pg35 & ng1521;
  assign new_n9291_ = ng1500 & new_n7195_;
  assign new_n9292_ = ng1306 & ~new_n9291_;
  assign new_n9293_ = ng1339 & new_n9291_;
  assign new_n9294_ = ~new_n9292_ & ~new_n9293_;
  assign new_n9295_ = pg35 & ~new_n9294_;
  assign n2495 = new_n9290_ | new_n9295_;
  assign new_n9297_ = pg35 & ng1322;
  assign new_n9298_ = ~pg35 & new_n9297_;
  assign new_n9299_ = ng1514 & new_n6843_;
  assign new_n9300_ = ng1500 & ~new_n9299_;
  assign new_n9301_ = ~ng1514 & new_n6843_;
  assign new_n9302_ = ~ng1500 & ~new_n9301_;
  assign new_n9303_ = ~new_n9300_ & ~new_n9302_;
  assign new_n9304_ = pg35 & ~new_n9303_;
  assign n2500 = new_n9298_ | new_n9304_;
  assign new_n9306_ = pg35 & ng4669;
  assign new_n9307_ = ~pg35 & new_n9306_;
  assign new_n9308_ = ng12 & new_n4924_;
  assign new_n9309_ = ng4727 & ~new_n9308_;
  assign new_n9310_ = n4955 & new_n9308_;
  assign new_n9311_ = ~new_n9309_ & ~new_n9310_;
  assign new_n9312_ = pg35 & ~new_n9311_;
  assign n2505 = new_n9307_ | new_n9312_;
  assign new_n9314_ = ~pg35 & ng3191;
  assign new_n9315_ = ~ng3161 & ng3155;
  assign new_n9316_ = new_n5962_ & new_n9315_;
  assign new_n9317_ = ng3219 & ~new_n9316_;
  assign new_n9318_ = ~new_n5966_ & new_n9316_;
  assign new_n9319_ = ~new_n9317_ & ~new_n9318_;
  assign new_n9320_ = pg35 & ~new_n9319_;
  assign n2510 = new_n9314_ | new_n9320_;
  assign new_n9322_ = ~pg35 & ng6645;
  assign new_n9323_ = ng6561 & new_n7456_;
  assign new_n9324_ = ng6597 & ~new_n9323_;
  assign new_n9325_ = ~new_n5966_ & new_n9323_;
  assign new_n9326_ = ~new_n9324_ & ~new_n9325_;
  assign new_n9327_ = pg35 & ~new_n9326_;
  assign n2515 = new_n9322_ | new_n9327_;
  assign new_n9329_ = ~pg35 & ng5957;
  assign new_n9330_ = ng5881 & ~ng5873;
  assign new_n9331_ = ng5869 & new_n9330_;
  assign new_n9332_ = ng5913 & ~new_n9331_;
  assign new_n9333_ = ~new_n5966_ & new_n9331_;
  assign new_n9334_ = ~new_n9332_ & ~new_n9333_;
  assign new_n9335_ = pg35 & ~new_n9334_;
  assign n2520 = new_n9329_ | new_n9335_;
  assign new_n9337_ = ~pg35 & ng3243;
  assign new_n9338_ = ng3161 & ng3155;
  assign new_n9339_ = new_n7151_ & new_n9338_;
  assign new_n9340_ = ng3259 & ~new_n9339_;
  assign new_n9341_ = ~new_n5966_ & new_n9339_;
  assign new_n9342_ = ~new_n9340_ & ~new_n9341_;
  assign new_n9343_ = pg35 & ~new_n9342_;
  assign n2525 = new_n9337_ | new_n9343_;
  assign new_n9345_ = pg35 & ng117;
  assign new_n9346_ = ~pg35 & new_n9345_;
  assign new_n9347_ = ng12 & n3583;
  assign new_n9348_ = new_n4954_ & new_n9347_;
  assign new_n9349_ = ~ng2932 & ~ng2999;
  assign new_n9350_ = ~new_n9348_ & ~new_n9349_;
  assign new_n9351_ = pg35 & new_n9350_;
  assign n2530 = new_n9346_ | new_n9351_;
  assign new_n9353_ = ~pg35 & ng2421;
  assign new_n9354_ = ~pg113 & new_n5653_1_;
  assign new_n9355_ = ~new_n4724_ & new_n9354_;
  assign new_n9356_ = new_n7554_ & new_n9355_;
  assign new_n9357_ = ng2495 & ~ng2465;
  assign new_n9358_ = ng112 & new_n9357_;
  assign new_n9359_ = ng112 & ~new_n9358_;
  assign new_n9360_ = new_n9357_ & ~new_n9358_;
  assign new_n9361_ = ~new_n9359_ & ~new_n9360_;
  assign new_n9362_ = new_n9356_ & ~new_n9361_;
  assign new_n9363_ = ng2472 & ~new_n9356_;
  assign new_n9364_ = ~new_n9362_ & ~new_n9363_;
  assign new_n9365_ = pg35 & ~new_n9364_;
  assign n2535 = new_n9353_ | new_n9365_;
  assign new_n9367_ = ~pg35 & ng3247;
  assign new_n9368_ = ~ng3171 & ~ng3179;
  assign new_n9369_ = ng3167 & new_n9368_;
  assign new_n9370_ = ng3195 & ~new_n9369_;
  assign new_n9371_ = ~new_n5966_ & new_n9369_;
  assign new_n9372_ = ~new_n9370_ & ~new_n9371_;
  assign new_n9373_ = pg35 & ~new_n9372_;
  assign n2540 = new_n9367_ | new_n9373_;
  assign new_n9375_ = ~pg35 & ng4382;
  assign new_n9376_ = pg35 & new_n5870_;
  assign n2545 = new_n9375_ | new_n9376_;
  assign new_n9378_ = ~pg35 & ng2912;
  assign new_n9379_ = ng12 & new_n4942_;
  assign new_n9380_ = n5814 & new_n9379_;
  assign new_n9381_ = ng2922 & ~new_n9379_;
  assign new_n9382_ = ~new_n9380_ & ~new_n9381_;
  assign new_n9383_ = pg35 & ~new_n9382_;
  assign n2550 = new_n9378_ | new_n9383_;
  assign new_n9385_ = ~pg35 & ng3451;
  assign new_n9386_ = ng3443 & ~ng3451;
  assign new_n9387_ = ~ng3401 & ~new_n9386_;
  assign new_n9388_ = ~ng3447 & ~new_n9387_;
  assign new_n9389_ = pg35 & new_n9388_;
  assign n2555 = new_n9385_ | new_n9389_;
  assign new_n9391_ = ~pg35 & ng3115;
  assign new_n9392_ = ng3119 & ~new_n7152_;
  assign new_n9393_ = ~ng3119 & new_n7152_;
  assign new_n9394_ = ~new_n9392_ & ~new_n9393_;
  assign new_n9395_ = pg35 & ~new_n9394_;
  assign n2560 = new_n9391_ | new_n9395_;
  assign new_n9397_ = ~pg35 & ng3255;
  assign new_n9398_ = ng3167 & new_n8744_;
  assign new_n9399_ = ng3211 & ~new_n9398_;
  assign new_n9400_ = ~new_n5966_ & new_n9398_;
  assign new_n9401_ = ~new_n9399_ & ~new_n9400_;
  assign new_n9402_ = pg35 & ~new_n9401_;
  assign n2565 = new_n9397_ | new_n9402_;
  assign new_n9404_ = ~pg35 & ng3817;
  assign new_n9405_ = ng3821 & ~new_n7011_1_;
  assign new_n9406_ = ~ng3821 & new_n7011_1_;
  assign new_n9407_ = ~new_n9405_ & ~new_n9406_;
  assign new_n9408_ = pg35 & ~new_n9407_;
  assign n2570 = new_n9404_ | new_n9408_;
  assign new_n9410_ = ~pg35 & ng3195;
  assign new_n9411_ = ~ng3161 & ~ng3155;
  assign new_n9412_ = ~ng3167 & new_n9411_;
  assign new_n9413_ = new_n5962_ & new_n9412_;
  assign new_n9414_ = ng3191 & ~new_n9413_;
  assign new_n9415_ = ~new_n5966_ & new_n9413_;
  assign new_n9416_ = ~new_n9414_ & ~new_n9415_;
  assign new_n9417_ = pg35 & ~new_n9416_;
  assign n2575 = new_n9410_ | new_n9417_;
  assign new_n9419_ = ~pg35 & ng2523;
  assign new_n9420_ = ng2485 & ng2453;
  assign new_n9421_ = new_n5907_1_ & new_n9420_;
  assign new_n9422_ = ng2527 & ~new_n9421_;
  assign new_n9423_ = ~ng2527 & new_n9421_;
  assign new_n9424_ = ~new_n9422_ & ~new_n9423_;
  assign new_n9425_ = pg35 & ~new_n9424_;
  assign n2580 = new_n9419_ | new_n9425_;
  assign new_n9427_ = ~pg35 & ng3227;
  assign new_n9428_ = new_n5963_ & new_n7151_;
  assign new_n9429_ = ng3243 & ~new_n9428_;
  assign new_n9430_ = ~new_n5966_ & new_n9428_;
  assign new_n9431_ = ~new_n9429_ & ~new_n9430_;
  assign new_n9432_ = pg35 & ~new_n9431_;
  assign n2585 = new_n9427_ | new_n9432_;
  assign new_n9434_ = ~pg35 & ng5256;
  assign new_n9435_ = ng5176 & new_n8407_;
  assign new_n9436_ = ng5204 & ~new_n9435_;
  assign new_n9437_ = ~new_n5966_ & new_n9435_;
  assign new_n9438_ = ~new_n9436_ & ~new_n9437_;
  assign new_n9439_ = pg35 & ~new_n9438_;
  assign n2590 = new_n9434_ | new_n9439_;
  assign new_n9441_ = pg35 & ng1858;
  assign new_n9442_ = ~pg35 & new_n9441_;
  assign new_n9443_ = ~ng1936 & ng1862;
  assign new_n9444_ = ~ng1936 & ~ng1906;
  assign new_n9445_ = ~new_n9443_ & ~new_n9444_;
  assign new_n9446_ = ~new_n9006_ & ~new_n9445_;
  assign new_n9447_ = ~new_n6667_1_ & new_n9446_;
  assign new_n9448_ = ng1862 & new_n6667_1_;
  assign new_n9449_ = ~new_n9447_ & ~new_n9448_;
  assign new_n9450_ = pg35 & ~new_n9449_;
  assign n2595 = new_n9442_ | new_n9450_;
  assign new_n9452_ = ~pg35 & ng6052;
  assign new_n9453_ = ng6058 & ~ng6052;
  assign new_n9454_ = ng6052 & ng6098;
  assign new_n9455_ = ~new_n9453_ & ~new_n9454_;
  assign new_n9456_ = ~ng6065 & ~new_n9455_;
  assign new_n9457_ = ng6065 & new_n7527_;
  assign new_n9458_ = new_n9455_ & new_n9457_;
  assign new_n9459_ = ~new_n9456_ & ~new_n9458_;
  assign new_n9460_ = pg35 & ~new_n9459_;
  assign n2600 = new_n9452_ | new_n9460_;
  assign new_n9462_ = ~pg35 & ng1183;
  assign new_n9463_ = ng1157 & ng996;
  assign new_n9464_ = ~ng1157 & ng1178;
  assign new_n9465_ = ~new_n9463_ & ~new_n9464_;
  assign new_n9466_ = pg35 & ~new_n9465_;
  assign n2605 = new_n9462_ | new_n9466_;
  assign new_n9468_ = ~pg35 & ng3522;
  assign new_n9469_ = ng3518 & ng3522;
  assign new_n9470_ = ~pg113 & new_n5800_;
  assign new_n9471_ = ~new_n4724_ & new_n9470_;
  assign new_n9472_ = ng43 & new_n9471_;
  assign new_n9473_ = ~ng3530 & ~new_n9472_;
  assign new_n9474_ = new_n9469_ & new_n9473_;
  assign new_n9475_ = ng3530 & ~new_n9472_;
  assign new_n9476_ = ~new_n9469_ & new_n9475_;
  assign new_n9477_ = ~new_n9474_ & ~new_n9476_;
  assign new_n9478_ = pg35 & ~new_n9477_;
  assign n2614 = new_n9468_ | new_n9478_;
  assign new_n9480_ = ~pg35 & ng4269;
  assign new_n9481_ = ng4269 & new_n8773_;
  assign new_n9482_ = ~ng4273 & new_n9481_;
  assign new_n9483_ = ng4273 & ~new_n9481_;
  assign new_n9484_ = ~new_n9482_ & ~new_n9483_;
  assign new_n9485_ = pg35 & ~new_n9484_;
  assign n2619 = new_n9480_ | new_n9485_;
  assign new_n9487_ = pg35 & ng4932;
  assign new_n9488_ = ~pg35 & new_n9487_;
  assign new_n9489_ = ~ng4871 & ~ng4836;
  assign new_n9490_ = ~ng4864 & new_n9489_;
  assign new_n9491_ = ~ng4878 & new_n9490_;
  assign new_n9492_ = ~ng4966 & new_n5675_;
  assign new_n9493_ = ng4991 & ng4983;
  assign new_n9494_ = ~ng4966 & new_n9493_;
  assign new_n9495_ = ~new_n9492_ & ~new_n9494_;
  assign new_n9496_ = ~new_n5751_ & ~new_n9495_;
  assign new_n9497_ = ng4912 & new_n5742_1_;
  assign new_n9498_ = ng4922 & new_n5744_;
  assign new_n9499_ = ng4907 & new_n5746_;
  assign new_n9500_ = ng4917 & new_n5674_;
  assign new_n9501_ = ~new_n9497_ & ~new_n9498_;
  assign new_n9502_ = ~new_n9499_ & ~new_n9500_;
  assign new_n9503_ = new_n9501_ & new_n9502_;
  assign new_n9504_ = ~new_n5751_ & ~new_n9503_;
  assign new_n9505_ = ~new_n9503_ & ~new_n9504_;
  assign new_n9506_ = ~new_n5751_ & ~new_n9504_;
  assign new_n9507_ = ~new_n9505_ & ~new_n9506_;
  assign new_n9508_ = new_n6462_ & ~new_n9507_;
  assign new_n9509_ = ~ng4966 & new_n6461_;
  assign new_n9510_ = ~ng4927 & new_n5674_;
  assign new_n9511_ = ~new_n5744_ & ~new_n5746_;
  assign new_n9512_ = ~new_n9510_ & new_n9511_;
  assign new_n9513_ = new_n9509_ & ~new_n9512_;
  assign new_n9514_ = ~new_n5676_ & ~new_n9496_;
  assign new_n9515_ = ~new_n9508_ & ~new_n9513_;
  assign new_n9516_ = new_n9514_ & new_n9515_;
  assign new_n9517_ = new_n9491_ & ~new_n9516_;
  assign new_n9518_ = ng4836 & ng5011;
  assign new_n9519_ = ng4871 & ng3684;
  assign new_n9520_ = ~ng3333 & ng4864;
  assign new_n9521_ = ~ng4035 & ng4878;
  assign new_n9522_ = ~new_n9518_ & ~new_n9519_;
  assign new_n9523_ = ~new_n9520_ & ~new_n9521_;
  assign new_n9524_ = new_n9522_ & new_n9523_;
  assign new_n9525_ = ~new_n9491_ & ~new_n9524_;
  assign new_n9526_ = ~new_n9517_ & ~new_n9525_;
  assign new_n9527_ = pg35 & ~new_n9526_;
  assign n2624 = new_n9488_ | new_n9527_;
  assign new_n9529_ = ~pg35 & ng2255;
  assign new_n9530_ = ng2185 & ng2217;
  assign new_n9531_ = ~ng2803 & new_n5902_1_;
  assign new_n9532_ = new_n5904_ & ~new_n9531_;
  assign new_n9533_ = ~ng2715 & ~new_n9532_;
  assign new_n9534_ = ~ng2719 & new_n9533_;
  assign new_n9535_ = new_n9530_ & new_n9534_;
  assign new_n9536_ = ng2259 & ~new_n9535_;
  assign new_n9537_ = ~ng2259 & new_n9535_;
  assign new_n9538_ = ~new_n9536_ & ~new_n9537_;
  assign new_n9539_ = pg35 & ~new_n9538_;
  assign n2629 = new_n9529_ | new_n9539_;
  assign new_n9541_ = ~pg35 & ng6187;
  assign new_n9542_ = ng6191 & ~new_n7064_;
  assign new_n9543_ = ng6181 & ~ng6187;
  assign new_n9544_ = ng6181 & ~new_n9543_;
  assign new_n9545_ = ~ng6187 & ~new_n9543_;
  assign new_n9546_ = ~new_n9544_ & ~new_n9545_;
  assign new_n9547_ = new_n7064_ & ~new_n9546_;
  assign new_n9548_ = ~new_n9542_ & ~new_n9547_;
  assign new_n9549_ = pg35 & ~new_n9548_;
  assign n2634 = new_n9541_ | new_n9549_;
  assign new_n9551_ = ~pg35 & ng6291;
  assign new_n9552_ = new_n5849_ & new_n7063_;
  assign new_n9553_ = ng6307 & ~new_n9552_;
  assign new_n9554_ = ~new_n5966_ & new_n9552_;
  assign new_n9555_ = ~new_n9553_ & ~new_n9554_;
  assign new_n9556_ = pg35 & ~new_n9555_;
  assign n2639 = new_n9551_ | new_n9556_;
  assign new_n9558_ = pg35 & ng2932;
  assign new_n9559_ = ~pg35 & new_n9558_;
  assign new_n9560_ = ~ng4639 & new_n8339_;
  assign new_n9561_ = pg35 & new_n9560_;
  assign n2649 = new_n9559_ | new_n9561_;
  assign new_n9563_ = ~pg35 & ng5033;
  assign new_n9564_ = ~new_n8138_ & ~new_n8143_;
  assign new_n9565_ = ~ng5037 & ~new_n9564_;
  assign new_n9566_ = ng5037 & new_n8107_;
  assign new_n9567_ = new_n9564_ & new_n9566_;
  assign new_n9568_ = ~new_n9565_ & ~new_n9567_;
  assign new_n9569_ = pg35 & ~new_n9568_;
  assign n2654 = new_n9563_ | new_n9569_;
  assign new_n9571_ = ~pg35 & ng6263;
  assign new_n9572_ = ~ng6227 & ~ng6219;
  assign new_n9573_ = ng6209 & ~ng6203;
  assign new_n9574_ = new_n9572_ & new_n9573_;
  assign new_n9575_ = ng6279 & ~new_n9574_;
  assign new_n9576_ = ~new_n5966_ & new_n9574_;
  assign new_n9577_ = ~new_n9575_ & ~new_n9576_;
  assign new_n9578_ = pg35 & ~new_n9577_;
  assign n2659 = new_n9571_ | new_n9578_;
  assign new_n9580_ = ~pg35 & ng457;
  assign new_n9581_ = ng471 & ~new_n5994_;
  assign new_n9582_ = ng269 & new_n5994_;
  assign new_n9583_ = ~new_n9581_ & ~new_n9582_;
  assign new_n9584_ = pg35 & ~new_n9583_;
  assign n2664 = new_n9580_ | new_n9584_;
  assign new_n9586_ = ~pg35 & ng5357;
  assign new_n9587_ = ng5357 & pg33959;
  assign new_n9588_ = pg33959 & new_n9187_;
  assign new_n9589_ = new_n4734_ & new_n9588_;
  assign new_n9590_ = ng5297 & ~new_n9589_;
  assign new_n9591_ = ~new_n9587_ & new_n9590_;
  assign new_n9592_ = ~ng5297 & ~new_n9589_;
  assign new_n9593_ = new_n9587_ & new_n9592_;
  assign new_n9594_ = ~new_n9591_ & ~new_n9593_;
  assign new_n9595_ = pg35 & ~new_n9594_;
  assign n2669 = new_n9586_ | new_n9595_;
  assign new_n9597_ = ~pg35 & ng255;
  assign new_n9598_ = ng875 & new_n6112_;
  assign new_n9599_ = ng232 & ~new_n6112_;
  assign new_n9600_ = ~new_n9598_ & ~new_n9599_;
  assign new_n9601_ = pg35 & ~new_n9600_;
  assign n2678 = new_n9597_ | new_n9601_;
  assign new_n9603_ = ~pg35 & ng3747;
  assign new_n9604_ = ~new_n6089_ & ~new_n6097_;
  assign new_n9605_ = pg35 & new_n9604_;
  assign n2683 = new_n9603_ | new_n9605_;
  assign new_n9607_ = pg35 & ng3684;
  assign new_n9608_ = ~pg35 & new_n9607_;
  assign new_n9609_ = ng3498 & ~new_n6770_;
  assign new_n9610_ = ~new_n5966_ & new_n9609_;
  assign new_n9611_ = new_n9609_ & ~new_n9610_;
  assign new_n9612_ = ~new_n5966_ & ~new_n9610_;
  assign new_n9613_ = ~new_n9611_ & ~new_n9612_;
  assign new_n9614_ = pg35 & ~new_n9613_;
  assign n2688 = new_n9608_ | new_n9614_;
  assign new_n9616_ = ~pg35 & ng6549;
  assign new_n9617_ = ng6555 & ~new_n8536_;
  assign new_n9618_ = ~ng6549 & new_n9617_;
  assign new_n9619_ = ~ng6555 & ~new_n8536_;
  assign new_n9620_ = ng6549 & new_n9619_;
  assign new_n9621_ = ~new_n9618_ & ~new_n9620_;
  assign new_n9622_ = pg35 & ~new_n9621_;
  assign n2693 = new_n9616_ | new_n9622_;
  assign new_n9624_ = ~pg35 & ng1467;
  assign new_n9625_ = new_n7196_ & new_n7472_;
  assign new_n9626_ = ng1467 & ng1472;
  assign new_n9627_ = ng1472 & ~new_n9626_;
  assign new_n9628_ = ng1467 & ~new_n9626_;
  assign new_n9629_ = ~new_n9627_ & ~new_n9628_;
  assign new_n9630_ = new_n9625_ & ~new_n9629_;
  assign new_n9631_ = ng1472 & ~new_n9625_;
  assign new_n9632_ = ~new_n9630_ & ~new_n9631_;
  assign new_n9633_ = pg35 & ~new_n9632_;
  assign n2698 = new_n9624_ | new_n9633_;
  assign new_n9635_ = pg35 & ng4743;
  assign new_n9636_ = ~pg35 & new_n9635_;
  assign new_n9637_ = new_n5667_ & new_n5840_;
  assign new_n9638_ = ~ng5990 & ~ng6040;
  assign new_n9639_ = ~ng6049 & new_n9638_;
  assign new_n9640_ = ng5990 & ng6040;
  assign new_n9641_ = ~ng6049 & new_n9640_;
  assign new_n9642_ = ~ng6044 & ~ng5990;
  assign new_n9643_ = ng6049 & new_n9642_;
  assign new_n9644_ = ng6044 & ng5990;
  assign new_n9645_ = ng6049 & new_n9644_;
  assign new_n9646_ = ~new_n9639_ & ~new_n9641_;
  assign new_n9647_ = ~new_n9643_ & ~new_n9645_;
  assign new_n9648_ = new_n9646_ & new_n9647_;
  assign new_n9649_ = ~ng4760 & new_n9648_;
  assign new_n9650_ = new_n9637_ & ~new_n9649_;
  assign new_n9651_ = new_n6353_ & new_n9650_;
  assign new_n9652_ = ng4760 & ~new_n6353_;
  assign new_n9653_ = ~new_n9651_ & ~new_n9652_;
  assign new_n9654_ = pg35 & ~new_n9653_;
  assign n2703 = new_n9636_ | new_n9654_;
  assign new_n9656_ = ~pg35 & ng2153;
  assign new_n9657_ = ~pg113 & new_n5652_;
  assign new_n9658_ = ~new_n4724_ & new_n9657_;
  assign new_n9659_ = new_n6521_ & new_n9658_;
  assign new_n9660_ = ~ng2197 & ng2227;
  assign new_n9661_ = ng112 & new_n9660_;
  assign new_n9662_ = ng112 & ~new_n9661_;
  assign new_n9663_ = new_n9660_ & ~new_n9661_;
  assign new_n9664_ = ~new_n9662_ & ~new_n9663_;
  assign new_n9665_ = new_n9659_ & ~new_n9664_;
  assign new_n9666_ = ng2204 & ~new_n9659_;
  assign new_n9667_ = ~new_n9665_ & ~new_n9666_;
  assign new_n9668_ = pg35 & ~new_n9667_;
  assign n2708 = new_n9656_ | new_n9668_;
  assign new_n9670_ = ~pg35 & ng890;
  assign new_n9671_ = ng896 & ~ng890;
  assign new_n9672_ = ~ng896 & ng862;
  assign new_n9673_ = ~new_n9671_ & ~new_n9672_;
  assign new_n9674_ = pg35 & ~new_n9673_;
  assign n2713 = new_n9670_ | new_n9674_;
  assign new_n9676_ = ~pg35 & ng6732;
  assign new_n9677_ = ng6727 & new_n8611_;
  assign new_n9678_ = ng6732 & ~new_n9677_;
  assign new_n9679_ = pg35 & new_n9678_;
  assign n2718 = new_n9676_ | new_n9679_;
  assign new_n9681_ = ~pg35 & ng6505;
  assign new_n9682_ = ng6500 & ~new_n7213_1_;
  assign new_n9683_ = ~ng6741 & ~ng6682;
  assign new_n9684_ = ~ng6727 & new_n9683_;
  assign new_n9685_ = ng6715 & ng6633;
  assign new_n9686_ = new_n9684_ & new_n9685_;
  assign new_n9687_ = ~ng6741 & ng6682;
  assign new_n9688_ = ~ng6727 & new_n9687_;
  assign new_n9689_ = ng6605 & ng6723;
  assign new_n9690_ = new_n9688_ & new_n9689_;
  assign new_n9691_ = ng6741 & ~ng6682;
  assign new_n9692_ = ~ng6727 & new_n9691_;
  assign new_n9693_ = ng6649 & ng6719;
  assign new_n9694_ = new_n9692_ & new_n9693_;
  assign new_n9695_ = ~ng6727 & new_n4759_;
  assign new_n9696_ = ng6697 & ng6601;
  assign new_n9697_ = new_n9695_ & new_n9696_;
  assign new_n9698_ = ~new_n9686_ & ~new_n9690_;
  assign new_n9699_ = ~new_n9694_ & ~new_n9697_;
  assign new_n9700_ = new_n9698_ & new_n9699_;
  assign new_n9701_ = ng6727 & new_n9683_;
  assign new_n9702_ = ng6589 & ng6723;
  assign new_n9703_ = new_n9701_ & new_n9702_;
  assign new_n9704_ = ng6697 & ng6727;
  assign new_n9705_ = ng6697 & ~new_n9704_;
  assign new_n9706_ = ng6727 & ~new_n9704_;
  assign new_n9707_ = ~new_n9705_ & ~new_n9706_;
  assign new_n9708_ = new_n9687_ & new_n9707_;
  assign new_n9709_ = ng6613 & ng6675;
  assign new_n9710_ = new_n9708_ & new_n9709_;
  assign new_n9711_ = ng6727 & new_n9691_;
  assign new_n9712_ = ng6697 & ng6585;
  assign new_n9713_ = new_n9711_ & new_n9712_;
  assign new_n9714_ = new_n4759_ & new_n9707_;
  assign new_n9715_ = ng6704 & ng6629;
  assign new_n9716_ = new_n9714_ & new_n9715_;
  assign new_n9717_ = ~new_n9703_ & ~new_n9710_;
  assign new_n9718_ = ~new_n9713_ & ~new_n9716_;
  assign new_n9719_ = new_n9717_ & new_n9718_;
  assign new_n9720_ = ng6581 & ng6692;
  assign new_n9721_ = new_n9701_ & new_n9720_;
  assign new_n9722_ = ng6727 & new_n9687_;
  assign new_n9723_ = ng6625 & ng6715;
  assign new_n9724_ = new_n9722_ & new_n9723_;
  assign new_n9725_ = ng6711 & ng6609;
  assign new_n9726_ = new_n9711_ & new_n9725_;
  assign new_n9727_ = ng6727 & new_n4759_;
  assign new_n9728_ = ng6641 & ng6719;
  assign new_n9729_ = new_n9727_ & new_n9728_;
  assign new_n9730_ = ~new_n9721_ & ~new_n9724_;
  assign new_n9731_ = ~new_n9726_ & ~new_n9729_;
  assign new_n9732_ = new_n9730_ & new_n9731_;
  assign new_n9733_ = new_n9683_ & new_n9707_;
  assign new_n9734_ = ng6645 & ng6661;
  assign new_n9735_ = new_n9733_ & new_n9734_;
  assign new_n9736_ = ng6593 & ng6692;
  assign new_n9737_ = new_n9688_ & new_n9736_;
  assign new_n9738_ = ng6597 & ng6668;
  assign new_n9739_ = new_n9692_ & new_n9738_;
  assign new_n9740_ = ng6711 & ng6617;
  assign new_n9741_ = new_n9695_ & new_n9740_;
  assign new_n9742_ = ~new_n9735_ & ~new_n9737_;
  assign new_n9743_ = ~new_n9739_ & ~new_n9741_;
  assign new_n9744_ = new_n9742_ & new_n9743_;
  assign new_n9745_ = new_n9719_ & new_n9732_;
  assign new_n9746_ = new_n9744_ & new_n9745_;
  assign new_n9747_ = new_n9683_ & ~new_n9707_;
  assign new_n9748_ = ng6621 & ng6675;
  assign new_n9749_ = new_n9747_ & new_n9748_;
  assign new_n9750_ = new_n9687_ & ~new_n9707_;
  assign new_n9751_ = ng6653 & ng6661;
  assign new_n9752_ = new_n9750_ & new_n9751_;
  assign new_n9753_ = new_n9691_ & ~new_n9707_;
  assign new_n9754_ = ng6704 & ng6637;
  assign new_n9755_ = new_n9753_ & new_n9754_;
  assign new_n9756_ = ng6657 & ng6668;
  assign new_n9757_ = new_n9727_ & new_n9756_;
  assign new_n9758_ = ~new_n9749_ & ~new_n9752_;
  assign new_n9759_ = ~new_n9755_ & ~new_n9757_;
  assign new_n9760_ = new_n9758_ & new_n9759_;
  assign new_n9761_ = new_n9700_ & new_n9746_;
  assign new_n9762_ = new_n9760_ & new_n9761_;
  assign new_n9763_ = new_n9682_ & ~new_n9762_;
  assign new_n9764_ = new_n9682_ & ~new_n9763_;
  assign new_n9765_ = ~new_n9762_ & ~new_n9763_;
  assign new_n9766_ = ~new_n9764_ & ~new_n9765_;
  assign new_n9767_ = new_n7218_1_ & ~new_n9766_;
  assign new_n9768_ = ng6500 & ~new_n7218_1_;
  assign new_n9769_ = ~new_n9767_ & ~new_n9768_;
  assign new_n9770_ = pg35 & ~new_n9769_;
  assign n2723 = new_n9681_ | new_n9770_;
  assign new_n9772_ = ~pg35 & ng2719;
  assign new_n9773_ = ng2724 & ~new_n6639_;
  assign new_n9774_ = ~ng2724 & new_n6639_;
  assign new_n9775_ = ~new_n9773_ & ~new_n9774_;
  assign new_n9776_ = ng2841 & ~new_n9775_;
  assign new_n9777_ = pg35 & new_n9776_;
  assign n2728 = new_n9772_ | new_n9777_;
  assign new_n9779_ = ~pg35 & ng2898;
  assign new_n9780_ = n6079 & new_n7895_;
  assign new_n9781_ = ~ng2882 & new_n5037_;
  assign new_n9782_ = ~new_n9780_ & ~new_n9781_;
  assign new_n9783_ = pg35 & new_n9782_;
  assign n2733 = new_n9779_ | new_n9783_;
  assign new_n9785_ = ~pg35 & ng2537;
  assign new_n9786_ = ~ng2495 & ~ng2421;
  assign new_n9787_ = ~new_n7555_ & new_n9786_;
  assign new_n9788_ = ng2541 & ~new_n9787_;
  assign new_n9789_ = ~ng2541 & new_n9787_;
  assign new_n9790_ = ~new_n9788_ & ~new_n9789_;
  assign new_n9791_ = pg35 & ~new_n9790_;
  assign n2738 = new_n9785_ | new_n9791_;
  assign new_n9793_ = ~pg35 & ng6637;
  assign new_n9794_ = new_n6316_ & new_n7159_;
  assign new_n9795_ = ng6653 & ~new_n9794_;
  assign new_n9796_ = ~new_n5966_ & new_n9794_;
  assign new_n9797_ = ~new_n9795_ & ~new_n9796_;
  assign new_n9798_ = pg35 & ~new_n9797_;
  assign n2743 = new_n9793_ | new_n9798_;
  assign new_n9800_ = pg35 & ng4899;
  assign new_n9801_ = ~pg35 & new_n9800_;
  assign new_n9802_ = ~ng6682 & ~ng6732;
  assign new_n9803_ = ~ng6741 & new_n9802_;
  assign new_n9804_ = ng6682 & ng6732;
  assign new_n9805_ = ~ng6741 & new_n9804_;
  assign new_n9806_ = ~ng6736 & ~ng6682;
  assign new_n9807_ = ng6741 & new_n9806_;
  assign new_n9808_ = ng6736 & ng6682;
  assign new_n9809_ = ng6741 & new_n9808_;
  assign new_n9810_ = ~new_n9803_ & ~new_n9805_;
  assign new_n9811_ = ~new_n9807_ & ~new_n9809_;
  assign new_n9812_ = new_n9810_ & new_n9811_;
  assign new_n9813_ = ~ng4894 & new_n9812_;
  assign new_n9814_ = new_n6053_ & ~new_n9813_;
  assign new_n9815_ = new_n7218_1_ & new_n9814_;
  assign new_n9816_ = ng4894 & ~new_n7218_1_;
  assign new_n9817_ = ~new_n9815_ & ~new_n9816_;
  assign new_n9818_ = pg35 & ~new_n9817_;
  assign n2748 = new_n9801_ | new_n9818_;
  assign new_n9820_ = ~pg35 & ng2453;
  assign new_n9821_ = ~ng2453 & ~new_n5910_;
  assign new_n9822_ = new_n5907_1_ & ~new_n9821_;
  assign new_n9823_ = ng2476 & ~new_n5907_1_;
  assign new_n9824_ = ~new_n9822_ & ~new_n9823_;
  assign new_n9825_ = pg35 & ~new_n9824_;
  assign n2753 = new_n9820_ | new_n9825_;
  assign new_n9827_ = ~pg35 & ng2724;
  assign new_n9828_ = ~ng2729 & new_n6640_;
  assign new_n9829_ = ng2729 & ~new_n6640_;
  assign new_n9830_ = ~new_n9828_ & ~new_n9829_;
  assign new_n9831_ = ng2841 & ~new_n9830_;
  assign new_n9832_ = ng2841 & ~new_n9831_;
  assign new_n9833_ = pg35 & ~new_n9832_;
  assign n2758 = new_n9827_ | new_n9833_;
  assign new_n9835_ = ~pg35 & ng925;
  assign new_n9836_ = ng925 & new_n7079_;
  assign new_n9837_ = ng930 & ng1227;
  assign new_n9838_ = ~new_n9836_ & new_n9837_;
  assign new_n9839_ = ~ng930 & new_n9836_;
  assign new_n9840_ = ~new_n9838_ & ~new_n9839_;
  assign new_n9841_ = pg35 & ~new_n9840_;
  assign n2767 = new_n9835_ | new_n9841_;
  assign new_n9843_ = ~pg35 & ng6741;
  assign new_n9844_ = ng6741 & new_n7218_1_;
  assign new_n9845_ = ng6682 & ~new_n9189_;
  assign new_n9846_ = ~new_n9844_ & new_n9845_;
  assign new_n9847_ = ~ng6682 & ~new_n9189_;
  assign new_n9848_ = new_n9844_ & new_n9847_;
  assign new_n9849_ = ~new_n9846_ & ~new_n9848_;
  assign new_n9850_ = pg35 & ~new_n9849_;
  assign n2772 = new_n9843_ | new_n9850_;
  assign new_n9852_ = ~pg35 & ng2868;
  assign new_n9853_ = n4465 & new_n8526_;
  assign new_n9854_ = ng2873 & ~new_n8526_;
  assign new_n9855_ = ~new_n9853_ & ~new_n9854_;
  assign new_n9856_ = pg35 & ~new_n9855_;
  assign n2777 = new_n9852_ | new_n9856_;
  assign new_n9858_ = ~pg35 & ng4975;
  assign new_n9859_ = ng4975 & new_n7706_;
  assign new_n9860_ = ng4899 & ~new_n7708_;
  assign new_n9861_ = ~new_n9859_ & new_n9860_;
  assign new_n9862_ = ~ng4899 & ~new_n7708_;
  assign new_n9863_ = new_n9859_ & new_n9862_;
  assign new_n9864_ = ~new_n9861_ & ~new_n9863_;
  assign new_n9865_ = pg35 & ~new_n9864_;
  assign n2782 = new_n9858_ | new_n9865_;
  assign new_n9867_ = ~pg35 & ng3480;
  assign new_n9868_ = ng3484 & ~new_n7432_;
  assign new_n9869_ = ~ng3484 & new_n7432_;
  assign new_n9870_ = ~new_n9868_ & ~new_n9869_;
  assign new_n9871_ = pg35 & ~new_n9870_;
  assign n2792 = new_n9867_ | new_n9871_;
  assign new_n9873_ = ~pg35 & ng599;
  assign new_n9874_ = ng604 & ~new_n6545_;
  assign new_n9875_ = ~new_n9114_ & new_n9874_;
  assign new_n9876_ = ~ng604 & new_n9114_;
  assign new_n9877_ = ~new_n9875_ & ~new_n9876_;
  assign new_n9878_ = pg35 & ~new_n9877_;
  assign n2797 = new_n9873_ | new_n9878_;
  assign new_n9880_ = ~pg35 & ng1811;
  assign new_n9881_ = ng1825 & ~new_n6805_;
  assign new_n9882_ = ng1811 & new_n9881_;
  assign new_n9883_ = new_n9881_ & ~new_n9882_;
  assign new_n9884_ = ng1811 & ~new_n9882_;
  assign new_n9885_ = ~new_n9883_ & ~new_n9884_;
  assign new_n9886_ = new_n6683_ & ~new_n9885_;
  assign new_n9887_ = ng1825 & ~new_n6683_;
  assign new_n9888_ = ~new_n9886_ & ~new_n9887_;
  assign new_n9889_ = pg35 & ~new_n9888_;
  assign n2802 = new_n9880_ | new_n9889_;
  assign new_n9891_ = ~pg35 & ng4417;
  assign new_n9892_ = ~ng4417 & ng4392;
  assign new_n9893_ = ~ng4417 & ~new_n9892_;
  assign new_n9894_ = new_n7684_ & new_n9893_;
  assign new_n9895_ = ng4392 & ~new_n7684_;
  assign new_n9896_ = ~new_n9894_ & ~new_n9895_;
  assign new_n9897_ = pg35 & ~new_n9896_;
  assign n2807 = new_n9891_ | new_n9897_;
  assign new_n9899_ = pg35 & ng1413;
  assign new_n9900_ = ~pg35 & new_n9899_;
  assign new_n9901_ = ~ng1399 & ~ng1333;
  assign new_n9902_ = ~ng1500 & new_n9901_;
  assign new_n9903_ = ng1570 & ~new_n9902_;
  assign new_n9904_ = ng1395 & new_n9903_;
  assign new_n9905_ = ~ng1395 & ~new_n9903_;
  assign new_n9906_ = ~new_n9904_ & ~new_n9905_;
  assign new_n9907_ = ~ng1322 & new_n9906_;
  assign new_n9908_ = pg35 & new_n9907_;
  assign n2817 = new_n9900_ | new_n9908_;
  assign new_n9910_ = ~pg35 & ng676;
  assign new_n9911_ = ng499 & ~ng504;
  assign new_n9912_ = new_n6780_ & new_n9911_;
  assign new_n9913_ = new_n6067_ & new_n9912_;
  assign new_n9914_ = ng671 & new_n9913_;
  assign new_n9915_ = ng676 & new_n9914_;
  assign new_n9916_ = ~ng718 & ng655;
  assign new_n9917_ = ng655 & ~new_n9916_;
  assign new_n9918_ = ~ng718 & ~new_n9916_;
  assign new_n9919_ = ~new_n9917_ & ~new_n9918_;
  assign new_n9920_ = ng681 & ~ng645;
  assign new_n9921_ = ~ng650 & new_n9920_;
  assign new_n9922_ = ng661 & ~ng728;
  assign new_n9923_ = ng661 & ~new_n9922_;
  assign new_n9924_ = ~ng728 & ~new_n9922_;
  assign new_n9925_ = ~new_n9923_ & ~new_n9924_;
  assign new_n9926_ = ng699 & ~new_n9919_;
  assign new_n9927_ = new_n9921_ & new_n9926_;
  assign new_n9928_ = ~new_n9925_ & new_n9927_;
  assign new_n9929_ = new_n9913_ & new_n9928_;
  assign new_n9930_ = ng703 & ~new_n9929_;
  assign new_n9931_ = ~ng714 & new_n9930_;
  assign new_n9932_ = new_n9915_ & new_n9931_;
  assign new_n9933_ = ng714 & new_n9930_;
  assign new_n9934_ = ~new_n9915_ & new_n9933_;
  assign new_n9935_ = ~new_n9932_ & ~new_n9934_;
  assign new_n9936_ = pg35 & ~new_n9935_;
  assign n2822 = new_n9910_ | new_n9936_;
  assign new_n9938_ = ~pg35 & ng728;
  assign new_n9939_ = ~ng661 & ~ng728;
  assign new_n9940_ = new_n9913_ & ~new_n9939_;
  assign new_n9941_ = ng79 & ~new_n9913_;
  assign new_n9942_ = ~new_n9940_ & ~new_n9941_;
  assign new_n9943_ = pg35 & ~new_n9942_;
  assign n2827 = new_n9938_ | new_n9943_;
  assign new_n9945_ = ~pg35 & ng6541;
  assign new_n9946_ = ng6505 & ~new_n7390_;
  assign new_n9947_ = ng6541 & new_n7390_;
  assign new_n9948_ = ~new_n9946_ & ~new_n9947_;
  assign new_n9949_ = pg35 & ~new_n9948_;
  assign n2832 = new_n9945_ | new_n9949_;
  assign new_n9951_ = ~pg35 & ng5467;
  assign new_n9952_ = ng5462 & ~new_n8547_;
  assign new_n9953_ = ~ng5703 & ~ng5644;
  assign new_n9954_ = ~ng5689 & new_n9953_;
  assign new_n9955_ = ng5677 & ng5595;
  assign new_n9956_ = new_n9954_ & new_n9955_;
  assign new_n9957_ = ~ng5703 & ng5644;
  assign new_n9958_ = ~ng5689 & new_n9957_;
  assign new_n9959_ = ng5685 & ng5567;
  assign new_n9960_ = new_n9958_ & new_n9959_;
  assign new_n9961_ = ng5703 & ~ng5644;
  assign new_n9962_ = ~ng5689 & new_n9961_;
  assign new_n9963_ = ng5681 & ng5611;
  assign new_n9964_ = new_n9962_ & new_n9963_;
  assign new_n9965_ = ~ng5689 & new_n4749_;
  assign new_n9966_ = ng5563 & ng5659;
  assign new_n9967_ = new_n9965_ & new_n9966_;
  assign new_n9968_ = ~new_n9956_ & ~new_n9960_;
  assign new_n9969_ = ~new_n9964_ & ~new_n9967_;
  assign new_n9970_ = new_n9968_ & new_n9969_;
  assign new_n9971_ = ng5689 & new_n9953_;
  assign new_n9972_ = ng5685 & ng5551;
  assign new_n9973_ = new_n9971_ & new_n9972_;
  assign new_n9974_ = ng5689 & ng5659;
  assign new_n9975_ = ng5659 & ~new_n9974_;
  assign new_n9976_ = ng5689 & ~new_n9974_;
  assign new_n9977_ = ~new_n9975_ & ~new_n9976_;
  assign new_n9978_ = new_n9957_ & new_n9977_;
  assign new_n9979_ = ng5575 & ng5637;
  assign new_n9980_ = new_n9978_ & new_n9979_;
  assign new_n9981_ = ng5689 & new_n9961_;
  assign new_n9982_ = ng5547 & ng5659;
  assign new_n9983_ = new_n9981_ & new_n9982_;
  assign new_n9984_ = new_n4749_ & new_n9977_;
  assign new_n9985_ = ng5666 & ng5591;
  assign new_n9986_ = new_n9984_ & new_n9985_;
  assign new_n9987_ = ~new_n9973_ & ~new_n9980_;
  assign new_n9988_ = ~new_n9983_ & ~new_n9986_;
  assign new_n9989_ = new_n9987_ & new_n9988_;
  assign new_n9990_ = ng5543 & ng5654;
  assign new_n9991_ = new_n9971_ & new_n9990_;
  assign new_n9992_ = ng5689 & new_n9957_;
  assign new_n9993_ = ng5677 & ng5587;
  assign new_n9994_ = new_n9992_ & new_n9993_;
  assign new_n9995_ = ng5673 & ng5571;
  assign new_n9996_ = new_n9981_ & new_n9995_;
  assign new_n9997_ = ng5689 & new_n4749_;
  assign new_n9998_ = ng5681 & ng5603;
  assign new_n9999_ = new_n9997_ & new_n9998_;
  assign new_n10000_ = ~new_n9991_ & ~new_n9994_;
  assign new_n10001_ = ~new_n9996_ & ~new_n9999_;
  assign new_n10002_ = new_n10000_ & new_n10001_;
  assign new_n10003_ = new_n9953_ & new_n9977_;
  assign new_n10004_ = ng5623 & ng5607;
  assign new_n10005_ = new_n10003_ & new_n10004_;
  assign new_n10006_ = ng5654 & ng5555;
  assign new_n10007_ = new_n9958_ & new_n10006_;
  assign new_n10008_ = ng5630 & ng5559;
  assign new_n10009_ = new_n9962_ & new_n10008_;
  assign new_n10010_ = ng5673 & ng5579;
  assign new_n10011_ = new_n9965_ & new_n10010_;
  assign new_n10012_ = ~new_n10005_ & ~new_n10007_;
  assign new_n10013_ = ~new_n10009_ & ~new_n10011_;
  assign new_n10014_ = new_n10012_ & new_n10013_;
  assign new_n10015_ = new_n9989_ & new_n10002_;
  assign new_n10016_ = new_n10014_ & new_n10015_;
  assign new_n10017_ = new_n9953_ & ~new_n9977_;
  assign new_n10018_ = ng5583 & ng5637;
  assign new_n10019_ = new_n10017_ & new_n10018_;
  assign new_n10020_ = new_n9957_ & ~new_n9977_;
  assign new_n10021_ = ng5623 & ng5615;
  assign new_n10022_ = new_n10020_ & new_n10021_;
  assign new_n10023_ = new_n9961_ & ~new_n9977_;
  assign new_n10024_ = ng5599 & ng5666;
  assign new_n10025_ = new_n10023_ & new_n10024_;
  assign new_n10026_ = ng5630 & ng5619;
  assign new_n10027_ = new_n9997_ & new_n10026_;
  assign new_n10028_ = ~new_n10019_ & ~new_n10022_;
  assign new_n10029_ = ~new_n10025_ & ~new_n10027_;
  assign new_n10030_ = new_n10028_ & new_n10029_;
  assign new_n10031_ = new_n9970_ & new_n10016_;
  assign new_n10032_ = new_n10030_ & new_n10031_;
  assign new_n10033_ = new_n9952_ & ~new_n10032_;
  assign new_n10034_ = new_n9952_ & ~new_n10033_;
  assign new_n10035_ = ~new_n10032_ & ~new_n10033_;
  assign new_n10036_ = ~new_n10034_ & ~new_n10035_;
  assign new_n10037_ = new_n7745_ & ~new_n10036_;
  assign new_n10038_ = ng5462 & ~new_n7745_;
  assign new_n10039_ = ~new_n10037_ & ~new_n10038_;
  assign new_n10040_ = pg35 & ~new_n10039_;
  assign n2837 = new_n9951_ | new_n10040_;
  assign new_n10042_ = ~pg35 & ng3727;
  assign new_n10043_ = ~new_n6077_ & ~new_n6082_;
  assign new_n10044_ = ng3731 & new_n6104_;
  assign new_n10045_ = new_n10043_ & new_n10044_;
  assign new_n10046_ = ~ng3731 & ~new_n10043_;
  assign new_n10047_ = ~new_n10045_ & ~new_n10046_;
  assign new_n10048_ = pg35 & ~new_n10047_;
  assign n2842 = new_n10042_ | new_n10048_;
  assign new_n10050_ = ~pg35 & ng6419;
  assign new_n10051_ = ~new_n6605_ & ~new_n6610_;
  assign new_n10052_ = ng6423 & new_n6632_1_;
  assign new_n10053_ = new_n10051_ & new_n10052_;
  assign new_n10054_ = ~ng6423 & ~new_n10051_;
  assign new_n10055_ = ~new_n10053_ & ~new_n10054_;
  assign new_n10056_ = pg35 & ~new_n10055_;
  assign n2847 = new_n10050_ | new_n10056_;
  assign new_n10058_ = ~pg35 & ng5069;
  assign new_n10059_ = ~new_n8100_ & ~new_n8104_;
  assign new_n10060_ = pg35 & new_n10059_;
  assign n2852 = new_n10058_ | new_n10060_;
  assign new_n10062_ = ~pg35 & ng1644;
  assign new_n10063_ = ng1592 & ~new_n9016_;
  assign new_n10064_ = ~new_n7537_1_ & new_n10063_;
  assign new_n10065_ = ng1636 & new_n7537_1_;
  assign new_n10066_ = ~new_n10064_ & ~new_n10065_;
  assign new_n10067_ = pg35 & ~new_n10066_;
  assign n2857 = new_n10062_ | new_n10067_;
  assign new_n10069_ = pg35 & ng4831;
  assign new_n10070_ = ~pg35 & new_n10069_;
  assign new_n10071_ = ng5869 & new_n8432_;
  assign new_n10072_ = ng5849 & ~new_n10071_;
  assign new_n10073_ = ~new_n5966_ & new_n10072_;
  assign new_n10074_ = new_n10072_ & ~new_n10073_;
  assign new_n10075_ = ~new_n5966_ & ~new_n10073_;
  assign new_n10076_ = ~new_n10074_ & ~new_n10075_;
  assign new_n10077_ = pg35 & ~new_n10076_;
  assign n2862 = new_n10070_ | new_n10077_;
  assign new_n10079_ = ~pg35 & ng2204;
  assign new_n10080_ = ~new_n4724_ & new_n5652_;
  assign new_n10081_ = ~pg113 & new_n10080_;
  assign new_n10082_ = ng112 & new_n10081_;
  assign new_n10083_ = ng2153 & ~new_n10082_;
  assign new_n10084_ = ~new_n6522_ & new_n10083_;
  assign new_n10085_ = ng2197 & new_n6522_;
  assign new_n10086_ = ~new_n10084_ & ~new_n10085_;
  assign new_n10087_ = pg35 & ~new_n10086_;
  assign n2867 = new_n10079_ | new_n10087_;
  assign new_n10089_ = ~pg35 & ng4164;
  assign new_n10090_ = new_n4705_ & new_n4706_1_;
  assign new_n10091_ = new_n5980_ & new_n10090_;
  assign new_n10092_ = ng4129 & ~new_n10091_;
  assign new_n10093_ = ng4164 & new_n10091_;
  assign new_n10094_ = ~new_n10092_ & ~new_n10093_;
  assign new_n10095_ = pg35 & ~new_n10094_;
  assign n2872 = new_n10089_ | new_n10095_;
  assign new_n10097_ = ~pg35 & ng1854;
  assign new_n10098_ = ng1858 & ~new_n7735_;
  assign new_n10099_ = ~ng1854 & ng1848;
  assign new_n10100_ = ng1848 & ~new_n10099_;
  assign new_n10101_ = ~ng1854 & ~new_n10099_;
  assign new_n10102_ = ~new_n10100_ & ~new_n10101_;
  assign new_n10103_ = new_n7735_ & ~new_n10102_;
  assign new_n10104_ = ~new_n10098_ & ~new_n10103_;
  assign new_n10105_ = pg35 & ~new_n10104_;
  assign n2877 = new_n10097_ | new_n10105_;
  assign new_n10107_ = ~pg35 & ng6573;
  assign new_n10108_ = ~ng6573 & ~ng6565;
  assign new_n10109_ = new_n6336_ & new_n10108_;
  assign new_n10110_ = ng6581 & ~new_n10109_;
  assign new_n10111_ = ~new_n5966_ & new_n10109_;
  assign new_n10112_ = ~new_n10110_ & ~new_n10111_;
  assign new_n10113_ = pg35 & ~new_n10112_;
  assign n2882 = new_n10107_ | new_n10113_;
  assign new_n10115_ = ~pg35 & ng1882;
  assign new_n10116_ = new_n5204_ & new_n8171_;
  assign new_n10117_ = ng1902 & ~new_n10116_;
  assign new_n10118_ = ~ng1862 & ng1906;
  assign new_n10119_ = new_n10116_ & ~new_n10118_;
  assign new_n10120_ = ~new_n10117_ & ~new_n10119_;
  assign new_n10121_ = pg35 & ~new_n10120_;
  assign n2887 = new_n10115_ | new_n10121_;
  assign new_n10123_ = ~pg35 & ng2122;
  assign new_n10124_ = ng2126 & ~new_n9160_;
  assign new_n10125_ = ng2116 & ~ng2122;
  assign new_n10126_ = ng2116 & ~new_n10125_;
  assign new_n10127_ = ~ng2122 & ~new_n10125_;
  assign new_n10128_ = ~new_n10126_ & ~new_n10127_;
  assign new_n10129_ = new_n9160_ & ~new_n10128_;
  assign new_n10130_ = ~new_n10124_ & ~new_n10129_;
  assign new_n10131_ = pg35 & ~new_n10130_;
  assign n2892 = new_n10123_ | new_n10131_;
  assign new_n10133_ = ~pg35 & ng577;
  assign new_n10134_ = ng582 & ~new_n6545_;
  assign new_n10135_ = ~new_n6562_1_ & new_n10134_;
  assign new_n10136_ = ~ng582 & new_n6562_1_;
  assign new_n10137_ = ~new_n10135_ & ~new_n10136_;
  assign new_n10138_ = pg35 & ~new_n10137_;
  assign n2901 = new_n10133_ | new_n10138_;
  assign new_n10140_ = ~pg35 & ng3841;
  assign new_n10141_ = ng3845 & ~new_n7011_1_;
  assign new_n10142_ = ~ng3841 & ng3835;
  assign new_n10143_ = ng3835 & ~new_n10142_;
  assign new_n10144_ = ~ng3841 & ~new_n10142_;
  assign new_n10145_ = ~new_n10143_ & ~new_n10144_;
  assign new_n10146_ = new_n7011_1_ & ~new_n10145_;
  assign new_n10147_ = ~new_n10141_ & ~new_n10146_;
  assign new_n10148_ = pg35 & ~new_n10147_;
  assign n2906 = new_n10140_ | new_n10148_;
  assign new_n10150_ = ~pg35 & ng5742;
  assign new_n10151_ = ~ng5731 & new_n6708_;
  assign new_n10152_ = ~ng5736 & new_n10151_;
  assign new_n10153_ = ~ng5742 & new_n10152_;
  assign new_n10154_ = ng5731 & new_n6710_;
  assign new_n10155_ = ng5736 & new_n10154_;
  assign new_n10156_ = ng5742 & new_n10155_;
  assign new_n10157_ = ~new_n10153_ & ~new_n10156_;
  assign new_n10158_ = ~ng5747 & ~new_n10157_;
  assign new_n10159_ = ng5747 & new_n6424_;
  assign new_n10160_ = new_n10157_ & new_n10159_;
  assign new_n10161_ = ~new_n10158_ & ~new_n10160_;
  assign new_n10162_ = pg35 & ~new_n10161_;
  assign n2911 = new_n10150_ | new_n10162_;
  assign new_n10164_ = ~pg35 & ng2060;
  assign new_n10165_ = ~ng2051 & ng2028;
  assign new_n10166_ = ng2020 & new_n10165_;
  assign new_n10167_ = ~ng2060 & ~ng2028;
  assign new_n10168_ = ng2016 & new_n10167_;
  assign new_n10169_ = ng2024 & new_n5208_;
  assign new_n10170_ = ~new_n10166_ & ~new_n10168_;
  assign new_n10171_ = ~new_n10169_ & new_n10170_;
  assign new_n10172_ = ng2051 & ~ng2028;
  assign new_n10173_ = ng2004 & new_n10172_;
  assign new_n10174_ = ng2008 & new_n9159_;
  assign new_n10175_ = ~ng2051 & ng2060;
  assign new_n10176_ = ng2012 & new_n10175_;
  assign new_n10177_ = new_n10171_ & ~new_n10173_;
  assign new_n10178_ = ~new_n10174_ & ~new_n10176_;
  assign new_n10179_ = new_n10177_ & new_n10178_;
  assign new_n10180_ = new_n9143_ & ~new_n10179_;
  assign new_n10181_ = ng2079 & ~new_n9143_;
  assign new_n10182_ = ~new_n10180_ & ~new_n10181_;
  assign new_n10183_ = pg35 & ~new_n10182_;
  assign n2916 = new_n10164_ | new_n10183_;
  assign new_n10185_ = ~pg35 & ng6077;
  assign new_n10186_ = ~ng6065 & new_n9453_;
  assign new_n10187_ = ~ng6069 & new_n10186_;
  assign new_n10188_ = ~ng6073 & new_n10187_;
  assign new_n10189_ = ~ng6077 & new_n10188_;
  assign new_n10190_ = ng6065 & new_n9454_;
  assign new_n10191_ = ng6069 & new_n10190_;
  assign new_n10192_ = ng6073 & new_n10191_;
  assign new_n10193_ = ng6077 & new_n10192_;
  assign new_n10194_ = ~new_n10189_ & ~new_n10193_;
  assign new_n10195_ = ~ng6082 & ~new_n10194_;
  assign new_n10196_ = ng6082 & new_n7527_;
  assign new_n10197_ = new_n10194_ & new_n10196_;
  assign new_n10198_ = ~new_n10195_ & ~new_n10197_;
  assign new_n10199_ = pg35 & ~new_n10198_;
  assign n2921 = new_n10185_ | new_n10199_;
  assign new_n10201_ = ~pg35 & ng5835;
  assign new_n10202_ = ng5841 & ~new_n10071_;
  assign new_n10203_ = ng5835 & new_n10071_;
  assign new_n10204_ = ~new_n10202_ & ~new_n10203_;
  assign new_n10205_ = pg35 & ~new_n10204_;
  assign n2926 = new_n10201_ | new_n10205_;
  assign new_n10207_ = ~pg35 & ng4273;
  assign new_n10208_ = pg35 & ~ng4239;
  assign n2931 = new_n10207_ | new_n10208_;
  assign new_n10210_ = ~pg35 & ng5142;
  assign new_n10211_ = ng5148 & ~pg26801;
  assign new_n10212_ = ng5142 & pg26801;
  assign new_n10213_ = ~new_n10211_ & ~new_n10212_;
  assign new_n10214_ = pg35 & ~new_n10213_;
  assign n2936 = new_n10210_ | new_n10214_;
  assign new_n10216_ = ~pg35 & ng5272;
  assign new_n10217_ = ~ng5297 & ~ng5357;
  assign new_n10218_ = ~ng5343 & new_n10217_;
  assign new_n10219_ = ng5248 & ng5331;
  assign new_n10220_ = new_n10218_ & new_n10219_;
  assign new_n10221_ = ng5297 & ~ng5357;
  assign new_n10222_ = ~ng5343 & new_n10221_;
  assign new_n10223_ = ng5339 & ng5220;
  assign new_n10224_ = new_n10222_ & new_n10223_;
  assign new_n10225_ = ~ng5297 & ng5357;
  assign new_n10226_ = ~ng5343 & new_n10225_;
  assign new_n10227_ = ng5335 & ng5264;
  assign new_n10228_ = new_n10226_ & new_n10227_;
  assign new_n10229_ = ~ng5343 & pg25114;
  assign new_n10230_ = ng5216 & ng5313;
  assign new_n10231_ = new_n10229_ & new_n10230_;
  assign new_n10232_ = ~new_n10220_ & ~new_n10224_;
  assign new_n10233_ = ~new_n10228_ & ~new_n10231_;
  assign new_n10234_ = new_n10232_ & new_n10233_;
  assign new_n10235_ = ng5343 & new_n10217_;
  assign new_n10236_ = ng5204 & ng5339;
  assign new_n10237_ = new_n10235_ & new_n10236_;
  assign new_n10238_ = ng5343 & ng5313;
  assign new_n10239_ = ng5313 & ~new_n10238_;
  assign new_n10240_ = ng5343 & ~new_n10238_;
  assign new_n10241_ = ~new_n10239_ & ~new_n10240_;
  assign new_n10242_ = new_n10221_ & new_n10241_;
  assign new_n10243_ = ng5290 & ng5228;
  assign new_n10244_ = new_n10242_ & new_n10243_;
  assign new_n10245_ = ng5343 & new_n10225_;
  assign new_n10246_ = ng5200 & ng5313;
  assign new_n10247_ = new_n10245_ & new_n10246_;
  assign new_n10248_ = pg25114 & new_n10241_;
  assign new_n10249_ = ng5244 & ng5320;
  assign new_n10250_ = new_n10248_ & new_n10249_;
  assign new_n10251_ = ~new_n10237_ & ~new_n10244_;
  assign new_n10252_ = ~new_n10247_ & ~new_n10250_;
  assign new_n10253_ = new_n10251_ & new_n10252_;
  assign new_n10254_ = ng5196 & ng5308;
  assign new_n10255_ = new_n10235_ & new_n10254_;
  assign new_n10256_ = ng5343 & new_n10221_;
  assign new_n10257_ = ng5240 & ng5331;
  assign new_n10258_ = new_n10256_ & new_n10257_;
  assign new_n10259_ = ng5327 & ng5224;
  assign new_n10260_ = new_n10245_ & new_n10259_;
  assign new_n10261_ = ng5343 & pg25114;
  assign new_n10262_ = ng5256 & ng5335;
  assign new_n10263_ = new_n10261_ & new_n10262_;
  assign new_n10264_ = ~new_n10255_ & ~new_n10258_;
  assign new_n10265_ = ~new_n10260_ & ~new_n10263_;
  assign new_n10266_ = new_n10264_ & new_n10265_;
  assign new_n10267_ = new_n10217_ & new_n10241_;
  assign new_n10268_ = ng5276 & ng5260;
  assign new_n10269_ = new_n10267_ & new_n10268_;
  assign new_n10270_ = ng5308 & ng5208;
  assign new_n10271_ = new_n10222_ & new_n10270_;
  assign new_n10272_ = ng5283 & ng5212;
  assign new_n10273_ = new_n10226_ & new_n10272_;
  assign new_n10274_ = ng5327 & ng5232;
  assign new_n10275_ = new_n10229_ & new_n10274_;
  assign new_n10276_ = ~new_n10269_ & ~new_n10271_;
  assign new_n10277_ = ~new_n10273_ & ~new_n10275_;
  assign new_n10278_ = new_n10276_ & new_n10277_;
  assign new_n10279_ = new_n10253_ & new_n10266_;
  assign new_n10280_ = new_n10278_ & new_n10279_;
  assign new_n10281_ = new_n10217_ & ~new_n10241_;
  assign new_n10282_ = ng5290 & ng5236;
  assign new_n10283_ = new_n10281_ & new_n10282_;
  assign new_n10284_ = new_n10221_ & ~new_n10241_;
  assign new_n10285_ = ng5268 & ng5276;
  assign new_n10286_ = new_n10284_ & new_n10285_;
  assign new_n10287_ = new_n10225_ & ~new_n10241_;
  assign new_n10288_ = ng5252 & ng5320;
  assign new_n10289_ = new_n10287_ & new_n10288_;
  assign new_n10290_ = ng5283 & ng5272;
  assign new_n10291_ = new_n10261_ & new_n10290_;
  assign new_n10292_ = ~new_n10283_ & ~new_n10286_;
  assign new_n10293_ = ~new_n10289_ & ~new_n10291_;
  assign new_n10294_ = new_n10292_ & new_n10293_;
  assign new_n10295_ = new_n10234_ & new_n10280_;
  assign new_n10296_ = new_n10294_ & new_n10295_;
  assign new_n10297_ = pg33959 & ~new_n10296_;
  assign new_n10298_ = ng128 & ~pg33959;
  assign new_n10299_ = ~new_n10297_ & ~new_n10298_;
  assign new_n10300_ = pg35 & ~new_n10299_;
  assign n2953 = new_n10216_ | new_n10300_;
  assign new_n10302_ = ~pg35 & ng2587;
  assign new_n10303_ = ~ng2819 & new_n5902_1_;
  assign new_n10304_ = new_n5904_ & ~new_n10303_;
  assign new_n10305_ = ng2715 & ~new_n10304_;
  assign new_n10306_ = ng2719 & new_n10305_;
  assign new_n10307_ = ~pg113 & new_n5195_;
  assign new_n10308_ = new_n5909_ & new_n10307_;
  assign new_n10309_ = ~ng2587 & ~new_n10308_;
  assign new_n10310_ = new_n10306_ & ~new_n10309_;
  assign new_n10311_ = ng2610 & ~new_n10306_;
  assign new_n10312_ = ~new_n10310_ & ~new_n10311_;
  assign new_n10313_ = pg35 & ~new_n10312_;
  assign n2958 = new_n10302_ | new_n10313_;
  assign new_n10315_ = ~pg35 & ng6723;
  assign new_n10316_ = ng6727 & ~new_n8611_;
  assign new_n10317_ = ~ng6727 & new_n8611_;
  assign new_n10318_ = ~new_n10316_ & ~new_n10317_;
  assign new_n10319_ = pg35 & ~new_n10318_;
  assign n2963 = new_n10315_ | new_n10319_;
  assign n2968 = ~pg35 & ng4741;
  assign new_n10322_ = ~pg35 & ng3139;
  assign new_n10323_ = ng3143 & ~new_n7152_;
  assign new_n10324_ = ~ng3139 & ng3133;
  assign new_n10325_ = ng3133 & ~new_n10324_;
  assign new_n10326_ = ~ng3139 & ~new_n10324_;
  assign new_n10327_ = ~new_n10325_ & ~new_n10326_;
  assign new_n10328_ = new_n7152_ & ~new_n10327_;
  assign new_n10329_ = ~new_n10323_ & ~new_n10328_;
  assign new_n10330_ = pg35 & ~new_n10329_;
  assign n2973 = new_n10322_ | new_n10330_;
  assign new_n10332_ = ~pg35 & ng4912;
  assign new_n10333_ = ng4927 & ~new_n7449_;
  assign new_n10334_ = ~n6079 & new_n7449_;
  assign new_n10335_ = ~new_n10333_ & ~new_n10334_;
  assign new_n10336_ = pg35 & ~new_n10335_;
  assign n2978 = new_n10332_ | new_n10336_;
  assign new_n10338_ = ~pg35 & ng5073;
  assign new_n10339_ = ng5069 & ng5073;
  assign new_n10340_ = pg35 & new_n10339_;
  assign n2983 = new_n10338_ | new_n10340_;
  assign new_n10342_ = ~pg35 & ng2319;
  assign new_n10343_ = ~pg113 & new_n5193_;
  assign new_n10344_ = new_n5909_ & new_n10343_;
  assign new_n10345_ = ~ng2319 & ~new_n10344_;
  assign new_n10346_ = new_n7259_ & ~new_n10345_;
  assign new_n10347_ = ng2342 & ~new_n7259_;
  assign new_n10348_ = ~new_n10346_ & ~new_n10347_;
  assign new_n10349_ = pg35 & ~new_n10348_;
  assign n2988 = new_n10342_ | new_n10349_;
  assign new_n10351_ = ~pg35 & ng3550;
  assign new_n10352_ = ng3530 & ~ng3522;
  assign new_n10353_ = ng3506 & ~ng3512;
  assign new_n10354_ = new_n10352_ & new_n10353_;
  assign new_n10355_ = ng3574 & ~new_n10354_;
  assign new_n10356_ = ~new_n5966_ & new_n10354_;
  assign new_n10357_ = ~new_n10355_ & ~new_n10356_;
  assign new_n10358_ = pg35 & ~new_n10357_;
  assign n2993 = new_n10351_ | new_n10358_;
  assign new_n10360_ = ~pg35 & ng4135;
  assign new_n10361_ = new_n4706_1_ & new_n6904_;
  assign new_n10362_ = new_n5980_ & new_n10361_;
  assign new_n10363_ = ng4138 & ~new_n10362_;
  assign new_n10364_ = ng4164 & new_n10362_;
  assign new_n10365_ = ~new_n10363_ & ~new_n10364_;
  assign new_n10366_ = pg35 & ~new_n10365_;
  assign n2998 = new_n10360_ | new_n10366_;
  assign new_n10368_ = ~pg35 & ng2327;
  assign new_n10369_ = ng2319 & ~ng2351;
  assign new_n10370_ = ~ng2342 & ~ng2351;
  assign new_n10371_ = ~new_n10369_ & ~new_n10370_;
  assign new_n10372_ = ~new_n10344_ & new_n10371_;
  assign new_n10373_ = new_n7259_ & ~new_n10372_;
  assign new_n10374_ = ng2319 & ~new_n7259_;
  assign new_n10375_ = ~new_n10373_ & ~new_n10374_;
  assign new_n10376_ = pg35 & ~new_n10375_;
  assign n3003 = new_n10368_ | new_n10376_;
  assign new_n10378_ = ~pg35 & ng5802;
  assign new_n10379_ = ~ng5802 & ng5794;
  assign new_n10380_ = ~ng5752 & ~new_n10379_;
  assign new_n10381_ = ~ng5798 & ~new_n10380_;
  assign new_n10382_ = pg35 & new_n10381_;
  assign n3008 = new_n10378_ | new_n10382_;
  assign new_n10384_ = ng22 & pg34927;
  assign new_n10385_ = ~ng22 & n5005;
  assign n3013 = new_n10384_ | new_n10385_;
  assign new_n10387_ = ~pg35 & ng5787;
  assign new_n10388_ = ng5774 & ng5782;
  assign new_n10389_ = ng5787 & new_n10388_;
  assign new_n10390_ = ~ng5791 & new_n10389_;
  assign new_n10391_ = ng5791 & ~new_n10389_;
  assign new_n10392_ = ~new_n10390_ & ~new_n10391_;
  assign new_n10393_ = pg35 & ~new_n10392_;
  assign n3018 = new_n10387_ | new_n10393_;
  assign new_n10395_ = ~pg35 & ng1036;
  assign new_n10396_ = ~new_n5939_ & ~new_n5940_1_;
  assign new_n10397_ = ng1041 & ~new_n10396_;
  assign new_n10398_ = ~ng1041 & ng1008;
  assign new_n10399_ = new_n10396_ & new_n10398_;
  assign new_n10400_ = ~new_n10397_ & ~new_n10399_;
  assign new_n10401_ = pg35 & ~new_n10400_;
  assign n3023 = new_n10395_ | new_n10401_;
  assign new_n10403_ = ~pg35 & ng3767;
  assign new_n10404_ = ng3774 & new_n9043_;
  assign new_n10405_ = ~ng3774 & new_n9047_;
  assign new_n10406_ = ~new_n10404_ & ~new_n10405_;
  assign new_n10407_ = pg35 & ~new_n10406_;
  assign n3028 = new_n10403_ | new_n10407_;
  assign new_n10409_ = pg35 & ~ng4581;
  assign new_n10410_ = ~pg35 & ~new_n10409_;
  assign new_n10411_ = ng4473 & ng4467;
  assign new_n10412_ = ~ng4462 & ~new_n10411_;
  assign new_n10413_ = ~new_n9232_ & new_n10412_;
  assign new_n10414_ = pg35 & ~new_n10413_;
  assign n3033 = new_n10410_ | new_n10414_;
  assign new_n10416_ = ~pg35 & ng2273;
  assign new_n10417_ = ng2279 & ~new_n9535_;
  assign new_n10418_ = ng2273 & new_n9535_;
  assign new_n10419_ = ~new_n10417_ & ~new_n10418_;
  assign new_n10420_ = pg35 & ~new_n10419_;
  assign n3038 = new_n10416_ | new_n10420_;
  assign new_n10422_ = pg35 & ng632;
  assign new_n10423_ = ~pg35 & new_n10422_;
  assign new_n10424_ = pg35 & ng106;
  assign n3043 = new_n10423_ | new_n10424_;
  assign new_n10426_ = ~pg35 & ng2555;
  assign new_n10427_ = ~pg113 & new_n5655_;
  assign new_n10428_ = ~new_n4724_ & new_n10427_;
  assign new_n10429_ = new_n7173_1_ & new_n10428_;
  assign new_n10430_ = ~ng2599 & ng2629;
  assign new_n10431_ = ng112 & new_n10430_;
  assign new_n10432_ = ng112 & ~new_n10431_;
  assign new_n10433_ = new_n10430_ & ~new_n10431_;
  assign new_n10434_ = ~new_n10432_ & ~new_n10433_;
  assign new_n10435_ = new_n10429_ & ~new_n10434_;
  assign new_n10436_ = ng2606 & ~new_n10429_;
  assign new_n10437_ = ~new_n10435_ & ~new_n10436_;
  assign new_n10438_ = pg35 & ~new_n10437_;
  assign n3048 = new_n10426_ | new_n10438_;
  assign new_n10440_ = ~pg35 & ng232;
  assign new_n10441_ = ng878 & new_n6112_;
  assign new_n10442_ = ng262 & ~new_n6112_;
  assign new_n10443_ = ~new_n10441_ & ~new_n10442_;
  assign new_n10444_ = pg35 & ~new_n10443_;
  assign n3053 = new_n10440_ | new_n10444_;
  assign new_n10446_ = pg35 & ng3494;
  assign new_n10447_ = ~pg35 & new_n10446_;
  assign new_n10448_ = ng12 & new_n5059_;
  assign new_n10449_ = n3583 & new_n10448_;
  assign new_n10450_ = ng3502 & ~new_n10448_;
  assign new_n10451_ = ~new_n10449_ & ~new_n10450_;
  assign new_n10452_ = pg35 & ~new_n10451_;
  assign n3058 = new_n10447_ | new_n10452_;
  assign new_n10454_ = ~pg35 & ng5808;
  assign new_n10455_ = ng5817 & ~new_n6354_;
  assign new_n10456_ = ng5808 & ng5813;
  assign new_n10457_ = ng5813 & ~new_n10456_;
  assign new_n10458_ = ng5808 & ~new_n10456_;
  assign new_n10459_ = ~new_n10457_ & ~new_n10458_;
  assign new_n10460_ = new_n6354_ & ~new_n10459_;
  assign new_n10461_ = ~new_n10455_ & ~new_n10460_;
  assign new_n10462_ = pg35 & ~new_n10461_;
  assign n3063 = new_n10454_ | new_n10462_;
  assign new_n10464_ = ~pg35 & ng4950;
  assign new_n10465_ = ~new_n6055_1_ & ~new_n8974_;
  assign new_n10466_ = ng4950 & ~new_n6055_1_;
  assign new_n10467_ = ~new_n6058_ & ~new_n10466_;
  assign new_n10468_ = ~new_n10465_ & ~new_n10467_;
  assign new_n10469_ = ng4944 & new_n10465_;
  assign new_n10470_ = ~new_n10468_ & ~new_n10469_;
  assign new_n10471_ = pg35 & ~new_n10470_;
  assign n3068 = new_n10464_ | new_n10471_;
  assign new_n10473_ = ~pg35 & ng3821;
  assign new_n10474_ = ng3827 & ~new_n6468_;
  assign new_n10475_ = ng3821 & new_n6468_;
  assign new_n10476_ = ~new_n10474_ & ~new_n10475_;
  assign new_n10477_ = pg35 & ~new_n10476_;
  assign n3073 = new_n10473_ | new_n10477_;
  assign new_n10479_ = pg35 & ng4709;
  assign new_n10480_ = ~pg35 & new_n10479_;
  assign new_n10481_ = new_n5665_ & new_n5667_;
  assign new_n10482_ = ~ng5297 & ~ng5348;
  assign new_n10483_ = ~ng5357 & new_n10482_;
  assign new_n10484_ = ng5297 & ng5348;
  assign new_n10485_ = ~ng5357 & new_n10484_;
  assign new_n10486_ = ~ng5297 & ~ng5352;
  assign new_n10487_ = ng5357 & new_n10486_;
  assign new_n10488_ = ng5297 & ng5352;
  assign new_n10489_ = ng5357 & new_n10488_;
  assign new_n10490_ = ~new_n10483_ & ~new_n10485_;
  assign new_n10491_ = ~new_n10487_ & ~new_n10489_;
  assign new_n10492_ = new_n10490_ & new_n10491_;
  assign new_n10493_ = ~ng4704 & new_n10492_;
  assign new_n10494_ = new_n10481_ & ~new_n10493_;
  assign new_n10495_ = pg33959 & new_n10494_;
  assign new_n10496_ = ng4704 & ~pg33959;
  assign new_n10497_ = ~new_n10495_ & ~new_n10496_;
  assign new_n10498_ = pg35 & ~new_n10497_;
  assign n3078 = new_n10480_ | new_n10498_;
  assign new_n10500_ = ~pg35 & ng311;
  assign new_n10501_ = ng336 & new_n6481_;
  assign new_n10502_ = ~new_n7286_ & ~new_n10501_;
  assign new_n10503_ = pg35 & ~new_n10502_;
  assign n3083 = new_n10500_ | new_n10503_;
  assign new_n10505_ = pg35 & ng2152;
  assign new_n10506_ = ~pg35 & new_n10505_;
  assign new_n10507_ = ng2153 & ~ng2227;
  assign new_n10508_ = ~ng2197 & ~ng2227;
  assign new_n10509_ = ~new_n10507_ & ~new_n10508_;
  assign new_n10510_ = ~new_n10082_ & ~new_n10509_;
  assign new_n10511_ = ~new_n6522_ & new_n10510_;
  assign new_n10512_ = ng2153 & new_n6522_;
  assign new_n10513_ = ~new_n10511_ & ~new_n10512_;
  assign new_n10514_ = pg35 & ~new_n10513_;
  assign n3088 = new_n10506_ | new_n10514_;
  assign new_n10516_ = ~pg35 & ng3476;
  assign new_n10517_ = ng3480 & ~new_n7432_;
  assign new_n10518_ = ng3470 & ~ng3476;
  assign new_n10519_ = ng3470 & ~new_n10518_;
  assign new_n10520_ = ~ng3476 & ~new_n10518_;
  assign new_n10521_ = ~new_n10519_ & ~new_n10520_;
  assign new_n10522_ = new_n7432_ & ~new_n10521_;
  assign new_n10523_ = ~new_n10517_ & ~new_n10522_;
  assign new_n10524_ = pg35 & ~new_n10523_;
  assign n3093 = new_n10516_ | new_n10524_;
  assign new_n10526_ = pg35 & ng4955;
  assign new_n10527_ = ~pg35 & new_n10526_;
  assign new_n10528_ = ~new_n5670_ & ~new_n8716_;
  assign new_n10529_ = ~ng4674 & ~ng4646;
  assign new_n10530_ = ~new_n8716_ & new_n10529_;
  assign new_n10531_ = new_n10528_ & new_n10530_;
  assign new_n10532_ = ~ng4681 & new_n10531_;
  assign new_n10533_ = pg35 & new_n10532_;
  assign n3101 = new_n10527_ | new_n10533_;
  assign new_n10535_ = ~pg35 & ng5352;
  assign new_n10536_ = ~ng5357 & ~new_n9589_;
  assign new_n10537_ = pg33959 & new_n10536_;
  assign new_n10538_ = ng5357 & ~pg33959;
  assign new_n10539_ = ~new_n10537_ & ~new_n10538_;
  assign new_n10540_ = pg35 & ~new_n10539_;
  assign n3106 = new_n10535_ | new_n10540_;
  assign new_n10542_ = ~pg35 & ng4922;
  assign new_n10543_ = ng4907 & ~new_n7449_;
  assign new_n10544_ = n5814 & new_n7449_;
  assign new_n10545_ = ~new_n10543_ & ~new_n10544_;
  assign new_n10546_ = pg35 & ~new_n10545_;
  assign n3111 = new_n10542_ | new_n10546_;
  assign new_n10548_ = ~pg35 & ng3921;
  assign new_n10549_ = new_n6894_ & new_n7125_;
  assign new_n10550_ = ng3937 & ~new_n10549_;
  assign new_n10551_ = ~new_n5966_ & new_n10549_;
  assign new_n10552_ = ~new_n10550_ & ~new_n10551_;
  assign new_n10553_ = pg35 & ~new_n10552_;
  assign n3116 = new_n10548_ | new_n10553_;
  assign new_n10555_ = ~pg35 & ng5933;
  assign new_n10556_ = new_n7995_ & new_n8646_;
  assign new_n10557_ = ng5949 & ~new_n10556_;
  assign new_n10558_ = ~new_n5966_ & new_n10556_;
  assign new_n10559_ = ~new_n10557_ & ~new_n10558_;
  assign new_n10560_ = pg35 & ~new_n10559_;
  assign n3121 = new_n10555_ | new_n10560_;
  assign new_n10562_ = ~pg35 & ng1848;
  assign new_n10563_ = ng1854 & ~new_n7735_;
  assign new_n10564_ = ng1848 & new_n7735_;
  assign new_n10565_ = ~new_n10563_ & ~new_n10564_;
  assign new_n10566_ = pg35 & ~new_n10565_;
  assign n3126 = new_n10562_ | new_n10566_;
  assign new_n10568_ = ~pg35 & ng4072;
  assign new_n10569_ = ng4169 & ~ng4064;
  assign new_n10570_ = ng4169 & ~new_n10569_;
  assign new_n10571_ = pg35 & ~new_n10570_;
  assign n3131 = new_n10568_ | new_n10571_;
  assign new_n10573_ = ~pg35 & ng6251;
  assign new_n10574_ = new_n6761_1_ & new_n7088_;
  assign new_n10575_ = ng6247 & ~new_n10574_;
  assign new_n10576_ = ~new_n5966_ & new_n10574_;
  assign new_n10577_ = ~new_n10575_ & ~new_n10576_;
  assign new_n10578_ = pg35 & ~new_n10577_;
  assign n3136 = new_n10573_ | new_n10578_;
  assign new_n10580_ = ~pg35 & ng1256;
  assign new_n10581_ = ~ng1259 & new_n9069_;
  assign new_n10582_ = ng1570 & ng1259;
  assign new_n10583_ = ~new_n9069_ & new_n10582_;
  assign new_n10584_ = ~new_n10581_ & ~new_n10583_;
  assign new_n10585_ = pg35 & ~new_n10584_;
  assign n3141 = new_n10580_ | new_n10585_;
  assign new_n10587_ = ~pg35 & ng6641;
  assign new_n10588_ = ng6561 & new_n10108_;
  assign new_n10589_ = ng6589 & ~new_n10588_;
  assign new_n10590_ = ~new_n5966_ & new_n10588_;
  assign new_n10591_ = ~new_n10589_ & ~new_n10590_;
  assign new_n10592_ = pg35 & ~new_n10591_;
  assign n3146 = new_n10587_ | new_n10592_;
  assign new_n10594_ = ~pg35 & ng3010;
  assign new_n10595_ = ~ng3010 & ~ng3050;
  assign new_n10596_ = ng3004 & new_n10595_;
  assign new_n10597_ = ~ng3004 & new_n8954_;
  assign new_n10598_ = ~new_n10595_ & new_n10597_;
  assign new_n10599_ = ~new_n10596_ & ~new_n10598_;
  assign new_n10600_ = pg35 & ~new_n10599_;
  assign n3151 = new_n10594_ | new_n10600_;
  assign new_n10602_ = ~pg35 & ng1862;
  assign new_n10603_ = ~pg113 & new_n5642_;
  assign new_n10604_ = ~new_n4724_ & new_n10603_;
  assign new_n10605_ = new_n6666_ & new_n10604_;
  assign new_n10606_ = ng1936 & ~ng1906;
  assign new_n10607_ = ng112 & new_n10606_;
  assign new_n10608_ = ng112 & ~new_n10607_;
  assign new_n10609_ = new_n10606_ & ~new_n10607_;
  assign new_n10610_ = ~new_n10608_ & ~new_n10609_;
  assign new_n10611_ = new_n10605_ & ~new_n10610_;
  assign new_n10612_ = ng1913 & ~new_n10605_;
  assign new_n10613_ = ~new_n10611_ & ~new_n10612_;
  assign new_n10614_ = pg35 & ~new_n10613_;
  assign n3166 = new_n10602_ | new_n10614_;
  assign new_n10616_ = ~pg35 & ng5485;
  assign new_n10617_ = ng5489 & ~new_n8548_;
  assign new_n10618_ = ~ng5489 & new_n8548_;
  assign new_n10619_ = ~new_n10617_ & ~new_n10618_;
  assign new_n10620_ = pg35 & ~new_n10619_;
  assign n3171 = new_n10616_ | new_n10620_;
  assign new_n10622_ = ~pg35 & ng405;
  assign new_n10623_ = ng182 & ~new_n5994_;
  assign new_n10624_ = ng446 & new_n5994_;
  assign new_n10625_ = ~new_n10623_ & ~new_n10624_;
  assign new_n10626_ = pg35 & ~new_n10625_;
  assign n3176 = new_n10622_ | new_n10626_;
  assign new_n10628_ = pg35 & ng968;
  assign new_n10629_ = ~pg35 & new_n10628_;
  assign new_n10630_ = ~ng1668 & ng1592;
  assign new_n10631_ = ~ng1668 & ~ng1636;
  assign new_n10632_ = ~new_n10630_ & ~new_n10631_;
  assign new_n10633_ = ~new_n9016_ & ~new_n10632_;
  assign new_n10634_ = ~new_n7537_1_ & new_n10633_;
  assign new_n10635_ = ng1592 & new_n7537_1_;
  assign new_n10636_ = ~new_n10634_ & ~new_n10635_;
  assign new_n10637_ = pg35 & ~new_n10636_;
  assign n3181 = new_n10629_ | new_n10637_;
  assign new_n10639_ = pg35 & ng2685;
  assign new_n10640_ = ~pg35 & new_n10639_;
  assign new_n10641_ = n4465 & new_n10448_;
  assign new_n10642_ = ng2689 & ~new_n10448_;
  assign new_n10643_ = ~new_n10641_ & ~new_n10642_;
  assign new_n10644_ = pg35 & ~new_n10643_;
  assign n3186 = new_n10640_ | new_n10644_;
  assign new_n10646_ = ~pg35 & ng3085;
  assign new_n10647_ = ng3085 & new_n6791_1_;
  assign new_n10648_ = ~ng3089 & new_n10647_;
  assign new_n10649_ = ng3089 & ~new_n10647_;
  assign new_n10650_ = ~new_n10648_ & ~new_n10649_;
  assign new_n10651_ = pg35 & ~new_n10650_;
  assign n3191 = new_n10646_ | new_n10651_;
  assign new_n10653_ = ~pg35 & ng2495;
  assign new_n10654_ = ng2509 & ~new_n9786_;
  assign new_n10655_ = ng1589 & new_n7551_1_;
  assign new_n10656_ = ~new_n8463_ & ~new_n10655_;
  assign new_n10657_ = new_n10654_ & ~new_n10656_;
  assign new_n10658_ = new_n10654_ & ~new_n10657_;
  assign new_n10659_ = ~new_n10656_ & ~new_n10657_;
  assign new_n10660_ = ~new_n10658_ & ~new_n10659_;
  assign new_n10661_ = ~new_n7555_ & ~new_n10660_;
  assign new_n10662_ = ng2509 & new_n7555_;
  assign new_n10663_ = ~new_n10661_ & ~new_n10662_;
  assign new_n10664_ = pg35 & ~new_n10663_;
  assign n3201 = new_n10653_ | new_n10664_;
  assign new_n10666_ = ~pg35 & ng3893;
  assign new_n10667_ = new_n6894_ & new_n8490_;
  assign new_n10668_ = ng3921 & ~new_n10667_;
  assign new_n10669_ = ~new_n5966_ & new_n10667_;
  assign new_n10670_ = ~new_n10668_ & ~new_n10669_;
  assign new_n10671_ = pg35 & ~new_n10670_;
  assign n3206 = new_n10666_ | new_n10671_;
  assign new_n10673_ = ~pg35 & ng1744;
  assign new_n10674_ = ~new_n6236_ & new_n7322_;
  assign new_n10675_ = ng1756 & ~new_n10674_;
  assign new_n10676_ = ng4180 & new_n6231_;
  assign new_n10677_ = ~new_n6232_ & ~new_n10676_;
  assign new_n10678_ = ~ng1242 & new_n6232_;
  assign new_n10679_ = ~new_n10677_ & ~new_n10678_;
  assign new_n10680_ = new_n10674_ & ~new_n10679_;
  assign new_n10681_ = ~new_n10675_ & ~new_n10680_;
  assign new_n10682_ = pg35 & ~new_n10681_;
  assign n3211 = new_n10673_ | new_n10682_;
  assign new_n10684_ = ~pg35 & ng6113;
  assign new_n10685_ = ng6120 & new_n7789_;
  assign new_n10686_ = ~ng6120 & new_n7793_;
  assign new_n10687_ = ~new_n10685_ & ~new_n10686_;
  assign new_n10688_ = pg35 & ~new_n10687_;
  assign n3216 = new_n10684_ | new_n10688_;
  assign new_n10690_ = ~pg35 & ng2936;
  assign new_n10691_ = n6079 & new_n9379_;
  assign new_n10692_ = ng2950 & ~new_n9379_;
  assign new_n10693_ = ~new_n10691_ & ~new_n10692_;
  assign new_n10694_ = pg35 & ~new_n10693_;
  assign n3221 = new_n10690_ | new_n10694_;
  assign new_n10696_ = ~pg35 & ng246;
  assign new_n10697_ = ng872 & new_n6112_;
  assign new_n10698_ = ng446 & ~new_n6112_;
  assign new_n10699_ = ~new_n10697_ & ~new_n10698_;
  assign new_n10700_ = pg35 & ~new_n10699_;
  assign n3226 = new_n10696_ | new_n10700_;
  assign new_n10702_ = ~pg35 & ng4340;
  assign new_n10703_ = ng4340 & new_n5862_;
  assign new_n10704_ = ng4349 & ~new_n5873_1_;
  assign new_n10705_ = ~new_n10703_ & new_n10704_;
  assign new_n10706_ = ~ng4349 & ~new_n5873_1_;
  assign new_n10707_ = new_n10703_ & new_n10706_;
  assign new_n10708_ = ~new_n10705_ & ~new_n10707_;
  assign new_n10709_ = pg35 & ~new_n10708_;
  assign n3231 = new_n10702_ | new_n10709_;
  assign new_n10711_ = ~pg35 & ng6154;
  assign new_n10712_ = ng6163 & ~new_n6700_;
  assign new_n10713_ = ng6159 & ng6154;
  assign new_n10714_ = ng6159 & ~new_n10713_;
  assign new_n10715_ = ng6154 & ~new_n10713_;
  assign new_n10716_ = ~new_n10714_ & ~new_n10715_;
  assign new_n10717_ = new_n6700_ & ~new_n10716_;
  assign new_n10718_ = ~new_n10712_ & ~new_n10717_;
  assign new_n10719_ = pg35 & ~new_n10718_;
  assign n3236 = new_n10711_ | new_n10719_;
  assign new_n10721_ = ~pg35 & ng5232;
  assign new_n10722_ = ng5188 & ~ng5180;
  assign new_n10723_ = new_n7581_ & new_n10722_;
  assign new_n10724_ = ng5248 & ~new_n10723_;
  assign new_n10725_ = ~new_n5966_ & new_n10723_;
  assign new_n10726_ = ~new_n10724_ & ~new_n10725_;
  assign new_n10727_ = pg35 & ~new_n10726_;
  assign n3241 = new_n10721_ | new_n10727_;
  assign new_n10729_ = ~pg35 & ng4443;
  assign new_n10730_ = ~ng4392 & new_n8046_;
  assign new_n10731_ = ~ng4382 & ng4438;
  assign new_n10732_ = ~new_n8046_ & new_n10731_;
  assign new_n10733_ = ~new_n10730_ & ~new_n10732_;
  assign new_n10734_ = pg35 & ~new_n10733_;
  assign n3246 = new_n10729_ | new_n10734_;
  assign new_n10736_ = ~pg35 & ng2946;
  assign new_n10737_ = ng4200 & ng4180;
  assign new_n10738_ = ng4180 & ~new_n10737_;
  assign new_n10739_ = ng4200 & ~new_n10737_;
  assign new_n10740_ = ~new_n10738_ & ~new_n10739_;
  assign new_n10741_ = ~ng4207 & ~ng4180;
  assign new_n10742_ = ~ng4210 & ~ng4204;
  assign new_n10743_ = new_n10741_ & new_n10742_;
  assign new_n10744_ = ~ng4200 & ~ng4194;
  assign new_n10745_ = ~ng4197 & ~ng4188;
  assign new_n10746_ = new_n10744_ & new_n10745_;
  assign new_n10747_ = new_n10743_ & new_n10746_;
  assign new_n10748_ = ~ng4191 & new_n10747_;
  assign new_n10749_ = new_n10740_ & ~new_n10748_;
  assign new_n10750_ = pg35 & ~new_n10749_;
  assign n3251 = new_n10736_ | new_n10750_;
  assign new_n10752_ = ~pg35 & ng2112;
  assign new_n10753_ = ng2116 & ~new_n8022_;
  assign new_n10754_ = ~ng2116 & new_n8022_;
  assign new_n10755_ = ~new_n10753_ & ~new_n10754_;
  assign new_n10756_ = pg35 & ~new_n10755_;
  assign n3256 = new_n10752_ | new_n10756_;
  assign new_n10758_ = ~pg35 & ng2689;
  assign new_n10759_ = n5005 & new_n10448_;
  assign new_n10760_ = ng2697 & ~new_n10448_;
  assign new_n10761_ = ~new_n10759_ & ~new_n10760_;
  assign new_n10762_ = pg35 & ~new_n10761_;
  assign n3261 = new_n10758_ | new_n10762_;
  assign new_n10764_ = ng22 & pg34923;
  assign new_n10765_ = ~ng22 & n6079;
  assign n3270 = new_n10764_ | new_n10765_;
  assign new_n10767_ = ~pg35 & ng2461;
  assign new_n10768_ = ~ng2485 & ng2453;
  assign new_n10769_ = ~ng2485 & ~ng2476;
  assign new_n10770_ = ~new_n10768_ & ~new_n10769_;
  assign new_n10771_ = ~new_n5910_ & new_n10770_;
  assign new_n10772_ = new_n5907_1_ & ~new_n10771_;
  assign new_n10773_ = ng2453 & ~new_n5907_1_;
  assign new_n10774_ = ~new_n10772_ & ~new_n10773_;
  assign new_n10775_ = pg35 & ~new_n10774_;
  assign n3275 = new_n10767_ | new_n10775_;
  assign new_n10777_ = ~pg35 & ng3385;
  assign new_n10778_ = ~ng3368 & new_n8386_;
  assign new_n10779_ = ~ng3372 & new_n10778_;
  assign new_n10780_ = ~ng3376 & new_n10779_;
  assign new_n10781_ = ~ng3380 & new_n10780_;
  assign new_n10782_ = ~ng3385 & new_n10781_;
  assign new_n10783_ = ng3368 & new_n8387_;
  assign new_n10784_ = ng3372 & new_n10783_;
  assign new_n10785_ = ng3376 & new_n10784_;
  assign new_n10786_ = ng3380 & new_n10785_;
  assign new_n10787_ = ng3385 & new_n10786_;
  assign new_n10788_ = ~new_n10782_ & ~new_n10787_;
  assign new_n10789_ = ng3391 & new_n8400_;
  assign new_n10790_ = new_n10788_ & new_n10789_;
  assign new_n10791_ = ~ng3391 & ~new_n10788_;
  assign new_n10792_ = ~new_n10790_ & ~new_n10791_;
  assign new_n10793_ = pg35 & ~new_n10792_;
  assign n3280 = new_n10777_ | new_n10793_;
  assign new_n10795_ = ~pg35 & ng4534;
  assign new_n10796_ = ng4537 & ng4534;
  assign new_n10797_ = ng4537 & ~new_n10796_;
  assign new_n10798_ = ng4534 & ~new_n10796_;
  assign new_n10799_ = ~new_n10797_ & ~new_n10798_;
  assign new_n10800_ = pg35 & ~new_n10799_;
  assign n3285 = new_n10795_ | new_n10800_;
  assign new_n10802_ = ~pg35 & ng3590;
  assign new_n10803_ = new_n7697_ & new_n10352_;
  assign new_n10804_ = ng3606 & ~new_n10803_;
  assign new_n10805_ = ~new_n5966_ & new_n10803_;
  assign new_n10806_ = ~new_n10804_ & ~new_n10805_;
  assign new_n10807_ = pg35 & ~new_n10806_;
  assign n3290 = new_n10802_ | new_n10807_;
  assign new_n10809_ = ~pg35 & ng837;
  assign new_n10810_ = ng847 & new_n6067_;
  assign new_n10811_ = ng837 & ng843;
  assign new_n10812_ = ~new_n10810_ & new_n10811_;
  assign new_n10813_ = ng837 & ~ng843;
  assign new_n10814_ = new_n10810_ & new_n10813_;
  assign new_n10815_ = ~new_n10812_ & ~new_n10814_;
  assign new_n10816_ = pg35 & ~new_n10815_;
  assign n3295 = new_n10809_ | new_n10816_;
  assign new_n10818_ = pg35 & ng3440;
  assign new_n10819_ = ~pg35 & new_n10818_;
  assign new_n10820_ = ~ng3518 & ~new_n9472_;
  assign new_n10821_ = ~ng3506 & new_n10820_;
  assign new_n10822_ = pg35 & new_n10821_;
  assign n3300 = new_n10819_ | new_n10822_;
  assign new_n10824_ = ~pg35 & ng1030;
  assign new_n10825_ = new_n6144_1_ & ~new_n6146_;
  assign new_n10826_ = ng1036 & ~new_n10825_;
  assign new_n10827_ = ~ng1036 & new_n6138_;
  assign new_n10828_ = new_n10825_ & new_n10827_;
  assign new_n10829_ = ~new_n10826_ & ~new_n10828_;
  assign new_n10830_ = pg35 & ~new_n10829_;
  assign n3305 = new_n10824_ | new_n10830_;
  assign new_n10832_ = ~pg35 & ng4108;
  assign new_n10833_ = ng4087 & new_n7187_;
  assign new_n10834_ = ng4093 & new_n10833_;
  assign new_n10835_ = ng4098 & new_n10834_;
  assign new_n10836_ = ng4108 & new_n10835_;
  assign new_n10837_ = ~ng4104 & new_n10836_;
  assign new_n10838_ = ng4104 & ~new_n10836_;
  assign new_n10839_ = ~new_n10837_ & ~new_n10838_;
  assign new_n10840_ = ng4169 & ~new_n10839_;
  assign new_n10841_ = ng4169 & ~new_n10840_;
  assign new_n10842_ = pg35 & ~new_n10841_;
  assign n3310 = new_n10832_ | new_n10842_;
  assign new_n10844_ = ~pg35 & ng1700;
  assign new_n10845_ = ~ng1668 & ~ng1592;
  assign new_n10846_ = ~new_n7537_1_ & new_n10845_;
  assign new_n10847_ = ng1706 & ~new_n10846_;
  assign new_n10848_ = ng1700 & new_n10846_;
  assign new_n10849_ = ~new_n10847_ & ~new_n10848_;
  assign new_n10850_ = pg35 & ~new_n10849_;
  assign n3315 = new_n10844_ | new_n10850_;
  assign new_n10852_ = ~pg35 & ng6404;
  assign new_n10853_ = ~ng6404 & ~ng6444;
  assign new_n10854_ = ng6398 & new_n10853_;
  assign new_n10855_ = ~ng6398 & new_n6632_1_;
  assign new_n10856_ = ~new_n10853_ & new_n10855_;
  assign new_n10857_ = ~new_n10854_ & ~new_n10856_;
  assign new_n10858_ = pg35 & ~new_n10857_;
  assign n3320 = new_n10852_ | new_n10858_;
  assign new_n10860_ = ~pg35 & ng5517;
  assign new_n10861_ = ng5511 & ng5517;
  assign new_n10862_ = ~ng5523 & ~new_n8302_;
  assign new_n10863_ = new_n10861_ & new_n10862_;
  assign new_n10864_ = ng5523 & new_n10862_;
  assign new_n10865_ = ~new_n10861_ & new_n10864_;
  assign new_n10866_ = ~new_n10863_ & ~new_n10865_;
  assign new_n10867_ = pg35 & ~new_n10866_;
  assign n3325 = new_n10860_ | new_n10867_;
  assign new_n10869_ = ~pg35 & ng6195;
  assign new_n10870_ = ng6159 & ~new_n7064_;
  assign new_n10871_ = ng6195 & new_n7064_;
  assign new_n10872_ = ~new_n10870_ & ~new_n10871_;
  assign new_n10873_ = pg35 & ~new_n10872_;
  assign n3330 = new_n10869_ | new_n10873_;
  assign new_n10875_ = ~pg35 & ng2950;
  assign new_n10876_ = n4465 & new_n9379_;
  assign new_n10877_ = ng2960 & ~new_n9379_;
  assign new_n10878_ = ~new_n10876_ & ~new_n10877_;
  assign new_n10879_ = pg35 & ~new_n10878_;
  assign n3335 = new_n10875_ | new_n10879_;
  assign new_n10881_ = ~pg35 & ng5489;
  assign new_n10882_ = ng5523 & new_n6885_;
  assign new_n10883_ = ng5495 & ~new_n10882_;
  assign new_n10884_ = ng5489 & new_n10882_;
  assign new_n10885_ = ~new_n10883_ & ~new_n10884_;
  assign new_n10886_ = pg35 & ~new_n10885_;
  assign n3340 = new_n10881_ | new_n10886_;
  assign new_n10888_ = ~pg35 & ng2965;
  assign new_n10889_ = ng12 & n5005;
  assign new_n10890_ = new_n4937_ & new_n10889_;
  assign new_n10891_ = ~ng2975 & new_n5112_1_;
  assign new_n10892_ = ~new_n10890_ & ~new_n10891_;
  assign new_n10893_ = pg35 & new_n10892_;
  assign n3345 = new_n10888_ | new_n10893_;
  assign new_n10895_ = pg35 & ng6483;
  assign new_n10896_ = ~pg35 & new_n10895_;
  assign new_n10897_ = ~ng6549 & new_n8654_;
  assign new_n10898_ = pg35 & new_n10897_;
  assign n3350 = new_n10896_ | new_n10898_;
  assign new_n10900_ = ~pg35 & ng2303;
  assign new_n10901_ = ~new_n7886_ & new_n9176_;
  assign new_n10902_ = ng2315 & ~new_n10901_;
  assign new_n10903_ = ~new_n8906_ & new_n10901_;
  assign new_n10904_ = ~new_n10902_ & ~new_n10903_;
  assign new_n10905_ = pg35 & ~new_n10904_;
  assign n3355 = new_n10900_ | new_n10905_;
  assign new_n10907_ = ~pg35 & ng2575;
  assign new_n10908_ = new_n5219_ & new_n10306_;
  assign new_n10909_ = ng2595 & ~new_n10908_;
  assign new_n10910_ = ng2599 & ~ng2555;
  assign new_n10911_ = new_n10908_ & ~new_n10910_;
  assign new_n10912_ = ~new_n10909_ & ~new_n10911_;
  assign new_n10913_ = pg35 & ~new_n10912_;
  assign n3360 = new_n10907_ | new_n10913_;
  assign new_n10915_ = pg35 & ng6537;
  assign new_n10916_ = ~pg35 & new_n10915_;
  assign new_n10917_ = n2287 & new_n10448_;
  assign new_n10918_ = ng6545 & ~new_n10448_;
  assign new_n10919_ = ~new_n10917_ & ~new_n10918_;
  assign new_n10920_ = pg35 & ~new_n10919_;
  assign n3365 = new_n10916_ | new_n10920_;
  assign new_n10922_ = ~pg35 & ng2638;
  assign new_n10923_ = ng2610 & ~ng2587;
  assign new_n10924_ = ng2652 & ~new_n10923_;
  assign new_n10925_ = ng2638 & new_n10924_;
  assign new_n10926_ = new_n10924_ & ~new_n10925_;
  assign new_n10927_ = ng2638 & ~new_n10925_;
  assign new_n10928_ = ~new_n10926_ & ~new_n10927_;
  assign new_n10929_ = new_n10306_ & ~new_n10928_;
  assign new_n10930_ = ng2652 & ~new_n10306_;
  assign new_n10931_ = ~new_n10929_ & ~new_n10930_;
  assign new_n10932_ = pg35 & ~new_n10931_;
  assign n3370 = new_n10922_ | new_n10932_;
  assign new_n10934_ = ~pg35 & ng6227;
  assign new_n10935_ = new_n7088_ & new_n9572_;
  assign new_n10936_ = ng6235 & ~new_n10935_;
  assign new_n10937_ = ~new_n5966_ & new_n10935_;
  assign new_n10938_ = ~new_n10936_ & ~new_n10937_;
  assign new_n10939_ = pg35 & ~new_n10938_;
  assign n3375 = new_n10934_ | new_n10939_;
  assign new_n10941_ = ~pg35 & ng3380;
  assign new_n10942_ = ~new_n10781_ & ~new_n10786_;
  assign new_n10943_ = ~ng3385 & ~new_n10942_;
  assign new_n10944_ = ng3385 & new_n8400_;
  assign new_n10945_ = new_n10942_ & new_n10944_;
  assign new_n10946_ = ~new_n10943_ & ~new_n10945_;
  assign new_n10947_ = pg35 & ~new_n10946_;
  assign n3380 = new_n10941_ | new_n10947_;
  assign new_n10949_ = ~pg35 & ng546;
  assign new_n10950_ = ~ng542 & ng691;
  assign new_n10951_ = ~new_n6578_ & ~new_n10950_;
  assign new_n10952_ = pg35 & new_n10951_;
  assign n3385 = new_n10949_ | new_n10952_;
  assign new_n10954_ = ~pg35 & ng1834;
  assign new_n10955_ = ng1840 & ~new_n8571_;
  assign new_n10956_ = ng1834 & new_n8571_;
  assign new_n10957_ = ~new_n10955_ & ~new_n10956_;
  assign new_n10958_ = pg35 & ~new_n10957_;
  assign n3390 = new_n10954_ | new_n10958_;
  assign new_n10960_ = ~pg35 & ng847;
  assign new_n10961_ = ng703 & ~new_n6067_;
  assign new_n10962_ = ng822 & ng817;
  assign new_n10963_ = ng723 & new_n10962_;
  assign new_n10964_ = ~ng847 & new_n10963_;
  assign new_n10965_ = ng703 & ~ng812;
  assign new_n10966_ = ~ng837 & ng703;
  assign new_n10967_ = ng703 & ~ng847;
  assign new_n10968_ = ~new_n10964_ & ~new_n10965_;
  assign new_n10969_ = ~new_n10966_ & ~new_n10967_;
  assign new_n10970_ = new_n10968_ & new_n10969_;
  assign new_n10971_ = new_n6067_ & ~new_n10970_;
  assign new_n10972_ = ~new_n10961_ & ~new_n10971_;
  assign new_n10973_ = pg35 & ~new_n10972_;
  assign n3395 = new_n10960_ | new_n10973_;
  assign new_n10975_ = pg35 & ng5297;
  assign new_n10976_ = ~pg35 & new_n10975_;
  assign new_n10977_ = pg35 & ng5188;
  assign n3400 = new_n10976_ | new_n10977_;
  assign new_n10979_ = ~pg35 & ng4125;
  assign new_n10980_ = ~ng4141 & ~ng4064;
  assign new_n10981_ = ~ng4057 & new_n10980_;
  assign new_n10982_ = ~ng4082 & new_n10981_;
  assign new_n10983_ = ng4076 & new_n5805_;
  assign new_n10984_ = new_n10982_ & new_n10983_;
  assign new_n10985_ = ~ng4169 & ~new_n10984_;
  assign new_n10986_ = pg35 & new_n10985_;
  assign n3404 = new_n10979_ | new_n10986_;
  assign new_n10988_ = ~pg35 & ng3129;
  assign new_n10989_ = new_n6915_ & new_n6918_;
  assign new_n10990_ = ng3133 & ~new_n10989_;
  assign new_n10991_ = ~ng3133 & new_n10989_;
  assign new_n10992_ = ~new_n10990_ & ~new_n10991_;
  assign new_n10993_ = pg35 & ~new_n10992_;
  assign n3409 = new_n10988_ | new_n10993_;
  assign new_n10995_ = ~pg35 & ng1913;
  assign new_n10996_ = ng1862 & ~new_n9006_;
  assign new_n10997_ = ~new_n6667_1_ & new_n10996_;
  assign new_n10998_ = ng1906 & new_n6667_1_;
  assign new_n10999_ = ~new_n10997_ & ~new_n10998_;
  assign new_n11000_ = pg35 & ~new_n10999_;
  assign n3419 = new_n10995_ | new_n11000_;
  assign new_n11002_ = ~pg35 & ng4907;
  assign new_n11003_ = ng4912 & ~new_n7449_;
  assign new_n11004_ = n2287 & new_n7449_;
  assign new_n11005_ = ~new_n11003_ & ~new_n11004_;
  assign new_n11006_ = pg35 & ~new_n11005_;
  assign n3424 = new_n11002_ | new_n11006_;
  assign new_n11008_ = ~pg35 & ng1945;
  assign new_n11009_ = ng1959 & ~new_n9091_;
  assign new_n11010_ = ng1945 & new_n11009_;
  assign new_n11011_ = new_n11009_ & ~new_n11010_;
  assign new_n11012_ = ng1945 & ~new_n11010_;
  assign new_n11013_ = ~new_n11011_ & ~new_n11012_;
  assign new_n11014_ = new_n8171_ & ~new_n11013_;
  assign new_n11015_ = ng1959 & ~new_n8171_;
  assign new_n11016_ = ~new_n11014_ & ~new_n11015_;
  assign new_n11017_ = pg35 & ~new_n11016_;
  assign n3429 = new_n11008_ | new_n11017_;
  assign new_n11019_ = pg35 & ng3791;
  assign new_n11020_ = ~pg35 & new_n11019_;
  assign new_n11021_ = ~ng3869 & ~new_n6204_;
  assign new_n11022_ = ~ng3857 & new_n11021_;
  assign new_n11023_ = pg35 & new_n11022_;
  assign n3434 = new_n11020_ | new_n11023_;
  assign new_n11025_ = ~pg35 & ng2361;
  assign new_n11026_ = ng2375 & ~new_n7887_;
  assign new_n11027_ = ~ng1589 & new_n7882_;
  assign new_n11028_ = ~new_n8904_ & ~new_n11027_;
  assign new_n11029_ = new_n11026_ & ~new_n11028_;
  assign new_n11030_ = new_n11026_ & ~new_n11029_;
  assign new_n11031_ = ~new_n11028_ & ~new_n11029_;
  assign new_n11032_ = ~new_n11030_ & ~new_n11031_;
  assign new_n11033_ = ~new_n7886_ & ~new_n11032_;
  assign new_n11034_ = ng2375 & new_n7886_;
  assign new_n11035_ = ~new_n11033_ & ~new_n11034_;
  assign new_n11036_ = pg35 & ~new_n11035_;
  assign n3439 = new_n11025_ | new_n11036_;
  assign new_n11038_ = ~pg35 & ng4983;
  assign new_n11039_ = ng4983 & new_n5679_;
  assign new_n11040_ = ~new_n7706_ & ~new_n7708_;
  assign new_n11041_ = ng4991 & new_n11040_;
  assign new_n11042_ = ~new_n11039_ & new_n11041_;
  assign new_n11043_ = ~ng4991 & new_n11040_;
  assign new_n11044_ = new_n11039_ & new_n11043_;
  assign new_n11045_ = ~new_n11042_ & ~new_n11044_;
  assign new_n11046_ = pg35 & ~new_n11045_;
  assign n3444 = new_n11038_ | new_n11046_;
  assign new_n11048_ = ~pg35 & ng4291;
  assign new_n11049_ = pg35 & ~new_n7631_;
  assign n3449 = new_n11048_ | new_n11049_;
  assign new_n11051_ = ~pg35 & ng2771;
  assign new_n11052_ = ng2715 & ~ng2787;
  assign new_n11053_ = ~ng2715 & ~ng2783;
  assign new_n11054_ = ~new_n11052_ & ~new_n11053_;
  assign new_n11055_ = ng2719 & new_n11054_;
  assign new_n11056_ = ng2715 & ~ng2775;
  assign new_n11057_ = ~ng2715 & ~ng2771;
  assign new_n11058_ = ~new_n11056_ & ~new_n11057_;
  assign new_n11059_ = ~ng2719 & new_n11058_;
  assign new_n11060_ = ~new_n11055_ & ~new_n11059_;
  assign new_n11061_ = new_n7335_ & new_n11060_;
  assign new_n11062_ = ng2715 & ng2079;
  assign new_n11063_ = ~ng2715 & ng1945;
  assign new_n11064_ = ~new_n11062_ & ~new_n11063_;
  assign new_n11065_ = ng2719 & new_n11064_;
  assign new_n11066_ = ng2715 & ng1811;
  assign new_n11067_ = ~ng2715 & ng1677;
  assign new_n11068_ = ~new_n11066_ & ~new_n11067_;
  assign new_n11069_ = ~ng2719 & new_n11068_;
  assign new_n11070_ = ~new_n11065_ & ~new_n11069_;
  assign new_n11071_ = ~new_n7335_ & new_n11070_;
  assign new_n11072_ = ~new_n11061_ & ~new_n11071_;
  assign new_n11073_ = pg35 & ~new_n11072_;
  assign n3454 = new_n11051_ | new_n11073_;
  assign new_n11075_ = ~pg35 & ng736;
  assign new_n11076_ = ng739 & ~new_n6578_;
  assign new_n11077_ = ~new_n6577_ & new_n11076_;
  assign new_n11078_ = ~ng739 & ~new_n6578_;
  assign new_n11079_ = new_n6577_ & new_n11078_;
  assign new_n11080_ = ~new_n11077_ & ~new_n11079_;
  assign new_n11081_ = pg35 & ~new_n11080_;
  assign n3459 = new_n11075_ | new_n11081_;
  assign new_n11083_ = ~pg35 & ng5080;
  assign new_n11084_ = ~ng5069 & ng5077;
  assign new_n11085_ = ~ng5080 & ~new_n11084_;
  assign new_n11086_ = ~ng5084 & new_n11085_;
  assign new_n11087_ = ng5084 & ng5080;
  assign new_n11088_ = ~ng5073 & ng5077;
  assign new_n11089_ = ~new_n11086_ & ~new_n11087_;
  assign new_n11090_ = ~new_n11088_ & new_n11089_;
  assign new_n11091_ = pg35 & ~new_n11090_;
  assign n3464 = new_n11083_ | new_n11091_;
  assign new_n11093_ = ~pg35 & ng4776;
  assign new_n11094_ = ng4785 & ~new_n6160_;
  assign new_n11095_ = ~new_n6157_ & new_n11094_;
  assign new_n11096_ = ~ng4785 & ~new_n6160_;
  assign new_n11097_ = new_n6157_ & new_n11096_;
  assign new_n11098_ = ~new_n11095_ & ~new_n11097_;
  assign new_n11099_ = pg35 & ~new_n11098_;
  assign n3469 = new_n11093_ | new_n11099_;
  assign new_n11101_ = ~pg35 & ng2779;
  assign new_n11102_ = ~ng1902 & new_n7642_;
  assign new_n11103_ = ~ng2791 & ~new_n11102_;
  assign new_n11104_ = ~new_n7640_ & ~new_n11103_;
  assign new_n11105_ = pg35 & new_n11104_;
  assign n3474 = new_n11101_ | new_n11105_;
  assign new_n11107_ = ~pg35 & ng6581;
  assign new_n11108_ = new_n6317_ & new_n10108_;
  assign new_n11109_ = ng6609 & ~new_n11108_;
  assign new_n11110_ = ~new_n5966_ & new_n11108_;
  assign new_n11111_ = ~new_n11109_ & ~new_n11110_;
  assign new_n11112_ = pg35 & ~new_n11111_;
  assign n3479 = new_n11107_ | new_n11112_;
  assign new_n11114_ = ~pg35 & ng2093;
  assign new_n11115_ = new_n9143_ & new_n10172_;
  assign new_n11116_ = ng2098 & ~new_n11115_;
  assign new_n11117_ = ng2093 & ng2089;
  assign new_n11118_ = ng2093 & ~new_n11117_;
  assign new_n11119_ = ng2089 & ~new_n11117_;
  assign new_n11120_ = ~new_n11118_ & ~new_n11119_;
  assign new_n11121_ = new_n11115_ & ~new_n11120_;
  assign new_n11122_ = ~new_n11116_ & ~new_n11121_;
  assign new_n11123_ = pg35 & ~new_n11122_;
  assign n3484 = new_n11114_ | new_n11123_;
  assign new_n11125_ = ~pg35 & ng6451;
  assign new_n11126_ = ~new_n6621_ & ~new_n6629_;
  assign new_n11127_ = pg35 & new_n11126_;
  assign n3489 = new_n11125_ | new_n11127_;
  assign new_n11129_ = ~pg35 & ng3598;
  assign new_n11130_ = ~ng3530 & ~ng3522;
  assign new_n11131_ = ng3518 & new_n11130_;
  assign new_n11132_ = ng3546 & ~new_n11131_;
  assign new_n11133_ = ~new_n5966_ & new_n11131_;
  assign new_n11134_ = ~new_n11132_ & ~new_n11133_;
  assign new_n11135_ = pg35 & ~new_n11134_;
  assign n3494 = new_n11129_ | new_n11135_;
  assign new_n11137_ = ~pg35 & ng2193;
  assign new_n11138_ = ng2185 & ~ng2217;
  assign new_n11139_ = ~ng2217 & ~ng2208;
  assign new_n11140_ = ~new_n11138_ & ~new_n11139_;
  assign new_n11141_ = ~pg113 & new_n5188_;
  assign new_n11142_ = new_n5909_ & new_n11141_;
  assign new_n11143_ = new_n11140_ & ~new_n11142_;
  assign new_n11144_ = new_n9534_ & ~new_n11143_;
  assign new_n11145_ = ng2185 & ~new_n9534_;
  assign new_n11146_ = ~new_n11144_ & ~new_n11145_;
  assign new_n11147_ = pg35 & ~new_n11146_;
  assign n3499 = new_n11137_ | new_n11147_;
  assign new_n11149_ = ~pg35 & ng2476;
  assign new_n11150_ = ~new_n4724_ & new_n5908_;
  assign new_n11151_ = new_n5907_1_ & new_n11150_;
  assign new_n11152_ = ng2485 & ~ng2476;
  assign new_n11153_ = ng110 & new_n11152_;
  assign new_n11154_ = ng110 & ~new_n11153_;
  assign new_n11155_ = new_n11152_ & ~new_n11153_;
  assign new_n11156_ = ~new_n11154_ & ~new_n11155_;
  assign new_n11157_ = new_n11151_ & ~new_n11156_;
  assign new_n11158_ = ng2491 & ~new_n11151_;
  assign new_n11159_ = ~new_n11157_ & ~new_n11158_;
  assign new_n11160_ = pg35 & ~new_n11159_;
  assign n3504 = new_n11149_ | new_n11160_;
  assign new_n11162_ = pg35 & ng1319;
  assign new_n11163_ = ~pg35 & new_n11162_;
  assign new_n11164_ = ng1312 & new_n6294_;
  assign new_n11165_ = new_n6298_ & new_n6833_;
  assign new_n11166_ = ~ng1351 & new_n11165_;
  assign new_n11167_ = ~ng1389 & new_n6300_1_;
  assign new_n11168_ = ng1351 & new_n11167_;
  assign new_n11169_ = ng1312 & new_n6298_;
  assign new_n11170_ = ~new_n11166_ & ~new_n11168_;
  assign new_n11171_ = ~new_n6302_ & ~new_n11169_;
  assign new_n11172_ = new_n11170_ & new_n11171_;
  assign new_n11173_ = ~new_n6294_ & ~new_n11172_;
  assign new_n11174_ = ~new_n11164_ & ~new_n11173_;
  assign new_n11175_ = pg35 & ~new_n11174_;
  assign n3509 = new_n11163_ | new_n11175_;
  assign new_n11177_ = ~pg35 & ng1124;
  assign new_n11178_ = ng1116 & new_n6663_;
  assign new_n11179_ = new_n5888_1_ & new_n11178_;
  assign new_n11180_ = ng1129 & ng1124;
  assign new_n11181_ = ng1129 & ~new_n11180_;
  assign new_n11182_ = ng1124 & ~new_n11180_;
  assign new_n11183_ = ~new_n11181_ & ~new_n11182_;
  assign new_n11184_ = new_n11179_ & ~new_n11183_;
  assign new_n11185_ = ng1129 & ~new_n11179_;
  assign new_n11186_ = ~new_n11184_ & ~new_n11185_;
  assign new_n11187_ = pg35 & ~new_n11186_;
  assign n3514 = new_n11177_ | new_n11187_;
  assign new_n11189_ = ~pg35 & ng1205;
  assign new_n11190_ = ~ng1221 & new_n8559_;
  assign new_n11191_ = ng1221 & ~new_n8559_;
  assign new_n11192_ = ~new_n11190_ & ~new_n11191_;
  assign new_n11193_ = pg35 & ~new_n11192_;
  assign n3519 = new_n11189_ | new_n11193_;
  assign new_n11195_ = ~pg35 & ng1632;
  assign new_n11196_ = ng1624 & ~ng1657;
  assign new_n11197_ = ~ng1657 & ~ng1648;
  assign new_n11198_ = ~new_n11196_ & ~new_n11197_;
  assign new_n11199_ = ~pg113 & new_n5173_;
  assign new_n11200_ = new_n5909_ & new_n11199_;
  assign new_n11201_ = new_n11198_ & ~new_n11200_;
  assign new_n11202_ = new_n7230_ & ~new_n11201_;
  assign new_n11203_ = ng1624 & ~new_n7230_;
  assign new_n11204_ = ~new_n11202_ & ~new_n11203_;
  assign new_n11205_ = pg35 & ~new_n11204_;
  assign n3524 = new_n11195_ | new_n11205_;
  assign new_n11207_ = ~pg35 & ng1844;
  assign new_n11208_ = ng1848 & ~new_n8571_;
  assign new_n11209_ = ~ng1848 & new_n8571_;
  assign new_n11210_ = ~new_n11208_ & ~new_n11209_;
  assign new_n11211_ = pg35 & ~new_n11210_;
  assign n3529 = new_n11207_ | new_n11211_;
  assign new_n11213_ = ~pg35 & ng4854;
  assign new_n11214_ = ng4854 & new_n7603_1_;
  assign new_n11215_ = ng4859 & new_n7606_;
  assign new_n11216_ = ~new_n11214_ & new_n11215_;
  assign new_n11217_ = ~ng4859 & new_n7606_;
  assign new_n11218_ = new_n11214_ & new_n11217_;
  assign new_n11219_ = ~new_n11216_ & ~new_n11218_;
  assign new_n11220_ = pg35 & ~new_n11219_;
  assign n3534 = new_n11213_ | new_n11220_;
  assign new_n11222_ = ~pg35 & ng2999;
  assign new_n11223_ = ~n5814 & new_n8526_;
  assign new_n11224_ = ng2994 & ~new_n8526_;
  assign new_n11225_ = ~new_n11223_ & ~new_n11224_;
  assign new_n11226_ = pg35 & ~new_n11225_;
  assign n3543 = new_n11222_ | new_n11226_;
  assign new_n11228_ = ~pg35 & ng1141;
  assign new_n11229_ = new_n5888_1_ & new_n7772_;
  assign new_n11230_ = ng1141 & ng956;
  assign new_n11231_ = ng956 & ~new_n11230_;
  assign new_n11232_ = ng1141 & ~new_n11230_;
  assign new_n11233_ = ~new_n11231_ & ~new_n11232_;
  assign new_n11234_ = new_n11229_ & ~new_n11233_;
  assign new_n11235_ = ng956 & ~new_n11229_;
  assign new_n11236_ = ~new_n11234_ & ~new_n11235_;
  assign new_n11237_ = pg35 & ~new_n11236_;
  assign n3548 = new_n11228_ | new_n11237_;
  assign new_n11239_ = pg35 & ng2417;
  assign new_n11240_ = ~pg35 & new_n11239_;
  assign new_n11241_ = ~ng2495 & ng2421;
  assign new_n11242_ = ~ng2495 & ~ng2465;
  assign new_n11243_ = ~new_n11241_ & ~new_n11242_;
  assign new_n11244_ = ~new_n7558_ & ~new_n11243_;
  assign new_n11245_ = ~new_n7555_ & new_n11244_;
  assign new_n11246_ = ng2421 & new_n7555_;
  assign new_n11247_ = ~new_n11245_ & ~new_n11246_;
  assign new_n11248_ = pg35 & ~new_n11247_;
  assign n3553 = new_n11240_ | new_n11248_;
  assign new_n11250_ = ~pg35 & ng6527;
  assign new_n11251_ = ng6533 & ~new_n7390_;
  assign new_n11252_ = ng6527 & new_n7390_;
  assign new_n11253_ = ~new_n11251_ & ~new_n11252_;
  assign new_n11254_ = pg35 & ~new_n11253_;
  assign n3558 = new_n11250_ | new_n11254_;
  assign new_n11256_ = ~pg35 & ng358;
  assign new_n11257_ = ng365 & ng376;
  assign new_n11258_ = ng385 & new_n11257_;
  assign new_n11259_ = ng370 & new_n11258_;
  assign new_n11260_ = new_n11258_ & ~new_n11259_;
  assign new_n11261_ = ng370 & ~new_n11259_;
  assign new_n11262_ = ~new_n11260_ & ~new_n11261_;
  assign new_n11263_ = pg35 & ~new_n11262_;
  assign n3563 = new_n11256_ | new_n11263_;
  assign new_n11265_ = ~pg35 & ng1955;
  assign new_n11266_ = ~new_n6667_1_ & new_n7238_;
  assign new_n11267_ = ng1874 & ~new_n11266_;
  assign new_n11268_ = ~new_n6674_ & new_n11266_;
  assign new_n11269_ = ~new_n11267_ & ~new_n11268_;
  assign new_n11270_ = pg35 & ~new_n11269_;
  assign n3568 = new_n11265_ | new_n11270_;
  assign new_n11272_ = ~pg35 & ng4169;
  assign new_n11273_ = ~ng4125 & ng4165;
  assign new_n11274_ = pg35 & new_n11273_;
  assign n3573 = new_n11272_ | new_n11274_;
  assign new_n11276_ = ~pg35 & ng5475;
  assign new_n11277_ = ng5481 & ~new_n8548_;
  assign new_n11278_ = ng5475 & new_n8548_;
  assign new_n11279_ = ~new_n11277_ & ~new_n11278_;
  assign new_n11280_ = pg35 & ~new_n11279_;
  assign n3578 = new_n11276_ | new_n11280_;
  assign new_n11282_ = ~pg35 & ng2331;
  assign new_n11283_ = ~new_n4724_ & new_n5654_;
  assign new_n11284_ = ~pg113 & new_n11283_;
  assign new_n11285_ = ng112 & new_n11284_;
  assign new_n11286_ = ng2331 & ~new_n11285_;
  assign new_n11287_ = ~new_n7886_ & new_n11286_;
  assign new_n11288_ = ng2361 & new_n7886_;
  assign new_n11289_ = ~new_n11287_ & ~new_n11288_;
  assign new_n11290_ = pg35 & ~new_n11289_;
  assign n3588 = new_n11282_ | new_n11290_;
  assign new_n11292_ = ~pg35 & ng2307;
  assign new_n11293_ = new_n5217_ & new_n7259_;
  assign new_n11294_ = ng2327 & ~new_n11293_;
  assign new_n11295_ = ~ng2287 & ng2331;
  assign new_n11296_ = new_n11293_ & ~new_n11295_;
  assign new_n11297_ = ~new_n11294_ & ~new_n11296_;
  assign new_n11298_ = pg35 & ~new_n11297_;
  assign n3593 = new_n11292_ | new_n11298_;
  assign new_n11300_ = ~pg35 & ng827;
  assign new_n11301_ = ng827 & new_n9053_;
  assign new_n11302_ = ng723 & new_n8009_;
  assign new_n11303_ = ~new_n11301_ & new_n11302_;
  assign new_n11304_ = ~ng723 & new_n8009_;
  assign new_n11305_ = new_n11301_ & new_n11304_;
  assign new_n11306_ = ~new_n11303_ & ~new_n11305_;
  assign new_n11307_ = pg35 & ~new_n11306_;
  assign n3598 = new_n11300_ | new_n11307_;
  assign new_n11309_ = ~pg35 & ng37;
  assign new_n11310_ = n4465 & new_n7615_;
  assign new_n11311_ = ng94 & ~new_n7615_;
  assign new_n11312_ = ~new_n11310_ & ~new_n11311_;
  assign new_n11313_ = pg35 & ~new_n11312_;
  assign n3603 = new_n11309_ | new_n11313_;
  assign new_n11315_ = ~pg35 & ng3698;
  assign new_n11316_ = new_n4743_ & new_n7747_;
  assign new_n11317_ = new_n7431_ & new_n11316_;
  assign new_n11318_ = new_n4735_ & new_n11317_;
  assign new_n11319_ = ~ng3703 & ~new_n11318_;
  assign new_n11320_ = new_n7431_ & new_n11319_;
  assign new_n11321_ = ng3703 & ~new_n7431_;
  assign new_n11322_ = ~new_n11320_ & ~new_n11321_;
  assign new_n11323_ = pg35 & ~new_n11322_;
  assign n3608 = new_n11315_ | new_n11323_;
  assign new_n11325_ = ~pg35 & ng4546;
  assign new_n11326_ = ~ng4575 & new_n8372_;
  assign new_n11327_ = ng4581 & ~new_n11326_;
  assign new_n11328_ = ng4546 & ~ng4581;
  assign new_n11329_ = ~new_n11327_ & ~new_n11328_;
  assign new_n11330_ = pg35 & ~new_n11329_;
  assign n3613 = new_n11325_ | new_n11330_;
  assign new_n11332_ = ~pg35 & ng1932;
  assign new_n11333_ = ~pg113 & new_n5175_;
  assign new_n11334_ = new_n5909_ & new_n11333_;
  assign new_n11335_ = ~ng1917 & ~new_n11334_;
  assign new_n11336_ = new_n8171_ & ~new_n11335_;
  assign new_n11337_ = ng1926 & ~new_n8171_;
  assign new_n11338_ = ~new_n11336_ & ~new_n11337_;
  assign new_n11339_ = pg35 & ~new_n11338_;
  assign n3623 = new_n11332_ | new_n11339_;
  assign new_n11341_ = ~pg35 & ng671;
  assign new_n11342_ = ~ng676 & new_n9930_;
  assign new_n11343_ = new_n9914_ & new_n11342_;
  assign new_n11344_ = ng676 & new_n9930_;
  assign new_n11345_ = ~new_n9914_ & new_n11344_;
  assign new_n11346_ = ~new_n11343_ & ~new_n11345_;
  assign new_n11347_ = pg35 & ~new_n11346_;
  assign n3628 = new_n11341_ | new_n11347_;
  assign new_n11349_ = ~pg35 & ng4555;
  assign new_n11350_ = pg6748 & pg35;
  assign n3633 = new_n11349_ | new_n11350_;
  assign new_n11352_ = ~pg35 & ng4836;
  assign new_n11353_ = ng4836 & ~new_n7605_;
  assign new_n11354_ = pg35 & new_n11353_;
  assign n3638 = new_n11352_ | new_n11354_;
  assign new_n11356_ = ~pg35 & ng1306;
  assign new_n11357_ = ng1521 & ng1500;
  assign new_n11358_ = ng1532 & ~ng1500;
  assign new_n11359_ = ~new_n11357_ & ~new_n11358_;
  assign new_n11360_ = pg35 & ~new_n11359_;
  assign n3643 = new_n11356_ | new_n11360_;
  assign new_n11362_ = ~pg35 & ng1384;
  assign new_n11363_ = ~new_n6294_ & ~new_n6298_;
  assign new_n11364_ = ng1351 & ~ng1384;
  assign new_n11365_ = new_n11363_ & ~new_n11364_;
  assign new_n11366_ = ng1389 & ~new_n11365_;
  assign new_n11367_ = ~ng1389 & ng1351;
  assign new_n11368_ = new_n11365_ & new_n11367_;
  assign new_n11369_ = ~new_n11366_ & ~new_n11368_;
  assign new_n11370_ = pg35 & ~new_n11369_;
  assign n3648 = new_n11362_ | new_n11370_;
  assign new_n11372_ = ~pg35 & ng2250;
  assign new_n11373_ = ~ng2185 & ng2208;
  assign new_n11374_ = new_n9534_ & new_n11373_;
  assign new_n11375_ = ng2255 & ~new_n11374_;
  assign new_n11376_ = ng2250 & ng2246;
  assign new_n11377_ = ng2250 & ~new_n11376_;
  assign new_n11378_ = ng2246 & ~new_n11376_;
  assign new_n11379_ = ~new_n11377_ & ~new_n11378_;
  assign new_n11380_ = new_n11374_ & ~new_n11379_;
  assign new_n11381_ = ~new_n11375_ & ~new_n11380_;
  assign new_n11382_ = pg35 & ~new_n11381_;
  assign n3662 = new_n11372_ | new_n11382_;
  assign new_n11384_ = ~pg35 & ng5495;
  assign new_n11385_ = ng5499 & ~new_n10882_;
  assign new_n11386_ = ng5489 & ~ng5495;
  assign new_n11387_ = ng5489 & ~new_n11386_;
  assign new_n11388_ = ~ng5495 & ~new_n11386_;
  assign new_n11389_ = ~new_n11387_ & ~new_n11388_;
  assign new_n11390_ = new_n10882_ & ~new_n11389_;
  assign new_n11391_ = ~new_n11385_ & ~new_n11390_;
  assign new_n11392_ = pg35 & ~new_n11391_;
  assign n3667 = new_n11384_ | new_n11392_;
  assign new_n11394_ = ~pg35 & ng4180;
  assign new_n11395_ = ng4253 & ng4164;
  assign new_n11396_ = ng4145 & ~ng4253;
  assign new_n11397_ = ~new_n11395_ & ~new_n11396_;
  assign new_n11398_ = pg35 & new_n11397_;
  assign n3672 = new_n11394_ | new_n11398_;
  assign new_n11400_ = ~pg35 & ng5889;
  assign new_n11401_ = new_n7650_ & new_n7995_;
  assign new_n11402_ = ng5917 & ~new_n11401_;
  assign new_n11403_ = ~new_n5966_ & new_n11401_;
  assign new_n11404_ = ~new_n11402_ & ~new_n11403_;
  assign new_n11405_ = pg35 & ~new_n11404_;
  assign n3676 = new_n11400_ | new_n11405_;
  assign new_n11407_ = ~pg35 & ng6163;
  assign new_n11408_ = ng6167 & ~new_n7064_;
  assign new_n11409_ = ~ng6167 & new_n7064_;
  assign new_n11410_ = ~new_n11408_ & ~new_n11409_;
  assign new_n11411_ = pg35 & ~new_n11410_;
  assign n3681 = new_n11407_ | new_n11411_;
  assign new_n11413_ = ~pg35 & ng3889;
  assign new_n11414_ = new_n7124_ & new_n8490_;
  assign new_n11415_ = ng3917 & ~new_n11414_;
  assign new_n11416_ = ~new_n5966_ & new_n11414_;
  assign new_n11417_ = ~new_n11415_ & ~new_n11416_;
  assign new_n11418_ = pg35 & ~new_n11417_;
  assign n3686 = new_n11413_ | new_n11418_;
  assign new_n11420_ = ~pg35 & ng2533;
  assign new_n11421_ = ng2537 & ~new_n9787_;
  assign new_n11422_ = ng2527 & ~ng2533;
  assign new_n11423_ = ng2527 & ~new_n11422_;
  assign new_n11424_ = ~ng2533 & ~new_n11422_;
  assign new_n11425_ = ~new_n11423_ & ~new_n11424_;
  assign new_n11426_ = new_n9787_ & ~new_n11425_;
  assign new_n11427_ = ~new_n11421_ & ~new_n11426_;
  assign new_n11428_ = pg35 & ~new_n11427_;
  assign n3691 = new_n11420_ | new_n11428_;
  assign new_n11430_ = ~pg35 & ng5252;
  assign new_n11431_ = ng5170 & ng5164;
  assign new_n11432_ = new_n5053_ & new_n11431_;
  assign new_n11433_ = ng5268 & ~new_n11432_;
  assign new_n11434_ = ~new_n5966_ & new_n11432_;
  assign new_n11435_ = ~new_n11433_ & ~new_n11434_;
  assign new_n11436_ = pg35 & ~new_n11435_;
  assign n3696 = new_n11430_ | new_n11436_;
  assign new_n11438_ = ~pg35 & ng3416;
  assign new_n11439_ = ~ng3408 & ng3416;
  assign new_n11440_ = ng3423 & new_n11439_;
  assign new_n11441_ = ~ng3412 & ng3416;
  assign new_n11442_ = ~ng3423 & new_n11441_;
  assign new_n11443_ = ~new_n11440_ & ~new_n11442_;
  assign new_n11444_ = pg35 & ~new_n11443_;
  assign n3705 = new_n11438_ | new_n11444_;
  assign new_n11446_ = ~pg35 & ng3873;
  assign new_n11447_ = ng3873 & ng3869;
  assign new_n11448_ = ~ng3881 & ~new_n6204_;
  assign new_n11449_ = new_n11447_ & new_n11448_;
  assign new_n11450_ = ng3881 & ~new_n6204_;
  assign new_n11451_ = ~new_n11447_ & new_n11450_;
  assign new_n11452_ = ~new_n11449_ & ~new_n11451_;
  assign new_n11453_ = pg35 & ~new_n11452_;
  assign n3710 = new_n11446_ | new_n11453_;
  assign new_n11455_ = ~pg35 & ng6109;
  assign new_n11456_ = ng6109 & ng6105;
  assign new_n11457_ = pg35 & new_n11456_;
  assign n3715 = new_n11455_ | new_n11457_;
  assign new_n11459_ = ~pg35 & ng5240;
  assign new_n11460_ = new_n8407_ & new_n11431_;
  assign new_n11461_ = ng5256 & ~new_n11460_;
  assign new_n11462_ = ~new_n5966_ & new_n11460_;
  assign new_n11463_ = ~new_n11461_ & ~new_n11462_;
  assign new_n11464_ = pg35 & ~new_n11463_;
  assign n3720 = new_n11459_ | new_n11464_;
  assign new_n11466_ = ~pg35 & ng5417;
  assign new_n11467_ = ng5413 & ng5417;
  assign new_n11468_ = pg35 & new_n11467_;
  assign n3725 = new_n11466_ | new_n11468_;
  assign new_n11470_ = ~pg35 & ng4727;
  assign new_n11471_ = ng4732 & ~new_n9308_;
  assign new_n11472_ = n3583 & new_n9308_;
  assign new_n11473_ = ~new_n11471_ & ~new_n11472_;
  assign new_n11474_ = pg35 & ~new_n11473_;
  assign n3730 = new_n11470_ | new_n11474_;
  assign new_n11476_ = ~pg35 & ng333;
  assign new_n11477_ = pg35 & ~ng347;
  assign n3735 = new_n11476_ | new_n11477_;
  assign new_n11479_ = ~pg35 & ng2882;
  assign new_n11480_ = n4465 & new_n7895_;
  assign new_n11481_ = pg91 & ~ng2878;
  assign new_n11482_ = ~new_n11480_ & ~new_n11481_;
  assign new_n11483_ = pg35 & new_n11482_;
  assign n3742 = new_n11479_ | new_n11483_;
  assign new_n11485_ = ~pg35 & ng930;
  assign new_n11486_ = ng930 & new_n9836_;
  assign new_n11487_ = ~new_n4686_ & new_n11486_;
  assign new_n11488_ = pg35 & new_n11487_;
  assign n3747 = new_n11485_ | new_n11488_;
  assign new_n11490_ = ~pg35 & ng4146;
  assign new_n11491_ = n2272 & new_n5972_;
  assign new_n11492_ = ng4157 & ~new_n5972_;
  assign new_n11493_ = ~new_n11491_ & ~new_n11492_;
  assign new_n11494_ = pg35 & ~new_n11493_;
  assign n3752 = new_n11490_ | new_n11494_;
  assign new_n11496_ = ~pg35 & ng3857;
  assign new_n11497_ = ng3863 & ~new_n6204_;
  assign new_n11498_ = ~ng3857 & new_n11497_;
  assign new_n11499_ = ~ng3863 & ~new_n6204_;
  assign new_n11500_ = ng3857 & new_n11499_;
  assign new_n11501_ = ~new_n11498_ & ~new_n11500_;
  assign new_n11502_ = pg35 & ~new_n11501_;
  assign n3757 = new_n11496_ | new_n11502_;
  assign new_n11504_ = ~pg35 & ng1664;
  assign new_n11505_ = ~ng1648 & ~new_n11200_;
  assign new_n11506_ = new_n7230_ & ~new_n11505_;
  assign new_n11507_ = ng1657 & ~new_n7230_;
  assign new_n11508_ = ~new_n11506_ & ~new_n11507_;
  assign new_n11509_ = pg35 & ~new_n11508_;
  assign n3767 = new_n11504_ | new_n11509_;
  assign new_n11511_ = ~pg35 & ng3965;
  assign new_n11512_ = new_n6467_ & ~new_n8272_;
  assign new_n11513_ = ng4035 & ~new_n6467_;
  assign new_n11514_ = ~new_n11512_ & ~new_n11513_;
  assign new_n11515_ = pg35 & ~new_n11514_;
  assign n3776 = new_n11511_ | new_n11515_;
  assign new_n11517_ = ~pg35 & ng686;
  assign new_n11518_ = ng686 & new_n6493_1_;
  assign new_n11519_ = ng667 & ~new_n6493_1_;
  assign new_n11520_ = ~new_n11518_ & ~new_n11519_;
  assign new_n11521_ = pg35 & ~new_n11520_;
  assign n3781 = new_n11517_ | new_n11521_;
  assign new_n11523_ = ~pg35 & ng5471;
  assign new_n11524_ = ng5475 & ~new_n10882_;
  assign new_n11525_ = ~ng5475 & new_n10882_;
  assign new_n11526_ = ~new_n11524_ & ~new_n11525_;
  assign new_n11527_ = pg35 & ~new_n11526_;
  assign n3786 = new_n11523_ | new_n11527_;
  assign new_n11529_ = ~pg35 & ng5587;
  assign new_n11530_ = new_n8033_ & new_n10861_;
  assign new_n11531_ = ng5603 & ~new_n11530_;
  assign new_n11532_ = ~new_n5966_ & new_n11530_;
  assign new_n11533_ = ~new_n11531_ & ~new_n11532_;
  assign new_n11534_ = pg35 & ~new_n11533_;
  assign n3791 = new_n11529_ | new_n11534_;
  assign new_n11536_ = ~pg35 & ng2715;
  assign new_n11537_ = ng2715 & ~ng2719;
  assign new_n11538_ = ~ng2715 & ng2719;
  assign new_n11539_ = ~new_n11537_ & ~new_n11538_;
  assign new_n11540_ = ng2841 & ~new_n11539_;
  assign new_n11541_ = ng2841 & ~new_n11540_;
  assign new_n11542_ = pg35 & ~new_n11541_;
  assign n3796 = new_n11536_ | new_n11542_;
  assign new_n11544_ = ~pg35 & ng3933;
  assign new_n11545_ = new_n7124_ & new_n8079_;
  assign new_n11546_ = ng3949 & ~new_n11545_;
  assign new_n11547_ = ~new_n5966_ & new_n11545_;
  assign new_n11548_ = ~new_n11546_ & ~new_n11547_;
  assign new_n11549_ = pg35 & ~new_n11548_;
  assign n3801 = new_n11544_ | new_n11549_;
  assign new_n11551_ = ~pg35 & ng191;
  assign new_n11552_ = ng215 & ng218;
  assign new_n11553_ = ng209 & ~new_n11552_;
  assign new_n11554_ = ng191 & ng194;
  assign new_n11555_ = ng194 & ~new_n11554_;
  assign new_n11556_ = ng191 & ~new_n11554_;
  assign new_n11557_ = ~new_n11555_ & ~new_n11556_;
  assign new_n11558_ = new_n11552_ & ~new_n11557_;
  assign new_n11559_ = ~new_n11553_ & ~new_n11558_;
  assign new_n11560_ = pg35 & ~new_n11559_;
  assign n3806 = new_n11551_ | new_n11560_;
  assign new_n11562_ = ~pg35 & ng4473;
  assign new_n11563_ = ng4473 & ng4462;
  assign new_n11564_ = ~ng4643 & new_n11563_;
  assign new_n11565_ = ~new_n10411_ & ~new_n11564_;
  assign new_n11566_ = ~new_n9227_ & ~new_n9232_;
  assign new_n11567_ = new_n11565_ & new_n11566_;
  assign new_n11568_ = pg35 & ~new_n11567_;
  assign n3811 = new_n11562_ | new_n11568_;
  assign new_n11570_ = ~pg35 & ng4253;
  assign new_n11571_ = n5005 & new_n7806_;
  assign new_n11572_ = ng4249 & ~new_n7806_;
  assign new_n11573_ = ~new_n11571_ & ~new_n11572_;
  assign new_n11574_ = pg35 & ~new_n11573_;
  assign n3816 = new_n11570_ | new_n11574_;
  assign new_n11576_ = ~pg35 & ng5216;
  assign new_n11577_ = ~ng5170 & ng5164;
  assign new_n11578_ = new_n5053_ & new_n11577_;
  assign new_n11579_ = ng5236 & ~new_n11578_;
  assign new_n11580_ = ~new_n5966_ & new_n11578_;
  assign new_n11581_ = ~new_n11579_ & ~new_n11580_;
  assign new_n11582_ = pg35 & ~new_n11581_;
  assign n3821 = new_n11576_ | new_n11582_;
  assign new_n11584_ = ~pg35 & ng4843;
  assign new_n11585_ = ng4849 & new_n7606_;
  assign new_n11586_ = ~new_n7602_ & new_n11585_;
  assign new_n11587_ = ~ng4849 & new_n7606_;
  assign new_n11588_ = new_n7602_ & new_n11587_;
  assign new_n11589_ = ~new_n11586_ & ~new_n11588_;
  assign new_n11590_ = pg35 & ~new_n11589_;
  assign n3829 = new_n11584_ | new_n11590_;
  assign new_n11592_ = ~pg35 & ng2197;
  assign new_n11593_ = ng2197 & ~new_n10082_;
  assign new_n11594_ = ~new_n6522_ & new_n11593_;
  assign new_n11595_ = ng2227 & new_n6522_;
  assign new_n11596_ = ~new_n11594_ & ~new_n11595_;
  assign new_n11597_ = pg35 & ~new_n11596_;
  assign n3839 = new_n11592_ | new_n11597_;
  assign new_n11599_ = ~pg35 & ng6398;
  assign new_n11600_ = ~new_n6602_ & ~new_n6607_;
  assign new_n11601_ = ~ng6411 & ~new_n11600_;
  assign new_n11602_ = ng6411 & new_n6632_1_;
  assign new_n11603_ = new_n11600_ & new_n11602_;
  assign new_n11604_ = ~new_n11601_ & ~new_n11603_;
  assign new_n11605_ = pg35 & ~new_n11604_;
  assign n3844 = new_n11599_ | new_n11605_;
  assign new_n11607_ = ~pg35 & ng5109;
  assign new_n11608_ = ~ng5109 & ng5101;
  assign new_n11609_ = ~ng5062 & ~new_n11608_;
  assign new_n11610_ = ~ng5105 & ~new_n11609_;
  assign new_n11611_ = pg35 & new_n11610_;
  assign n3849 = new_n11607_ | new_n11611_;
  assign new_n11613_ = ~pg35 & ng411;
  assign new_n11614_ = ng424 & ~new_n6067_;
  assign new_n11615_ = ng411 & new_n6067_;
  assign new_n11616_ = ~new_n11614_ & ~new_n11615_;
  assign new_n11617_ = pg35 & ~new_n11616_;
  assign n3859 = new_n11613_ | new_n11617_;
  assign new_n11619_ = ~pg35 & ng1266;
  assign new_n11620_ = ng1570 & ng1280;
  assign new_n11621_ = ~new_n8887_ & new_n11620_;
  assign new_n11622_ = ~ng1280 & new_n8887_;
  assign new_n11623_ = ~new_n11621_ & ~new_n11622_;
  assign new_n11624_ = pg35 & ~new_n11623_;
  assign n3864 = new_n11619_ | new_n11624_;
  assign new_n11626_ = ~pg35 & ng699;
  assign new_n11627_ = ng650 & ~new_n7858_;
  assign new_n11628_ = ng681 & new_n7858_;
  assign new_n11629_ = ~new_n11627_ & ~new_n11628_;
  assign new_n11630_ = pg35 & ~new_n11629_;
  assign n3869 = new_n11626_ | new_n11630_;
  assign new_n11632_ = ~pg35 & ng2169;
  assign new_n11633_ = ~new_n6522_ & new_n9660_;
  assign new_n11634_ = ng2181 & ~new_n11633_;
  assign new_n11635_ = ~new_n6725_ & new_n11633_;
  assign new_n11636_ = ~new_n11634_ & ~new_n11635_;
  assign new_n11637_ = pg35 & ~new_n11636_;
  assign n3874 = new_n11632_ | new_n11637_;
  assign new_n11639_ = ~pg35 & ng1041;
  assign new_n11640_ = new_n10396_ & ~new_n10398_;
  assign new_n11641_ = ng1046 & ~new_n11640_;
  assign new_n11642_ = ~ng1046 & ng1008;
  assign new_n11643_ = new_n11640_ & new_n11642_;
  assign new_n11644_ = ~new_n11641_ & ~new_n11643_;
  assign new_n11645_ = pg35 & ~new_n11644_;
  assign n3879 = new_n11639_ | new_n11645_;
  assign new_n11647_ = ~pg35 & ng1351;
  assign new_n11648_ = ng1345 & new_n6294_;
  assign new_n11649_ = ~new_n6294_ & new_n6307_;
  assign new_n11650_ = ~new_n11648_ & ~new_n11649_;
  assign new_n11651_ = pg35 & ~new_n11650_;
  assign n3884 = new_n11647_ | new_n11651_;
  assign new_n11653_ = ~pg35 & ng5689;
  assign new_n11654_ = ng5689 & new_n6327_;
  assign new_n11655_ = ~ng5698 & ~new_n11654_;
  assign new_n11656_ = pg35 & new_n11655_;
  assign n3889 = new_n11653_ | new_n11656_;
  assign new_n11658_ = ~pg35 & ng2445;
  assign new_n11659_ = ng2495 & ng2421;
  assign new_n11660_ = ~new_n7555_ & new_n11659_;
  assign new_n11661_ = ng2441 & ~new_n11660_;
  assign new_n11662_ = ~new_n8465_ & new_n11660_;
  assign new_n11663_ = ~new_n11661_ & ~new_n11662_;
  assign new_n11664_ = pg35 & ~new_n11663_;
  assign n3894 = new_n11658_ | new_n11664_;
  assign new_n11666_ = ~pg35 & ng5619;
  assign new_n11667_ = new_n7745_ & ~new_n10032_;
  assign new_n11668_ = ng4821 & ~new_n7745_;
  assign new_n11669_ = ~new_n11667_ & ~new_n11668_;
  assign new_n11670_ = pg35 & ~new_n11669_;
  assign n3899 = new_n11666_ | new_n11670_;
  assign new_n11672_ = ~pg35 & ng3689;
  assign new_n11673_ = ng3689 & new_n9026_;
  assign new_n11674_ = ~ng3698 & ~new_n11673_;
  assign new_n11675_ = pg35 & new_n11674_;
  assign n3904 = new_n11672_ | new_n11675_;
  assign new_n11677_ = ~pg35 & ng2767;
  assign new_n11678_ = ~ng1768 & new_n7642_;
  assign new_n11679_ = ~ng2779 & ~new_n11678_;
  assign new_n11680_ = ~new_n7640_ & ~new_n11679_;
  assign new_n11681_ = pg35 & new_n11680_;
  assign n3909 = new_n11677_ | new_n11681_;
  assign new_n11683_ = ~pg35 & ng370;
  assign new_n11684_ = ~ng358 & ~ng376;
  assign new_n11685_ = ~ng358 & ~new_n11684_;
  assign new_n11686_ = ~ng376 & ~new_n11684_;
  assign new_n11687_ = ~new_n11685_ & ~new_n11686_;
  assign new_n11688_ = pg35 & ~new_n11687_;
  assign n3914 = new_n11683_ | new_n11688_;
  assign new_n11690_ = ~pg35 & ng936;
  assign new_n11691_ = ~ng907 & new_n7075_1_;
  assign new_n11692_ = ng907 & ng1227;
  assign new_n11693_ = ~new_n7075_1_ & new_n11692_;
  assign new_n11694_ = ~new_n11691_ & ~new_n11693_;
  assign new_n11695_ = pg35 & ~new_n11694_;
  assign n3919 = new_n11690_ | new_n11695_;
  assign new_n11697_ = ~pg35 & ng681;
  assign new_n11698_ = ng699 & ~new_n6067_;
  assign new_n11699_ = ~new_n7858_ & new_n11698_;
  assign new_n11700_ = ~new_n7858_ & ~new_n11699_;
  assign new_n11701_ = pg35 & ~new_n11700_;
  assign n3924 = new_n11697_ | new_n11701_;
  assign new_n11703_ = ~pg35 & ng3125;
  assign new_n11704_ = ng3129 & ~new_n10989_;
  assign new_n11705_ = ng3119 & ~ng3125;
  assign new_n11706_ = ng3119 & ~new_n11705_;
  assign new_n11707_ = ~ng3125 & ~new_n11705_;
  assign new_n11708_ = ~new_n11706_ & ~new_n11707_;
  assign new_n11709_ = new_n10989_ & ~new_n11708_;
  assign new_n11710_ = ~new_n11704_ & ~new_n11709_;
  assign new_n11711_ = pg35 & ~new_n11710_;
  assign n3929 = new_n11703_ | new_n11711_;
  assign new_n11713_ = ~pg35 & ng4704;
  assign new_n11714_ = ~new_n8500_ & ~new_n10481_;
  assign new_n11715_ = ng4704 & ~new_n8500_;
  assign new_n11716_ = ~new_n8503_ & ~new_n11715_;
  assign new_n11717_ = ~new_n11714_ & ~new_n11716_;
  assign new_n11718_ = ng4698 & new_n11714_;
  assign new_n11719_ = ~new_n11717_ & ~new_n11718_;
  assign new_n11720_ = pg35 & ~new_n11719_;
  assign n3934 = new_n11713_ | new_n11720_;
  assign new_n11722_ = ~pg35 & ng6031;
  assign new_n11723_ = ng6035 & ~new_n6452_;
  assign new_n11724_ = ~ng6035 & new_n6452_;
  assign new_n11725_ = ~new_n11723_ & ~new_n11724_;
  assign new_n11726_ = pg35 & ~new_n11725_;
  assign n3939 = new_n11722_ | new_n11726_;
  assign new_n11728_ = pg35 & ~ng70;
  assign new_n11729_ = ~pg35 & ~new_n11728_;
  assign new_n11730_ = ng4473 & ~ng4459;
  assign new_n11731_ = ng4507 & ~new_n11730_;
  assign new_n11732_ = pg113 & new_n11730_;
  assign new_n11733_ = ~new_n11731_ & ~new_n11732_;
  assign new_n11734_ = pg35 & ~new_n11733_;
  assign n3944 = new_n11729_ | new_n11734_;
  assign new_n11736_ = ~pg35 & ng4031;
  assign new_n11737_ = ng4040 & ~new_n6172_;
  assign new_n11738_ = ~ng4040 & new_n6172_;
  assign new_n11739_ = ~new_n11737_ & ~new_n11738_;
  assign new_n11740_ = pg35 & ~new_n11739_;
  assign n3949 = new_n11736_ | new_n11740_;
  assign new_n11742_ = ~pg35 & ng3376;
  assign new_n11743_ = ~new_n10780_ & ~new_n10785_;
  assign new_n11744_ = ng3380 & new_n8400_;
  assign new_n11745_ = new_n11743_ & new_n11744_;
  assign new_n11746_ = ~ng3380 & ~new_n11743_;
  assign new_n11747_ = ~new_n11745_ & ~new_n11746_;
  assign new_n11748_ = pg35 & ~new_n11747_;
  assign n3954 = new_n11742_ | new_n11748_;
  assign new_n11750_ = ~pg35 & ng5559;
  assign new_n11751_ = ng5535 & ~ng5527;
  assign new_n11752_ = new_n8035_ & new_n11751_;
  assign new_n11753_ = ng5555 & ~new_n11752_;
  assign new_n11754_ = ~new_n5966_ & new_n11752_;
  assign new_n11755_ = ~new_n11753_ & ~new_n11754_;
  assign new_n11756_ = pg35 & ~new_n11755_;
  assign n3959 = new_n11750_ | new_n11756_;
  assign new_n11758_ = ~pg35 & ng582;
  assign new_n11759_ = ~ng590 & new_n6564_;
  assign new_n11760_ = ng590 & ~new_n6545_;
  assign new_n11761_ = ~new_n6564_ & new_n11760_;
  assign new_n11762_ = ~new_n11759_ & ~new_n11761_;
  assign new_n11763_ = pg35 & ~new_n11762_;
  assign n3964 = new_n11758_ | new_n11763_;
  assign new_n11765_ = ~pg35 & ng1756;
  assign new_n11766_ = ~new_n6236_ & new_n6686_;
  assign new_n11767_ = ng1752 & ~new_n11766_;
  assign new_n11768_ = ~new_n10679_ & new_n11766_;
  assign new_n11769_ = ~new_n11767_ & ~new_n11768_;
  assign new_n11770_ = pg35 & ~new_n11769_;
  assign n3969 = new_n11765_ | new_n11770_;
  assign new_n11772_ = ~pg35 & ng4474;
  assign new_n11773_ = pg35 & ng4474;
  assign n3974 = new_n11772_ | new_n11773_;
  assign new_n11775_ = ~pg35 & ng1291;
  assign new_n11776_ = n4465 & new_n8829_;
  assign new_n11777_ = ng1306 & ~ng1296;
  assign new_n11778_ = ~new_n11776_ & ~new_n11777_;
  assign new_n11779_ = pg35 & new_n11778_;
  assign n3979 = new_n11775_ | new_n11779_;
  assign new_n11781_ = ~pg35 & ng4388;
  assign new_n11782_ = ng4375 & ~ng4382;
  assign new_n11783_ = ~ng4375 & ng4382;
  assign new_n11784_ = ~new_n11782_ & ~new_n11783_;
  assign new_n11785_ = ~new_n7684_ & ~new_n11784_;
  assign new_n11786_ = ~new_n9894_ & ~new_n11785_;
  assign new_n11787_ = pg35 & ~new_n11786_;
  assign n3984 = new_n11781_ | new_n11787_;
  assign new_n11789_ = pg35 & ng1070;
  assign new_n11790_ = ~pg35 & new_n11789_;
  assign new_n11791_ = ~ng1052 & ~new_n7672_;
  assign new_n11792_ = ~new_n7673_ & ~new_n11791_;
  assign new_n11793_ = ~ng979 & new_n11792_;
  assign new_n11794_ = pg35 & new_n11793_;
  assign n3989 = new_n11790_ | new_n11794_;
  assign new_n11796_ = pg35 & ng1724;
  assign new_n11797_ = ~pg35 & new_n11796_;
  assign new_n11798_ = ng1728 & ~ng1802;
  assign new_n11799_ = ~ng1772 & ~ng1802;
  assign new_n11800_ = ~new_n11798_ & ~new_n11799_;
  assign new_n11801_ = ~new_n6239_ & ~new_n11800_;
  assign new_n11802_ = ~new_n6236_ & new_n11801_;
  assign new_n11803_ = ng1728 & new_n6236_;
  assign new_n11804_ = ~new_n11802_ & ~new_n11803_;
  assign new_n11805_ = pg35 & ~new_n11804_;
  assign n3994 = new_n11797_ | new_n11805_;
  assign new_n11807_ = pg35 & ng976;
  assign new_n11808_ = ~pg35 & new_n11807_;
  assign new_n11809_ = ng969 & new_n5940_1_;
  assign new_n11810_ = new_n5939_ & new_n5942_;
  assign new_n11811_ = ~ng1008 & new_n11810_;
  assign new_n11812_ = ~ng1046 & new_n6132_;
  assign new_n11813_ = ng1008 & new_n11812_;
  assign new_n11814_ = ng969 & new_n5939_;
  assign new_n11815_ = ~new_n11811_ & ~new_n11813_;
  assign new_n11816_ = ~new_n6134_1_ & ~new_n11814_;
  assign new_n11817_ = new_n11815_ & new_n11816_;
  assign new_n11818_ = ~new_n5940_1_ & ~new_n11817_;
  assign new_n11819_ = ~new_n11809_ & ~new_n11818_;
  assign new_n11820_ = pg35 & ~new_n11819_;
  assign n3999 = new_n11808_ | new_n11820_;
  assign new_n11822_ = ~pg35 & ng351;
  assign new_n11823_ = ~ng351 & ~new_n6361_;
  assign new_n11824_ = pg35 & new_n11823_;
  assign n4004 = new_n11822_ | new_n11824_;
  assign new_n11826_ = ~pg35 & ng6444;
  assign new_n11827_ = pg35 & ng6727;
  assign n4014 = new_n11826_ | new_n11827_;
  assign new_n11829_ = ~pg35 & ng872;
  assign new_n11830_ = ng859 & new_n6112_;
  assign new_n11831_ = ng225 & ~new_n6112_;
  assign new_n11832_ = ~new_n11830_ & ~new_n11831_;
  assign new_n11833_ = pg35 & ~new_n11832_;
  assign n4018 = new_n11829_ | new_n11833_;
  assign new_n11835_ = ~pg35 & ng5863;
  assign new_n11836_ = ~pg113 & new_n5775_;
  assign new_n11837_ = ~new_n4724_ & new_n11836_;
  assign new_n11838_ = ng43 & new_n11837_;
  assign new_n11839_ = ~ng5869 & ~new_n11838_;
  assign new_n11840_ = new_n8646_ & new_n11839_;
  assign new_n11841_ = ng5869 & new_n11839_;
  assign new_n11842_ = ~new_n8646_ & new_n11841_;
  assign new_n11843_ = ~new_n11840_ & ~new_n11842_;
  assign new_n11844_ = pg35 & ~new_n11843_;
  assign n4023 = new_n11835_ | new_n11844_;
  assign new_n11846_ = ~pg35 & ng150;
  assign new_n11847_ = ~ng153 & new_n6282_;
  assign new_n11848_ = ng153 & new_n6276_;
  assign new_n11849_ = ~new_n6282_ & new_n11848_;
  assign new_n11850_ = ~new_n11847_ & ~new_n11849_;
  assign new_n11851_ = pg35 & ~new_n11850_;
  assign n4028 = new_n11846_ | new_n11851_;
  assign new_n11853_ = ~pg35 & ng2799;
  assign new_n11854_ = ~ng2327 & new_n7642_;
  assign new_n11855_ = ~ng2811 & ~new_n11854_;
  assign new_n11856_ = ~new_n7640_ & ~new_n11855_;
  assign new_n11857_ = pg35 & new_n11856_;
  assign n4033 = new_n11853_ | new_n11857_;
  assign new_n11859_ = ~pg35 & ng4098;
  assign new_n11860_ = ng4108 & ~new_n10835_;
  assign new_n11861_ = ~ng4108 & new_n10835_;
  assign new_n11862_ = ~new_n11860_ & ~new_n11861_;
  assign new_n11863_ = ng4169 & ~new_n11862_;
  assign new_n11864_ = ng4169 & ~new_n11863_;
  assign new_n11865_ = pg35 & ~new_n11864_;
  assign n4047 = new_n11859_ | new_n11865_;
  assign new_n11867_ = ~pg35 & ng5873;
  assign new_n11868_ = ng5869 & ng5873;
  assign new_n11869_ = ~ng5881 & ~new_n11838_;
  assign new_n11870_ = new_n11868_ & new_n11869_;
  assign new_n11871_ = ng5881 & ~new_n11838_;
  assign new_n11872_ = ~new_n11868_ & new_n11871_;
  assign new_n11873_ = ~new_n11870_ & ~new_n11872_;
  assign new_n11874_ = pg35 & ~new_n11873_;
  assign n4052 = new_n11867_ | new_n11874_;
  assign new_n11876_ = pg35 & ng1046;
  assign new_n11877_ = ~pg35 & new_n11876_;
  assign new_n11878_ = ng1146 & ~new_n7772_;
  assign new_n11879_ = ng1146 & ~ng1152;
  assign new_n11880_ = ng1099 & ~new_n11879_;
  assign new_n11881_ = new_n7772_ & ~new_n11880_;
  assign new_n11882_ = ~new_n11878_ & ~new_n11881_;
  assign new_n11883_ = pg35 & ~new_n11882_;
  assign n4057 = new_n11877_ | new_n11883_;
  assign new_n11885_ = ~pg35 & ng513;
  assign new_n11886_ = ng513 & ~new_n6494_;
  assign new_n11887_ = new_n6493_1_ & new_n11886_;
  assign new_n11888_ = ng518 & ~new_n6493_1_;
  assign new_n11889_ = ~new_n11887_ & ~new_n11888_;
  assign new_n11890_ = pg35 & ~new_n11889_;
  assign n4062 = new_n11885_ | new_n11890_;
  assign new_n11892_ = ~pg35 & ng66;
  assign new_n11893_ = ~ng4340 & ~ng4349;
  assign new_n11894_ = ~ng4358 & new_n11893_;
  assign new_n11895_ = ng4643 & new_n5621_;
  assign new_n11896_ = new_n11894_ & new_n11895_;
  assign new_n11897_ = pg35 & new_n11896_;
  assign n4067 = new_n11892_ | new_n11897_;
  assign new_n11899_ = ~pg35 & ng3040;
  assign new_n11900_ = ~ng3029 & new_n8930_;
  assign new_n11901_ = ~ng3034 & new_n11900_;
  assign new_n11902_ = ~ng3040 & new_n11901_;
  assign new_n11903_ = ng3029 & new_n8934_;
  assign new_n11904_ = ng3034 & new_n11903_;
  assign new_n11905_ = ng3040 & new_n11904_;
  assign new_n11906_ = ~new_n11902_ & ~new_n11905_;
  assign new_n11907_ = ~ng3045 & ~new_n11906_;
  assign new_n11908_ = ng3045 & new_n8954_;
  assign new_n11909_ = new_n11906_ & new_n11908_;
  assign new_n11910_ = ~new_n11907_ & ~new_n11909_;
  assign new_n11911_ = pg35 & ~new_n11910_;
  assign n4072 = new_n11899_ | new_n11911_;
  assign new_n11913_ = ~pg35 & ng464;
  assign new_n11914_ = ng468 & ~new_n5994_;
  assign new_n11915_ = ng464 & new_n5994_;
  assign new_n11916_ = ~new_n11914_ & ~new_n11915_;
  assign new_n11917_ = pg35 & ~new_n11916_;
  assign n4077 = new_n11913_ | new_n11917_;
  assign new_n11919_ = ~pg35 & ng5037;
  assign new_n11920_ = ~new_n8139_ & ~new_n8144_;
  assign new_n11921_ = ng5041 & new_n8107_;
  assign new_n11922_ = new_n11920_ & new_n11921_;
  assign new_n11923_ = ~ng5041 & ~new_n11920_;
  assign new_n11924_ = ~new_n11922_ & ~new_n11923_;
  assign new_n11925_ = pg35 & ~new_n11924_;
  assign n4082 = new_n11919_ | new_n11925_;
  assign new_n11927_ = ~pg35 & ng2994;
  assign new_n11928_ = n2287 & new_n8526_;
  assign new_n11929_ = ng2988 & ~new_n8526_;
  assign new_n11930_ = ~new_n11928_ & ~new_n11929_;
  assign new_n11931_ = pg35 & ~new_n11930_;
  assign n4087 = new_n11927_ | new_n11931_;
  assign new_n11933_ = ~pg35 & ng1514;
  assign new_n11934_ = ng1514 & ng1500;
  assign new_n11935_ = ~ng1526 & new_n6843_;
  assign new_n11936_ = ~new_n11934_ & ~new_n11935_;
  assign new_n11937_ = ng1526 & new_n6843_;
  assign new_n11938_ = new_n11934_ & ~new_n11937_;
  assign new_n11939_ = ~new_n11936_ & ~new_n11938_;
  assign new_n11940_ = pg35 & ~new_n11939_;
  assign n4092 = new_n11933_ | new_n11940_;
  assign new_n11942_ = ~pg35 & ng562;
  assign new_n11943_ = ng568 & ~new_n6545_;
  assign new_n11944_ = ~new_n6547_1_ & new_n11943_;
  assign new_n11945_ = ~ng568 & new_n6547_1_;
  assign new_n11946_ = ~new_n11944_ & ~new_n11945_;
  assign new_n11947_ = pg35 & ~new_n11946_;
  assign n4097 = new_n11942_ | new_n11947_;
  assign new_n11949_ = ~pg35 & ng4239;
  assign new_n11950_ = ~ng4297 & ~ng4294;
  assign new_n11951_ = pg35 & new_n11950_;
  assign n4102 = new_n11949_ | new_n11951_;
  assign new_n11953_ = ~pg35 & ng3454;
  assign new_n11954_ = ~ng3454 & ng3447;
  assign new_n11955_ = ~ng3361 & ~new_n11954_;
  assign new_n11956_ = ~ng3443 & ~new_n11955_;
  assign new_n11957_ = pg35 & new_n11956_;
  assign n4106 = new_n11953_ | new_n11957_;
  assign new_n11959_ = ~pg35 & ng4567;
  assign new_n11960_ = ~ng4578 & new_n8372_;
  assign new_n11961_ = ng4581 & ~new_n11960_;
  assign new_n11962_ = ~ng4581 & ng4567;
  assign new_n11963_ = ~new_n11961_ & ~new_n11962_;
  assign new_n11964_ = pg35 & ~new_n11963_;
  assign n4111 = new_n11959_ | new_n11964_;
  assign new_n11966_ = ~pg35 & ng3068;
  assign new_n11967_ = ng3065 & ~ng3057;
  assign new_n11968_ = ~ng3068 & ~new_n11967_;
  assign new_n11969_ = ~ng3072 & new_n11968_;
  assign new_n11970_ = ng3072 & ng3068;
  assign new_n11971_ = ~ng3061 & ng3065;
  assign new_n11972_ = ~new_n11969_ & ~new_n11970_;
  assign new_n11973_ = ~new_n11971_ & new_n11972_;
  assign new_n11974_ = pg35 & ~new_n11973_;
  assign n4116 = new_n11966_ | new_n11974_;
  assign new_n11976_ = ~pg35 & ng6148;
  assign new_n11977_ = ~ng6148 & ng6140;
  assign new_n11978_ = ~ng6098 & ~new_n11977_;
  assign new_n11979_ = ~ng6144 & ~new_n11978_;
  assign new_n11980_ = pg35 & new_n11979_;
  assign n4121 = new_n11976_ | new_n11980_;
  assign new_n11982_ = ~pg35 & ng6267;
  assign new_n11983_ = new_n7865_ & new_n9573_;
  assign new_n11984_ = ng6283 & ~new_n11983_;
  assign new_n11985_ = ~new_n5966_ & new_n11983_;
  assign new_n11986_ = ~new_n11984_ & ~new_n11985_;
  assign new_n11987_ = pg35 & ~new_n11986_;
  assign n4126 = new_n11982_ | new_n11987_;
  assign new_n11989_ = ~pg35 & ng6411;
  assign new_n11990_ = ~new_n6603_ & ~new_n6608_;
  assign new_n11991_ = ng6415 & new_n6632_1_;
  assign new_n11992_ = new_n11990_ & new_n11991_;
  assign new_n11993_ = ~ng6415 & ~new_n11990_;
  assign new_n11994_ = ~new_n11992_ & ~new_n11993_;
  assign new_n11995_ = pg35 & ~new_n11994_;
  assign n4131 = new_n11989_ | new_n11995_;
  assign new_n11997_ = ~pg35 & ng5156;
  assign new_n11998_ = ng5120 & ~pg26801;
  assign new_n11999_ = ng5156 & pg26801;
  assign new_n12000_ = ~new_n11998_ & ~new_n11999_;
  assign new_n12001_ = pg35 & ~new_n12000_;
  assign n4136 = new_n11997_ | new_n12001_;
  assign new_n12003_ = ~pg35 & ng1333;
  assign new_n12004_ = ng1322 & ~ng1579;
  assign new_n12005_ = ~ng1579 & ~new_n12004_;
  assign new_n12006_ = ng1322 & ~new_n12004_;
  assign new_n12007_ = ~new_n12005_ & ~new_n12006_;
  assign new_n12008_ = new_n8879_ & new_n12007_;
  assign new_n12009_ = ng1333 & new_n12008_;
  assign new_n12010_ = ng1333 & ~new_n12009_;
  assign new_n12011_ = new_n12008_ & ~new_n12009_;
  assign new_n12012_ = ~new_n12010_ & ~new_n12011_;
  assign new_n12013_ = pg35 & ~new_n12012_;
  assign n4141 = new_n12003_ | new_n12013_;
  assign new_n12015_ = ~pg35 & ng4311;
  assign new_n12016_ = ~ng4322 & new_n5874_;
  assign new_n12017_ = new_n5866_ & new_n12016_;
  assign new_n12018_ = ng4322 & new_n5874_;
  assign new_n12019_ = ~new_n5866_ & new_n12018_;
  assign new_n12020_ = ~new_n12017_ & ~new_n12019_;
  assign new_n12021_ = pg35 & ~new_n12020_;
  assign n4146 = new_n12015_ | new_n12021_;
  assign new_n12023_ = ~pg35 & ng5236;
  assign new_n12024_ = new_n5053_ & new_n7581_;
  assign new_n12025_ = ng5252 & ~new_n12024_;
  assign new_n12026_ = ~new_n5966_ & new_n12024_;
  assign new_n12027_ = ~new_n12025_ & ~new_n12026_;
  assign new_n12028_ = pg35 & ~new_n12027_;
  assign n4151 = new_n12023_ | new_n12028_;
  assign new_n12030_ = ~pg35 & ng1270;
  assign new_n12031_ = ng1570 & ng1274;
  assign new_n12032_ = ~new_n9072_ & new_n12031_;
  assign new_n12033_ = ~ng1274 & new_n9072_;
  assign new_n12034_ = ~new_n12032_ & ~new_n12033_;
  assign new_n12035_ = pg35 & ~new_n12034_;
  assign n4156 = new_n12030_ | new_n12035_;
  assign new_n12037_ = ~new_n5661_ & pg34383;
  assign new_n12038_ = new_n5661_ & ~new_n5726_;
  assign n4161 = new_n12037_ | new_n12038_;
  assign new_n12040_ = ~pg35 & ng5029;
  assign new_n12041_ = ~new_n8137_ & ~new_n8142_;
  assign new_n12042_ = ng5033 & new_n8107_;
  assign new_n12043_ = new_n12041_ & new_n12042_;
  assign new_n12044_ = ~ng5033 & ~new_n12041_;
  assign new_n12045_ = ~new_n12043_ & ~new_n12044_;
  assign new_n12046_ = pg35 & ~new_n12045_;
  assign n4166 = new_n12040_ | new_n12046_;
  assign new_n12048_ = pg35 & ng4888;
  assign new_n12049_ = ~pg35 & new_n12048_;
  assign new_n12050_ = new_n5676_ & new_n5742_1_;
  assign new_n12051_ = ~ng3343 & ~ng3288;
  assign new_n12052_ = ~ng3352 & new_n12051_;
  assign new_n12053_ = ng3343 & ng3288;
  assign new_n12054_ = ~ng3352 & new_n12053_;
  assign new_n12055_ = ~ng3288 & ~ng3347;
  assign new_n12056_ = ng3352 & new_n12055_;
  assign new_n12057_ = ng3288 & ng3347;
  assign new_n12058_ = ng3352 & new_n12057_;
  assign new_n12059_ = ~new_n12052_ & ~new_n12054_;
  assign new_n12060_ = ~new_n12056_ & ~new_n12058_;
  assign new_n12061_ = new_n12059_ & new_n12060_;
  assign new_n12062_ = ~ng4939 & new_n12061_;
  assign new_n12063_ = new_n12050_ & ~new_n12062_;
  assign new_n12064_ = new_n6915_ & new_n12063_;
  assign new_n12065_ = ng4939 & ~new_n6915_;
  assign new_n12066_ = ~new_n12064_ & ~new_n12065_;
  assign new_n12067_ = pg35 & ~new_n12066_;
  assign n4171 = new_n12049_ | new_n12067_;
  assign new_n12069_ = ~pg35 & ng5092;
  assign new_n12070_ = ng5097 & ~new_n9273_;
  assign new_n12071_ = ~ng5097 & new_n9273_;
  assign new_n12072_ = ~new_n12070_ & ~new_n12071_;
  assign new_n12073_ = pg35 & ~new_n12072_;
  assign n4176 = new_n12069_ | new_n12073_;
  assign new_n12075_ = ~pg35 & ng3396;
  assign new_n12076_ = ~new_n8393_ & ~new_n8397_;
  assign new_n12077_ = pg35 & new_n12076_;
  assign n4185 = new_n12075_ | new_n12077_;
  assign new_n12079_ = ~pg35 & ng939;
  assign new_n12080_ = n2272 & new_n6861_;
  assign new_n12081_ = ~ng943 & new_n4686_;
  assign new_n12082_ = ~new_n12080_ & ~new_n12081_;
  assign new_n12083_ = pg35 & new_n12082_;
  assign n4195 = new_n12079_ | new_n12083_;
  assign new_n12085_ = ~pg35 & ng5204;
  assign new_n12086_ = new_n7580_1_ & new_n8995_;
  assign new_n12087_ = ng5200 & ~new_n12086_;
  assign new_n12088_ = ~new_n5966_ & new_n12086_;
  assign new_n12089_ = ~new_n12087_ & ~new_n12088_;
  assign new_n12090_ = pg35 & ~new_n12089_;
  assign n4200 = new_n12085_ | new_n12090_;
  assign new_n12092_ = ~pg35 & ng2907;
  assign new_n12093_ = n3583 & new_n9379_;
  assign new_n12094_ = ng2912 & ~new_n9379_;
  assign new_n12095_ = ~new_n12093_ & ~new_n12094_;
  assign new_n12096_ = pg35 & ~new_n12095_;
  assign n4205 = new_n12092_ | new_n12096_;
  assign new_n12098_ = ~pg35 & ng3347;
  assign new_n12099_ = new_n6915_ & new_n7748_;
  assign new_n12100_ = new_n4735_ & new_n12099_;
  assign new_n12101_ = ~ng3352 & ~new_n12100_;
  assign new_n12102_ = new_n6915_ & new_n12101_;
  assign new_n12103_ = ng3352 & ~new_n6915_;
  assign new_n12104_ = ~new_n12102_ & ~new_n12103_;
  assign new_n12105_ = pg35 & ~new_n12104_;
  assign n4210 = new_n12098_ | new_n12105_;
  assign new_n12107_ = ~pg35 & ng3119;
  assign new_n12108_ = ng3125 & ~new_n10989_;
  assign new_n12109_ = ng3119 & new_n10989_;
  assign new_n12110_ = ~new_n12108_ & ~new_n12109_;
  assign new_n12111_ = pg35 & ~new_n12110_;
  assign n4215 = new_n12107_ | new_n12111_;
  assign new_n12113_ = ~pg35 & ng1982;
  assign new_n12114_ = ng1988 & ~new_n8172_;
  assign new_n12115_ = ng1982 & new_n8172_;
  assign new_n12116_ = ~new_n12114_ & ~new_n12115_;
  assign new_n12117_ = pg35 & ~new_n12116_;
  assign n4220 = new_n12113_ | new_n12117_;
  assign new_n12119_ = ~pg35 & ng5343;
  assign new_n12120_ = ng5320 & ng5313;
  assign new_n12121_ = ng5290 & ng5276;
  assign new_n12122_ = new_n12120_ & new_n12121_;
  assign new_n12123_ = ng5343 & new_n12122_;
  assign new_n12124_ = ~ng5352 & ~new_n12123_;
  assign new_n12125_ = pg35 & new_n12124_;
  assign n4225 = new_n12119_ | new_n12125_;
  assign new_n12127_ = ~pg35 & ng4455;
  assign n4230 = new_n9897_ | new_n12127_;
  assign new_n12129_ = ~pg35 & ng1870;
  assign new_n12130_ = ~ng1936 & ng1906;
  assign new_n12131_ = ~new_n6667_1_ & new_n12130_;
  assign new_n12132_ = ng1878 & ~new_n12131_;
  assign new_n12133_ = ~new_n6674_ & new_n12131_;
  assign new_n12134_ = ~new_n12132_ & ~new_n12133_;
  assign new_n12135_ = pg35 & ~new_n12134_;
  assign n4235 = new_n12129_ | new_n12135_;
  assign new_n12137_ = ~pg35 & ng2541;
  assign new_n12138_ = ng2547 & ~new_n9421_;
  assign new_n12139_ = ng2541 & new_n9421_;
  assign new_n12140_ = ~new_n12138_ & ~new_n12139_;
  assign new_n12141_ = pg35 & ~new_n12140_;
  assign n4240 = new_n12137_ | new_n12141_;
  assign new_n12143_ = ~pg35 & ng5339;
  assign new_n12144_ = ng5343 & ~new_n12122_;
  assign new_n12145_ = ~ng5343 & new_n12122_;
  assign new_n12146_ = ~new_n12144_ & ~new_n12145_;
  assign new_n12147_ = pg35 & ~new_n12146_;
  assign n4245 = new_n12143_ | new_n12147_;
  assign new_n12149_ = ng22 & pg34921;
  assign new_n12150_ = ~ng22 & n2287;
  assign n4250 = new_n12149_ | new_n12150_;
  assign new_n12152_ = ~pg35 & ng5611;
  assign new_n12153_ = ng5523 & new_n11751_;
  assign new_n12154_ = ng5567 & ~new_n12153_;
  assign new_n12155_ = ~new_n5966_ & new_n12153_;
  assign new_n12156_ = ~new_n12154_ & ~new_n12155_;
  assign new_n12157_ = pg35 & ~new_n12156_;
  assign n4259 = new_n12152_ | new_n12157_;
  assign new_n12159_ = ~pg35 & ng1246;
  assign new_n12160_ = ~ng1083 & ng1233;
  assign new_n12161_ = ng1083 & ng1227;
  assign new_n12162_ = ~new_n12160_ & ~new_n12161_;
  assign new_n12163_ = pg35 & ~new_n12162_;
  assign n4264 = new_n12159_ | new_n12163_;
  assign new_n12165_ = ~pg35 & ng732;
  assign new_n12166_ = ng732 & new_n5996_;
  assign new_n12167_ = ng753 & ~new_n5996_;
  assign new_n12168_ = ~new_n12166_ & ~new_n12167_;
  assign new_n12169_ = pg35 & ~new_n12168_;
  assign n4269 = new_n12165_ | new_n12169_;
  assign new_n12171_ = ~pg35 & ng347;
  assign new_n12172_ = ~ng347 & ng344;
  assign new_n12173_ = pg35 & new_n12172_;
  assign n4274 = new_n12171_ | new_n12173_;
  assign new_n12175_ = ~pg35 & ng3171;
  assign new_n12176_ = ng3171 & ng3167;
  assign new_n12177_ = ~ng3179 & ~new_n6249_;
  assign new_n12178_ = new_n12176_ & new_n12177_;
  assign new_n12179_ = ng3179 & ~new_n6249_;
  assign new_n12180_ = ~new_n12176_ & new_n12179_;
  assign new_n12181_ = ~new_n12178_ & ~new_n12180_;
  assign new_n12182_ = pg35 & ~new_n12181_;
  assign n4284 = new_n12175_ | new_n12182_;
  assign new_n12184_ = ~pg35 & ng2815;
  assign new_n12185_ = ng2807 & ~new_n8663_;
  assign new_n12186_ = ng2811 & ~new_n5870_;
  assign new_n12187_ = ~new_n6045_1_ & ~new_n12186_;
  assign new_n12188_ = new_n8663_ & new_n12187_;
  assign new_n12189_ = ~new_n12185_ & ~new_n12188_;
  assign new_n12190_ = pg35 & ~new_n12189_;
  assign n4289 = new_n12184_ | new_n12190_;
  assign new_n12192_ = ~pg35 & ng1668;
  assign new_n12193_ = ng1682 & ~new_n10845_;
  assign new_n12194_ = ng1246 & new_n7536_;
  assign new_n12195_ = ~new_n7541_ & ~new_n12194_;
  assign new_n12196_ = new_n12193_ & ~new_n12195_;
  assign new_n12197_ = new_n12193_ & ~new_n12196_;
  assign new_n12198_ = ~new_n12195_ & ~new_n12196_;
  assign new_n12199_ = ~new_n12197_ & ~new_n12198_;
  assign new_n12200_ = ~new_n7537_1_ & ~new_n12199_;
  assign new_n12201_ = ng1682 & new_n7537_1_;
  assign new_n12202_ = ~new_n12200_ & ~new_n12201_;
  assign new_n12203_ = pg35 & ~new_n12202_;
  assign n4294 = new_n12192_ | new_n12203_;
  assign new_n12205_ = ~pg35 & ng5827;
  assign new_n12206_ = ng5831 & ~new_n6354_;
  assign new_n12207_ = ~ng5827 & ng5821;
  assign new_n12208_ = ng5821 & ~new_n12207_;
  assign new_n12209_ = ~ng5827 & ~new_n12207_;
  assign new_n12210_ = ~new_n12208_ & ~new_n12209_;
  assign new_n12211_ = new_n6354_ & ~new_n12210_;
  assign new_n12212_ = ~new_n12206_ & ~new_n12211_;
  assign new_n12213_ = pg35 & ~new_n12212_;
  assign n4299 = new_n12205_ | new_n12213_;
  assign new_n12215_ = ~pg35 & ng3215;
  assign new_n12216_ = new_n5963_ & new_n9368_;
  assign new_n12217_ = ng3231 & ~new_n12216_;
  assign new_n12218_ = ~new_n5966_ & new_n12216_;
  assign new_n12219_ = ~new_n12217_ & ~new_n12218_;
  assign new_n12220_ = pg35 & ~new_n12219_;
  assign n4304 = new_n12215_ | new_n12220_;
  assign new_n12222_ = ~pg35 & ng4483;
  assign n4309 = new_n11350_ | new_n12222_;
  assign new_n12224_ = ~pg35 & ng5555;
  assign new_n12225_ = new_n7566_1_ & new_n11751_;
  assign new_n12226_ = ng5579 & ~new_n12225_;
  assign new_n12227_ = ~new_n5966_ & new_n12225_;
  assign new_n12228_ = ~new_n12226_ & ~new_n12227_;
  assign new_n12229_ = pg35 & ~new_n12228_;
  assign n4314 = new_n12224_ | new_n12229_;
  assign new_n12231_ = ~pg35 & ng6609;
  assign new_n12232_ = ng6555 & ~ng6549;
  assign new_n12233_ = new_n10108_ & new_n12232_;
  assign new_n12234_ = ng6625 & ~new_n12233_;
  assign new_n12235_ = ~new_n5966_ & new_n12233_;
  assign new_n12236_ = ~new_n12234_ & ~new_n12235_;
  assign new_n12237_ = pg35 & ~new_n12236_;
  assign n4319 = new_n12231_ | new_n12237_;
  assign new_n12239_ = ~pg35 & ng3752;
  assign new_n12240_ = pg35 & ng4040;
  assign n4324 = new_n12239_ | new_n12240_;
  assign new_n12242_ = ~pg35 & ng4401;
  assign new_n12243_ = ng4401 & new_n7684_;
  assign new_n12244_ = ng4392 & new_n12243_;
  assign new_n12245_ = ~ng4411 & ~new_n12244_;
  assign new_n12246_ = pg35 & ~new_n12245_;
  assign n4329 = new_n12242_ | new_n12246_;
  assign new_n12248_ = ~pg35 & ng4561;
  assign new_n12249_ = pg6750 & pg35;
  assign n4334 = new_n12248_ | new_n12249_;
  assign new_n12251_ = ~pg35 & ng5381;
  assign new_n12252_ = ~ng5381 & new_n6370_;
  assign new_n12253_ = ng5381 & new_n6373_;
  assign new_n12254_ = ~new_n12252_ & ~new_n12253_;
  assign new_n12255_ = ng5385 & new_n6394_;
  assign new_n12256_ = new_n12254_ & new_n12255_;
  assign new_n12257_ = ~ng5385 & ~new_n12254_;
  assign new_n12258_ = ~new_n12256_ & ~new_n12257_;
  assign new_n12259_ = pg35 & ~new_n12258_;
  assign n4343 = new_n12251_ | new_n12259_;
  assign new_n12261_ = ~pg35 & ng2610;
  assign new_n12262_ = ~new_n4724_ & new_n10307_;
  assign new_n12263_ = new_n10306_ & new_n12262_;
  assign new_n12264_ = ~ng2610 & ng2619;
  assign new_n12265_ = ng110 & new_n12264_;
  assign new_n12266_ = ng110 & ~new_n12265_;
  assign new_n12267_ = new_n12264_ & ~new_n12265_;
  assign new_n12268_ = ~new_n12266_ & ~new_n12267_;
  assign new_n12269_ = new_n12263_ & ~new_n12268_;
  assign new_n12270_ = ng2625 & ~new_n12263_;
  assign new_n12271_ = ~new_n12269_ & ~new_n12270_;
  assign new_n12272_ = pg35 & ~new_n12271_;
  assign n4348 = new_n12261_ | new_n12272_;
  assign new_n12274_ = ~pg35 & ng3949;
  assign new_n12275_ = ng3869 & new_n7124_;
  assign new_n12276_ = ng3897 & ~new_n12275_;
  assign new_n12277_ = ~new_n5966_ & new_n12275_;
  assign new_n12278_ = ~new_n12276_ & ~new_n12277_;
  assign new_n12279_ = pg35 & ~new_n12278_;
  assign n4353 = new_n12274_ | new_n12279_;
  assign new_n12281_ = ~pg35 & ng2852;
  assign new_n12282_ = n5814 & new_n5972_;
  assign new_n12283_ = ng2860 & ~new_n5972_;
  assign new_n12284_ = ~new_n12282_ & ~new_n12283_;
  assign new_n12285_ = pg35 & ~new_n12284_;
  assign n4358 = new_n12281_ | new_n12285_;
  assign new_n12287_ = ~pg35 & ng6625;
  assign new_n12288_ = new_n7159_ & new_n10108_;
  assign new_n12289_ = ng6641 & ~new_n12288_;
  assign new_n12290_ = ~new_n5966_ & new_n12288_;
  assign new_n12291_ = ~new_n12289_ & ~new_n12290_;
  assign new_n12292_ = pg35 & ~new_n12291_;
  assign n4363 = new_n12287_ | new_n12292_;
  assign new_n12294_ = ~pg35 & ng5390;
  assign new_n12295_ = ~ng5385 & new_n12252_;
  assign new_n12296_ = ~ng5390 & new_n12295_;
  assign new_n12297_ = ng5385 & new_n12253_;
  assign new_n12298_ = ng5390 & new_n12297_;
  assign new_n12299_ = ~new_n12296_ & ~new_n12298_;
  assign new_n12300_ = ng5396 & new_n6394_;
  assign new_n12301_ = new_n12299_ & new_n12300_;
  assign new_n12302_ = ~ng5396 & ~new_n12299_;
  assign new_n12303_ = ~new_n12301_ & ~new_n12302_;
  assign new_n12304_ = pg35 & ~new_n12303_;
  assign n4368 = new_n12294_ | new_n12304_;
  assign n4373 = ~pg35 & ng2145;
  assign new_n12307_ = ~pg35 & ng3530;
  assign new_n12308_ = ~ng3506 & ~ng3512;
  assign new_n12309_ = ~ng3518 & new_n12308_;
  assign new_n12310_ = new_n11130_ & new_n12309_;
  assign new_n12311_ = ng3538 & ~new_n12310_;
  assign new_n12312_ = ~new_n5966_ & new_n12310_;
  assign new_n12313_ = ~new_n12311_ & ~new_n12312_;
  assign new_n12314_ = pg35 & ~new_n12313_;
  assign n4378 = new_n12307_ | new_n12314_;
  assign new_n12316_ = ~pg35 & ng6519;
  assign new_n12317_ = ng6523 & ~new_n7219_;
  assign new_n12318_ = ~ng6519 & ng6513;
  assign new_n12319_ = ng6513 & ~new_n12318_;
  assign new_n12320_ = ~ng6519 & ~new_n12318_;
  assign new_n12321_ = ~new_n12319_ & ~new_n12320_;
  assign new_n12322_ = new_n7219_ & ~new_n12321_;
  assign new_n12323_ = ~new_n12317_ & ~new_n12322_;
  assign new_n12324_ = pg35 & ~new_n12323_;
  assign n4383 = new_n12316_ | new_n12324_;
  assign new_n12326_ = ~pg35 & ng3259;
  assign new_n12327_ = ng3263 & ~new_n7152_;
  assign new_n12328_ = ~new_n5966_ & new_n7152_;
  assign new_n12329_ = ~new_n12327_ & ~new_n12328_;
  assign new_n12330_ = pg35 & ~new_n12329_;
  assign n4388 = new_n12326_ | new_n12330_;
  assign new_n12332_ = ~pg35 & ng3606;
  assign new_n12333_ = ng3518 & new_n10352_;
  assign new_n12334_ = ng3562 & ~new_n12333_;
  assign new_n12335_ = ~new_n5966_ & new_n12333_;
  assign new_n12336_ = ~new_n12334_ & ~new_n12335_;
  assign new_n12337_ = pg35 & ~new_n12336_;
  assign n4393 = new_n12332_ | new_n12337_;
  assign new_n12339_ = ~pg35 & ng5921;
  assign new_n12340_ = ~ng5857 & ng5863;
  assign new_n12341_ = new_n7649_ & new_n12340_;
  assign new_n12342_ = ng5937 & ~new_n12341_;
  assign new_n12343_ = ~new_n5966_ & new_n12341_;
  assign new_n12344_ = ~new_n12342_ & ~new_n12343_;
  assign new_n12345_ = pg35 & ~new_n12344_;
  assign n4402 = new_n12339_ | new_n12345_;
  assign new_n12347_ = pg35 & ng4754;
  assign new_n12348_ = ~pg35 & new_n12347_;
  assign new_n12349_ = ~ng6386 & ~ng6336;
  assign new_n12350_ = ~ng6395 & new_n12349_;
  assign new_n12351_ = ng6386 & ng6336;
  assign new_n12352_ = ~ng6395 & new_n12351_;
  assign new_n12353_ = ~ng6336 & ~ng6390;
  assign new_n12354_ = ng6395 & new_n12353_;
  assign new_n12355_ = ng6336 & ng6390;
  assign new_n12356_ = ng6395 & new_n12355_;
  assign new_n12357_ = ~new_n12350_ & ~new_n12352_;
  assign new_n12358_ = ~new_n12354_ & ~new_n12356_;
  assign new_n12359_ = new_n12357_ & new_n12358_;
  assign new_n12360_ = ~ng4771 & new_n12359_;
  assign new_n12361_ = new_n8498_ & ~new_n12360_;
  assign new_n12362_ = new_n6699_ & new_n12361_;
  assign new_n12363_ = ng4771 & ~new_n6699_;
  assign new_n12364_ = ~new_n12362_ & ~new_n12363_;
  assign new_n12365_ = pg35 & ~new_n12364_;
  assign n4412 = new_n12348_ | new_n12365_;
  assign new_n12367_ = ~pg35 & ng4991;
  assign new_n12368_ = ng4991 & new_n11039_;
  assign new_n12369_ = ng4966 & new_n11040_;
  assign new_n12370_ = ~new_n12368_ & new_n12369_;
  assign new_n12371_ = ~ng4966 & new_n11040_;
  assign new_n12372_ = new_n12368_ & new_n12371_;
  assign new_n12373_ = ~new_n12370_ & ~new_n12372_;
  assign new_n12374_ = pg35 & ~new_n12373_;
  assign n4420 = new_n12367_ | new_n12374_;
  assign new_n12376_ = ~pg35 & ng1193;
  assign new_n12377_ = ~ng1199 & new_n5953_;
  assign new_n12378_ = new_n8812_ & new_n12377_;
  assign new_n12379_ = ng1199 & new_n5953_;
  assign new_n12380_ = ~new_n8812_ & new_n12379_;
  assign new_n12381_ = ~new_n12378_ & ~new_n12380_;
  assign new_n12382_ = pg35 & ~new_n12381_;
  assign n4429 = new_n12376_ | new_n12382_;
  assign new_n12384_ = ~pg35 & ng5925;
  assign new_n12385_ = new_n9330_ & new_n12340_;
  assign new_n12386_ = ng5941 & ~new_n12385_;
  assign new_n12387_ = ~new_n5966_ & new_n12385_;
  assign new_n12388_ = ~new_n12386_ & ~new_n12387_;
  assign new_n12389_ = pg35 & ~new_n12388_;
  assign n4434 = new_n12384_ | new_n12389_;
  assign new_n12391_ = ~pg35 & ng1146;
  assign new_n12392_ = ng1152 & ~new_n7772_;
  assign new_n12393_ = ng1146 & new_n7772_;
  assign new_n12394_ = ~new_n12392_ & ~new_n12393_;
  assign new_n12395_ = pg35 & ~new_n12394_;
  assign n4439 = new_n12391_ | new_n12395_;
  assign new_n12397_ = ~pg35 & ng2848;
  assign new_n12398_ = n3583 & new_n7895_;
  assign new_n12399_ = ~ng2856 & new_n4867_1_;
  assign new_n12400_ = ~new_n12398_ & ~new_n12399_;
  assign new_n12401_ = pg35 & new_n12400_;
  assign n4447 = new_n12397_ | new_n12401_;
  assign new_n12403_ = ~pg35 & ng990;
  assign new_n12404_ = ng990 & new_n7417_1_;
  assign new_n12405_ = ng990 & ~new_n12404_;
  assign new_n12406_ = new_n7417_1_ & ~new_n12404_;
  assign new_n12407_ = ~new_n12405_ & ~new_n12406_;
  assign new_n12408_ = pg35 & ~new_n12407_;
  assign n4456 = new_n12403_ | new_n12408_;
  assign new_n12410_ = ~pg35 & ng1959;
  assign new_n12411_ = new_n8171_ & new_n9091_;
  assign new_n12412_ = ng1964 & ~new_n12411_;
  assign new_n12413_ = ng1959 & ng1955;
  assign new_n12414_ = ng1959 & ~new_n12413_;
  assign new_n12415_ = ng1955 & ~new_n12413_;
  assign new_n12416_ = ~new_n12414_ & ~new_n12415_;
  assign new_n12417_ = new_n12411_ & ~new_n12416_;
  assign new_n12418_ = ~new_n12412_ & ~new_n12417_;
  assign new_n12419_ = pg35 & ~new_n12418_;
  assign n4460 = new_n12410_ | new_n12419_;
  assign new_n12421_ = ~pg35 & ng5396;
  assign new_n12422_ = ~ng5396 & new_n12296_;
  assign new_n12423_ = ng5396 & new_n12298_;
  assign new_n12424_ = ~new_n12422_ & ~new_n12423_;
  assign new_n12425_ = ~ng5401 & ~new_n12424_;
  assign new_n12426_ = ng5401 & new_n6394_;
  assign new_n12427_ = new_n12424_ & new_n12426_;
  assign new_n12428_ = ~new_n12425_ & ~new_n12427_;
  assign new_n12429_ = pg35 & ~new_n12428_;
  assign n4470 = new_n12421_ | new_n12429_;
  assign new_n12431_ = ~pg35 & ng5164;
  assign new_n12432_ = ng5170 & ~new_n7369_1_;
  assign new_n12433_ = ~ng5164 & new_n12432_;
  assign new_n12434_ = ~ng5170 & ~new_n7369_1_;
  assign new_n12435_ = ng5164 & new_n12434_;
  assign new_n12436_ = ~new_n12433_ & ~new_n12435_;
  assign new_n12437_ = pg35 & ~new_n12436_;
  assign n4475 = new_n12431_ | new_n12437_;
  assign new_n12439_ = ~pg35 & ng1564;
  assign new_n12440_ = ng1548 & ng1430;
  assign new_n12441_ = ng1564 & new_n12440_;
  assign new_n12442_ = ng1559 & ~new_n8877_;
  assign new_n12443_ = ~new_n12441_ & new_n12442_;
  assign new_n12444_ = ~ng1559 & ~new_n8877_;
  assign new_n12445_ = new_n12441_ & new_n12444_;
  assign new_n12446_ = ~new_n12443_ & ~new_n12445_;
  assign new_n12447_ = pg35 & ~new_n12446_;
  assign n4480 = new_n12439_ | new_n12447_;
  assign new_n12449_ = ~pg35 & ng4878;
  assign new_n12450_ = ~ng4843 & new_n7606_;
  assign new_n12451_ = ng4878 & new_n12450_;
  assign new_n12452_ = ng4843 & new_n7606_;
  assign new_n12453_ = ~ng4878 & new_n12452_;
  assign new_n12454_ = ~new_n12451_ & ~new_n12453_;
  assign new_n12455_ = pg35 & ~new_n12454_;
  assign n4485 = new_n12449_ | new_n12455_;
  assign new_n12457_ = ~pg35 & ng6653;
  assign new_n12458_ = ng6657 & ~new_n7390_;
  assign new_n12459_ = ~new_n5966_ & new_n7390_;
  assign new_n12460_ = ~new_n12458_ & ~new_n12459_;
  assign new_n12461_ = pg35 & ~new_n12460_;
  assign n4494 = new_n12457_ | new_n12461_;
  assign new_n12463_ = ~pg35 & ng2860;
  assign new_n12464_ = n2287 & new_n5972_;
  assign new_n12465_ = ng2894 & ~new_n5972_;
  assign new_n12466_ = ~new_n12464_ & ~new_n12465_;
  assign new_n12467_ = pg35 & ~new_n12466_;
  assign n4499 = new_n12463_ | new_n12467_;
  assign new_n12469_ = pg35 & ng4531;
  assign new_n12470_ = ~pg35 & new_n12469_;
  assign new_n12471_ = ~ng4311 & new_n5874_;
  assign new_n12472_ = new_n5865_ & new_n12471_;
  assign new_n12473_ = ng4311 & new_n5874_;
  assign new_n12474_ = ~new_n5865_ & new_n12473_;
  assign new_n12475_ = ~new_n12472_ & ~new_n12474_;
  assign new_n12476_ = pg35 & ~new_n12475_;
  assign n4504 = new_n12470_ | new_n12476_;
  assign new_n12478_ = ~pg35 & ng3199;
  assign new_n12479_ = new_n8744_ & new_n9315_;
  assign new_n12480_ = ng3223 & ~new_n12479_;
  assign new_n12481_ = ~new_n5966_ & new_n12479_;
  assign new_n12482_ = ~new_n12480_ & ~new_n12481_;
  assign new_n12483_ = pg35 & ~new_n12482_;
  assign n4509 = new_n12478_ | new_n12483_;
  assign new_n12485_ = ~pg35 & ng3235;
  assign new_n12486_ = new_n5962_ & new_n9338_;
  assign new_n12487_ = ng3251 & ~new_n12486_;
  assign new_n12488_ = ~new_n5966_ & new_n12486_;
  assign new_n12489_ = ~new_n12487_ & ~new_n12488_;
  assign new_n12490_ = pg35 & ~new_n12489_;
  assign n4514 = new_n12485_ | new_n12490_;
  assign new_n12492_ = ~pg35 & ng5615;
  assign new_n12493_ = ng5619 & ~new_n10882_;
  assign new_n12494_ = ~new_n5966_ & new_n10882_;
  assign new_n12495_ = ~new_n12493_ & ~new_n12494_;
  assign new_n12496_ = pg35 & ~new_n12495_;
  assign n4519 = new_n12492_ | new_n12496_;
  assign new_n12498_ = ~pg35 & ng807;
  assign new_n12499_ = ~new_n6578_ & new_n8625_;
  assign new_n12500_ = ng790 & new_n12499_;
  assign new_n12501_ = ng794 & new_n12500_;
  assign new_n12502_ = ~new_n6578_ & new_n12501_;
  assign new_n12503_ = ~new_n6578_ & new_n12502_;
  assign new_n12504_ = ng807 & new_n12503_;
  assign new_n12505_ = ~ng554 & new_n12504_;
  assign new_n12506_ = ng554 & ~new_n6578_;
  assign new_n12507_ = ~new_n12504_ & new_n12506_;
  assign new_n12508_ = ~new_n12505_ & ~new_n12507_;
  assign new_n12509_ = pg35 & ~new_n12508_;
  assign n4529 = new_n12498_ | new_n12509_;
  assign new_n12511_ = ~pg35 & ng1783;
  assign new_n12512_ = ~new_n4724_ & new_n6731_1_;
  assign new_n12513_ = new_n6683_ & new_n12512_;
  assign new_n12514_ = ng110 & new_n6809_;
  assign new_n12515_ = ng110 & ~new_n12514_;
  assign new_n12516_ = new_n6809_ & ~new_n12514_;
  assign new_n12517_ = ~new_n12515_ & ~new_n12516_;
  assign new_n12518_ = new_n12513_ & ~new_n12517_;
  assign new_n12519_ = ng1798 & ~new_n12513_;
  assign new_n12520_ = ~new_n12518_ & ~new_n12519_;
  assign new_n12521_ = pg35 & ~new_n12520_;
  assign n4534 = new_n12511_ | new_n12521_;
  assign new_n12523_ = ~pg35 & ng4864;
  assign new_n12524_ = ng4864 & ~new_n7605_;
  assign new_n12525_ = pg35 & new_n12524_;
  assign n4539 = new_n12523_ | new_n12525_;
  assign new_n12527_ = ~pg35 & ng4633;
  assign new_n12528_ = ng4633 & ng4621;
  assign new_n12529_ = new_n8339_ & new_n12528_;
  assign new_n12530_ = ~ng4639 & new_n12529_;
  assign new_n12531_ = pg35 & new_n12530_;
  assign n4549 = new_n12527_ | new_n12531_;
  assign new_n12533_ = ~pg35 & ng2886;
  assign new_n12534_ = new_n4945_1_ & new_n10889_;
  assign new_n12535_ = ~ng34 & ~ng2980;
  assign new_n12536_ = ~new_n12534_ & ~new_n12535_;
  assign new_n12537_ = pg35 & new_n12536_;
  assign n4554 = new_n12533_ | new_n12537_;
  assign new_n12539_ = ~pg35 & ng5905;
  assign new_n12540_ = new_n7997_ & new_n9330_;
  assign new_n12541_ = ng5901 & ~new_n12540_;
  assign new_n12542_ = ~new_n5966_ & new_n12540_;
  assign new_n12543_ = ~new_n12541_ & ~new_n12542_;
  assign new_n12544_ = pg35 & ~new_n12543_;
  assign n4559 = new_n12539_ | new_n12544_;
  assign new_n12546_ = pg35 & ng468;
  assign new_n12547_ = ~pg35 & new_n12546_;
  assign new_n12548_ = ng174 & new_n6270_1_;
  assign new_n12549_ = ng182 & ng203;
  assign new_n12550_ = new_n12548_ & new_n12549_;
  assign new_n12551_ = ng168 & new_n6270_1_;
  assign new_n12552_ = new_n12549_ & new_n12551_;
  assign new_n12553_ = ng168 & ng174;
  assign new_n12554_ = new_n6271_ & new_n12553_;
  assign new_n12555_ = ~new_n12550_ & ~new_n12552_;
  assign new_n12556_ = ~new_n12554_ & new_n12555_;
  assign new_n12557_ = pg35 & ~new_n12556_;
  assign n4564 = new_n12547_ | new_n12557_;
  assign new_n12559_ = ~pg35 & ng4688;
  assign new_n12560_ = ~ng4653 & new_n10528_;
  assign new_n12561_ = ng4688 & new_n12560_;
  assign new_n12562_ = ng4653 & new_n10528_;
  assign new_n12563_ = ~ng4688 & new_n12562_;
  assign new_n12564_ = ~new_n12561_ & ~new_n12563_;
  assign new_n12565_ = pg35 & ~new_n12564_;
  assign n4569 = new_n12559_ | new_n12565_;
  assign new_n12567_ = ~pg35 & ng5421;
  assign new_n12568_ = ~ng5413 & ng5421;
  assign new_n12569_ = ng5428 & new_n12568_;
  assign new_n12570_ = ng5421 & ~ng5417;
  assign new_n12571_ = ~ng5428 & new_n12570_;
  assign new_n12572_ = ~new_n12569_ & ~new_n12571_;
  assign new_n12573_ = pg35 & ~new_n12572_;
  assign n4574 = new_n12567_ | new_n12573_;
  assign new_n12575_ = ~pg35 & ng1111;
  assign new_n12576_ = ng1116 & new_n5950_1_;
  assign new_n12577_ = new_n5888_1_ & new_n12576_;
  assign new_n12578_ = ng1105 & ng1111;
  assign new_n12579_ = ng1105 & ~new_n12578_;
  assign new_n12580_ = ng1111 & ~new_n12578_;
  assign new_n12581_ = ~new_n12579_ & ~new_n12580_;
  assign new_n12582_ = new_n12577_ & ~new_n12581_;
  assign new_n12583_ = ng1105 & ~new_n12577_;
  assign new_n12584_ = ~new_n12582_ & ~new_n12583_;
  assign new_n12585_ = pg35 & ~new_n12584_;
  assign n4579 = new_n12575_ | new_n12585_;
  assign new_n12587_ = ~pg35 & ng3881;
  assign new_n12588_ = new_n6896_ & new_n7124_;
  assign new_n12589_ = ng3889 & ~new_n12588_;
  assign new_n12590_ = ~new_n5966_ & new_n12588_;
  assign new_n12591_ = ~new_n12589_ & ~new_n12590_;
  assign new_n12592_ = pg35 & ~new_n12591_;
  assign n4584 = new_n12587_ | new_n12592_;
  assign new_n12594_ = ~pg35 & ng4093;
  assign new_n12595_ = ~ng4098 & new_n10834_;
  assign new_n12596_ = ng4098 & ~new_n10834_;
  assign new_n12597_ = ~new_n12595_ & ~new_n12596_;
  assign new_n12598_ = ng4169 & ~new_n12597_;
  assign new_n12599_ = ng4169 & ~new_n12598_;
  assign new_n12600_ = pg35 & ~new_n12599_;
  assign n4589 = new_n12594_ | new_n12600_;
  assign new_n12602_ = ~pg35 & ng4501;
  assign new_n12603_ = ~ng59 & new_n8372_;
  assign new_n12604_ = ng4581 & ~new_n12603_;
  assign new_n12605_ = ng4501 & ~ng4581;
  assign new_n12606_ = ~new_n12604_ & ~new_n12605_;
  assign new_n12607_ = pg35 & ~new_n12606_;
  assign n4594 = new_n12602_ | new_n12607_;
  assign new_n12609_ = ~pg35 & ng1585;
  assign new_n12610_ = pg35 & ng1570;
  assign n4599 = new_n12609_ | new_n12610_;
  assign new_n12612_ = ~pg35 & ng6049;
  assign new_n12613_ = ng6049 & new_n6353_;
  assign new_n12614_ = new_n6353_ & new_n11316_;
  assign new_n12615_ = new_n4734_ & new_n12614_;
  assign new_n12616_ = ng5990 & ~new_n12615_;
  assign new_n12617_ = ~new_n12613_ & new_n12616_;
  assign new_n12618_ = ~ng5990 & ~new_n12615_;
  assign new_n12619_ = new_n12613_ & new_n12618_;
  assign new_n12620_ = ~new_n12617_ & ~new_n12619_;
  assign new_n12621_ = pg35 & ~new_n12620_;
  assign n4604 = new_n12612_ | new_n12621_;
  assign new_n12623_ = ~pg35 & ng6255;
  assign new_n12624_ = new_n7063_ & new_n7866_;
  assign new_n12625_ = ng6275 & ~new_n12624_;
  assign new_n12626_ = ~new_n5966_ & new_n12624_;
  assign new_n12627_ = ~new_n12625_ & ~new_n12626_;
  assign new_n12628_ = pg35 & ~new_n12627_;
  assign n4613 = new_n12623_ | new_n12628_;
  assign new_n12630_ = ~pg35 & ng6243;
  assign new_n12631_ = new_n7088_ & new_n7865_;
  assign new_n12632_ = ng6239 & ~new_n12631_;
  assign new_n12633_ = ~new_n5966_ & new_n12631_;
  assign new_n12634_ = ~new_n12632_ & ~new_n12633_;
  assign new_n12635_ = pg35 & ~new_n12634_;
  assign n4618 = new_n12630_ | new_n12635_;
  assign new_n12637_ = ~pg35 & ng5456;
  assign new_n12638_ = ng5448 & ~ng5456;
  assign new_n12639_ = ~ng5406 & ~new_n12638_;
  assign new_n12640_ = ~ng5452 & ~new_n12639_;
  assign new_n12641_ = pg35 & new_n12640_;
  assign n4628 = new_n12637_ | new_n12641_;
  assign new_n12643_ = ~pg35 & ng164;
  assign new_n12644_ = ng150 & new_n6276_;
  assign new_n12645_ = ~new_n6280_1_ & new_n12644_;
  assign new_n12646_ = ~ng150 & new_n6280_1_;
  assign new_n12647_ = ~new_n12645_ & ~new_n12646_;
  assign new_n12648_ = pg35 & ~new_n12647_;
  assign n4633 = new_n12643_ | new_n12648_;
  assign new_n12650_ = pg35 & ng554;
  assign new_n12651_ = ~pg35 & new_n12650_;
  assign new_n12652_ = new_n4910_ & new_n8183_;
  assign new_n12653_ = ~ng209 & ~ng538;
  assign new_n12654_ = ~new_n12652_ & ~new_n12653_;
  assign new_n12655_ = pg35 & new_n12654_;
  assign n4638 = new_n12651_ | new_n12655_;
  assign new_n12657_ = ~pg35 & ng4749;
  assign new_n12658_ = new_n5667_ & new_n5836_;
  assign new_n12659_ = ~new_n8500_ & ~new_n12658_;
  assign new_n12660_ = ng4749 & ~new_n8500_;
  assign new_n12661_ = ~new_n8503_ & ~new_n12660_;
  assign new_n12662_ = ~new_n12659_ & ~new_n12661_;
  assign new_n12663_ = ng4743 & new_n12659_;
  assign new_n12664_ = ~new_n12662_ & ~new_n12663_;
  assign new_n12665_ = pg35 & ~new_n12664_;
  assign n4643 = new_n12657_ | new_n12665_;
  assign new_n12667_ = ~pg35 & ng5543;
  assign new_n12668_ = new_n7566_1_ & new_n8033_;
  assign new_n12669_ = ng5571 & ~new_n12668_;
  assign new_n12670_ = ~new_n5966_ & new_n12668_;
  assign new_n12671_ = ~new_n12669_ & ~new_n12670_;
  assign new_n12672_ = pg35 & ~new_n12671_;
  assign n4648 = new_n12667_ | new_n12672_;
  assign new_n12674_ = ~pg35 & ng5188;
  assign new_n12675_ = new_n8407_ & new_n8995_;
  assign new_n12676_ = ng5196 & ~new_n12675_;
  assign new_n12677_ = ~new_n5966_ & new_n12675_;
  assign new_n12678_ = ~new_n12676_ & ~new_n12677_;
  assign new_n12679_ = pg35 & ~new_n12678_;
  assign n4653 = new_n12674_ | new_n12679_;
  assign new_n12681_ = ~pg35 & ng2357;
  assign new_n12682_ = ~ng2342 & ~new_n10344_;
  assign new_n12683_ = new_n7259_ & ~new_n12682_;
  assign new_n12684_ = ng2351 & ~new_n7259_;
  assign new_n12685_ = ~new_n12683_ & ~new_n12684_;
  assign new_n12686_ = pg35 & ~new_n12685_;
  assign n4658 = new_n12681_ | new_n12686_;
  assign new_n12688_ = ~pg35 & ng4452;
  assign new_n12689_ = ng4430 & new_n10730_;
  assign new_n12690_ = ~ng4452 & ~new_n12689_;
  assign new_n12691_ = pg35 & ~new_n12690_;
  assign n4663 = new_n12688_ | new_n12691_;
  assign new_n12693_ = ~pg35 & ng160;
  assign new_n12694_ = ng160 & new_n6286_;
  assign new_n12695_ = pg35 & new_n12694_;
  assign n4668 = new_n12693_ | new_n12695_;
  assign new_n12697_ = pg35 & ng203;
  assign new_n12698_ = ~pg35 & new_n12697_;
  assign new_n12699_ = ng370 & ng376;
  assign new_n12700_ = ng365 & ~ng385;
  assign new_n12701_ = new_n12699_ & new_n12700_;
  assign new_n12702_ = ng854 & ~new_n12701_;
  assign new_n12703_ = ng174 & ~ng392;
  assign new_n12704_ = ng452 & ng392;
  assign new_n12705_ = ~new_n12703_ & ~new_n12704_;
  assign new_n12706_ = ng182 & ~new_n12705_;
  assign new_n12707_ = ~ng182 & new_n12705_;
  assign new_n12708_ = ~new_n12706_ & ~new_n12707_;
  assign new_n12709_ = ng411 & ~ng392;
  assign new_n12710_ = ng441 & ng392;
  assign new_n12711_ = ~new_n12709_ & ~new_n12710_;
  assign new_n12712_ = ~ng417 & new_n12711_;
  assign new_n12713_ = new_n12708_ & new_n12712_;
  assign new_n12714_ = ~ng691 & new_n12713_;
  assign new_n12715_ = ~ng405 & ~ng392;
  assign new_n12716_ = ng424 & new_n12715_;
  assign new_n12717_ = ng405 & ng392;
  assign new_n12718_ = ng392 & ~new_n12717_;
  assign new_n12719_ = ng405 & ~new_n12717_;
  assign new_n12720_ = ~new_n12718_ & ~new_n12719_;
  assign new_n12721_ = ng437 & ~new_n12720_;
  assign new_n12722_ = ~new_n12716_ & ~new_n12721_;
  assign new_n12723_ = ng401 & new_n12717_;
  assign new_n12724_ = new_n12722_ & ~new_n12723_;
  assign new_n12725_ = ng417 & ~new_n12724_;
  assign new_n12726_ = ng417 & ~new_n12725_;
  assign new_n12727_ = ~new_n12724_ & ~new_n12725_;
  assign new_n12728_ = ~new_n12726_ & ~new_n12727_;
  assign new_n12729_ = ~new_n12714_ & ~new_n12728_;
  assign new_n12730_ = new_n12701_ & ~new_n12729_;
  assign new_n12731_ = ~new_n12702_ & ~new_n12730_;
  assign new_n12732_ = pg35 & ~new_n12731_;
  assign n4673 = new_n12698_ | new_n12732_;
  assign new_n12734_ = ~pg35 & ng2504;
  assign new_n12735_ = ng2476 & ~ng2453;
  assign new_n12736_ = ng2518 & ~new_n12735_;
  assign new_n12737_ = ng2504 & new_n12736_;
  assign new_n12738_ = new_n12736_ & ~new_n12737_;
  assign new_n12739_ = ng2504 & ~new_n12737_;
  assign new_n12740_ = ~new_n12738_ & ~new_n12739_;
  assign new_n12741_ = new_n5907_1_ & ~new_n12740_;
  assign new_n12742_ = ng2518 & ~new_n5907_1_;
  assign new_n12743_ = ~new_n12741_ & ~new_n12742_;
  assign new_n12744_ = pg35 & ~new_n12743_;
  assign n4678 = new_n12734_ | new_n12744_;
  assign new_n12746_ = ~pg35 & ng4608;
  assign new_n12747_ = ng4584 & new_n8849_;
  assign new_n12748_ = ng4593 & new_n12747_;
  assign new_n12749_ = ng4601 & new_n12748_;
  assign new_n12750_ = ng4608 & new_n12749_;
  assign new_n12751_ = ~ng4616 & new_n8853_;
  assign new_n12752_ = new_n12750_ & new_n12751_;
  assign new_n12753_ = ng4616 & new_n8853_;
  assign new_n12754_ = ~new_n12750_ & new_n12753_;
  assign new_n12755_ = ~new_n12752_ & ~new_n12754_;
  assign new_n12756_ = pg35 & ~new_n12755_;
  assign n4696 = new_n12746_ | new_n12756_;
  assign new_n12758_ = ~pg35 & ng2518;
  assign new_n12759_ = new_n5907_1_ & new_n12735_;
  assign new_n12760_ = ng2523 & ~new_n12759_;
  assign new_n12761_ = ng2518 & ng2514;
  assign new_n12762_ = ng2518 & ~new_n12761_;
  assign new_n12763_ = ng2514 & ~new_n12761_;
  assign new_n12764_ = ~new_n12762_ & ~new_n12763_;
  assign new_n12765_ = new_n12759_ & ~new_n12764_;
  assign new_n12766_ = ~new_n12760_ & ~new_n12765_;
  assign new_n12767_ = pg35 & ~new_n12766_;
  assign n4701 = new_n12758_ | new_n12767_;
  assign new_n12769_ = ~pg35 & ng2547;
  assign new_n12770_ = ng2551 & ~new_n9421_;
  assign new_n12771_ = ng2541 & ~ng2547;
  assign new_n12772_ = ng2541 & ~new_n12771_;
  assign new_n12773_ = ~ng2547 & ~new_n12771_;
  assign new_n12774_ = ~new_n12772_ & ~new_n12773_;
  assign new_n12775_ = new_n9421_ & ~new_n12774_;
  assign new_n12776_ = ~new_n12770_ & ~new_n12775_;
  assign new_n12777_ = pg35 & ~new_n12776_;
  assign n4706 = new_n12769_ | new_n12777_;
  assign new_n12779_ = ~pg35 & ng2583;
  assign new_n12780_ = ~new_n7174_ & new_n10910_;
  assign new_n12781_ = ng2579 & ~new_n12780_;
  assign new_n12782_ = ~new_n8484_ & new_n12780_;
  assign new_n12783_ = ~new_n12781_ & ~new_n12782_;
  assign new_n12784_ = pg35 & ~new_n12783_;
  assign n4714 = new_n12779_ | new_n12784_;
  assign new_n12786_ = ~pg35 & ng3909;
  assign new_n12787_ = new_n7010_ & new_n8490_;
  assign new_n12788_ = ng3929 & ~new_n12787_;
  assign new_n12789_ = ~new_n5966_ & new_n12787_;
  assign new_n12790_ = ~new_n12788_ & ~new_n12789_;
  assign new_n12791_ = pg35 & ~new_n12790_;
  assign n4722 = new_n12786_ | new_n12791_;
  assign new_n12793_ = ~pg35 & ng2004;
  assign new_n12794_ = ~ng2070 & ng2040;
  assign new_n12795_ = ~new_n7025_ & new_n12794_;
  assign new_n12796_ = ng2012 & ~new_n12795_;
  assign new_n12797_ = ~new_n7032_ & new_n12795_;
  assign new_n12798_ = ~new_n12796_ & ~new_n12797_;
  assign new_n12799_ = pg35 & ~new_n12798_;
  assign n4727 = new_n12793_ | new_n12799_;
  assign new_n12801_ = pg35 & ng4372;
  assign new_n12802_ = ~pg35 & new_n12801_;
  assign new_n12803_ = ~ng4864 & ~ng4836;
  assign new_n12804_ = ~new_n7605_ & new_n12803_;
  assign new_n12805_ = new_n7606_ & new_n12804_;
  assign new_n12806_ = ~ng4871 & new_n12805_;
  assign new_n12807_ = pg35 & new_n12806_;
  assign n4732 = new_n12802_ | new_n12807_;
  assign new_n12809_ = ~pg35 & ng2102;
  assign new_n12810_ = ng2108 & ~new_n8022_;
  assign new_n12811_ = ng2102 & new_n8022_;
  assign new_n12812_ = ~new_n12810_ & ~new_n12811_;
  assign new_n12813_ = pg35 & ~new_n12812_;
  assign n4737 = new_n12809_ | new_n12813_;
  assign new_n12815_ = ~pg35 & ng2563;
  assign new_n12816_ = ng2599 & ~ng2629;
  assign new_n12817_ = ~new_n7174_ & new_n12816_;
  assign new_n12818_ = ng2571 & ~new_n12817_;
  assign new_n12819_ = ~new_n8484_ & new_n12817_;
  assign new_n12820_ = ~new_n12818_ & ~new_n12819_;
  assign new_n12821_ = pg35 & ~new_n12820_;
  assign n4742 = new_n12815_ | new_n12821_;
  assign new_n12823_ = ~pg35 & ng2079;
  assign new_n12824_ = ng2093 & ~new_n10172_;
  assign new_n12825_ = ng2079 & new_n12824_;
  assign new_n12826_ = new_n12824_ & ~new_n12825_;
  assign new_n12827_ = ng2079 & ~new_n12825_;
  assign new_n12828_ = ~new_n12826_ & ~new_n12827_;
  assign new_n12829_ = new_n9143_ & ~new_n12828_;
  assign new_n12830_ = ng2093 & ~new_n9143_;
  assign new_n12831_ = ~new_n12829_ & ~new_n12830_;
  assign new_n12832_ = pg35 & ~new_n12831_;
  assign n4747 = new_n12823_ | new_n12832_;
  assign new_n12834_ = ~pg35 & ng6474;
  assign new_n12835_ = ng6474 & ng6466;
  assign new_n12836_ = ng6479 & ~new_n12835_;
  assign new_n12837_ = ~ng6479 & new_n12835_;
  assign new_n12838_ = ~new_n12836_ & ~new_n12837_;
  assign new_n12839_ = pg35 & ~new_n12838_;
  assign n4752 = new_n12834_ | new_n12839_;
  assign new_n12841_ = ~pg35 & ng1559;
  assign new_n12842_ = ng1559 & new_n12441_;
  assign new_n12843_ = ng1554 & ~new_n8877_;
  assign new_n12844_ = ~new_n12842_ & new_n12843_;
  assign new_n12845_ = ~ng1554 & ~new_n8877_;
  assign new_n12846_ = new_n12842_ & new_n12845_;
  assign new_n12847_ = ~new_n12844_ & ~new_n12846_;
  assign new_n12848_ = pg35 & ~new_n12847_;
  assign n4757 = new_n12841_ | new_n12848_;
  assign new_n12850_ = ~pg35 & ng3211;
  assign new_n12851_ = new_n7151_ & new_n9412_;
  assign new_n12852_ = ng3207 & ~new_n12851_;
  assign new_n12853_ = ~new_n5966_ & new_n12851_;
  assign new_n12854_ = ~new_n12852_ & ~new_n12853_;
  assign new_n12855_ = pg35 & ~new_n12854_;
  assign n4762 = new_n12850_ | new_n12855_;
  assign new_n12857_ = ~pg35 & ng1714;
  assign new_n12858_ = ng1720 & ~new_n7231_;
  assign new_n12859_ = ng1714 & new_n7231_;
  assign new_n12860_ = ~new_n12858_ & ~new_n12859_;
  assign new_n12861_ = pg35 & ~new_n12860_;
  assign n4771 = new_n12857_ | new_n12861_;
  assign new_n12863_ = ~pg35 & ng1189;
  assign new_n12864_ = ng1070 & new_n8813_;
  assign new_n12865_ = ng1193 & ~new_n12864_;
  assign new_n12866_ = ~new_n5949_ & ~new_n12865_;
  assign new_n12867_ = pg35 & ~new_n12866_;
  assign n4776 = new_n12863_ | new_n12867_;
  assign new_n12869_ = ~pg35 & ng3239;
  assign new_n12870_ = new_n8744_ & new_n9338_;
  assign new_n12871_ = ng3255 & ~new_n12870_;
  assign new_n12872_ = ~new_n5966_ & new_n12870_;
  assign new_n12873_ = ~new_n12871_ & ~new_n12872_;
  assign new_n12874_ = pg35 & ~new_n12873_;
  assign n4781 = new_n12869_ | new_n12874_;
  assign new_n12876_ = ~pg35 & ng5897;
  assign new_n12877_ = new_n7649_ & new_n7997_;
  assign new_n12878_ = ng5893 & ~new_n12877_;
  assign new_n12879_ = ~new_n5966_ & new_n12877_;
  assign new_n12880_ = ~new_n12878_ & ~new_n12879_;
  assign new_n12881_ = pg35 & ~new_n12880_;
  assign n4786 = new_n12876_ | new_n12881_;
  assign n4791 = ~pg35 & ng4392;
  assign new_n12884_ = pg35 & ng6336;
  assign new_n12885_ = ~pg35 & new_n12884_;
  assign new_n12886_ = pg35 & ng6227;
  assign n4796 = new_n12885_ | new_n12886_;
  assign new_n12888_ = ~pg35 & ng1484;
  assign new_n12889_ = new_n6433_ & new_n7472_;
  assign new_n12890_ = ng1484 & ng1300;
  assign new_n12891_ = ng1300 & ~new_n12890_;
  assign new_n12892_ = ng1484 & ~new_n12890_;
  assign new_n12893_ = ~new_n12891_ & ~new_n12892_;
  assign new_n12894_ = new_n12889_ & ~new_n12893_;
  assign new_n12895_ = ng1300 & ~new_n12889_;
  assign new_n12896_ = ~new_n12894_ & ~new_n12895_;
  assign new_n12897_ = pg35 & ~new_n12896_;
  assign n4800 = new_n12888_ | new_n12897_;
  assign new_n12899_ = ~pg35 & ng3742;
  assign new_n12900_ = ~ng3736 & new_n6078_;
  assign new_n12901_ = ~ng3742 & new_n12900_;
  assign new_n12902_ = ng3736 & new_n6083_;
  assign new_n12903_ = ng3742 & new_n12902_;
  assign new_n12904_ = ~new_n12901_ & ~new_n12903_;
  assign new_n12905_ = ~ng3747 & ~new_n12904_;
  assign new_n12906_ = ng3747 & new_n6104_;
  assign new_n12907_ = new_n12904_ & new_n12906_;
  assign new_n12908_ = ~new_n12905_ & ~new_n12907_;
  assign new_n12909_ = pg35 & ~new_n12908_;
  assign n4805 = new_n12899_ | new_n12909_;
  assign new_n12911_ = ~pg35 & ng4549;
  assign new_n12912_ = ~ng4578 & new_n5871_;
  assign new_n12913_ = ng4581 & ~new_n12912_;
  assign new_n12914_ = ng4549 & ~ng4581;
  assign new_n12915_ = ~new_n12913_ & ~new_n12914_;
  assign new_n12916_ = pg35 & ~new_n12915_;
  assign n4810 = new_n12911_ | new_n12916_;
  assign new_n12918_ = ~pg35 & ng5413;
  assign new_n12919_ = ~new_n6383_ & ~new_n6391_;
  assign new_n12920_ = pg35 & new_n12919_;
  assign n4815 = new_n12918_ | new_n12920_;
  assign new_n12922_ = ~pg35 & ng3179;
  assign new_n12923_ = new_n9368_ & new_n9412_;
  assign new_n12924_ = ng3187 & ~new_n12923_;
  assign new_n12925_ = ~new_n5966_ & new_n12923_;
  assign new_n12926_ = ~new_n12924_ & ~new_n12925_;
  assign new_n12927_ = pg35 & ~new_n12926_;
  assign n4820 = new_n12922_ | new_n12927_;
  assign n4825 = ~pg35 & ng4927;
  assign new_n12930_ = pg35 & ng1992;
  assign new_n12931_ = ~pg35 & new_n12930_;
  assign new_n12932_ = ~ng2070 & ng1996;
  assign new_n12933_ = ~ng2070 & ~ng2040;
  assign new_n12934_ = ~new_n12932_ & ~new_n12933_;
  assign new_n12935_ = ~new_n9212_ & ~new_n12934_;
  assign new_n12936_ = ~new_n7025_ & new_n12935_;
  assign new_n12937_ = ng1996 & new_n7025_;
  assign new_n12938_ = ~new_n12936_ & ~new_n12937_;
  assign new_n12939_ = pg35 & ~new_n12938_;
  assign n4830 = new_n12931_ | new_n12939_;
  assign new_n12941_ = pg35 & ng3151;
  assign new_n12942_ = ~pg35 & new_n12941_;
  assign new_n12943_ = ~ng3625 & ng3649;
  assign new_n12944_ = ~ng3618 & ng3625;
  assign new_n12945_ = ~new_n12943_ & ~new_n12944_;
  assign new_n12946_ = ~new_n9026_ & new_n12945_;
  assign new_n12947_ = ~ng3632 & ng3661;
  assign new_n12948_ = ng3632 & ~ng3654;
  assign new_n12949_ = ~ng3661 & ng3618;
  assign new_n12950_ = new_n12946_ & ~new_n12947_;
  assign new_n12951_ = ~new_n12948_ & new_n12950_;
  assign new_n12952_ = ~new_n12949_ & new_n12951_;
  assign new_n12953_ = pg35 & new_n12952_;
  assign n4835 = new_n12942_ | new_n12953_;
  assign new_n12955_ = ~pg35 & ng3004;
  assign new_n12956_ = ~new_n8927_ & ~new_n8931_;
  assign new_n12957_ = ~ng3017 & ~new_n12956_;
  assign new_n12958_ = ng3017 & new_n8954_;
  assign new_n12959_ = new_n12956_ & new_n12958_;
  assign new_n12960_ = ~new_n12957_ & ~new_n12959_;
  assign new_n12961_ = pg35 & ~new_n12960_;
  assign n4839 = new_n12955_ | new_n12961_;
  assign new_n12963_ = ~pg35 & ng102;
  assign new_n12964_ = ~pg72 & ng255;
  assign new_n12965_ = pg73 & ~new_n12964_;
  assign new_n12966_ = pg72 & ng262;
  assign new_n12967_ = ~pg72 & ng269;
  assign new_n12968_ = ~new_n12966_ & ~new_n12967_;
  assign new_n12969_ = ~pg73 & new_n12968_;
  assign new_n12970_ = ~new_n12965_ & ~new_n12969_;
  assign new_n12971_ = pg35 & new_n12970_;
  assign n4844 = new_n12963_ | new_n12971_;
  assign new_n12973_ = ~pg35 & ng4717;
  assign new_n12974_ = ng4722 & ~new_n9308_;
  assign new_n12975_ = n2287 & new_n9308_;
  assign new_n12976_ = ~new_n12974_ & ~new_n12975_;
  assign new_n12977_ = pg35 & ~new_n12976_;
  assign n4852 = new_n12973_ | new_n12977_;
  assign new_n12979_ = ~pg35 & ng6159;
  assign new_n12980_ = ng6154 & ~new_n6694_;
  assign new_n12981_ = ~ng6336 & ~ng6395;
  assign new_n12982_ = ~ng6381 & new_n12981_;
  assign new_n12983_ = ng6369 & ng6287;
  assign new_n12984_ = new_n12982_ & new_n12983_;
  assign new_n12985_ = ng6336 & ~ng6395;
  assign new_n12986_ = ~ng6381 & new_n12985_;
  assign new_n12987_ = ng6377 & ng6259;
  assign new_n12988_ = new_n12986_ & new_n12987_;
  assign new_n12989_ = ~ng6336 & ng6395;
  assign new_n12990_ = ~ng6381 & new_n12989_;
  assign new_n12991_ = ng6303 & ng6373;
  assign new_n12992_ = new_n12990_ & new_n12991_;
  assign new_n12993_ = ~ng6381 & new_n4753_;
  assign new_n12994_ = ng6255 & ng6351;
  assign new_n12995_ = new_n12993_ & new_n12994_;
  assign new_n12996_ = ~new_n12984_ & ~new_n12988_;
  assign new_n12997_ = ~new_n12992_ & ~new_n12995_;
  assign new_n12998_ = new_n12996_ & new_n12997_;
  assign new_n12999_ = ng6381 & new_n12981_;
  assign new_n13000_ = ng6243 & ng6377;
  assign new_n13001_ = new_n12999_ & new_n13000_;
  assign new_n13002_ = ng6351 & ng6381;
  assign new_n13003_ = ng6351 & ~new_n13002_;
  assign new_n13004_ = ng6381 & ~new_n13002_;
  assign new_n13005_ = ~new_n13003_ & ~new_n13004_;
  assign new_n13006_ = new_n12985_ & new_n13005_;
  assign new_n13007_ = ng6267 & ng6329;
  assign new_n13008_ = new_n13006_ & new_n13007_;
  assign new_n13009_ = ng6381 & new_n12989_;
  assign new_n13010_ = ng6351 & ng6239;
  assign new_n13011_ = new_n13009_ & new_n13010_;
  assign new_n13012_ = new_n4753_ & new_n13005_;
  assign new_n13013_ = ng6283 & ng6358;
  assign new_n13014_ = new_n13012_ & new_n13013_;
  assign new_n13015_ = ~new_n13001_ & ~new_n13008_;
  assign new_n13016_ = ~new_n13011_ & ~new_n13014_;
  assign new_n13017_ = new_n13015_ & new_n13016_;
  assign new_n13018_ = ng6235 & ng6346;
  assign new_n13019_ = new_n12999_ & new_n13018_;
  assign new_n13020_ = ng6381 & new_n12985_;
  assign new_n13021_ = ng6279 & ng6369;
  assign new_n13022_ = new_n13020_ & new_n13021_;
  assign new_n13023_ = ng6365 & ng6263;
  assign new_n13024_ = new_n13009_ & new_n13023_;
  assign new_n13025_ = ng6381 & new_n4753_;
  assign new_n13026_ = ng6373 & ng6295;
  assign new_n13027_ = new_n13025_ & new_n13026_;
  assign new_n13028_ = ~new_n13019_ & ~new_n13022_;
  assign new_n13029_ = ~new_n13024_ & ~new_n13027_;
  assign new_n13030_ = new_n13028_ & new_n13029_;
  assign new_n13031_ = new_n12981_ & new_n13005_;
  assign new_n13032_ = ng6315 & ng6299;
  assign new_n13033_ = new_n13031_ & new_n13032_;
  assign new_n13034_ = ng6247 & ng6346;
  assign new_n13035_ = new_n12986_ & new_n13034_;
  assign new_n13036_ = ng6251 & ng6322;
  assign new_n13037_ = new_n12990_ & new_n13036_;
  assign new_n13038_ = ng6365 & ng6271;
  assign new_n13039_ = new_n12993_ & new_n13038_;
  assign new_n13040_ = ~new_n13033_ & ~new_n13035_;
  assign new_n13041_ = ~new_n13037_ & ~new_n13039_;
  assign new_n13042_ = new_n13040_ & new_n13041_;
  assign new_n13043_ = new_n13017_ & new_n13030_;
  assign new_n13044_ = new_n13042_ & new_n13043_;
  assign new_n13045_ = new_n12981_ & ~new_n13005_;
  assign new_n13046_ = ng6329 & ng6275;
  assign new_n13047_ = new_n13045_ & new_n13046_;
  assign new_n13048_ = new_n12985_ & ~new_n13005_;
  assign new_n13049_ = ng6315 & ng6307;
  assign new_n13050_ = new_n13048_ & new_n13049_;
  assign new_n13051_ = new_n12989_ & ~new_n13005_;
  assign new_n13052_ = ng6358 & ng6291;
  assign new_n13053_ = new_n13051_ & new_n13052_;
  assign new_n13054_ = ng6322 & ng6311;
  assign new_n13055_ = new_n13025_ & new_n13054_;
  assign new_n13056_ = ~new_n13047_ & ~new_n13050_;
  assign new_n13057_ = ~new_n13053_ & ~new_n13055_;
  assign new_n13058_ = new_n13056_ & new_n13057_;
  assign new_n13059_ = new_n12998_ & new_n13044_;
  assign new_n13060_ = new_n13058_ & new_n13059_;
  assign new_n13061_ = new_n12980_ & ~new_n13060_;
  assign new_n13062_ = new_n12980_ & ~new_n13061_;
  assign new_n13063_ = ~new_n13060_ & ~new_n13061_;
  assign new_n13064_ = ~new_n13062_ & ~new_n13063_;
  assign new_n13065_ = new_n6699_ & ~new_n13064_;
  assign new_n13066_ = ng6154 & ~new_n6699_;
  assign new_n13067_ = ~new_n13065_ & ~new_n13066_;
  assign new_n13068_ = pg35 & ~new_n13067_;
  assign n4857 = new_n12979_ | new_n13068_;
  assign new_n13070_ = ~pg35 & ng5248;
  assign new_n13071_ = new_n10722_ & new_n11431_;
  assign new_n13072_ = ng5264 & ~new_n13071_;
  assign new_n13073_ = ~new_n5966_ & new_n13071_;
  assign new_n13074_ = ~new_n13072_ & ~new_n13073_;
  assign new_n13075_ = pg35 & ~new_n13074_;
  assign n4862 = new_n13070_ | new_n13075_;
  assign new_n13077_ = pg35 & ng3143;
  assign new_n13078_ = ~pg35 & new_n13077_;
  assign new_n13079_ = n5814 & new_n10448_;
  assign new_n13080_ = ng3151 & ~new_n10448_;
  assign new_n13081_ = ~new_n13079_ & ~new_n13080_;
  assign new_n13082_ = pg35 & ~new_n13081_;
  assign n4867 = new_n13078_ | new_n13082_;
  assign new_n13084_ = ~pg35 & ng2878;
  assign new_n13085_ = n5005 & new_n7895_;
  assign new_n13086_ = ~ng2946 & ~ng2886;
  assign new_n13087_ = ~new_n13085_ & ~new_n13086_;
  assign new_n13088_ = pg35 & new_n13087_;
  assign n4872 = new_n13084_ | new_n13088_;
  assign new_n13090_ = ~pg35 & ng6381;
  assign new_n13091_ = ng6381 & new_n7307_;
  assign new_n13092_ = ~ng6390 & ~new_n13091_;
  assign new_n13093_ = pg35 & new_n13092_;
  assign n4877 = new_n13090_ | new_n13093_;
  assign new_n13095_ = ~pg35 & ng5731;
  assign new_n13096_ = ~new_n10151_ & ~new_n10154_;
  assign new_n13097_ = ~ng5736 & ~new_n13096_;
  assign new_n13098_ = ng5736 & new_n6424_;
  assign new_n13099_ = new_n13096_ & new_n13098_;
  assign new_n13100_ = ~new_n13097_ & ~new_n13099_;
  assign new_n13101_ = pg35 & ~new_n13100_;
  assign n4882 = new_n13095_ | new_n13101_;
  assign new_n13103_ = ~pg35 & ng4049;
  assign new_n13104_ = new_n4751_ & new_n7747_;
  assign new_n13105_ = new_n6467_ & new_n13104_;
  assign new_n13106_ = new_n4735_ & new_n13105_;
  assign new_n13107_ = ~ng4054 & ~new_n13106_;
  assign new_n13108_ = new_n6467_ & new_n13107_;
  assign new_n13109_ = ng4054 & ~new_n6467_;
  assign new_n13110_ = ~new_n13108_ & ~new_n13109_;
  assign new_n13111_ = pg35 & ~new_n13110_;
  assign n4887 = new_n13103_ | new_n13111_;
  assign new_n13113_ = ~pg35 & ng3470;
  assign new_n13114_ = ng3476 & ~new_n7432_;
  assign new_n13115_ = ng3470 & new_n7432_;
  assign new_n13116_ = ~new_n13114_ & ~new_n13115_;
  assign new_n13117_ = pg35 & ~new_n13116_;
  assign n4896 = new_n13113_ | new_n13117_;
  assign new_n13119_ = ~pg35 & ng59;
  assign new_n13120_ = ~ng4681 & ~ng4646;
  assign new_n13121_ = ~ng4674 & new_n13120_;
  assign new_n13122_ = ~ng4688 & new_n13121_;
  assign new_n13123_ = ~ng4776 & new_n5666_;
  assign new_n13124_ = ng4801 & ng4793;
  assign new_n13125_ = ~ng4776 & new_n13124_;
  assign new_n13126_ = ~new_n13123_ & ~new_n13125_;
  assign new_n13127_ = ~new_n5845_ & ~new_n13126_;
  assign new_n13128_ = ng4722 & new_n5836_;
  assign new_n13129_ = ng4732 & new_n5838_1_;
  assign new_n13130_ = ng4717 & new_n5840_;
  assign new_n13131_ = ng4727 & new_n5665_;
  assign new_n13132_ = ~new_n13128_ & ~new_n13129_;
  assign new_n13133_ = ~new_n13130_ & ~new_n13131_;
  assign new_n13134_ = new_n13132_ & new_n13133_;
  assign new_n13135_ = ~new_n5845_ & ~new_n13134_;
  assign new_n13136_ = ~new_n13134_ & ~new_n13135_;
  assign new_n13137_ = ~new_n5845_ & ~new_n13135_;
  assign new_n13138_ = ~new_n13136_ & ~new_n13137_;
  assign new_n13139_ = new_n5690_ & ~new_n13138_;
  assign new_n13140_ = ~ng4776 & new_n5689_;
  assign new_n13141_ = ~ng4737 & new_n5665_;
  assign new_n13142_ = ~new_n5838_1_ & ~new_n5840_;
  assign new_n13143_ = ~new_n13141_ & new_n13142_;
  assign new_n13144_ = new_n13140_ & ~new_n13143_;
  assign new_n13145_ = ~new_n5667_ & ~new_n13127_;
  assign new_n13146_ = ~new_n13139_ & ~new_n13144_;
  assign new_n13147_ = new_n13145_ & new_n13146_;
  assign new_n13148_ = new_n13122_ & ~new_n13147_;
  assign new_n13149_ = ng128 & ng4646;
  assign new_n13150_ = ng4831 & ng4681;
  assign new_n13151_ = ng4674 & ~ng4821;
  assign new_n13152_ = ~ng4826 & ng4688;
  assign new_n13153_ = ~new_n13149_ & ~new_n13150_;
  assign new_n13154_ = ~new_n13151_ & ~new_n13152_;
  assign new_n13155_ = new_n13153_ & new_n13154_;
  assign new_n13156_ = ~new_n13122_ & ~new_n13155_;
  assign new_n13157_ = ~new_n13148_ & ~new_n13156_;
  assign new_n13158_ = pg35 & ~new_n13157_;
  assign n4901 = new_n13119_ | new_n13158_;
  assign new_n13160_ = ~pg35 & ng5869;
  assign new_n13161_ = ng5873 & ~new_n11838_;
  assign new_n13162_ = ~ng5869 & new_n13161_;
  assign new_n13163_ = ~ng5873 & ~new_n11838_;
  assign new_n13164_ = ng5869 & new_n13163_;
  assign new_n13165_ = ~new_n13162_ & ~new_n13164_;
  assign new_n13166_ = pg35 & ~new_n13165_;
  assign n4906 = new_n13160_ | new_n13166_;
  assign new_n13168_ = ~pg35 & ng5706;
  assign new_n13169_ = ~new_n6401_ & ~new_n6403_;
  assign new_n13170_ = ~ng5719 & ~new_n13169_;
  assign new_n13171_ = ng5719 & new_n6424_;
  assign new_n13172_ = new_n13169_ & new_n13171_;
  assign new_n13173_ = ~new_n13170_ & ~new_n13172_;
  assign new_n13174_ = pg35 & ~new_n13173_;
  assign n4911 = new_n13168_ | new_n13174_;
  assign new_n13176_ = ~pg35 & ng4572;
  assign n4916 = new_n9527_ | new_n13176_;
  assign new_n13178_ = pg35 & ng4507;
  assign new_n13179_ = ~pg35 & new_n13178_;
  assign new_n13180_ = ng4467 & ng4462;
  assign new_n13181_ = ~new_n9232_ & new_n13180_;
  assign new_n13182_ = pg35 & ~new_n13181_;
  assign n4921 = new_n13179_ | new_n13182_;
  assign new_n13184_ = ~pg35 & ng6307;
  assign new_n13185_ = ng6311 & ~new_n7064_;
  assign new_n13186_ = ~new_n5966_ & new_n7064_;
  assign new_n13187_ = ~new_n13185_ & ~new_n13186_;
  assign new_n13188_ = pg35 & ~new_n13187_;
  assign n4926 = new_n13184_ | new_n13188_;
  assign new_n13190_ = ~pg35 & ng6311;
  assign new_n13191_ = new_n6699_ & ~new_n13060_;
  assign new_n13192_ = ng4826 & ~new_n6699_;
  assign new_n13193_ = ~new_n13191_ & ~new_n13192_;
  assign new_n13194_ = pg35 & ~new_n13193_;
  assign n4931 = new_n13190_ | new_n13194_;
  assign new_n13196_ = ~pg35 & ng3329;
  assign new_n13197_ = ng3338 & ~new_n8782_;
  assign new_n13198_ = ~ng3338 & new_n8782_;
  assign new_n13199_ = ~new_n13197_ & ~new_n13198_;
  assign new_n13200_ = pg35 & ~new_n13199_;
  assign n4940 = new_n13196_ | new_n13200_;
  assign new_n13202_ = ~pg35 & ng1691;
  assign new_n13203_ = new_n7230_ & new_n9259_;
  assign new_n13204_ = ng1696 & ~new_n13203_;
  assign new_n13205_ = ng1691 & ng1687;
  assign new_n13206_ = ng1691 & ~new_n13205_;
  assign new_n13207_ = ng1687 & ~new_n13205_;
  assign new_n13208_ = ~new_n13206_ & ~new_n13207_;
  assign new_n13209_ = new_n13203_ & ~new_n13208_;
  assign new_n13210_ = ~new_n13204_ & ~new_n13209_;
  assign new_n13211_ = pg35 & ~new_n13210_;
  assign n4945 = new_n13202_ | new_n13211_;
  assign new_n13213_ = ~pg35 & ng3021;
  assign new_n13214_ = ~new_n8929_ & ~new_n8933_;
  assign new_n13215_ = ~ng3025 & ~new_n13214_;
  assign new_n13216_ = ng3025 & new_n8954_;
  assign new_n13217_ = new_n13214_ & new_n13216_;
  assign new_n13218_ = ~new_n13215_ & ~new_n13217_;
  assign new_n13219_ = pg35 & ~new_n13218_;
  assign n4950 = new_n13213_ | new_n13219_;
  assign new_n13221_ = ~pg35 & ng3558;
  assign new_n13222_ = new_n6769_ & new_n10353_;
  assign new_n13223_ = ng3578 & ~new_n13222_;
  assign new_n13224_ = ~new_n5966_ & new_n13222_;
  assign new_n13225_ = ~new_n13223_ & ~new_n13224_;
  assign new_n13226_ = pg35 & ~new_n13225_;
  assign n4960 = new_n13221_ | new_n13226_;
  assign new_n13228_ = ~pg35 & ng2375;
  assign new_n13229_ = ng2380 & ~new_n7888_;
  assign new_n13230_ = ng2375 & new_n7888_;
  assign new_n13231_ = ~new_n13229_ & ~new_n13230_;
  assign new_n13232_ = pg35 & ~new_n13231_;
  assign n4965 = new_n13228_ | new_n13232_;
  assign new_n13234_ = ~pg35 & ng2643;
  assign new_n13235_ = ~new_n7174_ & new_n7491_;
  assign new_n13236_ = ng2648 & ~new_n13235_;
  assign new_n13237_ = ng2643 & new_n13235_;
  assign new_n13238_ = ~new_n13236_ & ~new_n13237_;
  assign new_n13239_ = pg35 & ~new_n13238_;
  assign n4970 = new_n13234_ | new_n13239_;
  assign new_n13241_ = ~pg35 & ng5436;
  assign new_n13242_ = ng5441 & ~new_n8965_;
  assign new_n13243_ = ~ng5441 & new_n8965_;
  assign new_n13244_ = ~new_n13242_ & ~new_n13243_;
  assign new_n13245_ = pg35 & ~new_n13244_;
  assign n4975 = new_n13241_ | new_n13245_;
  assign new_n13247_ = ~pg35 & ng106;
  assign new_n13248_ = pg35 & ng316;
  assign n4980 = new_n13247_ | new_n13248_;
  assign new_n13250_ = ~pg35 & ng4593;
  assign new_n13251_ = ~ng4601 & new_n8853_;
  assign new_n13252_ = new_n12748_ & new_n13251_;
  assign new_n13253_ = ng4601 & new_n8853_;
  assign new_n13254_ = ~new_n12748_ & new_n13253_;
  assign new_n13255_ = ~new_n13252_ & ~new_n13254_;
  assign new_n13256_ = pg35 & ~new_n13255_;
  assign n4985 = new_n13250_ | new_n13256_;
  assign new_n13258_ = ~pg35 & ng2648;
  assign new_n13259_ = ng2567 & ~new_n13235_;
  assign new_n13260_ = ~new_n8484_ & new_n13235_;
  assign new_n13261_ = ~new_n13259_ & ~new_n13260_;
  assign new_n13262_ = pg35 & ~new_n13261_;
  assign n4990 = new_n13258_ | new_n13262_;
  assign new_n13264_ = ~pg35 & ng446;
  assign new_n13265_ = ng896 & ng890;
  assign new_n13266_ = ~ng703 & ~new_n12729_;
  assign new_n13267_ = new_n12701_ & new_n13266_;
  assign new_n13268_ = ~new_n11258_ & ~new_n13267_;
  assign new_n13269_ = ng862 & new_n13268_;
  assign new_n13270_ = ~new_n9672_ & ~new_n13265_;
  assign new_n13271_ = ~new_n13269_ & new_n13270_;
  assign new_n13272_ = pg35 & ~new_n13271_;
  assign n4995 = new_n13264_ | new_n13272_;
  assign new_n13274_ = ~pg35 & ng2856;
  assign new_n13275_ = n5814 & new_n7895_;
  assign new_n13276_ = ~ng2864 & new_n4844_1_;
  assign new_n13277_ = ~new_n13275_ & ~new_n13276_;
  assign new_n13278_ = pg35 & new_n13277_;
  assign n5000 = new_n13274_ | new_n13278_;
  assign new_n13280_ = ~pg35 & ng4558;
  assign new_n13281_ = pg6749 & pg35;
  assign n5010 = new_n13280_ | new_n13281_;
  assign new_n13283_ = pg35 & ng128;
  assign new_n13284_ = ~pg35 & new_n13283_;
  assign new_n13285_ = ng5156 & ~pg26801;
  assign new_n13286_ = ~new_n5966_ & new_n13285_;
  assign new_n13287_ = new_n13285_ & ~new_n13286_;
  assign new_n13288_ = ~new_n5966_ & ~new_n13286_;
  assign new_n13289_ = ~new_n13287_ & ~new_n13288_;
  assign new_n13290_ = pg35 & ~new_n13289_;
  assign n5020 = new_n13284_ | new_n13290_;
  assign new_n13292_ = ~pg35 & ng2269;
  assign new_n13293_ = ng2273 & ~new_n6524_;
  assign new_n13294_ = ~ng2273 & new_n6524_;
  assign new_n13295_ = ~new_n13293_ & ~new_n13294_;
  assign new_n13296_ = pg35 & ~new_n13295_;
  assign n5025 = new_n13292_ | new_n13296_;
  assign new_n13298_ = pg35 & ng929;
  assign new_n13299_ = ~pg35 & new_n13298_;
  assign new_n13300_ = ~ng1227 & new_n7073_;
  assign new_n13301_ = ~ng904 & ng1227;
  assign new_n13302_ = ~new_n13300_ & ~new_n13301_;
  assign new_n13303_ = pg35 & ~new_n13302_;
  assign n5030 = new_n13299_ | new_n13303_;
  assign new_n13305_ = ~pg35 & ng6455;
  assign new_n13306_ = ng6451 & ng6455;
  assign new_n13307_ = pg35 & new_n13306_;
  assign n5035 = new_n13305_ | new_n13307_;
  assign new_n13309_ = ~pg35 & ng6219;
  assign new_n13310_ = ng6215 & ng6219;
  assign new_n13311_ = ~ng6227 & ~new_n5852_;
  assign new_n13312_ = new_n13310_ & new_n13311_;
  assign new_n13313_ = ng6227 & ~new_n5852_;
  assign new_n13314_ = ~new_n13310_ & new_n13313_;
  assign new_n13315_ = ~new_n13312_ & ~new_n13314_;
  assign new_n13316_ = pg35 & ~new_n13315_;
  assign n5040 = new_n13309_ | new_n13316_;
  assign new_n13318_ = pg35 & ng6137;
  assign new_n13319_ = ~pg35 & new_n13318_;
  assign new_n13320_ = ~ng6203 & new_n5853_1_;
  assign new_n13321_ = pg35 & new_n13320_;
  assign n5045 = new_n13319_ | new_n13321_;
  assign new_n13323_ = ~pg35 & ng4358;
  assign new_n13324_ = ~ng4332 & ~ng4311;
  assign new_n13325_ = ~ng4584 & ~ng4322;
  assign new_n13326_ = new_n13324_ & new_n13325_;
  assign new_n13327_ = ~ng4608 & ~ng4593;
  assign new_n13328_ = ~ng4616 & ~ng4601;
  assign new_n13329_ = new_n13327_ & new_n13328_;
  assign new_n13330_ = new_n13326_ & new_n13329_;
  assign new_n13331_ = ng4340 & ~ng4349;
  assign new_n13332_ = ~ng4358 & new_n13331_;
  assign new_n13333_ = new_n8692_ & new_n13330_;
  assign new_n13334_ = new_n13332_ & new_n13333_;
  assign new_n13335_ = pg35 & new_n13334_;
  assign n5050 = new_n13323_ | new_n13335_;
  assign new_n13337_ = ~pg35 & ng2246;
  assign new_n13338_ = ng2165 & ~new_n6524_;
  assign new_n13339_ = new_n6524_ & ~new_n6725_;
  assign new_n13340_ = ~new_n13338_ & ~new_n13339_;
  assign new_n13341_ = pg35 & ~new_n13340_;
  assign n5058 = new_n13337_ | new_n13341_;
  assign new_n13343_ = ~pg35 & ng4145;
  assign new_n13344_ = ng4112 & ~new_n10091_;
  assign new_n13345_ = ng4145 & new_n10091_;
  assign new_n13346_ = ~new_n13344_ & ~new_n13345_;
  assign new_n13347_ = pg35 & ~new_n13346_;
  assign n5063 = new_n13343_ | new_n13347_;
  assign new_n13349_ = ~pg35 & ng1978;
  assign new_n13350_ = ng1982 & ~new_n11266_;
  assign new_n13351_ = ~ng1982 & new_n11266_;
  assign new_n13352_ = ~new_n13350_ & ~new_n13351_;
  assign new_n13353_ = pg35 & ~new_n13352_;
  assign n5068 = new_n13349_ | new_n13353_;
  assign new_n13355_ = ~pg35 & ng4732;
  assign new_n13356_ = ng4717 & ~new_n9308_;
  assign new_n13357_ = n5814 & new_n9308_;
  assign new_n13358_ = ~new_n13356_ & ~new_n13357_;
  assign new_n13359_ = pg35 & ~new_n13358_;
  assign n5073 = new_n13355_ | new_n13359_;
  assign new_n13361_ = ~pg35 & ng3187;
  assign new_n13362_ = new_n9315_ & new_n9368_;
  assign new_n13363_ = ng3215 & ~new_n13362_;
  assign new_n13364_ = ~new_n5966_ & new_n13362_;
  assign new_n13365_ = ~new_n13363_ & ~new_n13364_;
  assign new_n13366_ = pg35 & ~new_n13365_;
  assign n5082 = new_n13361_ | new_n13366_;
  assign new_n13368_ = ~pg35 & ng1361;
  assign new_n13369_ = new_n6308_1_ & ~new_n6310_;
  assign new_n13370_ = ng1367 & ~new_n13369_;
  assign new_n13371_ = ~ng1367 & new_n6306_;
  assign new_n13372_ = new_n13369_ & new_n13371_;
  assign new_n13373_ = ~new_n13370_ & ~new_n13372_;
  assign new_n13374_ = pg35 & ~new_n13373_;
  assign n5087 = new_n13368_ | new_n13374_;
  assign new_n13376_ = ~pg35 & ng2028;
  assign new_n13377_ = ~pg113 & new_n5180_;
  assign new_n13378_ = new_n5909_ & new_n13377_;
  assign new_n13379_ = ~ng2028 & ~new_n13378_;
  assign new_n13380_ = new_n9143_ & ~new_n13379_;
  assign new_n13381_ = ng2051 & ~new_n9143_;
  assign new_n13382_ = ~new_n13380_ & ~new_n13381_;
  assign new_n13383_ = pg35 & ~new_n13382_;
  assign n5092 = new_n13376_ | new_n13383_;
  assign new_n13385_ = ~pg35 & ng1677;
  assign new_n13386_ = ng1691 & ~new_n9259_;
  assign new_n13387_ = ng1677 & new_n13386_;
  assign new_n13388_ = new_n13386_ & ~new_n13387_;
  assign new_n13389_ = ng1677 & ~new_n13387_;
  assign new_n13390_ = ~new_n13388_ & ~new_n13389_;
  assign new_n13391_ = new_n7230_ & ~new_n13390_;
  assign new_n13392_ = ng1691 & ~new_n7230_;
  assign new_n13393_ = ~new_n13391_ & ~new_n13392_;
  assign new_n13394_ = pg35 & ~new_n13393_;
  assign n5097 = new_n13385_ | new_n13394_;
  assign new_n13396_ = ~pg35 & ng1135;
  assign new_n13397_ = ng1111 & ~new_n12576_;
  assign new_n13398_ = ng1105 & new_n7775_;
  assign new_n13399_ = ng1105 & ~new_n13398_;
  assign new_n13400_ = new_n7775_ & ~new_n13398_;
  assign new_n13401_ = ~new_n13399_ & ~new_n13400_;
  assign new_n13402_ = ng1111 & ~new_n13401_;
  assign new_n13403_ = ~new_n7774_ & new_n13402_;
  assign new_n13404_ = new_n7774_ & ~new_n13401_;
  assign new_n13405_ = ~new_n13403_ & ~new_n13404_;
  assign new_n13406_ = new_n12576_ & ~new_n13405_;
  assign new_n13407_ = ~new_n13397_ & ~new_n13406_;
  assign new_n13408_ = pg35 & ~new_n13407_;
  assign n5102 = new_n13396_ | new_n13408_;
  assign new_n13410_ = ~pg35 & ng5817;
  assign new_n13411_ = ng5821 & ~new_n10071_;
  assign new_n13412_ = ~ng5821 & new_n10071_;
  assign new_n13413_ = ~new_n13411_ & ~new_n13412_;
  assign new_n13414_ = pg35 & ~new_n13413_;
  assign n5107 = new_n13410_ | new_n13414_;
  assign new_n13416_ = ~pg35 & ng417;
  assign new_n13417_ = ng411 & ~new_n6067_;
  assign new_n13418_ = ~ng417 & ~new_n12728_;
  assign new_n13419_ = ~ng417 & ~new_n13418_;
  assign new_n13420_ = ~new_n12728_ & ~new_n13418_;
  assign new_n13421_ = ~new_n13419_ & ~new_n13420_;
  assign new_n13422_ = new_n6067_ & ~new_n13421_;
  assign new_n13423_ = ~new_n13417_ & ~new_n13422_;
  assign new_n13424_ = pg35 & ~new_n13423_;
  assign n5112 = new_n13416_ | new_n13424_;
  assign new_n13426_ = ~pg35 & ng4064;
  assign new_n13427_ = ~new_n5979_1_ & ~new_n7047_;
  assign new_n13428_ = ng4169 & ~new_n13427_;
  assign new_n13429_ = pg35 & new_n13428_;
  assign n5117 = new_n13426_ | new_n13429_;
  assign new_n13431_ = ~pg35 & ng5759;
  assign new_n13432_ = ~new_n6413_ & ~new_n6421_;
  assign new_n13433_ = pg35 & new_n13432_;
  assign n5122 = new_n13431_ | new_n13433_;
  assign new_n13435_ = ~pg35 & ng2657;
  assign new_n13436_ = ng2619 & ng2587;
  assign new_n13437_ = new_n10306_ & new_n13436_;
  assign new_n13438_ = ng2661 & ~new_n13437_;
  assign new_n13439_ = ~ng2661 & new_n13437_;
  assign new_n13440_ = ~new_n13438_ & ~new_n13439_;
  assign new_n13441_ = pg35 & ~new_n13440_;
  assign n5131 = new_n13435_ | new_n13441_;
  assign new_n13443_ = ~pg35 & ng3057;
  assign new_n13444_ = ~new_n8943_ & ~new_n8951_;
  assign new_n13445_ = pg35 & new_n13444_;
  assign n5136 = new_n13443_ | new_n13445_;
  assign new_n13447_ = ~pg35 & ng2960;
  assign new_n13448_ = n5005 & new_n9379_;
  assign new_n13449_ = ng2970 & ~new_n9379_;
  assign new_n13450_ = ~new_n13448_ & ~new_n13449_;
  assign new_n13451_ = pg35 & ~new_n13450_;
  assign n5141 = new_n13447_ | new_n13451_;
  assign new_n13453_ = ~pg35 & ng4621;
  assign new_n13454_ = ng4628 & new_n8339_;
  assign new_n13455_ = ~new_n8337_ & new_n13454_;
  assign new_n13456_ = ~ng4628 & new_n8339_;
  assign new_n13457_ = new_n8337_ & new_n13456_;
  assign new_n13458_ = ~new_n13455_ & ~new_n13457_;
  assign new_n13459_ = pg35 & ~new_n13458_;
  assign n5146 = new_n13453_ | new_n13459_;
  assign new_n13461_ = ~pg56 & ng58;
  assign new_n13462_ = ~ng12 & new_n13461_;
  assign new_n13463_ = ~pg54 & new_n13462_;
  assign n5151 = new_n4890_ & new_n13463_;
  assign new_n13465_ = ~pg35 & ng2775;
  assign new_n13466_ = ng2771 & ~new_n6752_;
  assign new_n13467_ = ng2767 & ~new_n5870_;
  assign new_n13468_ = ~new_n8665_ & ~new_n13467_;
  assign new_n13469_ = new_n6752_ & new_n13468_;
  assign new_n13470_ = ~new_n13466_ & ~new_n13469_;
  assign new_n13471_ = pg35 & ~new_n13470_;
  assign n5156 = new_n13465_ | new_n13471_;
  assign new_n13473_ = ~pg35 & ng3542;
  assign new_n13474_ = new_n7038_ & new_n10353_;
  assign new_n13475_ = ng3570 & ~new_n13474_;
  assign new_n13476_ = ~new_n5966_ & new_n13474_;
  assign new_n13477_ = ~new_n13475_ & ~new_n13476_;
  assign new_n13478_ = pg35 & ~new_n13477_;
  assign n5161 = new_n13473_ | new_n13478_;
  assign new_n13480_ = ~pg35 & ng617;
  assign new_n13481_ = ng622 & ~new_n6545_;
  assign new_n13482_ = ~new_n9122_ & new_n13481_;
  assign new_n13483_ = ~ng622 & new_n9122_;
  assign new_n13484_ = ~new_n13482_ & ~new_n13483_;
  assign new_n13485_ = pg35 & ~new_n13484_;
  assign n5166 = new_n13480_ | new_n13485_;
  assign new_n13487_ = pg35 & ng3845;
  assign new_n13488_ = ~pg35 & new_n13487_;
  assign new_n13489_ = n4955 & new_n10448_;
  assign new_n13490_ = ng3853 & ~new_n10448_;
  assign new_n13491_ = ~new_n13489_ & ~new_n13490_;
  assign new_n13492_ = pg35 & ~new_n13491_;
  assign n5171 = new_n13488_ | new_n13492_;
  assign new_n13494_ = ~pg35 & ng2927;
  assign new_n13495_ = ng12 & n2287;
  assign new_n13496_ = new_n4937_ & new_n13495_;
  assign new_n13497_ = ~ng4153 & ~ng4072;
  assign new_n13498_ = ~ng2941 & new_n13497_;
  assign new_n13499_ = ~new_n13496_ & ~new_n13498_;
  assign new_n13500_ = pg35 & new_n13499_;
  assign n5176 = new_n13494_ | new_n13500_;
  assign new_n13502_ = ~pg35 & ng4722;
  assign new_n13503_ = ng4737 & ~new_n9308_;
  assign new_n13504_ = ~n6079 & new_n9308_;
  assign new_n13505_ = ~new_n13503_ & ~new_n13504_;
  assign new_n13506_ = pg35 & ~new_n13505_;
  assign n5186 = new_n13502_ | new_n13506_;
  assign new_n13508_ = ~pg35 & ng3436;
  assign new_n13509_ = ng3431 & ng3423;
  assign new_n13510_ = ng3436 & new_n13509_;
  assign new_n13511_ = ~ng3440 & new_n13510_;
  assign new_n13512_ = ng3440 & ~new_n13510_;
  assign new_n13513_ = ~new_n13511_ & ~new_n13512_;
  assign new_n13514_ = pg35 & ~new_n13513_;
  assign n5191 = new_n13508_ | new_n13514_;
  assign new_n13516_ = ~pg35 & ng5366;
  assign new_n13517_ = ~ng5406 & ~ng5366;
  assign new_n13518_ = ng5360 & new_n13517_;
  assign new_n13519_ = ~ng5360 & new_n6394_;
  assign new_n13520_ = ~new_n13517_ & new_n13519_;
  assign new_n13521_ = ~new_n13518_ & ~new_n13520_;
  assign new_n13522_ = pg35 & ~new_n13521_;
  assign n5196 = new_n13516_ | new_n13522_;
  assign new_n13524_ = ~pg35 & ng4760;
  assign new_n13525_ = ~new_n8500_ & ~new_n9637_;
  assign new_n13526_ = ng4760 & ~new_n8500_;
  assign new_n13527_ = ~new_n8503_ & ~new_n13526_;
  assign new_n13528_ = ~new_n13525_ & ~new_n13527_;
  assign new_n13529_ = ng4754 & new_n13525_;
  assign new_n13530_ = ~new_n13528_ & ~new_n13529_;
  assign new_n13531_ = pg35 & ~new_n13530_;
  assign n5201 = new_n13524_ | new_n13531_;
  assign new_n13533_ = ~pg35 & ng5008;
  assign new_n13534_ = ~ng4983 & new_n11040_;
  assign new_n13535_ = new_n5679_ & new_n13534_;
  assign new_n13536_ = ng4983 & new_n11040_;
  assign new_n13537_ = ~new_n5679_ & new_n13536_;
  assign new_n13538_ = ~new_n13535_ & ~new_n13537_;
  assign new_n13539_ = pg35 & ~new_n13538_;
  assign n5206 = new_n13533_ | new_n13539_;
  assign new_n13541_ = pg35 & ng4944;
  assign new_n13542_ = ~pg35 & new_n13541_;
  assign new_n13543_ = new_n5676_ & new_n5744_;
  assign new_n13544_ = ~ng4045 & ~ng3990;
  assign new_n13545_ = ~ng4054 & new_n13544_;
  assign new_n13546_ = ng4045 & ng3990;
  assign new_n13547_ = ~ng4054 & new_n13546_;
  assign new_n13548_ = ~ng4049 & ~ng3990;
  assign new_n13549_ = ng4054 & new_n13548_;
  assign new_n13550_ = ng4049 & ng3990;
  assign new_n13551_ = ng4054 & new_n13550_;
  assign new_n13552_ = ~new_n13545_ & ~new_n13547_;
  assign new_n13553_ = ~new_n13549_ & ~new_n13551_;
  assign new_n13554_ = new_n13552_ & new_n13553_;
  assign new_n13555_ = ~ng4961 & new_n13554_;
  assign new_n13556_ = new_n13543_ & ~new_n13555_;
  assign new_n13557_ = new_n6467_ & new_n13556_;
  assign new_n13558_ = ng4961 & ~new_n6467_;
  assign new_n13559_ = ~new_n13557_ & ~new_n13558_;
  assign new_n13560_ = pg35 & ~new_n13559_;
  assign n5211 = new_n13542_ | new_n13560_;
  assign new_n13562_ = ~pg35 & ng3490;
  assign new_n13563_ = ng3494 & ~new_n6770_;
  assign new_n13564_ = ng3484 & ~ng3490;
  assign new_n13565_ = ng3484 & ~new_n13564_;
  assign new_n13566_ = ~ng3490 & ~new_n13564_;
  assign new_n13567_ = ~new_n13565_ & ~new_n13566_;
  assign new_n13568_ = new_n6770_ & ~new_n13567_;
  assign new_n13569_ = ~new_n13563_ & ~new_n13568_;
  assign new_n13570_ = pg35 & ~new_n13569_;
  assign n5216 = new_n13562_ | new_n13570_;
  assign new_n13572_ = pg35 & ng4698;
  assign new_n13573_ = ~pg35 & new_n13572_;
  assign new_n13574_ = ~ng5694 & ~ng5644;
  assign new_n13575_ = ~ng5703 & new_n13574_;
  assign new_n13576_ = ng5694 & ng5644;
  assign new_n13577_ = ~ng5703 & new_n13576_;
  assign new_n13578_ = ~ng5698 & ~ng5644;
  assign new_n13579_ = ng5703 & new_n13578_;
  assign new_n13580_ = ng5698 & ng5644;
  assign new_n13581_ = ng5703 & new_n13580_;
  assign new_n13582_ = ~new_n13575_ & ~new_n13577_;
  assign new_n13583_ = ~new_n13579_ & ~new_n13581_;
  assign new_n13584_ = new_n13582_ & new_n13583_;
  assign new_n13585_ = ~ng4749 & new_n13584_;
  assign new_n13586_ = new_n12658_ & ~new_n13585_;
  assign new_n13587_ = new_n7745_ & new_n13586_;
  assign new_n13588_ = ng4749 & ~new_n7745_;
  assign new_n13589_ = ~new_n13587_ & ~new_n13588_;
  assign new_n13590_ = pg35 & ~new_n13589_;
  assign n5221 = new_n13573_ | new_n13590_;
  assign new_n13592_ = ~pg35 & ng2472;
  assign new_n13593_ = ng2421 & ~new_n7558_;
  assign new_n13594_ = ~new_n7555_ & new_n13593_;
  assign new_n13595_ = ng2465 & new_n7555_;
  assign new_n13596_ = ~new_n13594_ & ~new_n13595_;
  assign new_n13597_ = pg35 & ~new_n13596_;
  assign n5226 = new_n13592_ | new_n13597_;
  assign new_n13599_ = pg35 & ng4859;
  assign new_n13600_ = ~pg35 & new_n13599_;
  assign new_n13601_ = ng4917 & ~new_n7449_;
  assign new_n13602_ = n4955 & new_n7449_;
  assign new_n13603_ = ~new_n13601_ & ~new_n13602_;
  assign new_n13604_ = pg35 & ~new_n13603_;
  assign n5231 = new_n13600_ | new_n13604_;
  assign new_n13606_ = ~pg35 & ng1752;
  assign new_n13607_ = ng1728 & ng1802;
  assign new_n13608_ = ~new_n6236_ & new_n13607_;
  assign new_n13609_ = ng1748 & ~new_n13608_;
  assign new_n13610_ = ~new_n10679_ & new_n13608_;
  assign new_n13611_ = ~new_n13609_ & ~new_n13610_;
  assign new_n13612_ = pg35 & ~new_n13611_;
  assign n5240 = new_n13606_ | new_n13612_;
  assign new_n13614_ = pg35 & ng3288;
  assign new_n13615_ = ~pg35 & new_n13614_;
  assign new_n13616_ = pg35 & ng3179;
  assign n5245 = new_n13615_ | new_n13616_;
  assign new_n13618_ = ~pg35 & ng749;
  assign new_n13619_ = ~ng758 & new_n6584_;
  assign new_n13620_ = ng758 & ~new_n6578_;
  assign new_n13621_ = ~new_n6584_ & new_n13620_;
  assign new_n13622_ = ~new_n13619_ & ~new_n13621_;
  assign new_n13623_ = pg35 & ~new_n13622_;
  assign n5249 = new_n13618_ | new_n13623_;
  assign new_n13625_ = ~pg35 & ng1211;
  assign new_n13626_ = pg35 & ng102;
  assign n5254 = new_n13625_ | new_n13626_;
  assign new_n13628_ = ~pg35 & ng1648;
  assign new_n13629_ = ~new_n4724_ & new_n11199_;
  assign new_n13630_ = new_n7230_ & new_n13629_;
  assign new_n13631_ = ng110 & new_n9262_;
  assign new_n13632_ = ng110 & ~new_n13631_;
  assign new_n13633_ = new_n9262_ & ~new_n13631_;
  assign new_n13634_ = ~new_n13632_ & ~new_n13633_;
  assign new_n13635_ = new_n13630_ & ~new_n13634_;
  assign new_n13636_ = ng1664 & ~new_n13630_;
  assign new_n13637_ = ~new_n13635_ & ~new_n13636_;
  assign new_n13638_ = pg35 & ~new_n13637_;
  assign n5258 = new_n13628_ | new_n13638_;
  assign new_n13640_ = ~pg35 & ng518;
  assign new_n13641_ = ng528 & ~new_n6494_;
  assign new_n13642_ = ~new_n6778_ & new_n13641_;
  assign new_n13643_ = ~new_n6494_ & ~new_n6780_;
  assign new_n13644_ = ~ng528 & new_n13643_;
  assign new_n13645_ = new_n6778_ & new_n13644_;
  assign new_n13646_ = ~new_n13642_ & ~new_n13645_;
  assign new_n13647_ = pg35 & ~new_n13646_;
  assign n5263 = new_n13640_ | new_n13647_;
  assign new_n13649_ = ~pg35 & ng94;
  assign new_n13650_ = n4955 & new_n7895_;
  assign new_n13651_ = ~ng2848 & new_n5834_1_;
  assign new_n13652_ = ~new_n13650_ & ~new_n13651_;
  assign new_n13653_ = pg35 & new_n13652_;
  assign n5268 = new_n13649_ | new_n13653_;
  assign new_n13655_ = ~pg35 & ng1548;
  assign new_n13656_ = ~ng1564 & new_n12440_;
  assign new_n13657_ = ng1564 & ~new_n12440_;
  assign new_n13658_ = ~new_n13656_ & ~new_n13657_;
  assign new_n13659_ = pg35 & ~new_n13658_;
  assign n5273 = new_n13655_ | new_n13659_;
  assign new_n13661_ = ~pg35 & ng3805;
  assign new_n13662_ = ng3798 & ~ng3805;
  assign new_n13663_ = ~ng3712 & ~new_n13662_;
  assign new_n13664_ = ~ng3794 & ~new_n13663_;
  assign new_n13665_ = pg35 & new_n13664_;
  assign n5278 = new_n13661_ | new_n13665_;
  assign new_n13667_ = ~pg35 & ng1178;
  assign new_n13668_ = ng1157 & new_n6663_;
  assign new_n13669_ = ng962 & ~new_n13668_;
  assign new_n13670_ = ng996 & new_n13668_;
  assign new_n13671_ = ~new_n13669_ & ~new_n13670_;
  assign new_n13672_ = pg35 & ~new_n13671_;
  assign n5283 = new_n13667_ | new_n13672_;
  assign new_n13674_ = ~pg35 & ng452;
  assign new_n13675_ = ng457 & ~new_n5994_;
  assign new_n13676_ = ng452 & new_n5994_;
  assign new_n13677_ = ~new_n13675_ & ~new_n13676_;
  assign new_n13678_ = pg35 & ~new_n13677_;
  assign n5288 = new_n13674_ | new_n13678_;
  assign new_n13680_ = ~pg35 & ng5782;
  assign new_n13681_ = ng5787 & ~new_n10388_;
  assign new_n13682_ = ~ng5787 & new_n10388_;
  assign new_n13683_ = ~new_n13681_ & ~new_n13682_;
  assign new_n13684_ = pg35 & ~new_n13683_;
  assign n5293 = new_n13680_ | new_n13684_;
  assign new_n13686_ = ~pg35 & ng3827;
  assign new_n13687_ = ng3831 & ~new_n6468_;
  assign new_n13688_ = ng3821 & ~ng3827;
  assign new_n13689_ = ng3821 & ~new_n13688_;
  assign new_n13690_ = ~ng3827 & ~new_n13688_;
  assign new_n13691_ = ~new_n13689_ & ~new_n13690_;
  assign new_n13692_ = new_n6468_ & ~new_n13691_;
  assign new_n13693_ = ~new_n13687_ & ~new_n13692_;
  assign new_n13694_ = pg35 & ~new_n13693_;
  assign n5298 = new_n13686_ | new_n13694_;
  assign new_n13696_ = ~pg35 & ng4818;
  assign new_n13697_ = ~ng4793 & new_n6161_;
  assign new_n13698_ = new_n5670_ & new_n13697_;
  assign new_n13699_ = ng4793 & new_n6161_;
  assign new_n13700_ = ~new_n5670_ & new_n13699_;
  assign new_n13701_ = ~new_n13698_ & ~new_n13700_;
  assign new_n13702_ = pg35 & ~new_n13701_;
  assign n5303 = new_n13696_ | new_n13702_;
  assign new_n13704_ = ~pg35 & ng5813;
  assign new_n13705_ = ng5808 & ~new_n6349_;
  assign new_n13706_ = ~new_n7988_ & new_n13705_;
  assign new_n13707_ = new_n13705_ & ~new_n13706_;
  assign new_n13708_ = ~new_n7988_ & ~new_n13706_;
  assign new_n13709_ = ~new_n13707_ & ~new_n13708_;
  assign new_n13710_ = new_n6353_ & ~new_n13709_;
  assign new_n13711_ = ng5808 & ~new_n6353_;
  assign new_n13712_ = ~new_n13710_ & ~new_n13711_;
  assign new_n13713_ = pg35 & ~new_n13712_;
  assign n5308 = new_n13704_ | new_n13713_;
  assign new_n13715_ = ~pg35 & ng1878;
  assign new_n13716_ = ~new_n6667_1_ & new_n10606_;
  assign new_n13717_ = ng1890 & ~new_n13716_;
  assign new_n13718_ = ~new_n6674_ & new_n13716_;
  assign new_n13719_ = ~new_n13717_ & ~new_n13718_;
  assign new_n13720_ = pg35 & ~new_n13719_;
  assign n5316 = new_n13715_ | new_n13720_;
  assign new_n13722_ = ~pg35 & ng753;
  assign n5321 = new_n7468_ | new_n13722_;
  assign new_n13724_ = ~pg35 & ng5949;
  assign new_n13725_ = ng5869 & new_n7995_;
  assign new_n13726_ = ng5897 & ~new_n13725_;
  assign new_n13727_ = ~new_n5966_ & new_n13725_;
  assign new_n13728_ = ~new_n13726_ & ~new_n13727_;
  assign new_n13729_ = pg35 & ~new_n13728_;
  assign n5326 = new_n13724_ | new_n13729_;
  assign new_n13731_ = ~pg35 & ng3787;
  assign new_n13732_ = ng3787 & new_n7278_;
  assign new_n13733_ = ~ng3791 & new_n13732_;
  assign new_n13734_ = ng3791 & ~new_n13732_;
  assign new_n13735_ = ~new_n13733_ & ~new_n13734_;
  assign new_n13736_ = pg35 & ~new_n13735_;
  assign n5334 = new_n13731_ | new_n13736_;
  assign new_n13738_ = ~pg35 & ng4087;
  assign new_n13739_ = ng4093 & ~new_n10833_;
  assign new_n13740_ = ~ng4093 & new_n10833_;
  assign new_n13741_ = ~new_n13739_ & ~new_n13740_;
  assign new_n13742_ = ng4169 & ~new_n13741_;
  assign new_n13743_ = pg35 & new_n13742_;
  assign n5339 = new_n13738_ | new_n13743_;
  assign new_n13745_ = ~pg35 & ng2625;
  assign new_n13746_ = ~ng2610 & ~new_n10308_;
  assign new_n13747_ = new_n10306_ & ~new_n13746_;
  assign new_n13748_ = ng2619 & ~new_n10306_;
  assign new_n13749_ = ~new_n13747_ & ~new_n13748_;
  assign new_n13750_ = pg35 & ~new_n13749_;
  assign n5344 = new_n13745_ | new_n13750_;
  assign new_n13752_ = ~pg35 & ng718;
  assign new_n13753_ = ng661 & ~new_n7858_;
  assign new_n13754_ = ng718 & new_n7858_;
  assign new_n13755_ = ~new_n13753_ & ~new_n13754_;
  assign new_n13756_ = pg35 & ~new_n13755_;
  assign n5349 = new_n13752_ | new_n13756_;
  assign new_n13758_ = ~pg35 & ng1542;
  assign new_n13759_ = ng1542 & new_n6831_;
  assign new_n13760_ = ng1413 & new_n6843_;
  assign new_n13761_ = ~new_n13759_ & new_n13760_;
  assign new_n13762_ = ~ng1413 & new_n6843_;
  assign new_n13763_ = new_n13759_ & new_n13762_;
  assign new_n13764_ = ~new_n13761_ & ~new_n13763_;
  assign new_n13765_ = pg35 & ~new_n13764_;
  assign n5358 = new_n13758_ | new_n13765_;
  assign new_n13767_ = ~pg35 & ng2315;
  assign new_n13768_ = ~new_n7886_ & new_n11295_;
  assign new_n13769_ = ng2311 & ~new_n13768_;
  assign new_n13770_ = ~new_n8906_ & new_n13768_;
  assign new_n13771_ = ~new_n13769_ & ~new_n13770_;
  assign new_n13772_ = pg35 & ~new_n13771_;
  assign n5363 = new_n13767_ | new_n13772_;
  assign new_n13774_ = ~pg35 & ng5770;
  assign new_n13775_ = ~ng5759 & ng5767;
  assign new_n13776_ = ~ng5770 & ~new_n13775_;
  assign new_n13777_ = ~ng5774 & new_n13776_;
  assign new_n13778_ = ng5774 & ng5770;
  assign new_n13779_ = ~ng5763 & ng5767;
  assign new_n13780_ = ~new_n13777_ & ~new_n13778_;
  assign new_n13781_ = ~new_n13779_ & new_n13780_;
  assign new_n13782_ = pg35 & ~new_n13781_;
  assign n5368 = new_n13774_ | new_n13782_;
  assign new_n13784_ = ~pg35 & ng790;
  assign new_n13785_ = ~ng794 & new_n12500_;
  assign new_n13786_ = ng794 & ~new_n6578_;
  assign new_n13787_ = ~new_n12500_ & new_n13786_;
  assign new_n13788_ = ~new_n13785_ & ~new_n13787_;
  assign new_n13789_ = pg35 & ~new_n13788_;
  assign n5378 = new_n13784_ | new_n13789_;
  assign new_n13791_ = pg35 & ng4578;
  assign new_n13792_ = ~pg35 & new_n13791_;
  assign n5383 = new_n8767_ | new_n13792_;
  assign new_n13794_ = ~pg35 & ng2661;
  assign new_n13795_ = ng2667 & ~new_n13235_;
  assign new_n13796_ = ng2661 & new_n13235_;
  assign new_n13797_ = ~new_n13795_ & ~new_n13796_;
  assign new_n13798_ = pg35 & ~new_n13797_;
  assign n5387 = new_n13794_ | new_n13798_;
  assign new_n13800_ = pg35 & ng2551;
  assign new_n13801_ = ~pg35 & new_n13800_;
  assign new_n13802_ = ng2555 & ~ng2629;
  assign new_n13803_ = ~ng2599 & ~ng2629;
  assign new_n13804_ = ~new_n13802_ & ~new_n13803_;
  assign new_n13805_ = ~new_n7177_ & ~new_n13804_;
  assign new_n13806_ = ~new_n7174_ & new_n13805_;
  assign new_n13807_ = ng2555 & new_n7174_;
  assign new_n13808_ = ~new_n13806_ & ~new_n13807_;
  assign new_n13809_ = pg35 & ~new_n13808_;
  assign n5392 = new_n13801_ | new_n13809_;
  assign new_n13811_ = ~pg35 & ng4462;
  assign new_n13812_ = ~ng4473 & ~ng4467;
  assign new_n13813_ = pg35 & new_n13812_;
  assign n5397 = new_n13811_ | new_n13813_;
  assign new_n13815_ = ~pg35 & ng1620;
  assign new_n13816_ = ng1636 & ~ng1592;
  assign new_n13817_ = ~new_n7537_1_ & new_n13816_;
  assign new_n13818_ = ng1616 & ~new_n13817_;
  assign new_n13819_ = ~new_n7543_ & new_n13817_;
  assign new_n13820_ = ~new_n13818_ & ~new_n13819_;
  assign new_n13821_ = pg35 & ~new_n13820_;
  assign n5402 = new_n13815_ | new_n13821_;
  assign new_n13823_ = pg35 & ng4242;
  assign new_n13824_ = ~pg35 & new_n13823_;
  assign new_n13825_ = pg6745 & pg35;
  assign n5407 = new_n13824_ | new_n13825_;
  assign new_n13827_ = ~pg35 & ng225;
  assign new_n13828_ = ng869 & new_n6112_;
  assign new_n13829_ = ng255 & ~new_n6112_;
  assign new_n13830_ = ~new_n13828_ & ~new_n13829_;
  assign new_n13831_ = pg35 & ~new_n13830_;
  assign n5412 = new_n13827_ | new_n13831_;
  assign new_n13833_ = ~pg35 & ng3419;
  assign new_n13834_ = ~ng3419 & ~new_n11439_;
  assign new_n13835_ = ~ng3423 & new_n13834_;
  assign new_n13836_ = ng3419 & ng3423;
  assign new_n13837_ = ~new_n13835_ & ~new_n13836_;
  assign new_n13838_ = ~new_n11441_ & new_n13837_;
  assign new_n13839_ = pg35 & ~new_n13838_;
  assign n5417 = new_n13833_ | new_n13839_;
  assign new_n13841_ = ~pg35 & ng608;
  assign new_n13842_ = ng613 & ~new_n6545_;
  assign new_n13843_ = ~new_n9118_ & new_n13842_;
  assign new_n13844_ = ~ng613 & new_n9118_;
  assign new_n13845_ = ~new_n13843_ & ~new_n13844_;
  assign new_n13846_ = pg35 & ~new_n13845_;
  assign n5422 = new_n13841_ | new_n13846_;
  assign new_n13848_ = ~pg35 & ng5385;
  assign new_n13849_ = ~new_n12295_ & ~new_n12297_;
  assign new_n13850_ = ~ng5390 & ~new_n13849_;
  assign new_n13851_ = ng5390 & new_n6394_;
  assign new_n13852_ = new_n13849_ & new_n13851_;
  assign new_n13853_ = ~new_n13850_ & ~new_n13852_;
  assign new_n13854_ = pg35 & ~new_n13853_;
  assign n5427 = new_n13848_ | new_n13854_;
  assign new_n13856_ = ~pg35 & ng3029;
  assign new_n13857_ = ~new_n11900_ & ~new_n11903_;
  assign new_n13858_ = ~ng3034 & ~new_n13857_;
  assign new_n13859_ = ng3034 & new_n8954_;
  assign new_n13860_ = new_n13857_ & new_n13859_;
  assign new_n13861_ = ~new_n13858_ & ~new_n13860_;
  assign new_n13862_ = pg35 & ~new_n13861_;
  assign n5432 = new_n13856_ | new_n13862_;
  assign new_n13864_ = ~pg35 & ng812;
  assign new_n13865_ = ng817 & new_n8009_;
  assign new_n13866_ = ~new_n6067_ & new_n13865_;
  assign new_n13867_ = ~ng817 & new_n8009_;
  assign new_n13868_ = new_n6067_ & new_n13867_;
  assign new_n13869_ = ~new_n13866_ & ~new_n13868_;
  assign new_n13870_ = pg35 & ~new_n13869_;
  assign n5437 = new_n13864_ | new_n13870_;
  assign new_n13872_ = ~pg35 & ng691;
  assign new_n13873_ = ng703 & new_n9928_;
  assign new_n13874_ = ~ng691 & new_n13873_;
  assign new_n13875_ = new_n6493_1_ & ~new_n13874_;
  assign new_n13876_ = ng686 & ~new_n6493_1_;
  assign new_n13877_ = ~new_n13875_ & ~new_n13876_;
  assign new_n13878_ = pg35 & ~new_n13877_;
  assign n5442 = new_n13872_ | new_n13878_;
  assign new_n13880_ = ~pg35 & ng4486;
  assign n5447 = new_n13281_ | new_n13880_;
  assign new_n13882_ = ~pg35 & ng4961;
  assign new_n13883_ = ~new_n6055_1_ & ~new_n13543_;
  assign new_n13884_ = ng4961 & ~new_n6055_1_;
  assign new_n13885_ = ~new_n6058_ & ~new_n13884_;
  assign new_n13886_ = ~new_n13883_ & ~new_n13885_;
  assign new_n13887_ = ng4955 & new_n13883_;
  assign new_n13888_ = ~new_n13886_ & ~new_n13887_;
  assign new_n13889_ = pg35 & ~new_n13888_;
  assign n5452 = new_n13882_ | new_n13889_;
  assign new_n13891_ = ~pg35 & ng2671;
  assign new_n13892_ = ng2675 & ~new_n13235_;
  assign new_n13893_ = ~ng2675 & new_n13235_;
  assign new_n13894_ = ~new_n13892_ & ~new_n13893_;
  assign new_n13895_ = pg35 & ~new_n13894_;
  assign n5457 = new_n13891_ | new_n13895_;
  assign n5462 = ng12 | ng25;
  assign new_n13898_ = ~pg35 & ng901;
  assign new_n13899_ = pg35 & ng901;
  assign n5467 = new_n13898_ | new_n13899_;
  assign new_n13901_ = ~pg35 & ng319;
  assign new_n13902_ = pg35 & ng319;
  assign n5472 = new_n13901_ | new_n13902_;
  assign new_n13904_ = ~pg35 & ng5723;
  assign new_n13905_ = ~new_n6707_ & ~new_n6709_;
  assign new_n13906_ = ~ng5727 & ~new_n13905_;
  assign new_n13907_ = ng5727 & new_n6424_;
  assign new_n13908_ = new_n13905_ & new_n13907_;
  assign new_n13909_ = ~new_n13906_ & ~new_n13908_;
  assign new_n13910_ = pg35 & ~new_n13909_;
  assign n5485 = new_n13904_ | new_n13910_;
  assign new_n13912_ = ~pg35 & ng6434;
  assign new_n13913_ = ~ng6434 & new_n8596_;
  assign new_n13914_ = ng6434 & new_n8597_;
  assign new_n13915_ = ~new_n13913_ & ~new_n13914_;
  assign new_n13916_ = ~ng6439 & ~new_n13915_;
  assign new_n13917_ = ng6439 & new_n6632_1_;
  assign new_n13918_ = new_n13915_ & new_n13917_;
  assign new_n13919_ = ~new_n13916_ & ~new_n13918_;
  assign new_n13920_ = pg35 & ~new_n13919_;
  assign n5490 = new_n13912_ | new_n13920_;
  assign new_n13922_ = ~pg35 & ng2527;
  assign new_n13923_ = ng2533 & ~new_n9787_;
  assign new_n13924_ = ng2527 & new_n9787_;
  assign new_n13925_ = ~new_n13923_ & ~new_n13924_;
  assign new_n13926_ = pg35 & ~new_n13925_;
  assign n5495 = new_n13922_ | new_n13926_;
  assign new_n13928_ = ~pg35 & ng6497;
  assign new_n13929_ = ~ng6497 & ng6490;
  assign new_n13930_ = ~ng6404 & ~new_n13929_;
  assign new_n13931_ = ~ng6486 & ~new_n13930_;
  assign new_n13932_ = pg35 & new_n13931_;
  assign n5500 = new_n13928_ | new_n13932_;
  assign new_n13934_ = ~pg35 & ng2922;
  assign new_n13935_ = n2287 & new_n9379_;
  assign new_n13936_ = ng2936 & ~new_n9379_;
  assign new_n13937_ = ~new_n13935_ & ~new_n13936_;
  assign new_n13938_ = pg35 & ~new_n13937_;
  assign n5505 = new_n13934_ | new_n13938_;
  assign new_n13940_ = ~pg35 & ng6283;
  assign new_n13941_ = new_n5849_ & new_n7865_;
  assign new_n13942_ = ng6299 & ~new_n13941_;
  assign new_n13943_ = ~new_n5966_ & new_n13941_;
  assign new_n13944_ = ~new_n13942_ & ~new_n13943_;
  assign new_n13945_ = pg35 & ~new_n13944_;
  assign n5514 = new_n13940_ | new_n13945_;
  assign new_n13947_ = ~pg35 & ng3065;
  assign new_n13948_ = ng3072 & new_n11967_;
  assign new_n13949_ = ~ng3072 & new_n11971_;
  assign new_n13950_ = ~new_n13948_ & ~new_n13949_;
  assign new_n13951_ = pg35 & ~new_n13950_;
  assign n5519 = new_n13947_ | new_n13951_;
  assign new_n13953_ = ~pg35 & ng316;
  assign new_n13954_ = pg35 & ~new_n7288_;
  assign n5524 = new_n13953_ | new_n13954_;
  assign new_n13956_ = ~pg35 & ng1312;
  assign new_n13957_ = ng1351 & new_n6294_;
  assign new_n13958_ = ng1351 & ~new_n6300_1_;
  assign new_n13959_ = new_n6298_ & new_n13958_;
  assign new_n13960_ = ng1312 & ~new_n6298_;
  assign new_n13961_ = ng1351 & ~new_n6298_;
  assign new_n13962_ = ~ng1389 & ~new_n6300_1_;
  assign new_n13963_ = new_n13961_ & new_n13962_;
  assign new_n13964_ = ~new_n13959_ & ~new_n13960_;
  assign new_n13965_ = ~new_n13963_ & new_n13964_;
  assign new_n13966_ = ~new_n6294_ & ~new_n13965_;
  assign new_n13967_ = ~new_n13957_ & ~new_n13966_;
  assign new_n13968_ = pg35 & ~new_n13967_;
  assign n5529 = new_n13956_ | new_n13968_;
  assign new_n13970_ = ~pg35 & ng661;
  assign new_n13971_ = ng728 & ~new_n7858_;
  assign new_n13972_ = ng661 & new_n7858_;
  assign new_n13973_ = ~new_n13971_ & ~new_n13972_;
  assign new_n13974_ = pg35 & ~new_n13973_;
  assign n5537 = new_n13970_ | new_n13974_;
  assign new_n13976_ = ~pg35 & ng2070;
  assign new_n13977_ = ng2084 & ~new_n8021_;
  assign new_n13978_ = ~ng1246 & new_n7020_;
  assign new_n13979_ = ~new_n7030_ & ~new_n13978_;
  assign new_n13980_ = new_n13977_ & ~new_n13979_;
  assign new_n13981_ = new_n13977_ & ~new_n13980_;
  assign new_n13982_ = ~new_n13979_ & ~new_n13980_;
  assign new_n13983_ = ~new_n13981_ & ~new_n13982_;
  assign new_n13984_ = ~new_n7025_ & ~new_n13983_;
  assign new_n13985_ = ng2084 & new_n7025_;
  assign new_n13986_ = ~new_n13984_ & ~new_n13985_;
  assign new_n13987_ = pg35 & ~new_n13986_;
  assign n5542 = new_n13976_ | new_n13987_;
  assign new_n13989_ = ~pg35 & ng79;
  assign new_n13990_ = ~ng691 & new_n13874_;
  assign new_n13991_ = ng714 & ng691;
  assign new_n13992_ = ng703 & ~new_n13991_;
  assign new_n13993_ = ng691 & new_n13992_;
  assign new_n13994_ = ~new_n13990_ & ~new_n13993_;
  assign new_n13995_ = new_n6493_1_ & ~new_n13994_;
  assign new_n13996_ = ng691 & ~new_n6493_1_;
  assign new_n13997_ = ~new_n13995_ & ~new_n13996_;
  assign new_n13998_ = pg35 & ~new_n13997_;
  assign n5547 = new_n13989_ | new_n13998_;
  assign new_n14000_ = ~pg35 & ng5694;
  assign new_n14001_ = ng5694 & ~new_n11654_;
  assign new_n14002_ = pg35 & new_n14001_;
  assign n5552 = new_n14000_ | new_n14002_;
  assign new_n14004_ = ~pg35 & ng4527;
  assign new_n14005_ = ng4515 & ng4521;
  assign new_n14006_ = ~ng4527 & new_n7765_;
  assign new_n14007_ = ng4527 & ~new_n7765_;
  assign new_n14008_ = ~new_n14006_ & ~new_n14007_;
  assign new_n14009_ = ~ng4521 & ~new_n14008_;
  assign new_n14010_ = ~new_n14005_ & ~new_n14009_;
  assign new_n14011_ = pg35 & ~new_n14010_;
  assign n5557 = new_n14004_ | new_n14011_;
  assign new_n14013_ = ~pg35 & ng1886;
  assign new_n14014_ = ng1936 & ng1862;
  assign new_n14015_ = ~new_n6667_1_ & new_n14014_;
  assign new_n14016_ = ng1882 & ~new_n14015_;
  assign new_n14017_ = ~new_n6674_ & new_n14015_;
  assign new_n14018_ = ~new_n14016_ & ~new_n14017_;
  assign new_n14019_ = pg35 & ~new_n14018_;
  assign n5562 = new_n14013_ | new_n14019_;
  assign new_n14021_ = ~pg35 & ng6395;
  assign new_n14022_ = ng6395 & new_n6699_;
  assign new_n14023_ = new_n6699_ & new_n13104_;
  assign new_n14024_ = new_n4734_ & new_n14023_;
  assign new_n14025_ = ng6336 & ~new_n14024_;
  assign new_n14026_ = ~new_n14022_ & new_n14025_;
  assign new_n14027_ = ~ng6336 & ~new_n14024_;
  assign new_n14028_ = new_n14022_ & new_n14027_;
  assign new_n14029_ = ~new_n14026_ & ~new_n14028_;
  assign new_n14030_ = pg35 & ~new_n14029_;
  assign n5570 = new_n14021_ | new_n14030_;
  assign new_n14032_ = ~pg35 & ng5128;
  assign new_n14033_ = ng5134 & ~new_n6191_;
  assign new_n14034_ = ng5128 & new_n6191_;
  assign new_n14035_ = ~new_n14033_ & ~new_n14034_;
  assign new_n14036_ = pg35 & ~new_n14035_;
  assign n5575 = new_n14032_ | new_n14036_;
  assign new_n14038_ = ~pg35 & ng4082;
  assign new_n14039_ = ng4076 & ~new_n7186_;
  assign new_n14040_ = ~ng4076 & new_n7186_;
  assign new_n14041_ = ~new_n14039_ & ~new_n14040_;
  assign new_n14042_ = ng4169 & ~new_n14041_;
  assign new_n14043_ = ng4169 & ~new_n14042_;
  assign new_n14044_ = pg35 & ~new_n14043_;
  assign n5580 = new_n14038_ | new_n14044_;
  assign new_n14046_ = ~pg35 & ng1489;
  assign new_n14047_ = ng1495 & ~new_n6433_;
  assign new_n14048_ = ng1489 & new_n6433_;
  assign new_n14049_ = ~new_n14047_ & ~new_n14048_;
  assign new_n14050_ = pg35 & ~new_n14049_;
  assign n5585 = new_n14046_ | new_n14050_;
  assign new_n14052_ = ~pg35 & ng3034;
  assign new_n14053_ = ~new_n11901_ & ~new_n11904_;
  assign new_n14054_ = ng3040 & new_n8954_;
  assign new_n14055_ = new_n14053_ & new_n14054_;
  assign new_n14056_ = ~ng3040 & ~new_n14053_;
  assign new_n14057_ = ~new_n14055_ & ~new_n14056_;
  assign new_n14058_ = pg35 & ~new_n14057_;
  assign n5590 = new_n14052_ | new_n14058_;
  assign new_n14060_ = pg35 & ng5152;
  assign new_n14061_ = ~pg35 & new_n14060_;
  assign new_n14062_ = n2287 & new_n6181_;
  assign new_n14063_ = ng5160 & ~new_n6181_;
  assign new_n14064_ = ~new_n14062_ & ~new_n14063_;
  assign new_n14065_ = pg35 & ~new_n14064_;
  assign n5598 = new_n14061_ | new_n14065_;
  assign new_n14067_ = ~pg35 & ng962;
  assign new_n14068_ = ng1157 & ng1178;
  assign new_n14069_ = ~ng1157 & ng1189;
  assign new_n14070_ = ~new_n14068_ & ~new_n14069_;
  assign new_n14071_ = pg35 & ~new_n14070_;
  assign n5603 = new_n14067_ | new_n14071_;
  assign new_n14073_ = ~pg35 & ng3368;
  assign new_n14074_ = ~new_n10778_ & ~new_n10783_;
  assign new_n14075_ = ng3372 & new_n8400_;
  assign new_n14076_ = new_n14074_ & new_n14075_;
  assign new_n14077_ = ~ng3372 & ~new_n14074_;
  assign new_n14078_ = ~new_n14076_ & ~new_n14077_;
  assign new_n14079_ = pg35 & ~new_n14078_;
  assign n5608 = new_n14073_ | new_n14079_;
  assign new_n14081_ = ~pg35 & ng441;
  assign new_n14082_ = ng437 & ~new_n6067_;
  assign new_n14083_ = ng441 & new_n6067_;
  assign new_n14084_ = ~new_n14082_ & ~new_n14083_;
  assign new_n14085_ = pg35 & ~new_n14084_;
  assign n5613 = new_n14081_ | new_n14085_;
  assign new_n14087_ = pg35 & ng5445;
  assign new_n14088_ = ~pg35 & new_n14087_;
  assign new_n14089_ = ~ng5511 & new_n10862_;
  assign new_n14090_ = pg35 & new_n14089_;
  assign n5618 = new_n14088_ | new_n14090_;
  assign new_n14092_ = ~pg35 & ng3961;
  assign new_n14093_ = ng3965 & ~new_n7011_1_;
  assign new_n14094_ = ~new_n5966_ & new_n7011_1_;
  assign new_n14095_ = ~new_n14093_ & ~new_n14094_;
  assign new_n14096_ = pg35 & ~new_n14095_;
  assign n5623 = new_n14092_ | new_n14096_;
  assign new_n14098_ = ~pg35 & ng6479;
  assign new_n14099_ = ng6479 & new_n12835_;
  assign new_n14100_ = ~ng6483 & new_n14099_;
  assign new_n14101_ = ng6483 & ~new_n14099_;
  assign new_n14102_ = ~new_n14100_ & ~new_n14101_;
  assign new_n14103_ = pg35 & ~new_n14102_;
  assign n5628 = new_n14098_ | new_n14103_;
  assign new_n14105_ = ~pg35 & ng6181;
  assign new_n14106_ = ng6187 & ~new_n7064_;
  assign new_n14107_ = ng6181 & new_n7064_;
  assign new_n14108_ = ~new_n14106_ & ~new_n14107_;
  assign new_n14109_ = pg35 & ~new_n14108_;
  assign n5633 = new_n14105_ | new_n14109_;
  assign new_n14111_ = ~pg35 & ng911;
  assign new_n14112_ = ~ng914 & new_n7077_;
  assign new_n14113_ = ng1227 & ng914;
  assign new_n14114_ = ~new_n7077_ & new_n14113_;
  assign new_n14115_ = ~new_n14112_ & ~new_n14114_;
  assign new_n14116_ = pg35 & ~new_n14115_;
  assign n5638 = new_n14111_ | new_n14116_;
  assign new_n14118_ = ~pg35 & ng5603;
  assign new_n14119_ = ng5523 & new_n8033_;
  assign new_n14120_ = ng5551 & ~new_n14119_;
  assign new_n14121_ = ~new_n5966_ & new_n14119_;
  assign new_n14122_ = ~new_n14120_ & ~new_n14121_;
  assign new_n14123_ = pg35 & ~new_n14122_;
  assign n5643 = new_n14118_ | new_n14123_;
  assign new_n14125_ = ~pg35 & ng1367;
  assign new_n14126_ = new_n13369_ & ~new_n13371_;
  assign new_n14127_ = ng1373 & ~new_n14126_;
  assign new_n14128_ = ~ng1373 & new_n6306_;
  assign new_n14129_ = new_n14126_ & new_n14128_;
  assign new_n14130_ = ~new_n14127_ & ~new_n14129_;
  assign new_n14131_ = pg35 & ~new_n14130_;
  assign n5648 = new_n14125_ | new_n14131_;
  assign new_n14133_ = ~pg35 & ng5805;
  assign new_n14134_ = ng5798 & ~ng5805;
  assign new_n14135_ = ~ng5712 & ~new_n14134_;
  assign new_n14136_ = ~ng5794 & ~new_n14135_;
  assign new_n14137_ = pg35 & new_n14136_;
  assign n5653 = new_n14133_ | new_n14137_;
  assign new_n14139_ = ~pg35 & ng626;
  assign new_n14140_ = ~new_n6545_ & new_n9124_;
  assign new_n14141_ = ng626 & new_n14140_;
  assign new_n14142_ = ng632 & ~new_n6545_;
  assign new_n14143_ = ~new_n14141_ & new_n14142_;
  assign new_n14144_ = ~ng632 & new_n14141_;
  assign new_n14145_ = ~new_n14143_ & ~new_n14144_;
  assign new_n14146_ = pg35 & ~new_n14145_;
  assign n5658 = new_n14139_ | new_n14146_;
  assign new_n14148_ = ~pg35 & ng1242;
  assign new_n14149_ = pg35 & ng1227;
  assign n5663 = new_n14148_ | new_n14149_;
  assign new_n14151_ = ~pg35 & ng4495;
  assign new_n14152_ = ~ng59 & new_n7110_;
  assign new_n14153_ = ng4581 & ~new_n14152_;
  assign new_n14154_ = ng4495 & ~ng4581;
  assign new_n14155_ = ~new_n14153_ & ~new_n14154_;
  assign new_n14156_ = pg35 & ~new_n14155_;
  assign n5668 = new_n14151_ | new_n14156_;
  assign new_n14158_ = ~pg35 & ng2227;
  assign new_n14159_ = ng2241 & ~new_n6523_1_;
  assign new_n14160_ = ng1589 & new_n6513_1_;
  assign new_n14161_ = ~new_n6723_ & ~new_n14160_;
  assign new_n14162_ = new_n14159_ & ~new_n14161_;
  assign new_n14163_ = new_n14159_ & ~new_n14162_;
  assign new_n14164_ = ~new_n14161_ & ~new_n14162_;
  assign new_n14165_ = ~new_n14163_ & ~new_n14164_;
  assign new_n14166_ = ~new_n6522_ & ~new_n14165_;
  assign new_n14167_ = ng2241 & new_n6522_;
  assign new_n14168_ = ~new_n14166_ & ~new_n14167_;
  assign new_n14169_ = pg35 & ~new_n14168_;
  assign n5677 = new_n14158_ | new_n14169_;
  assign new_n14171_ = ~pg35 & ng2351;
  assign new_n14172_ = ~ng2342 & ng2319;
  assign new_n14173_ = ng2311 & new_n14172_;
  assign new_n14174_ = ~ng2319 & ~ng2351;
  assign new_n14175_ = ng2307 & new_n14174_;
  assign new_n14176_ = ng2315 & new_n5217_;
  assign new_n14177_ = ~new_n14173_ & ~new_n14175_;
  assign new_n14178_ = ~new_n14176_ & new_n14177_;
  assign new_n14179_ = ng2342 & ~ng2319;
  assign new_n14180_ = ng2295 & new_n14179_;
  assign new_n14181_ = ng2299 & new_n7255_;
  assign new_n14182_ = ~ng2342 & ng2351;
  assign new_n14183_ = ng2303 & new_n14182_;
  assign new_n14184_ = new_n14178_ & ~new_n14180_;
  assign new_n14185_ = ~new_n14181_ & ~new_n14183_;
  assign new_n14186_ = new_n14184_ & new_n14185_;
  assign new_n14187_ = new_n7259_ & ~new_n14186_;
  assign new_n14188_ = ng2370 & ~new_n7259_;
  assign new_n14189_ = ~new_n14187_ & ~new_n14188_;
  assign new_n14190_ = pg35 & ~new_n14189_;
  assign n5682 = new_n14171_ | new_n14190_;
  assign new_n14192_ = ~pg35 & ng5767;
  assign new_n14193_ = ng5774 & new_n13775_;
  assign new_n14194_ = ~ng5774 & new_n13779_;
  assign new_n14195_ = ~new_n14193_ & ~new_n14194_;
  assign new_n14196_ = pg35 & ~new_n14195_;
  assign n5687 = new_n14192_ | new_n14196_;
  assign new_n14198_ = ~pg35 & ng2748;
  assign new_n14199_ = ~ng2756 & new_n6644_;
  assign new_n14200_ = ng2756 & ~new_n6644_;
  assign new_n14201_ = ~new_n14199_ & ~new_n14200_;
  assign new_n14202_ = ng2841 & ~new_n14201_;
  assign new_n14203_ = ng2841 & ~new_n14202_;
  assign new_n14204_ = pg35 & ~new_n14203_;
  assign n5692 = new_n14198_ | new_n14204_;
  assign new_n14206_ = ~pg35 & ng3431;
  assign new_n14207_ = ng3436 & ~new_n13509_;
  assign new_n14208_ = ~ng3436 & new_n13509_;
  assign new_n14209_ = ~new_n14207_ & ~new_n14208_;
  assign new_n14210_ = pg35 & ~new_n14209_;
  assign n5697 = new_n14206_ | new_n14210_;
  assign new_n14212_ = ~pg35 & ng2509;
  assign new_n14213_ = ng2514 & ~new_n9787_;
  assign new_n14214_ = ng2509 & new_n9787_;
  assign new_n14215_ = ~new_n14213_ & ~new_n14214_;
  assign new_n14216_ = pg35 & ~new_n14215_;
  assign n5702 = new_n14212_ | new_n14216_;
  assign new_n14218_ = ~pg35 & ng2759;
  assign new_n14219_ = ng2759 & new_n6645_;
  assign new_n14220_ = ~ng2763 & new_n14219_;
  assign new_n14221_ = ng2763 & ~new_n14219_;
  assign new_n14222_ = ~new_n14220_ & ~new_n14221_;
  assign new_n14223_ = ng2841 & ~new_n14222_;
  assign new_n14224_ = ng2841 & ~new_n14223_;
  assign new_n14225_ = pg35 & ~new_n14224_;
  assign n5707 = new_n14218_ | new_n14225_;
  assign new_n14227_ = ~pg35 & ng6629;
  assign new_n14228_ = new_n7159_ & new_n7456_;
  assign new_n14229_ = ng6645 & ~new_n14228_;
  assign new_n14230_ = ~new_n5966_ & new_n14228_;
  assign new_n14231_ = ~new_n14229_ & ~new_n14230_;
  assign new_n14232_ = pg35 & ~new_n14231_;
  assign n5712 = new_n14227_ | new_n14232_;
  assign new_n14234_ = ~pg35 & ng3863;
  assign new_n14235_ = new_n8079_ & new_n11021_;
  assign new_n14236_ = ng3869 & new_n11021_;
  assign new_n14237_ = ~new_n8079_ & new_n14236_;
  assign new_n14238_ = ~new_n14235_ & ~new_n14237_;
  assign new_n14239_ = pg35 & ~new_n14238_;
  assign n5717 = new_n14234_ | new_n14239_;
  assign new_n14241_ = ~pg35 & ng2599;
  assign new_n14242_ = ng2599 & ~new_n7177_;
  assign new_n14243_ = ~new_n7174_ & new_n14242_;
  assign new_n14244_ = ng2629 & new_n7174_;
  assign new_n14245_ = ~new_n14243_ & ~new_n14244_;
  assign new_n14246_ = pg35 & ~new_n14245_;
  assign n5722 = new_n14241_ | new_n14246_;
  assign new_n14248_ = ng22 & pg34913;
  assign new_n14249_ = ~ng22 & n4955;
  assign n5727 = new_n14248_ | new_n14249_;
  assign new_n14251_ = pg35 & ng3853;
  assign new_n14252_ = ~pg35 & new_n14251_;
  assign n5732 = new_n5884_ | new_n14252_;
  assign new_n14254_ = ~pg35 & ng3703;
  assign new_n14255_ = ng3703 & new_n7431_;
  assign new_n14256_ = ng3639 & ~new_n11318_;
  assign new_n14257_ = ~new_n14255_ & new_n14256_;
  assign new_n14258_ = ~ng3639 & ~new_n11318_;
  assign new_n14259_ = new_n14255_ & new_n14258_;
  assign new_n14260_ = ~new_n14257_ & ~new_n14259_;
  assign new_n14261_ = pg35 & ~new_n14260_;
  assign n5737 = new_n14254_ | new_n14261_;
  assign new_n14263_ = ~pg35 & ng239;
  assign new_n14264_ = ng884 & new_n6112_;
  assign new_n14265_ = ng269 & ~new_n6112_;
  assign new_n14266_ = ~new_n14264_ & ~new_n14265_;
  assign new_n14267_ = pg35 & ~new_n14266_;
  assign n5742 = new_n14263_ | new_n14267_;
  assign new_n14269_ = ~pg35 & ng3941;
  assign new_n14270_ = new_n6874_ & new_n8079_;
  assign new_n14271_ = ng3957 & ~new_n14270_;
  assign new_n14272_ = ~new_n5966_ & new_n14270_;
  assign new_n14273_ = ~new_n14271_ & ~new_n14272_;
  assign new_n14274_ = pg35 & ~new_n14273_;
  assign n5747 = new_n14269_ | new_n14274_;
  assign new_n14276_ = ~pg35 & ng1171;
  assign new_n14277_ = ng1171 & ng1157;
  assign new_n14278_ = ~ng1183 & new_n5953_;
  assign new_n14279_ = ~new_n14277_ & ~new_n14278_;
  assign new_n14280_ = ng1183 & new_n5953_;
  assign new_n14281_ = new_n14277_ & ~new_n14280_;
  assign new_n14282_ = ~new_n14279_ & ~new_n14281_;
  assign new_n14283_ = pg35 & ~new_n14282_;
  assign n5752 = new_n14276_ | new_n14283_;
  assign new_n14285_ = ~pg35 & ng5763;
  assign new_n14286_ = ng5759 & ng5763;
  assign new_n14287_ = pg35 & new_n14286_;
  assign n5757 = new_n14285_ | new_n14287_;
  assign new_n14289_ = ~pg35 & ng4664;
  assign new_n14290_ = ng4653 & ng4688;
  assign new_n14291_ = ng4659 & new_n14290_;
  assign new_n14292_ = ng4664 & new_n14291_;
  assign new_n14293_ = ng4669 & new_n10528_;
  assign new_n14294_ = ~new_n14292_ & new_n14293_;
  assign new_n14295_ = ~ng4669 & new_n10528_;
  assign new_n14296_ = new_n14292_ & new_n14295_;
  assign new_n14297_ = ~new_n14294_ & ~new_n14296_;
  assign new_n14298_ = pg35 & ~new_n14297_;
  assign n5762 = new_n14289_ | new_n14298_;
  assign new_n14300_ = ~pg35 & ng3586;
  assign new_n14301_ = new_n7038_ & new_n7697_;
  assign new_n14302_ = ng3602 & ~new_n14301_;
  assign new_n14303_ = ~new_n5966_ & new_n14301_;
  assign new_n14304_ = ~new_n14302_ & ~new_n14303_;
  assign new_n14305_ = pg35 & ~new_n14304_;
  assign n5771 = new_n14300_ | new_n14305_;
  assign new_n14307_ = ~pg35 & ng4681;
  assign new_n14308_ = ng4681 & ~new_n8716_;
  assign new_n14309_ = pg35 & new_n14308_;
  assign n5776 = new_n14307_ | new_n14309_;
  assign new_n14311_ = ~pg35 & ng3207;
  assign new_n14312_ = new_n7151_ & new_n9315_;
  assign new_n14313_ = ng3227 & ~new_n14312_;
  assign new_n14314_ = ~new_n5966_ & new_n14312_;
  assign new_n14315_ = ~new_n14313_ & ~new_n14314_;
  assign new_n14316_ = pg35 & ~new_n14315_;
  assign n5781 = new_n14311_ | new_n14316_;
  assign new_n14318_ = ~pg35 & ng2047;
  assign new_n14319_ = ng1996 & ~new_n9212_;
  assign new_n14320_ = ~new_n7025_ & new_n14319_;
  assign new_n14321_ = ng2040 & new_n7025_;
  assign new_n14322_ = ~new_n14320_ & ~new_n14321_;
  assign new_n14323_ = pg35 & ~new_n14322_;
  assign n5789 = new_n14318_ | new_n14323_;
  assign new_n14325_ = ~pg35 & ng3391;
  assign new_n14326_ = ~ng3391 & new_n10782_;
  assign new_n14327_ = ng3391 & new_n10787_;
  assign new_n14328_ = ~new_n14326_ & ~new_n14327_;
  assign new_n14329_ = ~ng3396 & ~new_n14328_;
  assign new_n14330_ = ng3396 & new_n8400_;
  assign new_n14331_ = new_n14328_ & new_n14330_;
  assign new_n14332_ = ~new_n14329_ & ~new_n14331_;
  assign new_n14333_ = pg35 & ~new_n14332_;
  assign n5794 = new_n14325_ | new_n14333_;
  assign new_n14335_ = ~pg35 & ng6073;
  assign new_n14336_ = ~new_n10188_ & ~new_n10192_;
  assign new_n14337_ = ng6077 & new_n7527_;
  assign new_n14338_ = new_n14336_ & new_n14337_;
  assign new_n14339_ = ~ng6077 & ~new_n14336_;
  assign new_n14340_ = ~new_n14338_ & ~new_n14339_;
  assign new_n14341_ = pg35 & ~new_n14340_;
  assign n5799 = new_n14335_ | new_n14341_;
  assign new_n14343_ = ~pg35 & ng3017;
  assign new_n14344_ = ~new_n8928_ & ~new_n8932_;
  assign new_n14345_ = ng3021 & new_n8954_;
  assign new_n14346_ = new_n14344_ & new_n14345_;
  assign new_n14347_ = ~ng3021 & ~new_n14344_;
  assign new_n14348_ = ~new_n14346_ & ~new_n14347_;
  assign new_n14349_ = pg35 & ~new_n14348_;
  assign n5804 = new_n14343_ | new_n14349_;
  assign new_n14351_ = pg35 & ng5791;
  assign new_n14352_ = ~pg35 & new_n14351_;
  assign new_n14353_ = ~ng5857 & new_n11839_;
  assign new_n14354_ = pg35 & new_n14353_;
  assign n5809 = new_n14352_ | new_n14354_;
  assign new_n14356_ = ~pg35 & ng534;
  assign new_n14357_ = ng12 & n4465;
  assign new_n14358_ = new_n4910_ & new_n14357_;
  assign new_n14359_ = ng79 & ~ng550;
  assign new_n14360_ = ~new_n14358_ & ~new_n14359_;
  assign new_n14361_ = pg35 & new_n14360_;
  assign n5819 = new_n14356_ | new_n14361_;
  assign new_n14363_ = ~pg35 & ng278;
  assign new_n14364_ = ~ng283 & new_n6021_;
  assign new_n14365_ = pg35 & new_n14364_;
  assign n5824 = new_n14363_ | new_n14365_;
  assign new_n14367_ = ~pg35 & ng2791;
  assign new_n14368_ = ~ng2036 & new_n7642_;
  assign new_n14369_ = ~ng2795 & ~new_n14368_;
  assign new_n14370_ = ~new_n7640_ & ~new_n14369_;
  assign new_n14371_ = pg35 & new_n14370_;
  assign n5829 = new_n14367_ | new_n14371_;
  assign new_n14373_ = ~pg35 & ng222;
  assign new_n14374_ = new_n11552_ & new_n11557_;
  assign new_n14375_ = ng194 & ~new_n14374_;
  assign new_n14376_ = ~ng194 & new_n14374_;
  assign new_n14377_ = ~new_n14375_ & ~new_n14376_;
  assign new_n14378_ = pg35 & ~new_n14377_;
  assign n5834 = new_n14373_ | new_n14378_;
  assign new_n14380_ = ~pg35 & ng6044;
  assign new_n14381_ = ~ng6049 & ~new_n12615_;
  assign new_n14382_ = new_n6353_ & new_n14381_;
  assign new_n14383_ = ng6049 & ~new_n6353_;
  assign new_n14384_ = ~new_n14382_ & ~new_n14383_;
  assign new_n14385_ = pg35 & ~new_n14384_;
  assign n5838 = new_n14380_ | new_n14385_;
  assign new_n14387_ = ~pg35 & ng4141;
  assign new_n14388_ = ~ng4082 & new_n7185_;
  assign new_n14389_ = ng4082 & ~new_n7185_;
  assign new_n14390_ = ~new_n14388_ & ~new_n14389_;
  assign new_n14391_ = ng4169 & ~new_n14390_;
  assign new_n14392_ = ng4169 & ~new_n14391_;
  assign new_n14393_ = pg35 & ~new_n14392_;
  assign n5843 = new_n14387_ | new_n14393_;
  assign new_n14395_ = ~pg35 & ng1280;
  assign new_n14396_ = ~ng1252 & new_n8888_;
  assign new_n14397_ = ng1570 & ng1252;
  assign new_n14398_ = ~new_n8888_ & new_n14397_;
  assign new_n14399_ = ~new_n14396_ & ~new_n14398_;
  assign new_n14400_ = pg35 & ~new_n14399_;
  assign n5848 = new_n14395_ | new_n14400_;
  assign new_n14402_ = ~pg35 & ng5523;
  assign new_n14403_ = ng5527 & ~new_n8302_;
  assign new_n14404_ = ~ng5523 & new_n14403_;
  assign new_n14405_ = ~ng5527 & ~new_n8302_;
  assign new_n14406_ = ng5523 & new_n14405_;
  assign new_n14407_ = ~new_n14404_ & ~new_n14406_;
  assign new_n14408_ = pg35 & ~new_n14407_;
  assign n5853 = new_n14402_ | new_n14408_;
  assign new_n14410_ = ~pg35 & ng5196;
  assign new_n14411_ = new_n8407_ & new_n11577_;
  assign new_n14412_ = ng5224 & ~new_n14411_;
  assign new_n14413_ = ~new_n5966_ & new_n14411_;
  assign new_n14414_ = ~new_n14412_ & ~new_n14413_;
  assign new_n14415_ = pg35 & ~new_n14414_;
  assign n5858 = new_n14410_ | new_n14415_;
  assign new_n14417_ = ~pg35 & ng1283;
  assign new_n14418_ = n2272 & new_n8829_;
  assign new_n14419_ = ~ng1287 & new_n4689_;
  assign new_n14420_ = ~new_n14418_ & ~new_n14419_;
  assign new_n14421_ = pg35 & new_n14420_;
  assign n5863 = new_n14417_ | new_n14421_;
  assign new_n14423_ = ~pg35 & ng1592;
  assign new_n14424_ = ~pg113 & new_n5639_;
  assign new_n14425_ = ~new_n4724_ & new_n14424_;
  assign new_n14426_ = pg33533 & new_n14425_;
  assign new_n14427_ = ng112 & pg25259;
  assign new_n14428_ = ng112 & ~new_n14427_;
  assign new_n14429_ = pg25259 & ~new_n14427_;
  assign new_n14430_ = ~new_n14428_ & ~new_n14429_;
  assign new_n14431_ = new_n14426_ & ~new_n14430_;
  assign new_n14432_ = ng1644 & ~new_n14426_;
  assign new_n14433_ = ~new_n14431_ & ~new_n14432_;
  assign new_n14434_ = pg35 & ~new_n14433_;
  assign n5868 = new_n14423_ | new_n14434_;
  assign new_n14436_ = ~pg35 & ng5170;
  assign new_n14437_ = ~ng5176 & ~new_n7369_1_;
  assign new_n14438_ = new_n11431_ & new_n14437_;
  assign new_n14439_ = ng5176 & new_n14437_;
  assign new_n14440_ = ~new_n11431_ & new_n14439_;
  assign new_n14441_ = ~new_n14438_ & ~new_n14440_;
  assign new_n14442_ = pg35 & ~new_n14441_;
  assign n5873 = new_n14436_ | new_n14442_;
  assign new_n14444_ = ~pg35 & ng1532;
  assign new_n14445_ = ng1413 & new_n13759_;
  assign new_n14446_ = ng1536 & ~new_n14445_;
  assign new_n14447_ = ~new_n6840_ & ~new_n14446_;
  assign new_n14448_ = pg35 & ~new_n14447_;
  assign n5878 = new_n14444_ | new_n14448_;
  assign new_n14450_ = ~pg35 & ng5200;
  assign new_n14451_ = new_n7580_1_ & new_n11577_;
  assign new_n14452_ = ng5228 & ~new_n14451_;
  assign new_n14453_ = ~new_n5966_ & new_n14451_;
  assign new_n14454_ = ~new_n14452_ & ~new_n14453_;
  assign new_n14455_ = pg35 & ~new_n14454_;
  assign n5883 = new_n14450_ | new_n14455_;
  assign new_n14457_ = pg35 & ng4035;
  assign new_n14458_ = ~pg35 & new_n14457_;
  assign new_n14459_ = ng3849 & ~new_n7011_1_;
  assign new_n14460_ = ~new_n5966_ & new_n14459_;
  assign new_n14461_ = new_n14459_ & ~new_n14460_;
  assign new_n14462_ = ~new_n5966_ & ~new_n14460_;
  assign new_n14463_ = ~new_n14461_ & ~new_n14462_;
  assign new_n14464_ = pg35 & ~new_n14463_;
  assign n5888 = new_n14458_ | new_n14464_;
  assign new_n14466_ = ~pg35 & ng2295;
  assign new_n14467_ = ~ng2361 & ng2331;
  assign new_n14468_ = ~new_n7886_ & new_n14467_;
  assign new_n14469_ = ng2303 & ~new_n14468_;
  assign new_n14470_ = ~new_n8906_ & new_n14468_;
  assign new_n14471_ = ~new_n14469_ & ~new_n14470_;
  assign new_n14472_ = pg35 & ~new_n14471_;
  assign n5893 = new_n14466_ | new_n14472_;
  assign new_n14474_ = ~pg35 & ng3050;
  assign new_n14475_ = pg35 & ng3338;
  assign n5898 = new_n14474_ | new_n14475_;
  assign new_n14477_ = ~pg35 & ng336;
  assign new_n14478_ = ng324 & ~ng311;
  assign new_n14479_ = ~ng305 & ~new_n14478_;
  assign new_n14480_ = pg35 & ~new_n14479_;
  assign n5902 = new_n14477_ | new_n14480_;
  assign new_n14482_ = ~pg35 & ng6523;
  assign new_n14483_ = ng6527 & ~new_n7219_;
  assign new_n14484_ = ~ng6527 & new_n7219_;
  assign new_n14485_ = ~new_n14483_ & ~new_n14484_;
  assign new_n14486_ = pg35 & ~new_n14485_;
  assign n5907 = new_n14482_ | new_n14486_;
  assign new_n14488_ = ~pg35 & ng5703;
  assign new_n14489_ = ng5703 & new_n7745_;
  assign new_n14490_ = ng5644 & ~new_n7750_;
  assign new_n14491_ = ~new_n14489_ & new_n14490_;
  assign new_n14492_ = ~ng5644 & ~new_n7750_;
  assign new_n14493_ = new_n14489_ & new_n14492_;
  assign new_n14494_ = ~new_n14491_ & ~new_n14493_;
  assign new_n14495_ = pg35 & ~new_n14494_;
  assign n5912 = new_n14488_ | new_n14495_;
  assign n5917 = ~pg35 & ng1287;
  assign new_n14498_ = ~pg35 & ng3937;
  assign new_n14499_ = new_n6894_ & new_n8079_;
  assign new_n14500_ = ng3953 & ~new_n14499_;
  assign new_n14501_ = ~new_n5966_ & new_n14499_;
  assign new_n14502_ = ~new_n14500_ & ~new_n14501_;
  assign new_n14503_ = pg35 & ~new_n14502_;
  assign n5925 = new_n14498_ | new_n14503_;
  assign new_n14505_ = ~pg35 & ng146;
  assign new_n14506_ = ~ng164 & new_n6278_;
  assign new_n14507_ = ng164 & new_n6276_;
  assign new_n14508_ = ~new_n6278_ & new_n14507_;
  assign new_n14509_ = ~new_n14506_ & ~new_n14508_;
  assign new_n14510_ = pg35 & ~new_n14509_;
  assign n5930 = new_n14505_ | new_n14510_;
  assign new_n14512_ = ~pg35 & ng1624;
  assign new_n14513_ = ~ng1624 & ~new_n11200_;
  assign new_n14514_ = new_n7230_ & ~new_n14513_;
  assign new_n14515_ = ng1648 & ~new_n7230_;
  assign new_n14516_ = ~new_n14514_ & ~new_n14515_;
  assign new_n14517_ = pg35 & ~new_n14516_;
  assign n5935 = new_n14512_ | new_n14517_;
  assign n5940 = ~pg35 & ng1311;
  assign new_n14520_ = ~pg35 & ng6279;
  assign new_n14521_ = new_n5849_ & new_n9572_;
  assign new_n14522_ = ng6295 & ~new_n14521_;
  assign new_n14523_ = ~new_n5966_ & new_n14521_;
  assign new_n14524_ = ~new_n14522_ & ~new_n14523_;
  assign new_n14525_ = pg35 & ~new_n14524_;
  assign n5945 = new_n14520_ | new_n14525_;
  assign new_n14527_ = ~pg35 & ng1798;
  assign new_n14528_ = ~ng1783 & ~new_n6732_;
  assign new_n14529_ = new_n6683_ & ~new_n14528_;
  assign new_n14530_ = ng1792 & ~new_n6683_;
  assign new_n14531_ = ~new_n14529_ & ~new_n14530_;
  assign new_n14532_ = pg35 & ~new_n14531_;
  assign n5950 = new_n14527_ | new_n14532_;
  assign new_n14534_ = ~pg35 & ng2571;
  assign new_n14535_ = ~new_n7174_ & new_n10430_;
  assign new_n14536_ = ng2583 & ~new_n14535_;
  assign new_n14537_ = ~new_n8484_ & new_n14535_;
  assign new_n14538_ = ~new_n14536_ & ~new_n14537_;
  assign new_n14539_ = pg35 & ~new_n14538_;
  assign n5955 = new_n14534_ | new_n14539_;
  assign new_n14541_ = ~pg35 & ng3412;
  assign new_n14542_ = ng3412 & ng3408;
  assign new_n14543_ = pg35 & new_n14542_;
  assign n5960 = new_n14541_ | new_n14543_;
  assign new_n14545_ = ~pg35 & ng3401;
  assign new_n14546_ = pg35 & ng3689;
  assign n5965 = new_n14545_ | new_n14546_;
  assign new_n14548_ = ~pg35 & ng6459;
  assign new_n14549_ = ~ng6451 & ng6459;
  assign new_n14550_ = ng6466 & new_n14549_;
  assign new_n14551_ = ~ng6455 & ng6459;
  assign new_n14552_ = ~ng6466 & new_n14551_;
  assign new_n14553_ = ~new_n14550_ & ~new_n14552_;
  assign new_n14554_ = pg35 & ~new_n14553_;
  assign n5969 = new_n14548_ | new_n14554_;
  assign new_n14556_ = pg35 & ng199;
  assign new_n14557_ = ~pg35 & new_n14556_;
  assign new_n14558_ = ~ng278 & ~new_n6017_;
  assign new_n14559_ = ~new_n6010_ & ~new_n14558_;
  assign new_n14560_ = pg35 & new_n14559_;
  assign n5974 = new_n14557_ | new_n14560_;
  assign new_n14562_ = ~pg35 & ng6390;
  assign new_n14563_ = ~ng6395 & ~new_n14024_;
  assign new_n14564_ = new_n6699_ & new_n14563_;
  assign new_n14565_ = ng6395 & ~new_n6699_;
  assign new_n14566_ = ~new_n14564_ & ~new_n14565_;
  assign new_n14567_ = pg35 & ~new_n14566_;
  assign n5979 = new_n14562_ | new_n14567_;
  assign new_n14569_ = ~pg35 & ng758;
  assign new_n14570_ = ng763 & ~new_n6578_;
  assign new_n14571_ = ~new_n6586_1_ & new_n14570_;
  assign new_n14572_ = ~ng763 & new_n6586_1_;
  assign new_n14573_ = ~new_n14571_ & ~new_n14572_;
  assign new_n14574_ = pg35 & ~new_n14573_;
  assign n5988 = new_n14569_ | new_n14574_;
  assign new_n14576_ = ~pg35 & ng1612;
  assign new_n14577_ = pg25167 & new_n7230_;
  assign new_n14578_ = ng1632 & ~new_n14577_;
  assign new_n14579_ = ~new_n13816_ & new_n14577_;
  assign new_n14580_ = ~new_n14578_ & ~new_n14579_;
  assign new_n14581_ = pg35 & ~new_n14580_;
  assign n5993 = new_n14576_ | new_n14581_;
  assign new_n14583_ = ~pg35 & ng739;
  assign new_n14584_ = ~ng744 & new_n6580_;
  assign new_n14585_ = ng744 & ~new_n6578_;
  assign new_n14586_ = ~new_n6580_ & new_n14585_;
  assign new_n14587_ = ~new_n14584_ & ~new_n14586_;
  assign new_n14588_ = pg35 & ~new_n14587_;
  assign n5998 = new_n14583_ | new_n14588_;
  assign new_n14590_ = ~pg35 & ng1495;
  assign new_n14591_ = ng1442 & ~new_n6433_;
  assign new_n14592_ = ng1495 & new_n6433_;
  assign new_n14593_ = ~new_n14591_ & ~new_n14592_;
  assign new_n14594_ = pg35 & ~new_n14593_;
  assign n6003 = new_n14590_ | new_n14594_;
  assign new_n14596_ = ~pg35 & ng1478;
  assign new_n14597_ = ng1454 & ~new_n8067_;
  assign new_n14598_ = ng1448 & new_n6436_;
  assign new_n14599_ = ng1448 & ~new_n14598_;
  assign new_n14600_ = new_n6436_ & ~new_n14598_;
  assign new_n14601_ = ~new_n14599_ & ~new_n14600_;
  assign new_n14602_ = ng1454 & ~new_n14601_;
  assign new_n14603_ = ~new_n6435_1_ & new_n14602_;
  assign new_n14604_ = new_n6435_1_ & ~new_n14601_;
  assign new_n14605_ = ~new_n14603_ & ~new_n14604_;
  assign new_n14606_ = new_n8067_ & ~new_n14605_;
  assign new_n14607_ = ~new_n14597_ & ~new_n14606_;
  assign new_n14608_ = pg35 & ~new_n14607_;
  assign n6008 = new_n14596_ | new_n14608_;
  assign new_n14610_ = pg35 & ng2283;
  assign new_n14611_ = ~pg35 & new_n14610_;
  assign new_n14612_ = ~ng2361 & ng2287;
  assign new_n14613_ = ~ng2361 & ~ng2331;
  assign new_n14614_ = ~new_n14612_ & ~new_n14613_;
  assign new_n14615_ = ~new_n11285_ & ~new_n14614_;
  assign new_n14616_ = ~new_n7886_ & new_n14615_;
  assign new_n14617_ = ng2287 & new_n7886_;
  assign new_n14618_ = ~new_n14616_ & ~new_n14617_;
  assign new_n14619_ = pg35 & ~new_n14618_;
  assign n6013 = new_n14611_ | new_n14619_;
  assign new_n14621_ = ~pg35 & ng3538;
  assign new_n14622_ = new_n10353_ & new_n11130_;
  assign new_n14623_ = ng3566 & ~new_n14622_;
  assign new_n14624_ = ~new_n5966_ & new_n14622_;
  assign new_n14625_ = ~new_n14623_ & ~new_n14624_;
  assign new_n14626_ = pg35 & ~new_n14625_;
  assign n6018 = new_n14621_ | new_n14626_;
  assign new_n14628_ = ~pg35 & ng645;
  assign new_n14629_ = ng681 & ~new_n7858_;
  assign new_n14630_ = ng645 & new_n7858_;
  assign new_n14631_ = ~new_n14629_ & ~new_n14630_;
  assign new_n14632_ = pg35 & ~new_n14631_;
  assign n6023 = new_n14628_ | new_n14632_;
  assign new_n14634_ = ~pg35 & ng3512;
  assign new_n14635_ = new_n7697_ & new_n10820_;
  assign new_n14636_ = ng3518 & new_n10820_;
  assign new_n14637_ = ~new_n7697_ & new_n14636_;
  assign new_n14638_ = ~new_n14635_ & ~new_n14637_;
  assign new_n14639_ = pg35 & ~new_n14638_;
  assign n6028 = new_n14634_ | new_n14639_;
  assign new_n14641_ = ~pg35 & ng3831;
  assign new_n14642_ = ng3835 & ~new_n6468_;
  assign new_n14643_ = ~ng3835 & new_n6468_;
  assign new_n14644_ = ~new_n14642_ & ~new_n14643_;
  assign new_n14645_ = pg35 & ~new_n14644_;
  assign n6041 = new_n14641_ | new_n14645_;
  assign new_n14647_ = ~pg35 & ng182;
  assign new_n14648_ = ng174 & ~new_n5994_;
  assign new_n14649_ = ng182 & new_n5994_;
  assign new_n14650_ = ~new_n14648_ & ~new_n14649_;
  assign new_n14651_ = pg35 & ~new_n14650_;
  assign n6050 = new_n14647_ | new_n14651_;
  assign new_n14653_ = ~pg35 & ng5736;
  assign new_n14654_ = ~new_n10152_ & ~new_n10155_;
  assign new_n14655_ = ng5742 & new_n6424_;
  assign new_n14656_ = new_n14654_ & new_n14655_;
  assign new_n14657_ = ~ng5742 & ~new_n14654_;
  assign new_n14658_ = ~new_n14656_ & ~new_n14657_;
  assign new_n14659_ = pg35 & ~new_n14658_;
  assign n6055 = new_n14653_ | new_n14659_;
  assign new_n14661_ = ~pg35 & ng2787;
  assign new_n14662_ = ng2783 & ~new_n6043_;
  assign new_n14663_ = ng2791 & ~new_n5870_;
  assign new_n14664_ = ~new_n8665_ & ~new_n14663_;
  assign new_n14665_ = new_n6043_ & new_n14664_;
  assign new_n14666_ = ~new_n14662_ & ~new_n14665_;
  assign new_n14667_ = pg35 & ~new_n14666_;
  assign n6060 = new_n14661_ | new_n14667_;
  assign new_n14669_ = ~pg35 & ng6295;
  assign new_n14670_ = ng6215 & new_n9572_;
  assign new_n14671_ = ng6243 & ~new_n14670_;
  assign new_n14672_ = ~new_n5966_ & new_n14670_;
  assign new_n14673_ = ~new_n14671_ & ~new_n14672_;
  assign new_n14674_ = pg35 & ~new_n14673_;
  assign n6069 = new_n14669_ | new_n14674_;
  assign new_n14676_ = ~pg35 & ng6120;
  assign new_n14677_ = ng6120 & ~ng6128;
  assign new_n14678_ = ~ng6120 & ng6128;
  assign new_n14679_ = ~new_n14677_ & ~new_n14678_;
  assign new_n14680_ = pg35 & ~new_n14679_;
  assign n6074 = new_n14676_ | new_n14680_;
  assign new_n14682_ = ~pg35 & ng262;
  assign new_n14683_ = ng881 & new_n6112_;
  assign new_n14684_ = ng239 & ~new_n6112_;
  assign new_n14685_ = ~new_n14683_ & ~new_n14684_;
  assign new_n14686_ = pg35 & ~new_n14685_;
  assign n6084 = new_n14682_ | new_n14686_;
  assign n6096 = ~pg35 & ng2151;
  assign new_n14689_ = pg35 & ng86;
  assign new_n14690_ = ~pg35 & new_n14689_;
  assign new_n14691_ = ~ng5164 & new_n14437_;
  assign new_n14692_ = pg35 & new_n14691_;
  assign n6101 = new_n14690_ | new_n14692_;
  assign new_n14694_ = ~pg35 & ng2441;
  assign new_n14695_ = new_n5215_ & new_n5907_1_;
  assign new_n14696_ = ng2461 & ~new_n14695_;
  assign new_n14697_ = ~new_n9238_ & new_n14695_;
  assign new_n14698_ = ~new_n14696_ & ~new_n14697_;
  assign new_n14699_ = pg35 & ~new_n14698_;
  assign n6109 = new_n14694_ | new_n14699_;
  assign new_n14701_ = ~pg35 & ng4459;
  assign new_n14702_ = pg35 & ng4473;
  assign n6114 = new_n14701_ | new_n14702_;
  assign new_n14704_ = ~pg35 & ng3352;
  assign new_n14705_ = ng3352 & new_n6915_;
  assign new_n14706_ = ng3288 & ~new_n12100_;
  assign new_n14707_ = ~new_n14705_ & new_n14706_;
  assign new_n14708_ = ~ng3288 & ~new_n12100_;
  assign new_n14709_ = new_n14705_ & new_n14708_;
  assign new_n14710_ = ~new_n14707_ & ~new_n14709_;
  assign new_n14711_ = pg35 & ~new_n14710_;
  assign n6119 = new_n14704_ | new_n14711_;
  assign new_n14713_ = ~pg35 & ng1259;
  assign new_n14714_ = ng1570 & ng1263;
  assign new_n14715_ = ~new_n9070_ & new_n14714_;
  assign new_n14716_ = ~ng1263 & new_n9070_;
  assign new_n14717_ = ~new_n14715_ & ~new_n14716_;
  assign new_n14718_ = pg35 & ~new_n14717_;
  assign n6124 = new_n14713_ | new_n14718_;
  assign new_n14720_ = ~pg35 & ng4659;
  assign new_n14721_ = ~ng4664 & new_n10528_;
  assign new_n14722_ = new_n14291_ & new_n14721_;
  assign new_n14723_ = ng4664 & new_n10528_;
  assign new_n14724_ = ~new_n14291_ & new_n14723_;
  assign new_n14725_ = ~new_n14722_ & ~new_n14724_;
  assign new_n14726_ = pg35 & ~new_n14725_;
  assign n6129 = new_n14720_ | new_n14726_;
  assign new_n14728_ = ~pg35 & ng1996;
  assign new_n14729_ = ~pg113 & new_n5646_;
  assign new_n14730_ = ~new_n4724_ & new_n14729_;
  assign new_n14731_ = new_n7024_ & new_n14730_;
  assign new_n14732_ = ng2070 & ~ng2040;
  assign new_n14733_ = ng112 & new_n14732_;
  assign new_n14734_ = ng112 & ~new_n14733_;
  assign new_n14735_ = new_n14732_ & ~new_n14733_;
  assign new_n14736_ = ~new_n14734_ & ~new_n14735_;
  assign new_n14737_ = new_n14731_ & ~new_n14736_;
  assign new_n14738_ = ng2047 & ~new_n14731_;
  assign new_n14739_ = ~new_n14737_ & ~new_n14738_;
  assign new_n14740_ = pg35 & ~new_n14739_;
  assign n6134 = new_n14728_ | new_n14740_;
  assign new_n14742_ = ~pg35 & ng4434;
  assign new_n14743_ = ng4434 & new_n8046_;
  assign new_n14744_ = ng4392 & new_n14743_;
  assign new_n14745_ = ~ng4443 & ~new_n14744_;
  assign new_n14746_ = pg35 & ~new_n14745_;
  assign n6139 = new_n14742_ | new_n14746_;
  assign new_n14748_ = ~pg35 & ng568;
  assign new_n14749_ = ~ng572 & new_n6549_;
  assign new_n14750_ = ng572 & ~new_n6545_;
  assign new_n14751_ = ~new_n6549_ & new_n14750_;
  assign new_n14752_ = ~new_n14749_ & ~new_n14751_;
  assign new_n14753_ = pg35 & ~new_n14752_;
  assign n6144 = new_n14748_ | new_n14753_;
  assign new_n14755_ = ~pg35 & ng4054;
  assign new_n14756_ = ng4054 & new_n6467_;
  assign new_n14757_ = ng3990 & ~new_n13106_;
  assign new_n14758_ = ~new_n14756_ & new_n14757_;
  assign new_n14759_ = ~ng3990 & ~new_n13106_;
  assign new_n14760_ = new_n14756_ & new_n14759_;
  assign new_n14761_ = ~new_n14758_ & ~new_n14760_;
  assign new_n14762_ = pg35 & ~new_n14761_;
  assign n6149 = new_n14755_ | new_n14762_;
  assign new_n14764_ = ~pg35 & ng843;
  assign new_n14765_ = ng843 & new_n10810_;
  assign new_n14766_ = ng837 & ng812;
  assign new_n14767_ = ~new_n14765_ & new_n14766_;
  assign new_n14768_ = ng837 & ~ng812;
  assign new_n14769_ = new_n14765_ & new_n14768_;
  assign new_n14770_ = ~new_n14767_ & ~new_n14769_;
  assign new_n14771_ = pg35 & ~new_n14770_;
  assign n6154 = new_n14764_ | new_n14771_;
  assign new_n14773_ = ~pg35 & ng3614;
  assign new_n14774_ = ~ng3703 & ~ng3639;
  assign new_n14775_ = ~ng3689 & new_n14774_;
  assign new_n14776_ = ng3672 & ng3590;
  assign new_n14777_ = new_n14775_ & new_n14776_;
  assign new_n14778_ = ~ng3703 & ng3639;
  assign new_n14779_ = ~ng3689 & new_n14778_;
  assign new_n14780_ = ng3562 & ng3680;
  assign new_n14781_ = new_n14779_ & new_n14780_;
  assign new_n14782_ = ng3703 & ~ng3639;
  assign new_n14783_ = ~ng3689 & new_n14782_;
  assign new_n14784_ = ng3676 & ng3606;
  assign new_n14785_ = new_n14783_ & new_n14784_;
  assign new_n14786_ = ~ng3689 & new_n4762_1_;
  assign new_n14787_ = ng3654 & ng3558;
  assign new_n14788_ = new_n14786_ & new_n14787_;
  assign new_n14789_ = ~new_n14777_ & ~new_n14781_;
  assign new_n14790_ = ~new_n14785_ & ~new_n14788_;
  assign new_n14791_ = new_n14789_ & new_n14790_;
  assign new_n14792_ = ng3689 & new_n14774_;
  assign new_n14793_ = ng3546 & ng3680;
  assign new_n14794_ = new_n14792_ & new_n14793_;
  assign new_n14795_ = ng3689 & ng3654;
  assign new_n14796_ = ng3654 & ~new_n14795_;
  assign new_n14797_ = ng3689 & ~new_n14795_;
  assign new_n14798_ = ~new_n14796_ & ~new_n14797_;
  assign new_n14799_ = new_n14778_ & new_n14798_;
  assign new_n14800_ = ng3632 & ng3570;
  assign new_n14801_ = new_n14799_ & new_n14800_;
  assign new_n14802_ = ng3689 & new_n14782_;
  assign new_n14803_ = ng3654 & ng3542;
  assign new_n14804_ = new_n14802_ & new_n14803_;
  assign new_n14805_ = new_n4762_1_ & new_n14798_;
  assign new_n14806_ = ng3586 & ng3661;
  assign new_n14807_ = new_n14805_ & new_n14806_;
  assign new_n14808_ = ~new_n14794_ & ~new_n14801_;
  assign new_n14809_ = ~new_n14804_ & ~new_n14807_;
  assign new_n14810_ = new_n14808_ & new_n14809_;
  assign new_n14811_ = ng3538 & ng3649;
  assign new_n14812_ = new_n14792_ & new_n14811_;
  assign new_n14813_ = ng3689 & new_n14778_;
  assign new_n14814_ = ng3672 & ng3582;
  assign new_n14815_ = new_n14813_ & new_n14814_;
  assign new_n14816_ = ng3668 & ng3566;
  assign new_n14817_ = new_n14802_ & new_n14816_;
  assign new_n14818_ = ng3689 & new_n4762_1_;
  assign new_n14819_ = ng3676 & ng3598;
  assign new_n14820_ = new_n14818_ & new_n14819_;
  assign new_n14821_ = ~new_n14812_ & ~new_n14815_;
  assign new_n14822_ = ~new_n14817_ & ~new_n14820_;
  assign new_n14823_ = new_n14821_ & new_n14822_;
  assign new_n14824_ = new_n14774_ & new_n14798_;
  assign new_n14825_ = ng3618 & ng3602;
  assign new_n14826_ = new_n14824_ & new_n14825_;
  assign new_n14827_ = ng3550 & ng3649;
  assign new_n14828_ = new_n14779_ & new_n14827_;
  assign new_n14829_ = ng3625 & ng3554;
  assign new_n14830_ = new_n14783_ & new_n14829_;
  assign new_n14831_ = ng3668 & ng3574;
  assign new_n14832_ = new_n14786_ & new_n14831_;
  assign new_n14833_ = ~new_n14826_ & ~new_n14828_;
  assign new_n14834_ = ~new_n14830_ & ~new_n14832_;
  assign new_n14835_ = new_n14833_ & new_n14834_;
  assign new_n14836_ = new_n14810_ & new_n14823_;
  assign new_n14837_ = new_n14835_ & new_n14836_;
  assign new_n14838_ = new_n14774_ & ~new_n14798_;
  assign new_n14839_ = ng3632 & ng3578;
  assign new_n14840_ = new_n14838_ & new_n14839_;
  assign new_n14841_ = new_n14778_ & ~new_n14798_;
  assign new_n14842_ = ng3610 & ng3618;
  assign new_n14843_ = new_n14841_ & new_n14842_;
  assign new_n14844_ = new_n14782_ & ~new_n14798_;
  assign new_n14845_ = ng3661 & ng3594;
  assign new_n14846_ = new_n14844_ & new_n14845_;
  assign new_n14847_ = ng3614 & ng3625;
  assign new_n14848_ = new_n14818_ & new_n14847_;
  assign new_n14849_ = ~new_n14840_ & ~new_n14843_;
  assign new_n14850_ = ~new_n14846_ & ~new_n14848_;
  assign new_n14851_ = new_n14849_ & new_n14850_;
  assign new_n14852_ = new_n14791_ & new_n14837_;
  assign new_n14853_ = new_n14851_ & new_n14852_;
  assign new_n14854_ = new_n7431_ & ~new_n14853_;
  assign new_n14855_ = ng3684 & ~new_n7431_;
  assign new_n14856_ = ~new_n14854_ & ~new_n14855_;
  assign new_n14857_ = pg35 & ~new_n14856_;
  assign n6159 = new_n14773_ | new_n14857_;
  assign new_n14859_ = ~pg35 & ng429;
  assign new_n14860_ = ng401 & ~new_n6067_;
  assign new_n14861_ = ng429 & new_n6067_;
  assign new_n14862_ = ~new_n14860_ & ~new_n14861_;
  assign new_n14863_ = pg35 & ~new_n14862_;
  assign n6164 = new_n14859_ | new_n14863_;
  assign new_n14865_ = ~pg35 & ng572;
  assign new_n14866_ = ng586 & ~new_n6545_;
  assign new_n14867_ = ~new_n6551_ & new_n14866_;
  assign new_n14868_ = ~ng586 & new_n6551_;
  assign new_n14869_ = ~new_n14867_ & ~new_n14868_;
  assign new_n14870_ = pg35 & ~new_n14869_;
  assign n6174 = new_n14865_ | new_n14870_;
  assign new_n14872_ = ~pg35 & ng2389;
  assign new_n14873_ = ng2393 & ~new_n7260_;
  assign new_n14874_ = ~ng2393 & new_n7260_;
  assign new_n14875_ = ~new_n14873_ & ~new_n14874_;
  assign new_n14876_ = pg35 & ~new_n14875_;
  assign n6179 = new_n14872_ | new_n14876_;
  assign new_n14878_ = ~pg35 & ng5424;
  assign new_n14879_ = ~ng5424 & ~new_n12568_;
  assign new_n14880_ = ~ng5428 & new_n14879_;
  assign new_n14881_ = ng5424 & ng5428;
  assign new_n14882_ = ~new_n14880_ & ~new_n14881_;
  assign new_n14883_ = ~new_n12570_ & new_n14882_;
  assign new_n14884_ = pg35 & ~new_n14883_;
  assign n6184 = new_n14878_ | new_n14884_;
  assign new_n14886_ = ~pg35 & ng2595;
  assign new_n14887_ = ~ng2619 & ng2587;
  assign new_n14888_ = ~ng2610 & ~ng2619;
  assign new_n14889_ = ~new_n14887_ & ~new_n14888_;
  assign new_n14890_ = ~new_n10308_ & new_n14889_;
  assign new_n14891_ = new_n10306_ & ~new_n14890_;
  assign new_n14892_ = ng2587 & ~new_n10306_;
  assign new_n14893_ = ~new_n14891_ & ~new_n14892_;
  assign new_n14894_ = pg35 & ~new_n14893_;
  assign n6192 = new_n14886_ | new_n14894_;
  assign new_n14896_ = ~pg35 & ng6247;
  assign new_n14897_ = new_n6761_1_ & new_n7866_;
  assign new_n14898_ = ng6271 & ~new_n14897_;
  assign new_n14899_ = ~new_n5966_ & new_n14897_;
  assign new_n14900_ = ~new_n14898_ & ~new_n14899_;
  assign new_n14901_ = pg35 & ~new_n14900_;
  assign n6197 = new_n14896_ | new_n14901_;
  assign new_n14903_ = ~pg35 & ng2024;
  assign new_n14904_ = ~new_n7025_ & new_n9146_;
  assign new_n14905_ = ng2020 & ~new_n14904_;
  assign new_n14906_ = ~new_n7032_ & new_n14904_;
  assign new_n14907_ = ~new_n14905_ & ~new_n14906_;
  assign new_n14908_ = pg35 & ~new_n14907_;
  assign n6202 = new_n14903_ | new_n14908_;
  assign new_n14910_ = ~pg35 & ng168;
  assign new_n14911_ = ng460 & ~new_n5994_;
  assign new_n14912_ = ng246 & new_n5994_;
  assign new_n14913_ = ~new_n14911_ & ~new_n14912_;
  assign new_n14914_ = pg35 & ~new_n14913_;
  assign n6207 = new_n14910_ | new_n14914_;
  assign new_n14916_ = ~pg35 & ng3231;
  assign new_n14917_ = new_n9338_ & new_n9368_;
  assign new_n14918_ = ng3247 & ~new_n14917_;
  assign new_n14919_ = ~new_n5966_ & new_n14917_;
  assign new_n14920_ = ~new_n14918_ & ~new_n14919_;
  assign new_n14921_ = pg35 & ~new_n14920_;
  assign n6212 = new_n14916_ | new_n14921_;
  assign new_n14923_ = ~pg35 & ng136;
  assign new_n14924_ = new_n4910_ & new_n6820_;
  assign new_n14925_ = ~ng222 & ~ng199;
  assign new_n14926_ = ~new_n14924_ & ~new_n14925_;
  assign new_n14927_ = pg35 & new_n14926_;
  assign n6220 = new_n14923_ | new_n14927_;
  assign new_n14929_ = ~pg35 & ng5077;
  assign new_n14930_ = ng5084 & new_n11084_;
  assign new_n14931_ = ~ng5084 & new_n11088_;
  assign new_n14932_ = ~new_n14930_ & ~new_n14931_;
  assign new_n14933_ = pg35 & ~new_n14932_;
  assign n6225 = new_n14929_ | new_n14933_;
  assign new_n14935_ = ~pg35 & ng2955;
  assign new_n14936_ = new_n4937_ & new_n14357_;
  assign new_n14937_ = pg91 & new_n5037_;
  assign new_n14938_ = ~ng2965 & new_n14937_;
  assign new_n14939_ = ~new_n14936_ & ~new_n14938_;
  assign new_n14940_ = pg35 & new_n14939_;
  assign n6230 = new_n14935_ | new_n14940_;
  assign new_n14942_ = ~pg35 & ng1395;
  assign new_n14943_ = ng1404 & new_n9904_;
  assign new_n14944_ = ~ng1404 & ~new_n9904_;
  assign new_n14945_ = ~new_n14943_ & ~new_n14944_;
  assign new_n14946_ = ~ng1322 & new_n14945_;
  assign new_n14947_ = pg35 & new_n14946_;
  assign n6235 = new_n14942_ | new_n14947_;
  assign new_n14949_ = ~pg35 & ng613;
  assign new_n14950_ = ~ng617 & new_n9120_;
  assign new_n14951_ = ng617 & ~new_n6545_;
  assign new_n14952_ = ~new_n9120_ & new_n14951_;
  assign new_n14953_ = ~new_n14950_ & ~new_n14952_;
  assign new_n14954_ = pg35 & ~new_n14953_;
  assign n6240 = new_n14949_ | new_n14954_;
  assign new_n14956_ = ~pg35 & ng3155;
  assign new_n14957_ = ng3161 & ~new_n6249_;
  assign new_n14958_ = ~ng3155 & new_n14957_;
  assign new_n14959_ = ~ng3161 & ~new_n6249_;
  assign new_n14960_ = ng3155 & new_n14959_;
  assign new_n14961_ = ~new_n14958_ & ~new_n14960_;
  assign new_n14962_ = pg35 & ~new_n14961_;
  assign n6245 = new_n14956_ | new_n14962_;
  assign new_n14964_ = ~pg35 & ng1840;
  assign new_n14965_ = ng1844 & ~new_n8571_;
  assign new_n14966_ = ng1834 & ~ng1840;
  assign new_n14967_ = ng1834 & ~new_n14966_;
  assign new_n14968_ = ~ng1840 & ~new_n14966_;
  assign new_n14969_ = ~new_n14967_ & ~new_n14968_;
  assign new_n14970_ = new_n8571_ & ~new_n14969_;
  assign new_n14971_ = ~new_n14965_ & ~new_n14970_;
  assign new_n14972_ = pg35 & ~new_n14971_;
  assign n6250 = new_n14964_ | new_n14972_;
  assign new_n14974_ = ~pg35 & ng6105;
  assign new_n14975_ = ~new_n7516_ & ~new_n7524_1_;
  assign new_n14976_ = pg35 & new_n14975_;
  assign n6255 = new_n14974_ | new_n14976_;
  assign new_n14978_ = ~pg35 & ng1950;
  assign new_n14979_ = ng1955 & ~new_n11266_;
  assign new_n14980_ = ng1950 & new_n11266_;
  assign new_n14981_ = ~new_n14979_ & ~new_n14980_;
  assign new_n14982_ = pg35 & ~new_n14981_;
  assign n6260 = new_n14978_ | new_n14982_;
  assign new_n14984_ = ~pg35 & ng6415;
  assign new_n14985_ = ~new_n6604_1_ & ~new_n6609_1_;
  assign new_n14986_ = ~ng6419 & ~new_n14985_;
  assign new_n14987_ = ng6419 & new_n6632_1_;
  assign new_n14988_ = new_n14985_ & new_n14987_;
  assign new_n14989_ = ~new_n14986_ & ~new_n14988_;
  assign new_n14990_ = pg35 & ~new_n14989_;
  assign n6265 = new_n14984_ | new_n14990_;
  assign new_n14992_ = ~pg35 & ng667;
  assign new_n14993_ = ~ng671 & new_n9930_;
  assign new_n14994_ = new_n9913_ & new_n14993_;
  assign new_n14995_ = ng671 & new_n9930_;
  assign new_n14996_ = ~new_n9913_ & new_n14995_;
  assign new_n14997_ = ~new_n14994_ & ~new_n14996_;
  assign new_n14998_ = pg35 & ~new_n14997_;
  assign n6270 = new_n14992_ | new_n14998_;
  assign new_n15000_ = ~pg35 & ng1263;
  assign new_n15001_ = ~ng1270 & new_n9071_;
  assign new_n15002_ = ng1570 & ng1270;
  assign new_n15003_ = ~new_n9071_ & new_n15002_;
  assign new_n15004_ = ~new_n15001_ & ~new_n15003_;
  assign new_n15005_ = pg35 & ~new_n15004_;
  assign n6275 = new_n15000_ | new_n15005_;
  assign new_n15007_ = ~pg35 & ng5901;
  assign new_n15008_ = new_n7650_ & new_n9330_;
  assign new_n15009_ = ng5925 & ~new_n15008_;
  assign new_n15010_ = ~new_n5966_ & new_n15008_;
  assign new_n15011_ = ~new_n15009_ & ~new_n15010_;
  assign new_n15012_ = pg35 & ~new_n15011_;
  assign n6280 = new_n15007_ | new_n15012_;
  assign new_n15014_ = ~pg35 & ng2795;
  assign new_n15015_ = ng2787 & ~new_n8789_;
  assign new_n15016_ = ng2795 & ~new_n5870_;
  assign new_n15017_ = ~new_n8665_ & ~new_n15016_;
  assign new_n15018_ = new_n8789_ & new_n15017_;
  assign new_n15019_ = ~new_n15015_ & ~new_n15018_;
  assign new_n15020_ = pg35 & ~new_n15019_;
  assign n6285 = new_n15014_ | new_n15020_;
  assign new_n15022_ = ~pg35 & ng6605;
  assign new_n15023_ = new_n6316_ & new_n6336_;
  assign new_n15024_ = ng6601 & ~new_n15023_;
  assign new_n15025_ = ~new_n5966_ & new_n15023_;
  assign new_n15026_ = ~new_n15024_ & ~new_n15025_;
  assign new_n15027_ = pg35 & ~new_n15026_;
  assign n6290 = new_n15022_ | new_n15027_;
  assign new_n15029_ = ~pg35 & ng4116;
  assign new_n15030_ = ng4119 & ~new_n5982_;
  assign new_n15031_ = ng4145 & new_n5982_;
  assign new_n15032_ = ~new_n15030_ & ~new_n15031_;
  assign new_n15033_ = pg35 & ~new_n15032_;
  assign n6295 = new_n15029_ | new_n15033_;
  assign new_n15035_ = ~pg35 & ng5841;
  assign new_n15036_ = ng5845 & ~new_n10071_;
  assign new_n15037_ = ng5835 & ~ng5841;
  assign new_n15038_ = ng5835 & ~new_n15037_;
  assign new_n15039_ = ~ng5841 & ~new_n15037_;
  assign new_n15040_ = ~new_n15038_ & ~new_n15039_;
  assign new_n15041_ = new_n10071_ & ~new_n15040_;
  assign new_n15042_ = ~new_n15036_ & ~new_n15041_;
  assign new_n15043_ = pg35 & ~new_n15042_;
  assign n6300 = new_n15035_ | new_n15043_;
  assign new_n15045_ = ~pg35 & ng3554;
  assign new_n15046_ = new_n10352_ & new_n12309_;
  assign new_n15047_ = ng3550 & ~new_n15046_;
  assign new_n15048_ = ~new_n5966_ & new_n15046_;
  assign new_n15049_ = ~new_n15047_ & ~new_n15048_;
  assign new_n15050_ = pg35 & ~new_n15049_;
  assign n6308 = new_n15045_ | new_n15050_;
  assign new_n15052_ = ~pg35 & ng1682;
  assign new_n15053_ = ng1687 & ~new_n10846_;
  assign new_n15054_ = ng1682 & new_n10846_;
  assign new_n15055_ = ~new_n15053_ & ~new_n15054_;
  assign new_n15056_ = pg35 & ~new_n15055_;
  assign n6313 = new_n15052_ | new_n15056_;
  assign new_n15058_ = ~pg35 & ng1706;
  assign new_n15059_ = ng1710 & ~new_n10846_;
  assign new_n15060_ = ng1700 & ~ng1706;
  assign new_n15061_ = ng1700 & ~new_n15060_;
  assign new_n15062_ = ~ng1706 & ~new_n15060_;
  assign new_n15063_ = ~new_n15061_ & ~new_n15062_;
  assign new_n15064_ = new_n10846_ & ~new_n15063_;
  assign new_n15065_ = ~new_n15059_ & ~new_n15064_;
  assign new_n15066_ = pg35 & ~new_n15065_;
  assign n6318 = new_n15058_ | new_n15066_;
  assign new_n15068_ = ~pg35 & ng5148;
  assign new_n15069_ = ng5152 & ~pg26801;
  assign new_n15070_ = ng5142 & ~ng5148;
  assign new_n15071_ = ng5142 & ~new_n15070_;
  assign new_n15072_ = ~ng5148 & ~new_n15070_;
  assign new_n15073_ = ~new_n15071_ & ~new_n15072_;
  assign new_n15074_ = pg26801 & ~new_n15073_;
  assign new_n15075_ = ~new_n15069_ & ~new_n15074_;
  assign new_n15076_ = pg35 & ~new_n15075_;
  assign n6323 = new_n15068_ | new_n15076_;
  assign new_n15078_ = ~pg35 & ng2066;
  assign new_n15079_ = ~ng2051 & ~new_n13378_;
  assign new_n15080_ = new_n9143_ & ~new_n15079_;
  assign new_n15081_ = ng2060 & ~new_n9143_;
  assign new_n15082_ = ~new_n15080_ & ~new_n15081_;
  assign new_n15083_ = pg35 & ~new_n15082_;
  assign n6328 = new_n15078_ | new_n15083_;
  assign new_n15085_ = ~pg35 & ng3723;
  assign new_n15086_ = ~new_n6076_ & ~new_n6081_;
  assign new_n15087_ = ~ng3727 & ~new_n15086_;
  assign new_n15088_ = ng3727 & new_n6104_;
  assign new_n15089_ = new_n15086_ & new_n15088_;
  assign new_n15090_ = ~new_n15087_ & ~new_n15089_;
  assign new_n15091_ = pg35 & ~new_n15090_;
  assign n6333 = new_n15085_ | new_n15091_;
  assign new_n15093_ = ~pg35 & ng5041;
  assign new_n15094_ = ~new_n8140_ & ~new_n8145_;
  assign new_n15095_ = ~ng5046 & ~new_n15094_;
  assign new_n15096_ = ng5046 & new_n8107_;
  assign new_n15097_ = new_n15094_ & new_n15096_;
  assign new_n15098_ = ~new_n15095_ & ~new_n15097_;
  assign new_n15099_ = pg35 & ~new_n15098_;
  assign n6338 = new_n15093_ | new_n15099_;
  assign new_n15101_ = ~pg35 & ng4515;
  assign new_n15102_ = pg35 & ~new_n7761_;
  assign n6347 = new_n15101_ | new_n15102_;
  assign new_n15104_ = ~pg35 & ng3610;
  assign new_n15105_ = ng3614 & ~new_n6770_;
  assign new_n15106_ = ~new_n5966_ & new_n6770_;
  assign new_n15107_ = ~new_n15105_ & ~new_n15106_;
  assign new_n15108_ = pg35 & ~new_n15107_;
  assign n6352 = new_n15104_ | new_n15108_;
  assign new_n15110_ = ~pg35 & ng5268;
  assign new_n15111_ = ng5272 & ~pg26801;
  assign new_n15112_ = pg26801 & ~new_n5966_;
  assign new_n15113_ = ~new_n15111_ & ~new_n15112_;
  assign new_n15114_ = pg35 & ~new_n15113_;
  assign n6357 = new_n15110_ | new_n15114_;
  assign new_n15116_ = ~pg35 & ng4349;
  assign new_n15117_ = ng4349 & new_n10703_;
  assign new_n15118_ = ng4358 & ~new_n5873_1_;
  assign new_n15119_ = ~new_n15117_ & new_n15118_;
  assign new_n15120_ = ~ng4358 & ~new_n5873_1_;
  assign new_n15121_ = new_n15117_ & new_n15120_;
  assign new_n15122_ = ~new_n15119_ & ~new_n15121_;
  assign new_n15123_ = pg35 & ~new_n15122_;
  assign n6362 = new_n15116_ | new_n15123_;
  assign n6367 = ~pg35 & ng2975;
  assign new_n15126_ = ~pg35 & ng5459;
  assign new_n15127_ = ng5452 & ~ng5459;
  assign new_n15128_ = ~ng5366 & ~new_n15127_;
  assign new_n15129_ = ~ng5448 & ~new_n15128_;
  assign new_n15130_ = pg35 & new_n15129_;
  assign n6372 = new_n15126_ | new_n15130_;
  assign new_n15132_ = ~pg35 & ng5244;
  assign new_n15133_ = new_n7580_1_ & new_n11431_;
  assign new_n15134_ = ng5260 & ~new_n15133_;
  assign new_n15135_ = ~new_n5966_ & new_n15133_;
  assign new_n15136_ = ~new_n15134_ & ~new_n15135_;
  assign new_n15137_ = pg35 & ~new_n15136_;
  assign n6377 = new_n15132_ | new_n15137_;
  assign new_n15139_ = ~pg35 & ng4297;
  assign new_n15140_ = n6079 & new_n7806_;
  assign new_n15141_ = ~ng4300 & ~ng4242;
  assign new_n15142_ = ~new_n15140_ & ~new_n15141_;
  assign new_n15143_ = pg35 & new_n15142_;
  assign n6382 = new_n15139_ | new_n15143_;
  assign new_n15145_ = new_n5688_ & pg33935;
  assign new_n15146_ = ~new_n5688_ & ~new_n5751_;
  assign n6387 = new_n15145_ | new_n15146_;
  assign new_n15148_ = ~pg35 & ng2380;
  assign new_n15149_ = ng2299 & ~new_n7888_;
  assign new_n15150_ = new_n7888_ & ~new_n8906_;
  assign new_n15151_ = ~new_n15149_ & ~new_n15150_;
  assign new_n15152_ = pg35 & ~new_n15151_;
  assign n6392 = new_n15148_ | new_n15152_;
  assign new_n15154_ = ~pg35 & ng4489;
  assign n6397 = new_n12249_ | new_n15154_;
  assign new_n15156_ = ~pg35 & ng6133;
  assign new_n15157_ = ng6120 & ng6128;
  assign new_n15158_ = ng6133 & new_n15157_;
  assign new_n15159_ = ~ng6137 & new_n15158_;
  assign new_n15160_ = ng6137 & ~new_n15158_;
  assign new_n15161_ = ~new_n15159_ & ~new_n15160_;
  assign new_n15162_ = pg35 & ~new_n15161_;
  assign n6402 = new_n15156_ | new_n15162_;
  assign new_n15164_ = pg35 & ng3990;
  assign new_n15165_ = ~pg35 & new_n15164_;
  assign new_n15166_ = pg35 & ng3881;
  assign n6407 = new_n15165_ | new_n15166_;
  assign new_n15168_ = ~pg35 & ng3953;
  assign new_n15169_ = ng3869 & new_n6894_;
  assign new_n15170_ = ng3905 & ~new_n15169_;
  assign new_n15171_ = ~new_n5966_ & new_n15169_;
  assign new_n15172_ = ~new_n15170_ & ~new_n15171_;
  assign new_n15173_ = pg35 & ~new_n15172_;
  assign n6411 = new_n15168_ | new_n15173_;
  assign new_n15175_ = pg35 & ng4765;
  assign new_n15176_ = ~pg35 & new_n15175_;
  assign new_n15177_ = ~ng5283 & ng5308;
  assign new_n15178_ = ng5283 & ~ng5276;
  assign new_n15179_ = ~new_n15177_ & ~new_n15178_;
  assign new_n15180_ = ~new_n12122_ & new_n15179_;
  assign new_n15181_ = ~ng5290 & ng5320;
  assign new_n15182_ = ng5290 & ~ng5313;
  assign new_n15183_ = ~ng5320 & ng5276;
  assign new_n15184_ = new_n15180_ & ~new_n15181_;
  assign new_n15185_ = ~new_n15182_ & new_n15184_;
  assign new_n15186_ = ~new_n15183_ & new_n15185_;
  assign new_n15187_ = pg35 & new_n15186_;
  assign n6416 = new_n15176_ | new_n15187_;
  assign new_n15189_ = ~pg35 & ng1894;
  assign new_n15190_ = ~ng1894 & ~new_n11334_;
  assign new_n15191_ = new_n8171_ & ~new_n15190_;
  assign new_n15192_ = ng1917 & ~new_n8171_;
  assign new_n15193_ = ~new_n15191_ & ~new_n15192_;
  assign new_n15194_ = pg35 & ~new_n15193_;
  assign n6420 = new_n15189_ | new_n15194_;
  assign new_n15196_ = ~pg35 & ng5961;
  assign new_n15197_ = ng5965 & ~new_n10071_;
  assign new_n15198_ = ~new_n5966_ & new_n10071_;
  assign new_n15199_ = ~new_n15197_ & ~new_n15198_;
  assign new_n15200_ = pg35 & ~new_n15199_;
  assign n6425 = new_n15196_ | new_n15200_;
  assign new_n15202_ = ~pg35 & ng5917;
  assign new_n15203_ = new_n7995_ & new_n12340_;
  assign new_n15204_ = ng5933 & ~new_n15203_;
  assign new_n15205_ = ~new_n5966_ & new_n15203_;
  assign new_n15206_ = ~new_n15204_ & ~new_n15205_;
  assign new_n15207_ = pg35 & ~new_n15206_;
  assign n6430 = new_n15202_ | new_n15207_;
  assign new_n15209_ = ~pg35 & ng5595;
  assign new_n15210_ = new_n10861_ & new_n11751_;
  assign new_n15211_ = ng5611 & ~new_n15210_;
  assign new_n15212_ = ~new_n5966_ & new_n15210_;
  assign new_n15213_ = ~new_n15211_ & ~new_n15212_;
  assign new_n15214_ = pg35 & ~new_n15213_;
  assign n6435 = new_n15209_ | new_n15214_;
  assign new_n15216_ = ~pg35 & ng4564;
  assign new_n15217_ = ~new_n5871_ & new_n7816_;
  assign new_n15218_ = ng4561 & ng4555;
  assign new_n15219_ = ng4564 & new_n15218_;
  assign new_n15220_ = ng4558 & new_n15219_;
  assign new_n15221_ = ~ng2988 & ~new_n15220_;
  assign new_n15222_ = new_n5871_ & new_n15221_;
  assign new_n15223_ = ~new_n15217_ & ~new_n15222_;
  assign new_n15224_ = pg35 & new_n15223_;
  assign n6440 = new_n15216_ | new_n15224_;
  assign new_n15226_ = pg35 & ng490;
  assign new_n15227_ = ~pg35 & new_n15226_;
  assign new_n15228_ = ng417 & ~new_n6067_;
  assign new_n15229_ = ng446 & new_n6067_;
  assign new_n15230_ = ~new_n15228_ & ~new_n15229_;
  assign new_n15231_ = pg35 & ~new_n15230_;
  assign n6445 = new_n15227_ | new_n15231_;
  assign new_n15233_ = ~pg35 & ng1687;
  assign new_n15234_ = ng1604 & ~new_n10846_;
  assign new_n15235_ = ~new_n7543_ & new_n10846_;
  assign new_n15236_ = ~new_n15234_ & ~new_n15235_;
  assign new_n15237_ = pg35 & ~new_n15236_;
  assign n6450 = new_n15233_ | new_n15237_;
  assign new_n15239_ = ~pg35 & ng2089;
  assign new_n15240_ = ng2008 & ~new_n8022_;
  assign new_n15241_ = ~new_n7032_ & new_n8022_;
  assign new_n15242_ = ~new_n15240_ & ~new_n15241_;
  assign new_n15243_ = pg35 & ~new_n15242_;
  assign n6455 = new_n15239_ | new_n15243_;
  assign new_n15245_ = ~pg35 & ng2116;
  assign new_n15246_ = ng2122 & ~new_n9160_;
  assign new_n15247_ = ng2116 & new_n9160_;
  assign new_n15248_ = ~new_n15246_ & ~new_n15247_;
  assign new_n15249_ = pg35 & ~new_n15248_;
  assign n6460 = new_n15245_ | new_n15249_;
  assign new_n15251_ = ~pg35 & ng2514;
  assign new_n15252_ = ng2433 & ~new_n9787_;
  assign new_n15253_ = ~new_n8465_ & new_n9787_;
  assign new_n15254_ = ~new_n15252_ & ~new_n15253_;
  assign new_n15255_ = pg35 & ~new_n15254_;
  assign n6465 = new_n15251_ | new_n15255_;
  assign new_n15257_ = ~pg35 & ng4153;
  assign new_n15258_ = pg35 & ~new_n8730_;
  assign n6470 = new_n15257_ | new_n15258_;
  assign new_n15260_ = ~pg35 & ng6621;
  assign new_n15261_ = new_n6316_ & new_n12232_;
  assign new_n15262_ = ng6637 & ~new_n15261_;
  assign new_n15263_ = ~new_n5966_ & new_n15261_;
  assign new_n15264_ = ~new_n15262_ & ~new_n15263_;
  assign new_n15265_ = pg35 & ~new_n15264_;
  assign n6475 = new_n15260_ | new_n15265_;
  assign new_n15267_ = ~pg35 & ng3562;
  assign new_n15268_ = new_n6769_ & new_n12309_;
  assign new_n15269_ = ng3558 & ~new_n15268_;
  assign new_n15270_ = ~new_n5966_ & new_n15268_;
  assign new_n15271_ = ~new_n15269_ & ~new_n15270_;
  assign new_n15272_ = pg35 & ~new_n15271_;
  assign n6480 = new_n15267_ | new_n15272_;
  assign new_n15274_ = ~pg35 & ng153;
  assign new_n15275_ = ng157 & new_n6276_;
  assign new_n15276_ = ~new_n6284_ & new_n15275_;
  assign new_n15277_ = ~ng157 & new_n6284_;
  assign new_n15278_ = ~new_n15276_ & ~new_n15277_;
  assign new_n15279_ = pg35 & ~new_n15278_;
  assign n6485 = new_n15274_ | new_n15279_;
  assign new_n15281_ = ~pg35 & ng5945;
  assign new_n15282_ = new_n8432_ & new_n8646_;
  assign new_n15283_ = ng5961 & ~new_n15282_;
  assign new_n15284_ = ~new_n5966_ & new_n15282_;
  assign new_n15285_ = ~new_n15283_ & ~new_n15284_;
  assign new_n15286_ = pg35 & ~new_n15285_;
  assign n6493 = new_n15281_ | new_n15286_;
  assign new_n15288_ = ~pg35 & ng6613;
  assign new_n15289_ = new_n7456_ & new_n12232_;
  assign new_n15290_ = ng6629 & ~new_n15289_;
  assign new_n15291_ = ~new_n5966_ & new_n15289_;
  assign new_n15292_ = ~new_n15290_ & ~new_n15291_;
  assign new_n15293_ = pg35 & ~new_n15292_;
  assign n6498 = new_n15288_ | new_n15293_;
  assign new_n15295_ = ~pg35 & ng5428;
  assign new_n15296_ = ng5428 & ~ng5436;
  assign new_n15297_ = ~ng5428 & ng5436;
  assign new_n15298_ = ~new_n15296_ & ~new_n15297_;
  assign new_n15299_ = pg35 & ~new_n15298_;
  assign n6503 = new_n15295_ | new_n15299_;
  assign new_n15301_ = ~pg35 & ng1221;
  assign new_n15302_ = ng1216 & ~new_n8364_;
  assign new_n15303_ = ~new_n8560_ & new_n15302_;
  assign new_n15304_ = ~ng1216 & ~new_n8364_;
  assign new_n15305_ = new_n8560_ & new_n15304_;
  assign new_n15306_ = ~new_n15303_ & ~new_n15305_;
  assign new_n15307_ = pg35 & ~new_n15306_;
  assign n6508 = new_n15301_ | new_n15307_;
  assign new_n15309_ = ~pg35 & ng3736;
  assign new_n15310_ = ~new_n12900_ & ~new_n12902_;
  assign new_n15311_ = ng3742 & new_n6104_;
  assign new_n15312_ = new_n15310_ & new_n15311_;
  assign new_n15313_ = ~ng3742 & ~new_n15310_;
  assign new_n15314_ = ~new_n15312_ & ~new_n15313_;
  assign new_n15315_ = pg35 & ~new_n15314_;
  assign n6518 = new_n15309_ | new_n15315_;
  assign new_n15317_ = ~pg35 & ng5212;
  assign new_n15318_ = new_n8995_ & new_n10722_;
  assign new_n15319_ = ng5208 & ~new_n15318_;
  assign new_n15320_ = ~new_n5966_ & new_n15318_;
  assign new_n15321_ = ~new_n15319_ & ~new_n15320_;
  assign new_n15322_ = pg35 & ~new_n15321_;
  assign n6523 = new_n15317_ | new_n15322_;
  assign new_n15324_ = new_n5701_ & pg33636;
  assign new_n15325_ = ~new_n5701_ & ~new_n5845_;
  assign n6532 = new_n15324_ | new_n15325_;
  assign new_n15327_ = ~pg35 & ng5712;
  assign new_n15328_ = ~ng5752 & ~ng5712;
  assign new_n15329_ = ng5706 & new_n15328_;
  assign new_n15330_ = ~ng5706 & new_n6424_;
  assign new_n15331_ = ~new_n15328_ & new_n15330_;
  assign new_n15332_ = ~new_n15329_ & ~new_n15331_;
  assign new_n15333_ = pg35 & ~new_n15332_;
  assign n6537 = new_n15327_ | new_n15333_;
  assign new_n15335_ = ~pg35 & ng1802;
  assign new_n15336_ = ng1816 & ~new_n8570_;
  assign new_n15337_ = ~ng1246 & new_n6232_;
  assign new_n15338_ = ~new_n10677_ & ~new_n15337_;
  assign new_n15339_ = new_n15336_ & ~new_n15338_;
  assign new_n15340_ = new_n15336_ & ~new_n15339_;
  assign new_n15341_ = ~new_n15338_ & ~new_n15339_;
  assign new_n15342_ = ~new_n15340_ & ~new_n15341_;
  assign new_n15343_ = ~new_n6236_ & ~new_n15342_;
  assign new_n15344_ = ng1816 & new_n6236_;
  assign new_n15345_ = ~new_n15343_ & ~new_n15344_;
  assign new_n15346_ = pg35 & ~new_n15345_;
  assign n6542 = new_n15335_ | new_n15346_;
  assign new_n15348_ = ~pg35 & ng2399;
  assign new_n15349_ = ng2403 & ~new_n7888_;
  assign new_n15350_ = ~ng2399 & ng2393;
  assign new_n15351_ = ng2393 & ~new_n15350_;
  assign new_n15352_ = ~ng2399 & ~new_n15350_;
  assign new_n15353_ = ~new_n15351_ & ~new_n15352_;
  assign new_n15354_ = new_n7888_ & ~new_n15353_;
  assign new_n15355_ = ~new_n15349_ & ~new_n15354_;
  assign new_n15356_ = pg35 & ~new_n15355_;
  assign n6547 = new_n15348_ | new_n15356_;
  assign new_n15358_ = ~pg35 & ng947;
  assign new_n15359_ = n4465 & new_n6861_;
  assign new_n15360_ = ng962 & ~ng952;
  assign new_n15361_ = ~new_n15359_ & ~new_n15360_;
  assign new_n15362_ = pg35 & new_n15361_;
  assign n6552 = new_n15358_ | new_n15362_;
  assign new_n15364_ = ~pg35 & ng2208;
  assign new_n15365_ = ~new_n4724_ & new_n11141_;
  assign new_n15366_ = new_n9534_ & new_n15365_;
  assign new_n15367_ = ng2217 & ~ng2208;
  assign new_n15368_ = ng110 & new_n15367_;
  assign new_n15369_ = ng110 & ~new_n15368_;
  assign new_n15370_ = new_n15367_ & ~new_n15368_;
  assign new_n15371_ = ~new_n15369_ & ~new_n15370_;
  assign new_n15372_ = new_n15366_ & ~new_n15371_;
  assign new_n15373_ = ng2223 & ~new_n15366_;
  assign new_n15374_ = ~new_n15372_ & ~new_n15373_;
  assign new_n15375_ = pg35 & ~new_n15374_;
  assign n6557 = new_n15364_ | new_n15375_;
  assign new_n15377_ = ~pg35 & ng5941;
  assign new_n15378_ = new_n8646_ & new_n9330_;
  assign new_n15379_ = ng5957 & ~new_n15378_;
  assign new_n15380_ = ~new_n5966_ & new_n15378_;
  assign new_n15381_ = ~new_n15379_ & ~new_n15380_;
  assign new_n15382_ = pg35 & ~new_n15381_;
  assign n6562 = new_n15377_ | new_n15382_;
  assign new_n15384_ = pg35 & ng2126;
  assign new_n15385_ = ~pg35 & new_n15384_;
  assign new_n15386_ = n4465 & new_n6181_;
  assign new_n15387_ = ng2130 & ~new_n6181_;
  assign new_n15388_ = ~new_n15386_ & ~new_n15387_;
  assign new_n15389_ = pg35 & ~new_n15388_;
  assign n6571 = new_n15385_ | new_n15389_;
  assign new_n15391_ = ~pg35 & ng3712;
  assign new_n15392_ = ~ng3752 & ~ng3712;
  assign new_n15393_ = ng3706 & new_n15392_;
  assign new_n15394_ = ~ng3706 & new_n6104_;
  assign new_n15395_ = ~new_n15392_ & new_n15394_;
  assign new_n15396_ = ~new_n15393_ & ~new_n15395_;
  assign new_n15397_ = pg35 & ~new_n15396_;
  assign n6576 = new_n15391_ | new_n15397_;
  assign new_n15399_ = ~pg35 & ng817;
  assign new_n15400_ = ng832 & new_n8009_;
  assign new_n15401_ = ~new_n8005_ & new_n15400_;
  assign new_n15402_ = ~ng832 & new_n8009_;
  assign new_n15403_ = new_n8005_ & new_n15402_;
  assign new_n15404_ = ~new_n15401_ & ~new_n15403_;
  assign new_n15405_ = pg35 & ~new_n15404_;
  assign n6581 = new_n15399_ | new_n15405_;
  assign new_n15407_ = ~pg35 & ng2811;
  assign new_n15408_ = ~ng2461 & new_n7642_;
  assign new_n15409_ = ~ng2823 & ~new_n15408_;
  assign new_n15410_ = ~new_n7640_ & ~new_n15409_;
  assign new_n15411_ = pg35 & new_n15410_;
  assign n6586 = new_n15407_ | new_n15411_;
  assign new_n15413_ = ~pg35 & ng6035;
  assign new_n15414_ = ~ng6044 & ~new_n6453_;
  assign new_n15415_ = pg35 & new_n15414_;
  assign n6591 = new_n15413_ | new_n15415_;
  assign new_n15417_ = ~pg35 & ng1768;
  assign new_n15418_ = ~ng1792 & ng1760;
  assign new_n15419_ = ~ng1783 & ~ng1792;
  assign new_n15420_ = ~new_n15418_ & ~new_n15419_;
  assign new_n15421_ = ~new_n6732_ & new_n15420_;
  assign new_n15422_ = new_n6683_ & ~new_n15421_;
  assign new_n15423_ = ng1760 & ~new_n6683_;
  assign new_n15424_ = ~new_n15422_ & ~new_n15423_;
  assign new_n15425_ = pg35 & ~new_n15424_;
  assign n6596 = new_n15417_ | new_n15425_;
  assign new_n15427_ = ~pg35 & ng2173;
  assign new_n15428_ = new_n5213_ & new_n9534_;
  assign new_n15429_ = ng2193 & ~new_n15428_;
  assign new_n15430_ = ~new_n7096_ & new_n15428_;
  assign new_n15431_ = ~new_n15429_ & ~new_n15430_;
  assign new_n15432_ = pg35 & ~new_n15431_;
  assign n6604 = new_n15427_ | new_n15432_;
  assign new_n15434_ = ~pg35 & ng1236;
  assign n6609 = new_n14149_ | new_n15434_;
  assign new_n15436_ = ~pg35 & ng4477;
  assign new_n15437_ = pg73 & pg72;
  assign new_n15438_ = ~ng59 & new_n15437_;
  assign new_n15439_ = ng4581 & ~new_n15438_;
  assign new_n15440_ = ~ng4581 & ng4372;
  assign new_n15441_ = ~new_n15439_ & ~new_n15440_;
  assign new_n15442_ = pg35 & ~new_n15441_;
  assign n6619 = new_n15436_ | new_n15442_;
  assign new_n15444_ = ~pg35 & ng3566;
  assign new_n15445_ = new_n7039_ & new_n11130_;
  assign new_n15446_ = ng3582 & ~new_n15445_;
  assign new_n15447_ = ~new_n5966_ & new_n15445_;
  assign new_n15448_ = ~new_n15446_ & ~new_n15447_;
  assign new_n15449_ = pg35 & ~new_n15448_;
  assign n6624 = new_n15444_ | new_n15449_;
  assign new_n15451_ = ~pg35 & ng5503;
  assign new_n15452_ = ng5467 & ~new_n10882_;
  assign new_n15453_ = ng5503 & new_n10882_;
  assign new_n15454_ = ~new_n15452_ & ~new_n15453_;
  assign new_n15455_ = pg35 & ~new_n15454_;
  assign n6632 = new_n15451_ | new_n15455_;
  assign new_n15457_ = ~pg35 & ng4601;
  assign new_n15458_ = ~ng4608 & new_n8853_;
  assign new_n15459_ = new_n12749_ & new_n15458_;
  assign new_n15460_ = ng4608 & new_n8853_;
  assign new_n15461_ = ~new_n12749_ & new_n15460_;
  assign new_n15462_ = ~new_n15459_ & ~new_n15461_;
  assign new_n15463_ = pg35 & ~new_n15462_;
  assign n6637 = new_n15457_ | new_n15463_;
  assign new_n15465_ = ~pg35 & ng1902;
  assign new_n15466_ = ~ng1926 & ng1894;
  assign new_n15467_ = ~ng1926 & ~ng1917;
  assign new_n15468_ = ~new_n15466_ & ~new_n15467_;
  assign new_n15469_ = ~new_n11334_ & new_n15468_;
  assign new_n15470_ = new_n8171_ & ~new_n15469_;
  assign new_n15471_ = ng1894 & ~new_n8171_;
  assign new_n15472_ = ~new_n15470_ & ~new_n15471_;
  assign new_n15473_ = pg35 & ~new_n15472_;
  assign n6642 = new_n15465_ | new_n15473_;
  assign new_n15475_ = ~pg35 & ng6657;
  assign new_n15476_ = new_n7218_1_ & ~new_n9762_;
  assign new_n15477_ = ng5011 & ~new_n7218_1_;
  assign new_n15478_ = ~new_n15476_ & ~new_n15477_;
  assign new_n15479_ = pg35 & ~new_n15478_;
  assign n6647 = new_n15475_ | new_n15479_;
  assign new_n15481_ = ~pg35 & ng5857;
  assign new_n15482_ = ng5863 & ~new_n11838_;
  assign new_n15483_ = ~ng5857 & new_n15482_;
  assign new_n15484_ = ~ng5863 & ~new_n11838_;
  assign new_n15485_ = ng5857 & new_n15484_;
  assign new_n15486_ = ~new_n15483_ & ~new_n15485_;
  assign new_n15487_ = pg35 & ~new_n15486_;
  assign n6652 = new_n15481_ | new_n15487_;
  assign new_n15489_ = ~pg35 & ng6494;
  assign new_n15490_ = ng6486 & ~ng6494;
  assign new_n15491_ = ~ng6444 & ~new_n15490_;
  assign new_n15492_ = ~ng6490 & ~new_n15491_;
  assign new_n15493_ = pg35 & new_n15492_;
  assign n6657 = new_n15489_ | new_n15493_;
  assign new_n15495_ = ~pg35 & ng3719;
  assign new_n15496_ = ~new_n6075_ & ~new_n6080_;
  assign new_n15497_ = ng3723 & new_n6104_;
  assign new_n15498_ = new_n15496_ & new_n15497_;
  assign new_n15499_ = ~ng3723 & ~new_n15496_;
  assign new_n15500_ = ~new_n15498_ & ~new_n15499_;
  assign new_n15501_ = pg35 & ~new_n15500_;
  assign n6662 = new_n15495_ | new_n15501_;
  assign new_n15503_ = ~pg35 & ng5264;
  assign new_n15504_ = ng5176 & new_n10722_;
  assign new_n15505_ = ng5220 & ~new_n15504_;
  assign new_n15506_ = ~new_n5966_ & new_n15504_;
  assign new_n15507_ = ~new_n15505_ & ~new_n15506_;
  assign new_n15508_ = pg35 & ~new_n15507_;
  assign n6667 = new_n15503_ | new_n15508_;
  assign new_n15510_ = ~pg35 & ng2370;
  assign new_n15511_ = ng2384 & ~new_n14179_;
  assign new_n15512_ = ng2370 & new_n15511_;
  assign new_n15513_ = new_n15511_ & ~new_n15512_;
  assign new_n15514_ = ng2370 & ~new_n15512_;
  assign new_n15515_ = ~new_n15513_ & ~new_n15514_;
  assign new_n15516_ = new_n7259_ & ~new_n15515_;
  assign new_n15517_ = ng2384 & ~new_n7259_;
  assign new_n15518_ = ~new_n15516_ & ~new_n15517_;
  assign new_n15519_ = pg35 & ~new_n15518_;
  assign n6672 = new_n15510_ | new_n15519_;
  assign new_n15521_ = ~pg35 & ng4521;
  assign new_n15522_ = ng4521 & ~new_n14008_;
  assign new_n15523_ = ~ng4521 & new_n8691_;
  assign new_n15524_ = ~new_n15522_ & ~new_n15523_;
  assign new_n15525_ = pg35 & ~new_n15524_;
  assign n6677 = new_n15521_ | new_n15525_;
  assign new_n15527_ = pg35 & ng1389;
  assign new_n15528_ = ~pg35 & new_n15527_;
  assign new_n15529_ = ng1489 & ~new_n6433_;
  assign new_n15530_ = ~ng1495 & ng1489;
  assign new_n15531_ = ng1442 & ~new_n15530_;
  assign new_n15532_ = new_n6433_ & ~new_n15531_;
  assign new_n15533_ = ~new_n15529_ & ~new_n15532_;
  assign new_n15534_ = pg35 & ~new_n15533_;
  assign n6682 = new_n15528_ | new_n15534_;
  assign new_n15536_ = ~pg35 & ng4245;
  assign new_n15537_ = ~ng4277 & ~new_n7829_;
  assign new_n15538_ = ~new_n7829_ & ~new_n15537_;
  assign new_n15539_ = ~ng4277 & ~new_n15537_;
  assign new_n15540_ = ~new_n15538_ & ~new_n15539_;
  assign new_n15541_ = pg35 & ~new_n15540_;
  assign n6687 = new_n15536_ | new_n15541_;
  assign new_n15543_ = ~pg35 & ng3343;
  assign new_n15544_ = ng3343 & ~new_n8783_;
  assign new_n15545_ = pg35 & new_n15544_;
  assign n6691 = new_n15543_ | new_n15545_;
  assign new_n15547_ = ~pg35 & ng2259;
  assign new_n15548_ = ng2265 & ~new_n6524_;
  assign new_n15549_ = ng2259 & new_n6524_;
  assign new_n15550_ = ~new_n15548_ & ~new_n15549_;
  assign new_n15551_ = pg35 & ~new_n15550_;
  assign n6696 = new_n15547_ | new_n15551_;
  assign new_n15553_ = ~pg35 & ng1968;
  assign new_n15554_ = ng1974 & ~new_n11266_;
  assign new_n15555_ = ng1968 & new_n11266_;
  assign new_n15556_ = ~new_n15554_ & ~new_n15555_;
  assign new_n15557_ = pg35 & ~new_n15556_;
  assign n6701 = new_n15553_ | new_n15557_;
  assign new_n15559_ = ~pg35 & ng1105;
  assign new_n15560_ = ng1124 & ~new_n11178_;
  assign new_n15561_ = ng1129 & new_n7775_;
  assign new_n15562_ = ng1129 & ~new_n15561_;
  assign new_n15563_ = new_n7775_ & ~new_n15561_;
  assign new_n15564_ = ~new_n15562_ & ~new_n15563_;
  assign new_n15565_ = ng1124 & ~new_n15564_;
  assign new_n15566_ = ~new_n7774_ & new_n15565_;
  assign new_n15567_ = new_n7774_ & ~new_n15564_;
  assign new_n15568_ = ~new_n15566_ & ~new_n15567_;
  assign new_n15569_ = new_n11178_ & ~new_n15568_;
  assign new_n15570_ = ~new_n15560_ & ~new_n15569_;
  assign new_n15571_ = pg35 & ~new_n15570_;
  assign n6706 = new_n15559_ | new_n15571_;
  assign new_n15573_ = ~pg35 & ng2433;
  assign new_n15574_ = ng2421 & ~ng2465;
  assign new_n15575_ = ~new_n7555_ & new_n15574_;
  assign new_n15576_ = ng2429 & ~new_n15575_;
  assign new_n15577_ = ~new_n8465_ & new_n15575_;
  assign new_n15578_ = ~new_n15576_ & ~new_n15577_;
  assign new_n15579_ = pg35 & ~new_n15578_;
  assign n6711 = new_n15573_ | new_n15579_;
  assign new_n15581_ = ~pg35 & ng1974;
  assign new_n15582_ = ng1978 & ~new_n11266_;
  assign new_n15583_ = ~ng1974 & ng1968;
  assign new_n15584_ = ng1968 & ~new_n15583_;
  assign new_n15585_ = ~ng1974 & ~new_n15583_;
  assign new_n15586_ = ~new_n15584_ & ~new_n15585_;
  assign new_n15587_ = new_n11266_ & ~new_n15586_;
  assign new_n15588_ = ~new_n15582_ & ~new_n15587_;
  assign new_n15589_ = pg35 & ~new_n15588_;
  assign n6716 = new_n15581_ | new_n15589_;
  assign new_n15591_ = ~pg35 & ng6386;
  assign new_n15592_ = ng6386 & ~new_n13091_;
  assign new_n15593_ = pg35 & new_n15592_;
  assign n6721 = new_n15591_ | new_n15593_;
  assign new_n15595_ = ~pg35 & ng3203;
  assign new_n15596_ = new_n8744_ & new_n9412_;
  assign new_n15597_ = ng3199 & ~new_n15596_;
  assign new_n15598_ = ~new_n5966_ & new_n15596_;
  assign new_n15599_ = ~new_n15597_ & ~new_n15598_;
  assign new_n15600_ = pg35 & ~new_n15599_;
  assign n6726 = new_n15595_ | new_n15600_;
  assign new_n15602_ = ~pg35 & ng3061;
  assign new_n15603_ = ng3061 & ng3057;
  assign new_n15604_ = pg35 & new_n15603_;
  assign n6731 = new_n15602_ | new_n15604_;
  assign new_n15606_ = ~pg35 & ng1821;
  assign new_n15607_ = ng1740 & ~new_n8571_;
  assign new_n15608_ = new_n8571_ & ~new_n10679_;
  assign new_n15609_ = ~new_n15607_ & ~new_n15608_;
  assign new_n15610_ = pg35 & ~new_n15609_;
  assign n6736 = new_n15606_ | new_n15610_;
  assign new_n15612_ = ~pg35 & ng2675;
  assign new_n15613_ = ng2681 & ~new_n13437_;
  assign new_n15614_ = ng2675 & new_n13437_;
  assign new_n15615_ = ~new_n15613_ & ~new_n15614_;
  assign new_n15616_ = pg35 & ~new_n15615_;
  assign n6741 = new_n15612_ | new_n15616_;
  assign new_n15618_ = ~pg35 & ng2407;
  assign new_n15619_ = ng2413 & ~new_n7260_;
  assign new_n15620_ = ng2407 & new_n7260_;
  assign new_n15621_ = ~new_n15619_ & ~new_n15620_;
  assign new_n15622_ = pg35 & ~new_n15621_;
  assign n6746 = new_n15618_ | new_n15622_;
  assign new_n15624_ = ~pg35 & ng5348;
  assign new_n15625_ = ng5348 & ~new_n12123_;
  assign new_n15626_ = pg35 & new_n15625_;
  assign n6751 = new_n15624_ | new_n15626_;
  assign new_n15628_ = ~pg35 & ng6593;
  assign new_n15629_ = new_n6317_ & new_n6334_;
  assign new_n15630_ = ng6617 & ~new_n15629_;
  assign new_n15631_ = ~new_n5966_ & new_n15629_;
  assign new_n15632_ = ~new_n15630_ & ~new_n15631_;
  assign new_n15633_ = pg35 & ~new_n15632_;
  assign n6756 = new_n15628_ | new_n15633_;
  assign new_n15635_ = ~pg35 & ng2697;
  assign new_n15636_ = n2272 & new_n10448_;
  assign new_n15637_ = ng2704 & ~new_n10448_;
  assign new_n15638_ = ~new_n15636_ & ~new_n15637_;
  assign new_n15639_ = pg35 & ~new_n15638_;
  assign n6761 = new_n15635_ | new_n15639_;
  assign new_n15641_ = ~pg35 & ng2236;
  assign new_n15642_ = ng2250 & ~new_n11373_;
  assign new_n15643_ = ng2236 & new_n15642_;
  assign new_n15644_ = new_n15642_ & ~new_n15643_;
  assign new_n15645_ = ng2236 & ~new_n15643_;
  assign new_n15646_ = ~new_n15644_ & ~new_n15645_;
  assign new_n15647_ = new_n9534_ & ~new_n15646_;
  assign new_n15648_ = ng2250 & ~new_n9534_;
  assign new_n15649_ = ~new_n15647_ & ~new_n15648_;
  assign new_n15650_ = pg35 & ~new_n15649_;
  assign n6766 = new_n15641_ | new_n15650_;
  assign new_n15652_ = ~pg35 & ng2342;
  assign new_n15653_ = ~new_n4724_ & new_n10343_;
  assign new_n15654_ = new_n7259_ & new_n15653_;
  assign new_n15655_ = ng110 & new_n14182_;
  assign new_n15656_ = ng110 & ~new_n15655_;
  assign new_n15657_ = new_n14182_ & ~new_n15655_;
  assign new_n15658_ = ~new_n15656_ & ~new_n15657_;
  assign new_n15659_ = new_n15654_ & ~new_n15658_;
  assign new_n15660_ = ng2357 & ~new_n15654_;
  assign new_n15661_ = ~new_n15659_ & ~new_n15660_;
  assign new_n15662_ = pg35 & ~new_n15661_;
  assign n6771 = new_n15652_ | new_n15662_;
  assign new_n15664_ = ~pg35 & ng5120;
  assign new_n15665_ = ng5115 & ~new_n6190_;
  assign new_n15666_ = ~new_n10296_ & new_n15665_;
  assign new_n15667_ = new_n15665_ & ~new_n15666_;
  assign new_n15668_ = ~new_n10296_ & ~new_n15666_;
  assign new_n15669_ = ~new_n15667_ & ~new_n15668_;
  assign new_n15670_ = pg33959 & ~new_n15669_;
  assign new_n15671_ = ng5115 & ~pg33959;
  assign new_n15672_ = ~new_n15670_ & ~new_n15671_;
  assign new_n15673_ = pg35 & ~new_n15672_;
  assign n6776 = new_n15664_ | new_n15673_;
  assign new_n15675_ = ~pg35 & ng5579;
  assign new_n15676_ = new_n6886_ & new_n11751_;
  assign new_n15677_ = ng5595 & ~new_n15676_;
  assign new_n15678_ = ~new_n5966_ & new_n15676_;
  assign new_n15679_ = ~new_n15677_ & ~new_n15678_;
  assign new_n15680_ = pg35 & ~new_n15679_;
  assign n6781 = new_n15675_ | new_n15680_;
  assign new_n15682_ = ~pg35 & ng2729;
  assign new_n15683_ = ng2735 & ~new_n6641_;
  assign new_n15684_ = ~ng2735 & new_n6641_;
  assign new_n15685_ = ~new_n15683_ & ~new_n15684_;
  assign new_n15686_ = ng2841 & ~new_n15685_;
  assign new_n15687_ = ng2841 & ~new_n15686_;
  assign new_n15688_ = pg35 & ~new_n15687_;
  assign n6786 = new_n15682_ | new_n15688_;
  assign new_n15690_ = ~pg35 & ng4653;
  assign new_n15691_ = ng4659 & new_n10528_;
  assign new_n15692_ = ~new_n14290_ & new_n15691_;
  assign new_n15693_ = ~ng4659 & new_n10528_;
  assign new_n15694_ = new_n14290_ & new_n15693_;
  assign new_n15695_ = ~new_n15692_ & ~new_n15694_;
  assign new_n15696_ = pg35 & ~new_n15695_;
  assign n6791 = new_n15690_ | new_n15696_;
  assign new_n15698_ = ~pg35 & ng1099;
  assign new_n15699_ = ng1094 & ~new_n5887_;
  assign new_n15700_ = ng1135 & new_n7775_;
  assign new_n15701_ = ng1135 & ~new_n15700_;
  assign new_n15702_ = new_n7775_ & ~new_n15700_;
  assign new_n15703_ = ~new_n15701_ & ~new_n15702_;
  assign new_n15704_ = ng1094 & ~new_n15703_;
  assign new_n15705_ = ~new_n7774_ & new_n15704_;
  assign new_n15706_ = new_n7774_ & ~new_n15703_;
  assign new_n15707_ = ~new_n15705_ & ~new_n15706_;
  assign new_n15708_ = new_n5887_ & ~new_n15707_;
  assign new_n15709_ = ~new_n15699_ & ~new_n15708_;
  assign new_n15710_ = pg35 & ~new_n15709_;
  assign n6796 = new_n15698_ | new_n15710_;
  assign new_n15712_ = ~pg35 & ng542;
  assign new_n15713_ = ng12 & n6079;
  assign new_n15714_ = new_n4910_ & new_n15713_;
  assign new_n15715_ = ~ng301 & ~ng534;
  assign new_n15716_ = ~new_n15714_ & ~new_n15715_;
  assign new_n15717_ = pg35 & new_n15716_;
  assign n6801 = new_n15712_ | new_n15717_;
  assign new_n15719_ = ~pg35 & ng1526;
  assign new_n15720_ = ng1500 & ng1339;
  assign new_n15721_ = ng1521 & ~ng1500;
  assign new_n15722_ = ~new_n15720_ & ~new_n15721_;
  assign new_n15723_ = pg35 & ~new_n15722_;
  assign n6806 = new_n15719_ | new_n15723_;
  assign new_n15725_ = pg35 & ng4742;
  assign new_n15726_ = ~pg35 & new_n15725_;
  assign n6814 = new_n13158_ | new_n15726_;
  assign new_n15728_ = ~pg35 & ng767;
  assign new_n15729_ = ng772 & ~new_n6578_;
  assign new_n15730_ = ~new_n6590_ & new_n15729_;
  assign new_n15731_ = ~ng772 & new_n6590_;
  assign new_n15732_ = ~new_n15730_ & ~new_n15731_;
  assign new_n15733_ = pg35 & ~new_n15732_;
  assign n6819 = new_n15728_ | new_n15733_;
  assign new_n15735_ = ~pg35 & ng2567;
  assign new_n15736_ = ~ng2599 & ng2555;
  assign new_n15737_ = ~new_n7174_ & new_n15736_;
  assign new_n15738_ = ng2563 & ~new_n15737_;
  assign new_n15739_ = ~new_n8484_ & new_n15737_;
  assign new_n15740_ = ~new_n15738_ & ~new_n15739_;
  assign new_n15741_ = pg35 & ~new_n15740_;
  assign n6824 = new_n15735_ | new_n15741_;
  assign new_n15743_ = ~pg35 & ng3582;
  assign new_n15744_ = new_n7697_ & new_n11130_;
  assign new_n15745_ = ng3598 & ~new_n15744_;
  assign new_n15746_ = ~new_n5966_ & new_n15744_;
  assign new_n15747_ = ~new_n15745_ & ~new_n15746_;
  assign new_n15748_ = pg35 & ~new_n15747_;
  assign n6829 = new_n15743_ | new_n15748_;
  assign new_n15750_ = ~pg35 & ng291;
  assign new_n15751_ = ~ng294 & new_n6026_;
  assign new_n15752_ = ng294 & new_n6021_;
  assign new_n15753_ = ~new_n6026_ & new_n15752_;
  assign new_n15754_ = ~new_n15751_ & ~new_n15753_;
  assign new_n15755_ = pg35 & ~new_n15754_;
  assign n6834 = new_n15750_ | new_n15755_;
  assign new_n15757_ = ~pg35 & ng904;
  assign new_n15758_ = ~ng921 & new_n7073_;
  assign new_n15759_ = ng1227 & ng921;
  assign new_n15760_ = ~new_n7073_ & new_n15759_;
  assign new_n15761_ = ~new_n15758_ & ~new_n15760_;
  assign new_n15762_ = pg35 & ~new_n15761_;
  assign n6839 = new_n15757_ | new_n15762_;
  assign new_n15764_ = ~pg35 & ng3518;
  assign new_n15765_ = ng3522 & ~new_n9472_;
  assign new_n15766_ = ~ng3518 & new_n15765_;
  assign new_n15767_ = ~ng3522 & ~new_n9472_;
  assign new_n15768_ = ng3518 & new_n15767_;
  assign new_n15769_ = ~new_n15766_ & ~new_n15768_;
  assign new_n15770_ = pg35 & ~new_n15769_;
  assign n6844 = new_n15764_ | new_n15770_;
  assign new_n15772_ = ~pg35 & ng1373;
  assign new_n15773_ = new_n14126_ & ~new_n14128_;
  assign new_n15774_ = ng1379 & ~new_n15773_;
  assign new_n15775_ = ~ng1379 & new_n6306_;
  assign new_n15776_ = new_n15773_ & new_n15775_;
  assign new_n15777_ = ~new_n15774_ & ~new_n15776_;
  assign new_n15778_ = pg35 & ~new_n15777_;
  assign n6849 = new_n15772_ | new_n15778_;
  assign new_n15780_ = ~pg35 & ng5571;
  assign new_n15781_ = new_n6886_ & new_n8033_;
  assign new_n15782_ = ng5587 & ~new_n15781_;
  assign new_n15783_ = ~new_n5966_ & new_n15781_;
  assign new_n15784_ = ~new_n15782_ & ~new_n15783_;
  assign new_n15785_ = pg35 & ~new_n15784_;
  assign n6854 = new_n15780_ | new_n15785_;
  assign new_n15787_ = ~pg35 & ng1339;
  assign new_n15788_ = ~ng1582 & ~ng1333;
  assign new_n15789_ = ~ng1500 & new_n15788_;
  assign new_n15790_ = ~ng1459 & new_n15789_;
  assign new_n15791_ = ~ng1399 & new_n15790_;
  assign new_n15792_ = new_n12008_ & new_n15791_;
  assign new_n15793_ = new_n15791_ & ~new_n15792_;
  assign new_n15794_ = new_n12008_ & ~new_n15792_;
  assign new_n15795_ = ~new_n15793_ & ~new_n15794_;
  assign new_n15796_ = pg35 & ~new_n15795_;
  assign n6859 = new_n15787_ | new_n15796_;
  assign new_n15798_ = ~pg35 & ng4258;
  assign new_n15799_ = ~ng4264 & ng4258;
  assign new_n15800_ = ng4264 & ~ng4258;
  assign new_n15801_ = ~new_n15799_ & ~new_n15800_;
  assign new_n15802_ = pg35 & ~new_n15801_;
  assign n6863 = new_n15798_ | new_n15802_;
  assign new_n15804_ = ~pg35 & ng6275;
  assign new_n15805_ = new_n7063_ & new_n9573_;
  assign new_n15806_ = ng6291 & ~new_n15805_;
  assign new_n15807_ = ~new_n5966_ & new_n15805_;
  assign new_n15808_ = ~new_n15806_ & ~new_n15807_;
  assign new_n15809_ = pg35 & ~new_n15808_;
  assign n6868 = new_n15804_ | new_n15809_;
  assign new_n15811_ = ~pg35 & ng2941;
  assign new_n15812_ = new_n4937_ & new_n15713_;
  assign new_n15813_ = new_n4683_ & new_n4844_1_;
  assign new_n15814_ = ~ng2946 & new_n15813_;
  assign new_n15815_ = new_n5834_1_ & new_n15814_;
  assign new_n15816_ = new_n4867_1_ & new_n15815_;
  assign new_n15817_ = ~ng2955 & new_n15816_;
  assign new_n15818_ = ~new_n15812_ & ~new_n15817_;
  assign new_n15819_ = pg35 & new_n15818_;
  assign n6873 = new_n15811_ | new_n15819_;
  assign new_n15821_ = ~pg35 & ng3106;
  assign new_n15822_ = ng3115 & ~new_n10989_;
  assign new_n15823_ = ng3106 & ng3111;
  assign new_n15824_ = ng3111 & ~new_n15823_;
  assign new_n15825_ = ng3106 & ~new_n15823_;
  assign new_n15826_ = ~new_n15824_ & ~new_n15825_;
  assign new_n15827_ = new_n10989_ & ~new_n15826_;
  assign new_n15828_ = ~new_n15822_ & ~new_n15827_;
  assign new_n15829_ = pg35 & ~new_n15828_;
  assign n6878 = new_n15821_ | new_n15829_;
  assign new_n15831_ = ~pg35 & ng1720;
  assign new_n15832_ = ng1724 & ~new_n7231_;
  assign new_n15833_ = ~ng1720 & ng1714;
  assign new_n15834_ = ng1714 & ~new_n15833_;
  assign new_n15835_ = ~ng1720 & ~new_n15833_;
  assign new_n15836_ = ~new_n15834_ & ~new_n15835_;
  assign new_n15837_ = new_n7231_ & ~new_n15836_;
  assign new_n15838_ = ~new_n15832_ & ~new_n15837_;
  assign new_n15839_ = pg35 & ~new_n15838_;
  assign n6883 = new_n15831_ | new_n15839_;
  assign new_n15841_ = ~pg35 & ng6173;
  assign new_n15842_ = ng6177 & ~new_n6700_;
  assign new_n15843_ = ~ng6173 & ng6167;
  assign new_n15844_ = ng6167 & ~new_n15843_;
  assign new_n15845_ = ~ng6173 & ~new_n15843_;
  assign new_n15846_ = ~new_n15844_ & ~new_n15845_;
  assign new_n15847_ = new_n6700_ & ~new_n15846_;
  assign new_n15848_ = ~new_n15842_ & ~new_n15847_;
  assign new_n15849_ = pg35 & ~new_n15848_;
  assign n6888 = new_n15841_ | new_n15849_;
  assign new_n15851_ = ~pg35 & ng4584;
  assign new_n15852_ = ~ng4593 & new_n8853_;
  assign new_n15853_ = new_n12747_ & new_n15852_;
  assign new_n15854_ = ng4593 & new_n8853_;
  assign new_n15855_ = ~new_n12747_ & new_n15854_;
  assign new_n15856_ = ~new_n15853_ & ~new_n15855_;
  assign new_n15857_ = pg35 & ~new_n15856_;
  assign n6893 = new_n15851_ | new_n15857_;
  assign new_n15859_ = ~pg35 & ng1018;
  assign new_n15860_ = ng1024 & ~new_n6142_;
  assign new_n15861_ = new_n6142_ & new_n6143_;
  assign new_n15862_ = ~new_n15860_ & ~new_n15861_;
  assign new_n15863_ = pg35 & ~new_n15862_;
  assign n6898 = new_n15859_ | new_n15863_;
  assign new_n15865_ = ~pg35 & ng385;
  assign new_n15866_ = pg35 & new_n11258_;
  assign n6907 = new_n15865_ | new_n15866_;
  assign new_n15868_ = ~pg35 & ng5052;
  assign new_n15869_ = ~ng5052 & new_n8141_;
  assign new_n15870_ = ng5052 & new_n8146_;
  assign new_n15871_ = ~new_n15869_ & ~new_n15870_;
  assign new_n15872_ = ~ng5057 & ~new_n15871_;
  assign new_n15873_ = ng5057 & new_n8107_;
  assign new_n15874_ = new_n15871_ & new_n15873_;
  assign new_n15875_ = ~new_n15872_ & ~new_n15874_;
  assign new_n15876_ = pg35 & ~new_n15875_;
  assign n6912 = new_n15868_ | new_n15876_;
  assign new_n15878_ = ~pg35 & ng4801;
  assign new_n15879_ = ng4801 & new_n6155_;
  assign new_n15880_ = ng4776 & new_n6161_;
  assign new_n15881_ = ~new_n15879_ & new_n15880_;
  assign new_n15882_ = ~ng4776 & new_n6161_;
  assign new_n15883_ = new_n15879_ & new_n15882_;
  assign new_n15884_ = ~new_n15881_ & ~new_n15883_;
  assign new_n15885_ = pg35 & ~new_n15884_;
  assign n6921 = new_n15878_ | new_n15885_;
  assign new_n15887_ = ~pg35 & ng5575;
  assign new_n15888_ = new_n6886_ & new_n8129_;
  assign new_n15889_ = ng5591 & ~new_n15888_;
  assign new_n15890_ = ~new_n5966_ & new_n15888_;
  assign new_n15891_ = ~new_n15889_ & ~new_n15890_;
  assign new_n15892_ = pg35 & ~new_n15891_;
  assign n6926 = new_n15887_ | new_n15892_;
  assign new_n15894_ = pg35 & ng5499;
  assign new_n15895_ = ~pg35 & new_n15894_;
  assign new_n15896_ = n5814 & new_n6181_;
  assign new_n15897_ = ng5507 & ~new_n6181_;
  assign new_n15898_ = ~new_n15896_ & ~new_n15897_;
  assign new_n15899_ = pg35 & ~new_n15898_;
  assign n6931 = new_n15895_ | new_n15899_;
  assign new_n15901_ = ~pg35 & ng6082;
  assign new_n15902_ = ~ng6082 & new_n10189_;
  assign new_n15903_ = ng6082 & new_n10193_;
  assign new_n15904_ = ~new_n15902_ & ~new_n15903_;
  assign new_n15905_ = ng6088 & new_n7527_;
  assign new_n15906_ = new_n15904_ & new_n15905_;
  assign new_n15907_ = ~ng6088 & ~new_n15904_;
  assign new_n15908_ = ~new_n15906_ & ~new_n15907_;
  assign new_n15909_ = pg35 & ~new_n15908_;
  assign n6936 = new_n15901_ | new_n15909_;
  assign new_n15911_ = ~pg35 & ng460;
  assign new_n15912_ = ng452 & ~new_n5994_;
  assign new_n15913_ = ng460 & new_n5994_;
  assign new_n15914_ = ~new_n15912_ & ~new_n15913_;
  assign new_n15915_ = pg35 & ~new_n15914_;
  assign n6941 = new_n15911_ | new_n15915_;
  assign new_n15917_ = ~pg35 & ng794;
  assign new_n15918_ = ng807 & ~new_n6578_;
  assign new_n15919_ = ~new_n12502_ & new_n15918_;
  assign new_n15920_ = ~ng807 & new_n12502_;
  assign new_n15921_ = ~new_n15919_ & ~new_n15920_;
  assign new_n15922_ = pg35 & ~new_n15921_;
  assign n6946 = new_n15917_ | new_n15922_;
  assign new_n15924_ = ~pg35 & ng1604;
  assign new_n15925_ = ~ng1636 & ng1592;
  assign new_n15926_ = ~new_n7537_1_ & new_n15925_;
  assign new_n15927_ = ng1600 & ~new_n15926_;
  assign new_n15928_ = ~new_n7543_ & new_n15926_;
  assign new_n15929_ = ~new_n15927_ & ~new_n15928_;
  assign new_n15930_ = pg35 & ~new_n15929_;
  assign n6951 = new_n15924_ | new_n15930_;
  assign new_n15932_ = ~pg35 & ng4639;
  assign new_n15933_ = ng4621 & new_n8339_;
  assign new_n15934_ = ~ng4639 & new_n15933_;
  assign new_n15935_ = ~ng4621 & new_n8339_;
  assign new_n15936_ = ng4639 & new_n15935_;
  assign new_n15937_ = ~new_n15934_ & ~new_n15936_;
  assign new_n15938_ = pg35 & ~new_n15937_;
  assign n6956 = new_n15932_ | new_n15938_;
  assign new_n15940_ = ~pg35 & ng1152;
  assign new_n15941_ = ng1099 & ~new_n7772_;
  assign new_n15942_ = ng1152 & new_n7772_;
  assign new_n15943_ = ~new_n15941_ & ~new_n15942_;
  assign new_n15944_ = pg35 & ~new_n15943_;
  assign n6961 = new_n15940_ | new_n15944_;
  assign new_n15946_ = ~pg35 & ng2012;
  assign new_n15947_ = ~new_n7025_ & new_n14732_;
  assign new_n15948_ = ng2024 & ~new_n15947_;
  assign new_n15949_ = ~new_n7032_ & new_n15947_;
  assign new_n15950_ = ~new_n15948_ & ~new_n15949_;
  assign new_n15951_ = pg35 & ~new_n15950_;
  assign n6966 = new_n15946_ | new_n15951_;
  assign n6971 = ~pg35 & ng896;
  assign new_n15954_ = ~pg35 & ng4235;
  assign new_n15955_ = ~ng4213 & ~ng4219;
  assign new_n15956_ = ~ng4222 & ~ng4216;
  assign new_n15957_ = new_n15955_ & new_n15956_;
  assign new_n15958_ = ~ng4226 & ~ng4232;
  assign new_n15959_ = ~ng4229 & ~ng4235;
  assign new_n15960_ = new_n15958_ & new_n15959_;
  assign new_n15961_ = new_n15957_ & new_n15960_;
  assign new_n15962_ = ~ng4185 & new_n15961_;
  assign new_n15963_ = ng4222 & ng4235;
  assign new_n15964_ = ng4235 & ~new_n15963_;
  assign new_n15965_ = ng4222 & ~new_n15963_;
  assign new_n15966_ = ~new_n15964_ & ~new_n15965_;
  assign new_n15967_ = ~new_n15962_ & new_n15966_;
  assign new_n15968_ = new_n11397_ & ~new_n15967_;
  assign new_n15969_ = ~new_n15967_ & ~new_n15968_;
  assign new_n15970_ = new_n11397_ & ~new_n15968_;
  assign new_n15971_ = ~new_n15969_ & ~new_n15970_;
  assign new_n15972_ = pg35 & ~new_n15971_;
  assign n6976 = new_n15954_ | new_n15972_;
  assign new_n15974_ = ~pg35 & ng2735;
  assign new_n15975_ = ~ng2741 & new_n6642_1_;
  assign new_n15976_ = ng2741 & ~new_n6642_1_;
  assign new_n15977_ = ~new_n15975_ & ~new_n15976_;
  assign new_n15978_ = ng2841 & ~new_n15977_;
  assign new_n15979_ = pg35 & new_n15978_;
  assign n6981 = new_n15974_ | new_n15979_;
  assign new_n15981_ = ~pg35 & ng2223;
  assign new_n15982_ = ~ng2208 & ~new_n11142_;
  assign new_n15983_ = new_n9534_ & ~new_n15982_;
  assign new_n15984_ = ng2217 & ~new_n9534_;
  assign new_n15985_ = ~new_n15983_ & ~new_n15984_;
  assign new_n15986_ = pg35 & ~new_n15985_;
  assign n6986 = new_n15981_ | new_n15986_;
  assign new_n15988_ = ~pg35 & ng471;
  assign new_n15989_ = ng464 & ~new_n5994_;
  assign new_n15990_ = ng471 & new_n5994_;
  assign new_n15991_ = ~new_n15989_ & ~new_n15990_;
  assign new_n15992_ = pg35 & ~new_n15991_;
  assign n6991 = new_n15988_ | new_n15992_;
  assign new_n15994_ = ~pg35 & ng6215;
  assign new_n15995_ = ng6219 & ~new_n5852_;
  assign new_n15996_ = ~ng6215 & new_n15995_;
  assign new_n15997_ = ~ng6219 & ~new_n5852_;
  assign new_n15998_ = ng6215 & new_n15997_;
  assign new_n15999_ = ~new_n15996_ & ~new_n15998_;
  assign new_n16000_ = pg35 & ~new_n15999_;
  assign n6996 = new_n15994_ | new_n16000_;
  assign new_n16002_ = ~pg35 & ng1710;
  assign new_n16003_ = ng1714 & ~new_n10846_;
  assign new_n16004_ = ~ng1714 & new_n10846_;
  assign new_n16005_ = ~new_n16003_ & ~new_n16004_;
  assign new_n16006_ = pg35 & ~new_n16005_;
  assign n7001 = new_n16002_ | new_n16006_;
  assign new_n16008_ = ~pg35 & ng1964;
  assign new_n16009_ = ng1968 & ~new_n8172_;
  assign new_n16010_ = ~ng1968 & new_n8172_;
  assign new_n16011_ = ~new_n16009_ & ~new_n16010_;
  assign new_n16012_ = pg35 & ~new_n16011_;
  assign n7006 = new_n16008_ | new_n16012_;
  assign new_n16014_ = ~pg35 & ng4871;
  assign new_n16015_ = ng4871 & ~new_n7605_;
  assign new_n16016_ = pg35 & new_n16015_;
  assign n7011 = new_n16014_ | new_n16016_;
  assign new_n16018_ = pg35 & ng6545;
  assign new_n16019_ = ~pg35 & new_n16018_;
  assign new_n16020_ = ng3298 & ~ng3274;
  assign new_n16021_ = ~ng3267 & ng3274;
  assign new_n16022_ = ~new_n16020_ & ~new_n16021_;
  assign new_n16023_ = ~new_n8782_ & new_n16022_;
  assign new_n16024_ = ng3310 & ~ng3281;
  assign new_n16025_ = ng3281 & ~ng3303;
  assign new_n16026_ = ~ng3310 & ng3267;
  assign new_n16027_ = new_n16023_ & ~new_n16024_;
  assign new_n16028_ = ~new_n16025_ & new_n16027_;
  assign new_n16029_ = ~new_n16026_ & new_n16028_;
  assign new_n16030_ = pg35 & new_n16029_;
  assign n7016 = new_n16019_ | new_n16030_;
  assign new_n16032_ = pg35 & ng4821;
  assign new_n16033_ = ~pg35 & new_n16032_;
  assign new_n16034_ = ng5503 & ~new_n10882_;
  assign new_n16035_ = ~new_n5966_ & new_n16034_;
  assign new_n16036_ = new_n16034_ & ~new_n16035_;
  assign new_n16037_ = ~new_n5966_ & ~new_n16035_;
  assign new_n16038_ = ~new_n16036_ & ~new_n16037_;
  assign new_n16039_ = pg35 & ~new_n16038_;
  assign n7023 = new_n16033_ | new_n16039_;
  assign new_n16041_ = ~pg35 & ng590;
  assign new_n16042_ = ng595 & ~new_n6545_;
  assign new_n16043_ = ~new_n6566_1_ & new_n16042_;
  assign new_n16044_ = ~ng595 & new_n6566_1_;
  assign new_n16045_ = ~new_n16043_ & ~new_n16044_;
  assign new_n16046_ = pg35 & ~new_n16045_;
  assign n7031 = new_n16041_ | new_n16046_;
  assign new_n16048_ = ~pg35 & ng3546;
  assign new_n16049_ = new_n7038_ & new_n12309_;
  assign new_n16050_ = ng3542 & ~new_n16049_;
  assign new_n16051_ = ~new_n5966_ & new_n16049_;
  assign new_n16052_ = ~new_n16050_ & ~new_n16051_;
  assign new_n16053_ = pg35 & ~new_n16052_;
  assign n7036 = new_n16048_ | new_n16053_;
  assign new_n16055_ = ~pg35 & ng854;
  assign new_n16056_ = ng847 & ~new_n6067_;
  assign new_n16057_ = ng854 & new_n6067_;
  assign new_n16058_ = ~new_n16056_ & ~new_n16057_;
  assign new_n16059_ = pg35 & ~new_n16058_;
  assign n7041 = new_n16055_ | new_n16059_;
  assign new_n16061_ = pg35 & ng5507;
  assign new_n16062_ = ~pg35 & new_n16061_;
  assign new_n16063_ = ~ng5976 & ng6000;
  assign new_n16064_ = ~ng5969 & ng5976;
  assign new_n16065_ = ~new_n16063_ & ~new_n16064_;
  assign new_n16066_ = ~new_n6452_ & new_n16065_;
  assign new_n16067_ = ng6012 & ~ng5983;
  assign new_n16068_ = ng5983 & ~ng6005;
  assign new_n16069_ = ~ng6012 & ng5969;
  assign new_n16070_ = new_n16066_ & ~new_n16067_;
  assign new_n16071_ = ~new_n16068_ & new_n16070_;
  assign new_n16072_ = ~new_n16069_ & new_n16071_;
  assign new_n16073_ = pg35 & new_n16072_;
  assign n7046 = new_n16062_ | new_n16073_;
  assign new_n16075_ = ~pg35 & ng1740;
  assign new_n16076_ = ~ng1772 & ng1728;
  assign new_n16077_ = ~new_n6236_ & new_n16076_;
  assign new_n16078_ = ng1736 & ~new_n16077_;
  assign new_n16079_ = ~new_n10679_ & new_n16077_;
  assign new_n16080_ = ~new_n16078_ & ~new_n16079_;
  assign new_n16081_ = pg35 & ~new_n16080_;
  assign n7050 = new_n16075_ | new_n16081_;
  assign new_n16083_ = ng22 & pg34919;
  assign new_n16084_ = ~ng22 & n5814;
  assign n7055 = new_n16083_ | new_n16084_;
  assign new_n16086_ = ~pg35 & ng2384;
  assign new_n16087_ = new_n7259_ & new_n14179_;
  assign new_n16088_ = ng2389 & ~new_n16087_;
  assign new_n16089_ = ng2380 & ng2384;
  assign new_n16090_ = ng2384 & ~new_n16089_;
  assign new_n16091_ = ng2380 & ~new_n16089_;
  assign new_n16092_ = ~new_n16090_ & ~new_n16091_;
  assign new_n16093_ = new_n16087_ & ~new_n16092_;
  assign new_n16094_ = ~new_n16088_ & ~new_n16093_;
  assign new_n16095_ = pg35 & ~new_n16094_;
  assign n7060 = new_n16086_ | new_n16095_;
  assign new_n16097_ = ~pg35 & ng3774;
  assign new_n16098_ = ng3774 & ~ng3782;
  assign new_n16099_ = ~ng3774 & ng3782;
  assign new_n16100_ = ~new_n16098_ & ~new_n16099_;
  assign new_n16101_ = pg35 & ~new_n16100_;
  assign n7065 = new_n16097_ | new_n16101_;
  assign new_n16103_ = ~pg35 & ng2619;
  assign new_n16104_ = ~ng2610 & ng2587;
  assign new_n16105_ = ng2579 & new_n16104_;
  assign new_n16106_ = ~ng2619 & ~ng2587;
  assign new_n16107_ = ng2575 & new_n16106_;
  assign new_n16108_ = ng2583 & new_n5219_;
  assign new_n16109_ = ~new_n16105_ & ~new_n16107_;
  assign new_n16110_ = ~new_n16108_ & new_n16109_;
  assign new_n16111_ = ng2563 & new_n10923_;
  assign new_n16112_ = ng2567 & new_n13436_;
  assign new_n16113_ = ng2571 & new_n12264_;
  assign new_n16114_ = new_n16110_ & ~new_n16111_;
  assign new_n16115_ = ~new_n16112_ & ~new_n16113_;
  assign new_n16116_ = new_n16114_ & new_n16115_;
  assign new_n16117_ = new_n10306_ & ~new_n16116_;
  assign new_n16118_ = ng2638 & ~new_n10306_;
  assign new_n16119_ = ~new_n16117_ & ~new_n16118_;
  assign new_n16120_ = pg35 & ~new_n16119_;
  assign n7070 = new_n16103_ | new_n16120_;
  assign new_n16122_ = ~pg35 & ng2051;
  assign new_n16123_ = ~new_n4724_ & new_n13377_;
  assign new_n16124_ = new_n9143_ & new_n16123_;
  assign new_n16125_ = ng110 & new_n10175_;
  assign new_n16126_ = ng110 & ~new_n16125_;
  assign new_n16127_ = new_n10175_ & ~new_n16125_;
  assign new_n16128_ = ~new_n16126_ & ~new_n16127_;
  assign new_n16129_ = new_n16124_ & ~new_n16128_;
  assign new_n16130_ = ng2066 & ~new_n16124_;
  assign new_n16131_ = ~new_n16129_ & ~new_n16130_;
  assign new_n16132_ = pg35 & ~new_n16131_;
  assign n7075 = new_n16122_ | new_n16132_;
  assign new_n16134_ = pg35 & ng4157;
  assign new_n16135_ = ~pg35 & new_n16134_;
  assign new_n16136_ = pg35 & ~ng4258;
  assign n7080 = new_n16135_ | new_n16136_;
  assign new_n16138_ = ~pg35 & ng5208;
  assign new_n16139_ = new_n10722_ & new_n11577_;
  assign new_n16140_ = ng5232 & ~new_n16139_;
  assign new_n16141_ = ~new_n5966_ & new_n16139_;
  assign new_n16142_ = ~new_n16140_ & ~new_n16141_;
  assign new_n16143_ = pg35 & ~new_n16142_;
  assign n7085 = new_n16138_ | new_n16143_;
  assign new_n16145_ = ~pg35 & ng6069;
  assign new_n16146_ = ~new_n10187_ & ~new_n10191_;
  assign new_n16147_ = ~ng6073 & ~new_n16146_;
  assign new_n16148_ = ng6073 & new_n7527_;
  assign new_n16149_ = new_n16146_ & new_n16148_;
  assign new_n16150_ = ~new_n16147_ & ~new_n16149_;
  assign new_n16151_ = pg35 & ~new_n16150_;
  assign n7098 = new_n16145_ | new_n16151_;
  assign new_n16153_ = pg35 & ng3333;
  assign new_n16154_ = ~pg35 & new_n16153_;
  assign new_n16155_ = ng3147 & ~new_n7152_;
  assign new_n16156_ = ~new_n5966_ & new_n16155_;
  assign new_n16157_ = new_n16155_ & ~new_n16156_;
  assign new_n16158_ = ~new_n5966_ & ~new_n16156_;
  assign new_n16159_ = ~new_n16157_ & ~new_n16158_;
  assign new_n16160_ = pg35 & ~new_n16159_;
  assign n7103 = new_n16154_ | new_n16160_;
  assign new_n16162_ = ~pg35 & new_n4779_;
  assign n7108 = new_n5918_ | new_n16162_;
  assign new_n16164_ = ~pg35 & ng5551;
  assign new_n16165_ = new_n8035_ & new_n8129_;
  assign new_n16166_ = ng5547 & ~new_n16165_;
  assign new_n16167_ = ~new_n5966_ & new_n16165_;
  assign new_n16168_ = ~new_n16166_ & ~new_n16167_;
  assign new_n16169_ = pg35 & ~new_n16168_;
  assign n7113 = new_n16164_ | new_n16169_;
  assign new_n16171_ = ~pg35 & ng4119;
  assign new_n16172_ = ng4122 & ~new_n10362_;
  assign new_n16173_ = ng4145 & new_n10362_;
  assign new_n16174_ = ~new_n16172_ & ~new_n16173_;
  assign new_n16175_ = pg35 & ~new_n16174_;
  assign n7118 = new_n16171_ | new_n16175_;
  assign new_n16177_ = ~pg35 & ng1404;
  assign new_n16178_ = ~ng1570 & ng1404;
  assign new_n16179_ = ng1570 & ~ng1395;
  assign new_n16180_ = ~ng1404 & new_n16179_;
  assign new_n16181_ = ~new_n16178_ & ~new_n16180_;
  assign new_n16182_ = ng1399 & ~new_n16181_;
  assign new_n16183_ = pg35 & ~new_n16182_;
  assign n7123 = new_n16177_ | new_n16183_;
  assign new_n16185_ = ~pg35 & ng1616;
  assign new_n16186_ = ng1668 & ng1592;
  assign new_n16187_ = ~new_n7537_1_ & new_n16186_;
  assign new_n16188_ = ng1612 & ~new_n16187_;
  assign new_n16189_ = ~new_n7543_ & new_n16187_;
  assign new_n16190_ = ~new_n16188_ & ~new_n16189_;
  assign new_n16191_ = pg35 & ~new_n16190_;
  assign n7128 = new_n16185_ | new_n16191_;
  assign new_n16193_ = ~pg35 & ng5849;
  assign new_n16194_ = ng5813 & ~new_n10071_;
  assign new_n16195_ = ng5849 & new_n10071_;
  assign new_n16196_ = ~new_n16194_ & ~new_n16195_;
  assign new_n16197_ = pg35 & ~new_n16196_;
  assign n7133 = new_n16193_ | new_n16197_;
  assign new_n16199_ = pg35 & ng4138;
  assign new_n16200_ = ~pg35 & new_n16199_;
  assign new_n16201_ = new_n4927_ & new_n15713_;
  assign new_n16202_ = ~ng4153 & ~ng4172;
  assign new_n16203_ = ~new_n16201_ & ~new_n16202_;
  assign new_n16204_ = pg35 & new_n16203_;
  assign n7138 = new_n16200_ | new_n16204_;
  assign new_n16206_ = ~pg35 & ng3361;
  assign new_n16207_ = ~ng3401 & ~ng3361;
  assign new_n16208_ = ng3355 & new_n16207_;
  assign new_n16209_ = ~ng3355 & new_n8400_;
  assign new_n16210_ = ~new_n16207_ & new_n16209_;
  assign new_n16211_ = ~new_n16208_ & ~new_n16210_;
  assign new_n16212_ = pg35 & ~new_n16211_;
  assign n7143 = new_n16206_ | new_n16212_;
  assign new_n16214_ = ~pg35 & ng482;
  assign new_n16215_ = ng482 & new_n6782_;
  assign new_n16216_ = ~ng490 & ~new_n6494_;
  assign new_n16217_ = ~new_n16215_ & ~new_n16216_;
  assign new_n16218_ = ng490 & ~new_n6494_;
  assign new_n16219_ = new_n16215_ & ~new_n16218_;
  assign new_n16220_ = ~new_n16217_ & ~new_n16219_;
  assign new_n16221_ = pg35 & ~new_n16220_;
  assign n7148 = new_n16214_ | new_n16221_;
  assign new_n16223_ = ~pg35 & ng3462;
  assign new_n16224_ = ng3457 & ~new_n7427_;
  assign new_n16225_ = ~new_n14853_ & new_n16224_;
  assign new_n16226_ = new_n16224_ & ~new_n16225_;
  assign new_n16227_ = ~new_n14853_ & ~new_n16225_;
  assign new_n16228_ = ~new_n16226_ & ~new_n16227_;
  assign new_n16229_ = new_n7431_ & ~new_n16228_;
  assign new_n16230_ = ng3457 & ~new_n7431_;
  assign new_n16231_ = ~new_n16229_ & ~new_n16230_;
  assign new_n16232_ = pg35 & ~new_n16231_;
  assign n7153 = new_n16223_ | new_n16232_;
  assign new_n16234_ = ~pg35 & ng2890;
  assign new_n16235_ = n4955 & new_n5972_;
  assign new_n16236_ = ng2844 & ~new_n5972_;
  assign new_n16237_ = ~new_n16235_ & ~new_n16236_;
  assign new_n16238_ = pg35 & ~new_n16237_;
  assign n7158 = new_n16234_ | new_n16238_;
  assign new_n16240_ = ~pg35 & ng4785;
  assign new_n16241_ = ng4785 & new_n6157_;
  assign new_n16242_ = ng4709 & ~new_n6160_;
  assign new_n16243_ = ~new_n16241_ & new_n16242_;
  assign new_n16244_ = ~ng4709 & ~new_n6160_;
  assign new_n16245_ = new_n16241_ & new_n16244_;
  assign new_n16246_ = ~new_n16243_ & ~new_n16245_;
  assign new_n16247_ = pg35 & ~new_n16246_;
  assign n7163 = new_n16240_ | new_n16247_;
  assign new_n16249_ = pg35 & ng1300;
  assign new_n16250_ = ~pg35 & new_n16249_;
  assign new_n16251_ = n6079 & new_n8829_;
  assign new_n16252_ = ng1291 & ~new_n8829_;
  assign new_n16253_ = ~new_n16251_ & ~new_n16252_;
  assign new_n16254_ = pg35 & ~new_n16253_;
  assign n7168 = new_n16250_ | new_n16254_;
  assign new_n16256_ = ~pg35 & ng2437;
  assign new_n16257_ = ~new_n7555_ & new_n9357_;
  assign new_n16258_ = ng2449 & ~new_n16257_;
  assign new_n16259_ = ~new_n8465_ & new_n16257_;
  assign new_n16260_ = ~new_n16258_ & ~new_n16259_;
  assign new_n16261_ = pg35 & ~new_n16260_;
  assign n7173 = new_n16256_ | new_n16261_;
  assign new_n16263_ = ~pg35 & ng5260;
  assign new_n16264_ = ng5176 & new_n7580_1_;
  assign new_n16265_ = ng5212 & ~new_n16264_;
  assign new_n16266_ = ~new_n5966_ & new_n16264_;
  assign new_n16267_ = ~new_n16265_ & ~new_n16266_;
  assign new_n16268_ = pg35 & ~new_n16267_;
  assign n7178 = new_n16263_ | new_n16268_;
  assign new_n16270_ = ~pg35 & ng1825;
  assign new_n16271_ = new_n6683_ & new_n6805_;
  assign new_n16272_ = ng1830 & ~new_n16271_;
  assign new_n16273_ = ng1821 & ng1825;
  assign new_n16274_ = ng1825 & ~new_n16273_;
  assign new_n16275_ = ng1821 & ~new_n16273_;
  assign new_n16276_ = ~new_n16274_ & ~new_n16275_;
  assign new_n16277_ = new_n16271_ & ~new_n16276_;
  assign new_n16278_ = ~new_n16272_ & ~new_n16277_;
  assign new_n16279_ = pg35 & ~new_n16278_;
  assign n7183 = new_n16270_ | new_n16279_;
  assign new_n16281_ = ~pg35 & ng6466;
  assign new_n16282_ = ~ng6474 & ng6466;
  assign new_n16283_ = ng6474 & ~ng6466;
  assign new_n16284_ = ~new_n16282_ & ~new_n16283_;
  assign new_n16285_ = pg35 & ~new_n16284_;
  assign n7188 = new_n16281_ | new_n16285_;
  assign new_n16287_ = ~pg35 & ng4411;
  assign new_n16288_ = ~new_n7684_ & new_n11782_;
  assign new_n16289_ = ~new_n7685_ & ~new_n16288_;
  assign new_n16290_ = pg35 & ~new_n16289_;
  assign n7193 = new_n16287_ | new_n16290_;
  assign new_n16292_ = ~pg35 & ng3372;
  assign new_n16293_ = ~new_n10779_ & ~new_n10784_;
  assign new_n16294_ = ~ng3376 & ~new_n16293_;
  assign new_n16295_ = ng3376 & new_n8400_;
  assign new_n16296_ = new_n16293_ & new_n16295_;
  assign new_n16297_ = ~new_n16294_ & ~new_n16296_;
  assign new_n16298_ = pg35 & ~new_n16297_;
  assign n7198 = new_n16292_ | new_n16298_;
  assign new_n16300_ = ~pg35 & ng2984;
  assign new_n16301_ = n4955 & new_n9379_;
  assign new_n16302_ = ng2907 & ~new_n9379_;
  assign new_n16303_ = ~new_n16301_ & ~new_n16302_;
  assign new_n16304_ = pg35 & ~new_n16303_;
  assign n7203 = new_n16300_ | new_n16304_;
  assign new_n16306_ = ~pg35 & ng1061;
  assign new_n16307_ = ng1061 & ~ng1227;
  assign new_n16308_ = ~ng1052 & ng1227;
  assign new_n16309_ = ~ng1061 & new_n16308_;
  assign new_n16310_ = ~new_n16307_ & ~new_n16309_;
  assign new_n16311_ = ng1056 & ~new_n16310_;
  assign new_n16312_ = pg35 & ~new_n16311_;
  assign n7208 = new_n16306_ | new_n16312_;
  assign new_n16314_ = ~pg35 & ng2217;
  assign new_n16315_ = ng2185 & ~ng2208;
  assign new_n16316_ = ng2177 & new_n16315_;
  assign new_n16317_ = ~ng2185 & ~ng2217;
  assign new_n16318_ = ng2173 & new_n16317_;
  assign new_n16319_ = ng2181 & new_n5213_;
  assign new_n16320_ = ~new_n16316_ & ~new_n16318_;
  assign new_n16321_ = ~new_n16319_ & new_n16320_;
  assign new_n16322_ = ng2161 & new_n11373_;
  assign new_n16323_ = ng2165 & new_n9530_;
  assign new_n16324_ = ng2169 & new_n15367_;
  assign new_n16325_ = new_n16321_ & ~new_n16322_;
  assign new_n16326_ = ~new_n16323_ & ~new_n16324_;
  assign new_n16327_ = new_n16325_ & new_n16326_;
  assign new_n16328_ = new_n9534_ & ~new_n16327_;
  assign new_n16329_ = ng2236 & ~new_n9534_;
  assign new_n16330_ = ~new_n16328_ & ~new_n16329_;
  assign new_n16331_ = pg35 & ~new_n16330_;
  assign n7213 = new_n16314_ | new_n16331_;
  assign new_n16333_ = pg35 & ng5160;
  assign new_n16334_ = ~pg35 & new_n16333_;
  assign new_n16335_ = ng5654 & ~ng5630;
  assign new_n16336_ = ng5630 & ~ng5623;
  assign new_n16337_ = ~new_n16335_ & ~new_n16336_;
  assign new_n16338_ = ~new_n6327_ & new_n16337_;
  assign new_n16339_ = ng5666 & ~ng5637;
  assign new_n16340_ = ng5637 & ~ng5659;
  assign new_n16341_ = ~ng5666 & ng5623;
  assign new_n16342_ = new_n16338_ & ~new_n16339_;
  assign new_n16343_ = ~new_n16340_ & new_n16342_;
  assign new_n16344_ = ~new_n16341_ & new_n16343_;
  assign new_n16345_ = pg35 & new_n16344_;
  assign n7218 = new_n16334_ | new_n16345_;
  assign new_n16347_ = ~pg35 & ng6271;
  assign new_n16348_ = new_n6761_1_ & new_n9573_;
  assign new_n16349_ = ng6287 & ~new_n16348_;
  assign new_n16350_ = ~new_n5966_ & new_n16348_;
  assign new_n16351_ = ~new_n16349_ & ~new_n16350_;
  assign new_n16352_ = pg35 & ~new_n16351_;
  assign n7222 = new_n16347_ | new_n16352_;
  assign new_n16354_ = ~pg35 & ng5176;
  assign new_n16355_ = ng5180 & ~new_n7369_1_;
  assign new_n16356_ = ~ng5176 & new_n16355_;
  assign new_n16357_ = ~ng5180 & ~new_n7369_1_;
  assign new_n16358_ = ng5176 & new_n16357_;
  assign new_n16359_ = ~new_n16356_ & ~new_n16358_;
  assign new_n16360_ = pg35 & ~new_n16359_;
  assign n7227 = new_n16354_ | new_n16360_;
  assign new_n16362_ = ~pg35 & ng914;
  assign new_n16363_ = ng1227 & ng918;
  assign new_n16364_ = ~new_n7078_ & new_n16363_;
  assign new_n16365_ = ~ng918 & new_n7078_;
  assign new_n16366_ = ~new_n16364_ & ~new_n16365_;
  assign new_n16367_ = pg35 & ~new_n16366_;
  assign n7232 = new_n16362_ | new_n16367_;
  assign new_n16369_ = ~pg35 & ng5929;
  assign new_n16370_ = new_n8432_ & new_n12340_;
  assign new_n16371_ = ng5945 & ~new_n16370_;
  assign new_n16372_ = ~new_n5966_ & new_n16370_;
  assign new_n16373_ = ~new_n16371_ & ~new_n16372_;
  assign new_n16374_ = pg35 & ~new_n16373_;
  assign n7237 = new_n16369_ | new_n16374_;
  assign new_n16376_ = ~pg35 & ng5511;
  assign new_n16377_ = ng5517 & ~new_n8302_;
  assign new_n16378_ = ~ng5511 & new_n16377_;
  assign new_n16379_ = ~ng5517 & ~new_n8302_;
  assign new_n16380_ = ng5511 & new_n16379_;
  assign new_n16381_ = ~new_n16378_ & ~new_n16380_;
  assign new_n16382_ = pg35 & ~new_n16381_;
  assign n7242 = new_n16376_ | new_n16382_;
  assign new_n16384_ = ~pg35 & ng4249;
  assign new_n16385_ = n2272 & new_n7806_;
  assign new_n16386_ = ng4245 & ~new_n7806_;
  assign new_n16387_ = ~new_n16385_ & ~new_n16386_;
  assign new_n16388_ = pg35 & ~new_n16387_;
  assign n7247 = new_n16384_ | new_n16388_;
  assign new_n16390_ = ~pg35 & ng2241;
  assign new_n16391_ = ng2246 & ~new_n6524_;
  assign new_n16392_ = ng2241 & new_n6524_;
  assign new_n16393_ = ~new_n16391_ & ~new_n16392_;
  assign new_n16394_ = pg35 & ~new_n16393_;
  assign n7252 = new_n16390_ | new_n16394_;
  assign new_n16396_ = ~pg35 & ng1917;
  assign new_n16397_ = ~new_n4724_ & new_n11333_;
  assign new_n16398_ = new_n8171_ & new_n16397_;
  assign new_n16399_ = ng110 & new_n9094_;
  assign new_n16400_ = ng110 & ~new_n16399_;
  assign new_n16401_ = new_n9094_ & ~new_n16399_;
  assign new_n16402_ = ~new_n16400_ & ~new_n16401_;
  assign new_n16403_ = new_n16398_ & ~new_n16402_;
  assign new_n16404_ = ng1932 & ~new_n16398_;
  assign new_n16405_ = ~new_n16403_ & ~new_n16404_;
  assign new_n16406_ = pg35 & ~new_n16405_;
  assign n7257 = new_n16396_ | new_n16406_;
  assign new_n16408_ = ~pg35 & ng1589;
  assign new_n16409_ = ng1576 & ~ng1426;
  assign new_n16410_ = ng1570 & ng1426;
  assign new_n16411_ = ~new_n16409_ & ~new_n16410_;
  assign new_n16412_ = pg35 & ~new_n16411_;
  assign n7262 = new_n16408_ | new_n16412_;
  assign new_n16414_ = ~pg35 & ng3925;
  assign new_n16415_ = new_n6874_ & new_n7125_;
  assign new_n16416_ = ng3941 & ~new_n16415_;
  assign new_n16417_ = ~new_n5966_ & new_n16415_;
  assign new_n16418_ = ~new_n16416_ & ~new_n16417_;
  assign new_n16419_ = pg35 & ~new_n16418_;
  assign n7266 = new_n16414_ | new_n16419_;
  assign new_n16421_ = ~pg35 & ng1736;
  assign new_n16422_ = ng1772 & ~ng1802;
  assign new_n16423_ = ~new_n6236_ & new_n16422_;
  assign new_n16424_ = ng1744 & ~new_n16423_;
  assign new_n16425_ = ~new_n10679_ & new_n16423_;
  assign new_n16426_ = ~new_n16424_ & ~new_n16425_;
  assign new_n16427_ = pg35 & ~new_n16426_;
  assign n7271 = new_n16421_ | new_n16427_;
  assign new_n16429_ = ~pg35 & ng3506;
  assign new_n16430_ = ng3512 & ~new_n9472_;
  assign new_n16431_ = ~ng3506 & new_n16430_;
  assign new_n16432_ = ~ng3512 & ~new_n9472_;
  assign new_n16433_ = ng3506 & new_n16432_;
  assign new_n16434_ = ~new_n16431_ & ~new_n16433_;
  assign new_n16435_ = pg35 & ~new_n16434_;
  assign n7276 = new_n16429_ | new_n16435_;
  assign new_n16437_ = ~pg35 & ng2652;
  assign new_n16438_ = new_n10306_ & new_n10923_;
  assign new_n16439_ = ng2657 & ~new_n16438_;
  assign new_n16440_ = ng2652 & ng2648;
  assign new_n16441_ = ng2652 & ~new_n16440_;
  assign new_n16442_ = ng2648 & ~new_n16440_;
  assign new_n16443_ = ~new_n16441_ & ~new_n16442_;
  assign new_n16444_ = new_n16438_ & ~new_n16443_;
  assign new_n16445_ = ~new_n16439_ & ~new_n16444_;
  assign new_n16446_ = pg35 & ~new_n16445_;
  assign n7284 = new_n16437_ | new_n16446_;
  assign new_n16448_ = ~pg35 & ng4939;
  assign new_n16449_ = ~new_n6055_1_ & ~new_n12050_;
  assign new_n16450_ = ng4939 & ~new_n6055_1_;
  assign new_n16451_ = ~new_n6058_ & ~new_n16450_;
  assign new_n16452_ = ~new_n16449_ & ~new_n16451_;
  assign new_n16453_ = ng4933 & new_n16449_;
  assign new_n16454_ = ~new_n16452_ & ~new_n16453_;
  assign new_n16455_ = pg35 & ~new_n16454_;
  assign n7289 = new_n16448_ | new_n16455_;
  assign new_n16457_ = ~pg35 & ng604;
  assign new_n16458_ = ~ng608 & new_n9116_;
  assign new_n16459_ = ng608 & ~new_n6545_;
  assign new_n16460_ = ~new_n9116_ & new_n16459_;
  assign new_n16461_ = ~new_n16458_ & ~new_n16460_;
  assign new_n16462_ = pg35 & ~new_n16461_;
  assign n7294 = new_n16457_ | new_n16462_;
  assign new_n16464_ = ~pg35 & ng5774;
  assign new_n16465_ = ng5774 & ~ng5782;
  assign new_n16466_ = ~ng5774 & ng5782;
  assign new_n16467_ = ~new_n16465_ & ~new_n16466_;
  assign new_n16468_ = pg35 & ~new_n16467_;
  assign n7299 = new_n16464_ | new_n16468_;
  assign new_n16470_ = ~pg35 & ng1890;
  assign new_n16471_ = ~new_n6667_1_ & new_n10118_;
  assign new_n16472_ = ng1886 & ~new_n16471_;
  assign new_n16473_ = ~new_n6674_ & new_n16471_;
  assign new_n16474_ = ~new_n16472_ & ~new_n16473_;
  assign new_n16475_ = pg35 & ~new_n16474_;
  assign n7304 = new_n16470_ | new_n16475_;
  assign new_n16477_ = ~pg35 & ng969;
  assign new_n16478_ = ng1008 & new_n5940_1_;
  assign new_n16479_ = ng1008 & ~new_n6132_;
  assign new_n16480_ = new_n5939_ & new_n16479_;
  assign new_n16481_ = ng969 & ~new_n5939_;
  assign new_n16482_ = ng1008 & ~new_n5939_;
  assign new_n16483_ = ~ng1046 & ~new_n6132_;
  assign new_n16484_ = new_n16482_ & new_n16483_;
  assign new_n16485_ = ~new_n16480_ & ~new_n16481_;
  assign new_n16486_ = ~new_n16484_ & new_n16485_;
  assign new_n16487_ = ~new_n5940_1_ & ~new_n16486_;
  assign new_n16488_ = ~new_n16478_ & ~new_n16487_;
  assign new_n16489_ = pg35 & ~new_n16488_;
  assign n7309 = new_n16477_ | new_n16489_;
  assign new_n16491_ = pg35 & ng723;
  assign new_n16492_ = ~pg35 & new_n16491_;
  assign new_n16493_ = ng645 & ~new_n7858_;
  assign new_n16494_ = ng446 & new_n7858_;
  assign new_n16495_ = ~new_n16493_ & ~new_n16494_;
  assign new_n16496_ = pg35 & ~new_n16495_;
  assign n7314 = new_n16492_ | new_n16496_;
  assign new_n16498_ = ~pg35 & ng401;
  assign new_n16499_ = ng392 & ~new_n6067_;
  assign new_n16500_ = ~ng703 & ng854;
  assign new_n16501_ = new_n6067_ & new_n16500_;
  assign new_n16502_ = ~new_n16499_ & ~new_n16501_;
  assign new_n16503_ = pg35 & ~new_n16502_;
  assign n7319 = new_n16498_ | new_n16503_;
  assign new_n16505_ = ~pg35 & ng142;
  assign new_n16506_ = ng146 & new_n6276_;
  assign new_n16507_ = ~new_n6271_ & new_n16506_;
  assign new_n16508_ = ~ng146 & new_n6276_;
  assign new_n16509_ = new_n6271_ & new_n16508_;
  assign new_n16510_ = ~new_n16507_ & ~new_n16509_;
  assign new_n16511_ = pg35 & ~new_n16510_;
  assign n7324 = new_n16505_ | new_n16511_;
  assign new_n16513_ = ~pg35 & ng2667;
  assign new_n16514_ = ng2671 & ~new_n13235_;
  assign new_n16515_ = ng2661 & ~ng2667;
  assign new_n16516_ = ng2661 & ~new_n16515_;
  assign new_n16517_ = ~ng2667 & ~new_n16515_;
  assign new_n16518_ = ~new_n16516_ & ~new_n16517_;
  assign new_n16519_ = new_n13235_ & ~new_n16518_;
  assign new_n16520_ = ~new_n16514_ & ~new_n16519_;
  assign new_n16521_ = pg35 & ~new_n16520_;
  assign n7329 = new_n16513_ | new_n16521_;
  assign new_n16523_ = ~pg35 & ng6561;
  assign new_n16524_ = ng6565 & ~new_n8536_;
  assign new_n16525_ = ~ng6561 & new_n16524_;
  assign new_n16526_ = ~ng6565 & ~new_n8536_;
  assign new_n16527_ = ng6561 & new_n16526_;
  assign new_n16528_ = ~new_n16525_ & ~new_n16527_;
  assign new_n16529_ = pg35 & ~new_n16528_;
  assign n7334 = new_n16523_ | new_n16529_;
  assign new_n16531_ = ~pg35 & ng5913;
  assign new_n16532_ = new_n7997_ & new_n8432_;
  assign new_n16533_ = ng5909 & ~new_n16532_;
  assign new_n16534_ = ~new_n5966_ & new_n16532_;
  assign new_n16535_ = ~new_n16533_ & ~new_n16534_;
  assign new_n16536_ = pg35 & ~new_n16535_;
  assign n7339 = new_n16531_ | new_n16536_;
  assign new_n16538_ = ~pg35 & ng4366;
  assign new_n16539_ = ~ng4340 & new_n8691_;
  assign new_n16540_ = ~ng4340 & ~new_n16539_;
  assign new_n16541_ = ng4349 & new_n16540_;
  assign new_n16542_ = ~ng4349 & ~new_n16539_;
  assign new_n16543_ = ~new_n16541_ & ~new_n16542_;
  assign new_n16544_ = ng4358 & new_n16543_;
  assign new_n16545_ = ng4349 & ~new_n16539_;
  assign new_n16546_ = ~ng4322 & ~new_n5614_;
  assign new_n16547_ = ng4332 & new_n16546_;
  assign new_n16548_ = ~pg73 & ng4515;
  assign new_n16549_ = ~pg72 & new_n16548_;
  assign new_n16550_ = ng4311 & ~new_n16549_;
  assign new_n16551_ = ~ng4311 & ~new_n16549_;
  assign new_n16552_ = ~new_n16550_ & ~new_n16551_;
  assign new_n16553_ = ng4322 & new_n16552_;
  assign new_n16554_ = pg90 & ~ng2994;
  assign new_n16555_ = ~pg73 & ~new_n16554_;
  assign new_n16556_ = ~pg72 & new_n16555_;
  assign new_n16557_ = ng4311 & ~new_n16556_;
  assign new_n16558_ = ~ng4311 & ~new_n16556_;
  assign new_n16559_ = ~new_n16557_ & ~new_n16558_;
  assign new_n16560_ = ~ng4322 & new_n16559_;
  assign new_n16561_ = ~new_n16553_ & ~new_n16560_;
  assign new_n16562_ = ~ng4332 & new_n16561_;
  assign new_n16563_ = ~new_n16547_ & ~new_n16562_;
  assign new_n16564_ = ~ng4340 & ~new_n16563_;
  assign new_n16565_ = ~ng4340 & ~new_n16564_;
  assign new_n16566_ = ~ng4349 & new_n16565_;
  assign new_n16567_ = ~new_n16545_ & ~new_n16566_;
  assign new_n16568_ = ~ng4358 & new_n16567_;
  assign new_n16569_ = ~new_n16544_ & ~new_n16568_;
  assign new_n16570_ = pg35 & ~new_n16569_;
  assign n7344 = new_n16538_ | new_n16570_;
  assign new_n16572_ = pg35 & ng3089;
  assign new_n16573_ = ~pg35 & new_n16572_;
  assign new_n16574_ = ~ng3167 & ~new_n6249_;
  assign new_n16575_ = ~ng3155 & new_n16574_;
  assign new_n16576_ = pg35 & new_n16575_;
  assign n7349 = new_n16573_ | new_n16576_;
  assign new_n16578_ = ~pg35 & ng5591;
  assign new_n16579_ = new_n8129_ & new_n10861_;
  assign new_n16580_ = ng5607 & ~new_n16579_;
  assign new_n16581_ = ~new_n5966_ & new_n16579_;
  assign new_n16582_ = ~new_n16580_ & ~new_n16581_;
  assign new_n16583_ = pg35 & ~new_n16582_;
  assign n7354 = new_n16578_ | new_n16583_;
  assign new_n16585_ = ~pg35 & ng4512;
  assign new_n16586_ = ng4531 & ng4581;
  assign new_n16587_ = pg35 & ~new_n16586_;
  assign n7359 = new_n16585_ | new_n16587_;
  assign new_n16589_ = ~pg35 & ng559;
  assign new_n16590_ = ng626 & ng632;
  assign new_n16591_ = ~new_n6545_ & ~new_n16590_;
  assign new_n16592_ = ~ng562 & new_n16591_;
  assign new_n16593_ = new_n6544_ & new_n16592_;
  assign new_n16594_ = ng562 & new_n16591_;
  assign new_n16595_ = ~new_n6544_ & new_n16594_;
  assign new_n16596_ = ~new_n16593_ & ~new_n16595_;
  assign new_n16597_ = pg35 & ~new_n16596_;
  assign n7364 = new_n16589_ | new_n16597_;
  assign new_n16599_ = ~pg35 & ng6093;
  assign new_n16600_ = ~new_n7512_ & ~new_n7520_;
  assign new_n16601_ = pg35 & new_n16600_;
  assign n7369 = new_n16599_ | new_n16601_;
  assign new_n16603_ = ~pg35 & ng6462;
  assign new_n16604_ = ~ng6462 & ~new_n14549_;
  assign new_n16605_ = ~ng6466 & new_n16604_;
  assign new_n16606_ = ng6462 & ng6466;
  assign new_n16607_ = ~new_n16605_ & ~new_n16606_;
  assign new_n16608_ = ~new_n14551_ & new_n16607_;
  assign new_n16609_ = pg35 & ~new_n16608_;
  assign n7374 = new_n16603_ | new_n16609_;
  assign new_n16611_ = ~pg35 & ng6128;
  assign new_n16612_ = ng6133 & ~new_n15157_;
  assign new_n16613_ = ~ng6133 & new_n15157_;
  assign new_n16614_ = ~new_n16612_ & ~new_n16613_;
  assign new_n16615_ = pg35 & ~new_n16614_;
  assign n7379 = new_n16611_ | new_n16615_;
  assign new_n16617_ = ~pg35 & ng3574;
  assign new_n16618_ = new_n7039_ & new_n10352_;
  assign new_n16619_ = ng3590 & ~new_n16618_;
  assign new_n16620_ = ~new_n5966_ & new_n16618_;
  assign new_n16621_ = ~new_n16619_ & ~new_n16620_;
  assign new_n16622_ = pg35 & ~new_n16621_;
  assign n7388 = new_n16617_ | new_n16622_;
  assign new_n16624_ = ~pg35 & ng2036;
  assign new_n16625_ = ~ng2060 & ng2028;
  assign new_n16626_ = ~ng2051 & ~ng2060;
  assign new_n16627_ = ~new_n16625_ & ~new_n16626_;
  assign new_n16628_ = ~new_n13378_ & new_n16627_;
  assign new_n16629_ = new_n9143_ & ~new_n16628_;
  assign new_n16630_ = ng2028 & ~new_n9143_;
  assign new_n16631_ = ~new_n16629_ & ~new_n16630_;
  assign new_n16632_ = pg35 & ~new_n16631_;
  assign n7397 = new_n16624_ | new_n16632_;
  assign new_n16634_ = ~pg35 & ng2681;
  assign new_n16635_ = ng2685 & ~new_n13437_;
  assign new_n16636_ = ng2675 & ~ng2681;
  assign new_n16637_ = ng2675 & ~new_n16636_;
  assign new_n16638_ = ~ng2681 & ~new_n16636_;
  assign new_n16639_ = ~new_n16637_ & ~new_n16638_;
  assign new_n16640_ = new_n13437_ & ~new_n16639_;
  assign new_n16641_ = ~new_n16635_ & ~new_n16640_;
  assign new_n16642_ = pg35 & ~new_n16641_;
  assign n7402 = new_n16634_ | new_n16642_;
  assign new_n16644_ = ~pg35 & ng1772;
  assign new_n16645_ = ng1772 & ~new_n6239_;
  assign new_n16646_ = ~new_n6236_ & new_n16645_;
  assign new_n16647_ = ng1802 & new_n6236_;
  assign new_n16648_ = ~new_n16646_ & ~new_n16647_;
  assign new_n16649_ = pg35 & ~new_n16648_;
  assign n7407 = new_n16644_ | new_n16649_;
  assign new_n16651_ = ~pg35 & ng3484;
  assign new_n16652_ = ng3490 & ~new_n6770_;
  assign new_n16653_ = ng3484 & new_n6770_;
  assign new_n16654_ = ~new_n16652_ & ~new_n16653_;
  assign new_n16655_ = pg35 & ~new_n16654_;
  assign n7412 = new_n16651_ | new_n16655_;
  assign new_n16657_ = ~pg35 & ng3161;
  assign new_n16658_ = new_n9338_ & new_n16574_;
  assign new_n16659_ = ng3167 & new_n16574_;
  assign new_n16660_ = ~new_n9338_ & new_n16659_;
  assign new_n16661_ = ~new_n16658_ & ~new_n16660_;
  assign new_n16662_ = pg35 & ~new_n16661_;
  assign n7417 = new_n16657_ | new_n16662_;
  assign new_n16664_ = ~pg35 & ng2299;
  assign new_n16665_ = ng2287 & ~ng2331;
  assign new_n16666_ = ~new_n7886_ & new_n16665_;
  assign new_n16667_ = ng2295 & ~new_n16666_;
  assign new_n16668_ = ~new_n8906_ & new_n16666_;
  assign new_n16669_ = ~new_n16667_ & ~new_n16668_;
  assign new_n16670_ = pg35 & ~new_n16669_;
  assign n7422 = new_n16664_ | new_n16670_;
  assign new_n16672_ = ~pg35 & ng3849;
  assign new_n16673_ = ng3813 & ~new_n7011_1_;
  assign new_n16674_ = ng3849 & new_n7011_1_;
  assign new_n16675_ = ~new_n16673_ & ~new_n16674_;
  assign new_n16676_ = pg35 & ~new_n16675_;
  assign n7430 = new_n16672_ | new_n16676_;
  assign new_n16678_ = ~pg35 & ng1087;
  assign new_n16679_ = ng1087 & ~ng1205;
  assign new_n16680_ = ~ng1087 & ng1205;
  assign new_n16681_ = ~new_n16679_ & ~new_n16680_;
  assign new_n16682_ = pg35 & ~new_n16681_;
  assign n7435 = new_n16678_ | new_n16682_;
  assign new_n16684_ = ~pg35 & ng2185;
  assign new_n16685_ = ~ng2185 & ~new_n11142_;
  assign new_n16686_ = new_n9534_ & ~new_n16685_;
  assign new_n16687_ = ng2208 & ~new_n9534_;
  assign new_n16688_ = ~new_n16686_ & ~new_n16687_;
  assign new_n16689_ = pg35 & ~new_n16688_;
  assign n7440 = new_n16684_ | new_n16689_;
  assign new_n16691_ = ~pg35 & new_n6882_;
  assign new_n16692_ = ng732 & ~new_n5996_;
  assign new_n16693_ = ng246 & ng269;
  assign new_n16694_ = ng246 & ~new_n16693_;
  assign new_n16695_ = ng269 & ~new_n16693_;
  assign new_n16696_ = ~new_n16694_ & ~new_n16695_;
  assign new_n16697_ = ng262 & ng239;
  assign new_n16698_ = ng239 & ~new_n16697_;
  assign new_n16699_ = ng262 & ~new_n16697_;
  assign new_n16700_ = ~new_n16698_ & ~new_n16699_;
  assign new_n16701_ = ~new_n16696_ & ~new_n16700_;
  assign new_n16702_ = ~new_n16696_ & ~new_n16701_;
  assign new_n16703_ = ~new_n16700_ & ~new_n16701_;
  assign new_n16704_ = ~new_n16702_ & ~new_n16703_;
  assign new_n16705_ = ng232 & ng255;
  assign new_n16706_ = ng232 & ~new_n16705_;
  assign new_n16707_ = ng255 & ~new_n16705_;
  assign new_n16708_ = ~new_n16706_ & ~new_n16707_;
  assign new_n16709_ = ng225 & ~new_n16708_;
  assign new_n16710_ = ~new_n16708_ & ~new_n16709_;
  assign new_n16711_ = ng225 & ~new_n16709_;
  assign new_n16712_ = ~new_n16710_ & ~new_n16711_;
  assign new_n16713_ = ~new_n16704_ & ~new_n16712_;
  assign new_n16714_ = ~new_n16704_ & ~new_n16713_;
  assign new_n16715_ = ~new_n16712_ & ~new_n16713_;
  assign new_n16716_ = ~new_n16714_ & ~new_n16715_;
  assign new_n16717_ = new_n16692_ & ~new_n16716_;
  assign new_n16718_ = new_n16692_ & ~new_n16717_;
  assign new_n16719_ = ~new_n16716_ & ~new_n16717_;
  assign new_n16720_ = ~new_n16718_ & ~new_n16719_;
  assign new_n16721_ = pg35 & ~new_n16720_;
  assign n7445 = new_n16691_ | new_n16721_;
  assign n7450 = ~pg35 & ng967;
  assign new_n16724_ = ~pg35 & ng4172;
  assign new_n16725_ = new_n4927_ & new_n14357_;
  assign new_n16726_ = ~ng4072 & ~ng4176;
  assign new_n16727_ = ~new_n16725_ & ~new_n16726_;
  assign new_n16728_ = pg35 & new_n16727_;
  assign n7455 = new_n16724_ | new_n16728_;
  assign new_n16730_ = ~pg35 & ng6235;
  assign new_n16731_ = new_n7866_ & new_n9572_;
  assign new_n16732_ = ng6263 & ~new_n16731_;
  assign new_n16733_ = ~new_n5966_ & new_n16731_;
  assign new_n16734_ = ~new_n16732_ & ~new_n16733_;
  assign new_n16735_ = pg35 & ~new_n16734_;
  assign n7460 = new_n16730_ | new_n16735_;
  assign new_n16737_ = ~pg35 & ng4423;
  assign new_n16738_ = ~ng4575 & new_n15437_;
  assign new_n16739_ = ng4581 & ~new_n16738_;
  assign new_n16740_ = ~new_n15440_ & ~new_n16739_;
  assign new_n16741_ = pg35 & ~new_n16740_;
  assign n7465 = new_n16737_ | new_n16741_;
  assign new_n16743_ = ~pg35 & ng2831;
  assign n7470 = new_n11073_ | new_n16743_;
  assign new_n16745_ = ~pg35 & ng6727;
  assign new_n16746_ = ~ng6736 & ~new_n9677_;
  assign new_n16747_ = pg35 & new_n16746_;
  assign n7475 = new_n16745_ | new_n16747_;
  assign new_n16749_ = ~pg35 & ng3602;
  assign new_n16750_ = ng3518 & new_n7038_;
  assign new_n16751_ = ng3554 & ~new_n16750_;
  assign new_n16752_ = ~new_n5966_ & new_n16750_;
  assign new_n16753_ = ~new_n16751_ & ~new_n16752_;
  assign new_n16754_ = pg35 & ~new_n16753_;
  assign n7480 = new_n16749_ | new_n16754_;
  assign new_n16756_ = ~pg35 & ng744;
  assign new_n16757_ = ng749 & ~new_n6578_;
  assign new_n16758_ = ~new_n6582_ & new_n16757_;
  assign new_n16759_ = ~ng749 & new_n6582_;
  assign new_n16760_ = ~new_n16758_ & ~new_n16759_;
  assign new_n16761_ = pg35 & ~new_n16760_;
  assign n7485 = new_n16756_ | new_n16761_;
  assign new_n16763_ = ~pg35 & ng5599;
  assign new_n16764_ = new_n6885_ & new_n10861_;
  assign new_n16765_ = ng5615 & ~new_n16764_;
  assign new_n16766_ = ~new_n5966_ & new_n16764_;
  assign new_n16767_ = ~new_n16765_ & ~new_n16766_;
  assign new_n16768_ = pg35 & ~new_n16767_;
  assign n7490 = new_n16763_ | new_n16768_;
  assign new_n16770_ = pg35 & ng6191;
  assign new_n16771_ = ~pg35 & new_n16770_;
  assign new_n16772_ = n4955 & new_n6181_;
  assign new_n16773_ = ng6199 & ~new_n6181_;
  assign new_n16774_ = ~new_n16772_ & ~new_n16773_;
  assign new_n16775_ = pg35 & ~new_n16774_;
  assign n7495 = new_n16771_ | new_n16775_;
  assign new_n16777_ = ~pg35 & ng2084;
  assign new_n16778_ = ng2089 & ~new_n8022_;
  assign new_n16779_ = ng2084 & new_n8022_;
  assign new_n16780_ = ~new_n16778_ & ~new_n16779_;
  assign new_n16781_ = pg35 & ~new_n16780_;
  assign n7500 = new_n16777_ | new_n16781_;
  assign new_n16783_ = ~pg35 & ng6098;
  assign new_n16784_ = pg35 & ng6381;
  assign n7505 = new_n16783_ | new_n16784_;
  assign new_n16786_ = ~pg35 & ng3913;
  assign new_n16787_ = new_n6896_ & new_n7010_;
  assign new_n16788_ = ng3909 & ~new_n16787_;
  assign new_n16789_ = ~new_n5966_ & new_n16787_;
  assign new_n16790_ = ~new_n16788_ & ~new_n16789_;
  assign new_n16791_ = pg35 & ~new_n16790_;
  assign n7509 = new_n16786_ | new_n16791_;
  assign new_n16793_ = ~pg35 & ng2902;
  assign new_n16794_ = new_n4937_ & new_n9347_;
  assign new_n16795_ = ~ng2917 & new_n4694_;
  assign new_n16796_ = ~new_n16794_ & ~new_n16795_;
  assign new_n16797_ = pg35 & new_n16796_;
  assign n7514 = new_n16793_ | new_n16797_;
  assign new_n16799_ = ~pg35 & ng2485;
  assign new_n16800_ = ~ng2476 & ng2453;
  assign new_n16801_ = ng2445 & new_n16800_;
  assign new_n16802_ = ~ng2485 & ~ng2453;
  assign new_n16803_ = ng2441 & new_n16802_;
  assign new_n16804_ = ng2449 & new_n5215_;
  assign new_n16805_ = ~new_n16801_ & ~new_n16803_;
  assign new_n16806_ = ~new_n16804_ & new_n16805_;
  assign new_n16807_ = ng2429 & new_n12735_;
  assign new_n16808_ = ng2433 & new_n9420_;
  assign new_n16809_ = ng2437 & new_n11152_;
  assign new_n16810_ = new_n16806_ & ~new_n16807_;
  assign new_n16811_ = ~new_n16808_ & ~new_n16809_;
  assign new_n16812_ = new_n16810_ & new_n16811_;
  assign new_n16813_ = new_n5907_1_ & ~new_n16812_;
  assign new_n16814_ = ng2504 & ~new_n5907_1_;
  assign new_n16815_ = ~new_n16813_ & ~new_n16814_;
  assign new_n16816_ = pg35 & ~new_n16815_;
  assign n7519 = new_n16799_ | new_n16816_;
  assign new_n16818_ = ~pg35 & ng6088;
  assign new_n16819_ = ~ng6088 & new_n15902_;
  assign new_n16820_ = ng6088 & new_n15903_;
  assign new_n16821_ = ~new_n16819_ & ~new_n16820_;
  assign new_n16822_ = ~ng6093 & ~new_n16821_;
  assign new_n16823_ = ng6093 & new_n7527_;
  assign new_n16824_ = new_n16821_ & new_n16823_;
  assign new_n16825_ = ~new_n16822_ & ~new_n16824_;
  assign new_n16826_ = pg35 & ~new_n16825_;
  assign n7524 = new_n16818_ | new_n16826_;
  assign new_n16828_ = pg35 & ng3502;
  assign new_n16829_ = ~pg35 & new_n16828_;
  assign new_n16830_ = ~ng3976 & ng4000;
  assign new_n16831_ = ng3976 & ~ng3969;
  assign new_n16832_ = ~new_n16830_ & ~new_n16831_;
  assign new_n16833_ = ~new_n6172_ & new_n16832_;
  assign new_n16834_ = ~ng3983 & ng4012;
  assign new_n16835_ = ng3983 & ~ng4005;
  assign new_n16836_ = ~ng4012 & ng3969;
  assign new_n16837_ = new_n16833_ & ~new_n16834_;
  assign new_n16838_ = ~new_n16835_ & new_n16837_;
  assign new_n16839_ = ~new_n16836_ & new_n16838_;
  assign new_n16840_ = pg35 & new_n16839_;
  assign n7529 = new_n16829_ | new_n16840_;
  assign new_n16842_ = ~pg35 & ng2338;
  assign new_n16843_ = ng2287 & ~new_n11285_;
  assign new_n16844_ = ~new_n7886_ & new_n16843_;
  assign new_n16845_ = ng2331 & new_n7886_;
  assign new_n16846_ = ~new_n16844_ & ~new_n16845_;
  assign new_n16847_ = pg35 & ~new_n16846_;
  assign n7533 = new_n16842_ | new_n16847_;
  assign new_n16849_ = ~pg35 & ng6589;
  assign new_n16850_ = new_n6336_ & new_n7456_;
  assign new_n16851_ = ng6585 & ~new_n16850_;
  assign new_n16852_ = ~new_n5966_ & new_n16850_;
  assign new_n16853_ = ~new_n16851_ & ~new_n16852_;
  assign new_n16854_ = pg35 & ~new_n16853_;
  assign n7542 = new_n16849_ | new_n16854_;
  assign new_n16856_ = ~pg35 & ng6617;
  assign new_n16857_ = new_n6334_ & new_n12232_;
  assign new_n16858_ = ng6633 & ~new_n16857_;
  assign new_n16859_ = ~new_n5966_ & new_n16857_;
  assign new_n16860_ = ~new_n16858_ & ~new_n16859_;
  assign new_n16861_ = pg35 & ~new_n16860_;
  assign n7547 = new_n16856_ | new_n16861_;
  assign new_n16863_ = ~pg35 & ng6065;
  assign new_n16864_ = ~new_n10186_ & ~new_n10190_;
  assign new_n16865_ = ng6069 & new_n7527_;
  assign new_n16866_ = new_n16864_ & new_n16865_;
  assign new_n16867_ = ~ng6069 & ~new_n16864_;
  assign new_n16868_ = ~new_n16866_ & ~new_n16867_;
  assign new_n16869_ = pg35 & ~new_n16868_;
  assign n7556 = new_n16863_ | new_n16869_;
  assign new_n16871_ = ~pg35 & ng4543;
  assign new_n16872_ = ~ng4575 & new_n7110_;
  assign new_n16873_ = ng4581 & ~new_n16872_;
  assign new_n16874_ = ng4543 & ~ng4581;
  assign new_n16875_ = ~new_n16873_ & ~new_n16874_;
  assign new_n16876_ = pg35 & ~new_n16875_;
  assign n7561 = new_n16871_ | new_n16876_;
  assign new_n16878_ = ~pg35 & ng1579;
  assign n7566 = new_n12610_ | new_n16878_;
  assign new_n16880_ = ~pg35 & ng763;
  assign new_n16881_ = ~ng767 & new_n6588_;
  assign new_n16882_ = ng767 & ~new_n6578_;
  assign new_n16883_ = ~new_n6588_ & new_n16882_;
  assign new_n16884_ = ~new_n16881_ & ~new_n16883_;
  assign new_n16885_ = pg35 & ~new_n16884_;
  assign n7571 = new_n16880_ | new_n16885_;
  assign new_n16887_ = pg35 & ng5990;
  assign new_n16888_ = ~pg35 & new_n16887_;
  assign new_n16889_ = pg35 & ng5881;
  assign n7576 = new_n16888_ | new_n16889_;
  assign new_n16891_ = ~pg35 & ng6303;
  assign new_n16892_ = ng6215 & new_n6761_1_;
  assign new_n16893_ = ng6259 & ~new_n16892_;
  assign new_n16894_ = ~new_n5966_ & new_n16892_;
  assign new_n16895_ = ~new_n16893_ & ~new_n16894_;
  assign new_n16896_ = pg35 & ~new_n16895_;
  assign n7580 = new_n16891_ | new_n16896_;
  assign new_n16898_ = ~pg35 & ng3929;
  assign new_n16899_ = new_n7010_ & new_n7125_;
  assign new_n16900_ = ng3945 & ~new_n16899_;
  assign new_n16901_ = ~new_n5966_ & new_n16899_;
  assign new_n16902_ = ~new_n16900_ & ~new_n16901_;
  assign new_n16903_ = pg35 & ~new_n16902_;
  assign n7589 = new_n16898_ | new_n16903_;
  assign new_n16905_ = ~pg35 & ng2741;
  assign new_n16906_ = ng2748 & ~new_n6643_;
  assign new_n16907_ = ~ng2748 & new_n6643_;
  assign new_n16908_ = ~new_n16906_ & ~new_n16907_;
  assign new_n16909_ = ng2841 & ~new_n16908_;
  assign new_n16910_ = pg35 & new_n16909_;
  assign n7594 = new_n16905_ | new_n16910_;
  assign new_n16912_ = ~pg35 & ng2279;
  assign new_n16913_ = ng2283 & ~new_n9535_;
  assign new_n16914_ = ~ng2279 & ng2273;
  assign new_n16915_ = ng2273 & ~new_n16914_;
  assign new_n16916_ = ~ng2279 & ~new_n16914_;
  assign new_n16917_ = ~new_n16915_ & ~new_n16916_;
  assign new_n16918_ = new_n9535_ & ~new_n16917_;
  assign new_n16919_ = ~new_n16913_ & ~new_n16918_;
  assign new_n16920_ = pg35 & ~new_n16919_;
  assign n7599 = new_n16912_ | new_n16920_;
  assign new_n16922_ = ~pg35 & ng3694;
  assign new_n16923_ = ng3694 & ~new_n11673_;
  assign new_n16924_ = pg35 & new_n16923_;
  assign n7607 = new_n16922_ | new_n16924_;
  assign new_n16926_ = ~pg35 & ng305;
  assign new_n16927_ = pg6744 & pg35;
  assign n7612 = new_n16926_ | new_n16927_;
  assign new_n16929_ = ~pg35 & ng3045;
  assign new_n16930_ = ~new_n8939_ & ~new_n8947_;
  assign new_n16931_ = pg35 & new_n16930_;
  assign n7617 = new_n16929_ | new_n16931_;
  assign new_n16933_ = ~pg35 & ng1379;
  assign new_n16934_ = ng1384 & ~new_n11363_;
  assign new_n16935_ = new_n11363_ & new_n11364_;
  assign new_n16936_ = ~new_n16934_ & ~new_n16935_;
  assign new_n16937_ = pg35 & ~new_n16936_;
  assign n7622 = new_n16933_ | new_n16937_;
  assign new_n16939_ = pg35 & ng5845;
  assign new_n16940_ = ~pg35 & new_n16939_;
  assign new_n16941_ = n3583 & new_n6181_;
  assign new_n16942_ = ng5853 & ~new_n6181_;
  assign new_n16943_ = ~new_n16941_ & ~new_n16942_;
  assign new_n16944_ = pg35 & ~new_n16943_;
  assign n7627 = new_n16940_ | new_n16944_;
  assign new_n16946_ = ~pg35 & ng5607;
  assign new_n16947_ = ng5523 & new_n8129_;
  assign new_n16948_ = ng5559 & ~new_n16947_;
  assign new_n16949_ = ~new_n5966_ & new_n16947_;
  assign new_n16950_ = ~new_n16948_ & ~new_n16949_;
  assign new_n16951_ = pg35 & ~new_n16950_;
  assign n7632 = new_n16946_ | new_n16951_;
  assign new_n16953_ = ~pg35 & ng5953;
  assign new_n16954_ = ng5869 & new_n7649_;
  assign new_n16955_ = ng5905 & ~new_n16954_;
  assign new_n16956_ = ~new_n5966_ & new_n16954_;
  assign new_n16957_ = ~new_n16955_ & ~new_n16956_;
  assign new_n16958_ = pg35 & ~new_n16957_;
  assign n7637 = new_n16953_ | new_n16958_;
  assign new_n16960_ = ng22 & pg34925;
  assign new_n16961_ = ~ng22 & n4465;
  assign n7646 = new_n16960_ | new_n16961_;
  assign new_n16963_ = ~pg35 & ng5462;
  assign new_n16964_ = ng5471 & ~new_n8548_;
  assign new_n16965_ = ng5462 & ng5467;
  assign new_n16966_ = ng5467 & ~new_n16965_;
  assign new_n16967_ = ng5462 & ~new_n16965_;
  assign new_n16968_ = ~new_n16966_ & ~new_n16967_;
  assign new_n16969_ = new_n8548_ & ~new_n16968_;
  assign new_n16970_ = ~new_n16964_ & ~new_n16969_;
  assign new_n16971_ = pg35 & ~new_n16970_;
  assign n7651 = new_n16963_ | new_n16971_;
  assign new_n16973_ = ~pg35 & ng2161;
  assign new_n16974_ = ng2197 & ~ng2227;
  assign new_n16975_ = ~new_n6522_ & new_n16974_;
  assign new_n16976_ = ng2169 & ~new_n16975_;
  assign new_n16977_ = ~new_n6725_ & new_n16975_;
  assign new_n16978_ = ~new_n16976_ & ~new_n16977_;
  assign new_n16979_ = pg35 & ~new_n16978_;
  assign n7656 = new_n16973_ | new_n16979_;
  assign pg32454 = 1'b1;
  assign pg34597 = 1'b0;
  assign pg24151 = 1'b1;
  assign pg34232 = 1'b1;
  assign pg25583 = 1'b1;
  assign pg33948 = 1'b1;
  assign pg25584 = 1'b1;
  assign pg33949 = 1'b1;
  assign pg25585 = 1'b1;
  assign pg33946 = 1'b1;
  assign pg25586 = 1'b1;
  assign pg33947 = 1'b1;
  assign pg25590 = 1'b1;
  assign pg33945 = 1'b1;
  assign pg25582 = 1'b1;
  assign pg33950 = 1'b1;
  assign pg32429 = 1'b1;
  assign pg25587 = 1'b1;
  assign pg25588 = 1'b1;
  assign pg25589 = 1'b1;
  assign n4279 = 1'b0;
  assign pg30327 = ~ng37;
  assign pg30329 = ~ng136;
  assign pg12833 = ~pg5;
  assign pg23652 = ~ng2834;
  assign pg30331 = ~ng2831;
  assign pg8342 = ng3447;
  assign pg8353 = ng4815;
  assign pg8870 = ng4222;
  assign pg9048 = ng640;
  assign pg9741 = ng6144;
  assign pg13272 = ng1459;
  assign pg13906 = ng4023;
  assign pg8132 = ng4809;
  assign pg8783 = ng4188;
  assign pg9555 = ng5448;
  assign pg12184 = ng799;
  assign pg13068 = ng6000;
  assign pg13099 = ng6692;
  assign pg7260 = ng4449;
  assign pg8344 = ng3794;
  assign pg8784 = ng4194;
  assign pg14167 = ng887;
  assign pg17320 = ng1418;
  assign pg18101 = pg6746;
  assign pg34435 = pg31521;
  assign pg8398 = ng3798;
  assign pg8785 = ng4197;
  assign pg18100 = pg6751;
  assign pg20899 = ng79;
  assign pg8786 = ng4200;
  assign pg14828 = ng6675;
  assign pg20557 = ng86;
  assign pg20654 = ng121;
  assign pg24171 = pg92;
  assign pg24182 = pg127;
  assign pg7243 = ng4408;
  assign pg7540 = ng344;
  assign pg8235 = ng4812;
  assign pg8787 = ng4204;
  assign pg12470 = ng6697;
  assign pg17819 = ng6019;
  assign pg19334 = ng1056;
  assign pg24172 = pg99;
  assign pg24181 = pg126;
  assign pg8403 = ng5005;
  assign pg8788 = ng4207;
  assign pg9497 = ng5101;
  assign pg13926 = ng3632;
  assign pg14189 = ng859;
  assign pg14451 = ng3649;
  assign pg24162 = pg54;
  assign pg24180 = pg125;
  assign pg7245 = ng4446;
  assign pg8215 = ng3092;
  assign pg8789 = ng4210;
  assign pg10122 = ng4294;
  assign pg12919 = ng1227;
  assign pg16924 = ng3668;
  assign pg17291 = ng1075;
  assign pg20763 = ng74;
  assign pg24161 = pg53;
  assign pg24170 = pg91;
  assign pg34238 = pg34237;
  assign pg14705 = ng6369;
  assign pg14738 = ng5983;
  assign pg14749 = ng6715;
  assign pg16693 = ng3976;
  assign pg16718 = ng3310;
  assign pg17423 = ng1426;
  assign pg18097 = pg6747;
  assign pg24164 = pg57;
  assign pg24175 = pg114;
  assign pg29211 = ng74;
  assign pg18098 = pg6744;
  assign pg20901 = ng102;
  assign pg24163 = pg56;
  assign pg24176 = pg115;
  assign pg24185 = pg44;
  assign pg29210 = ng59;
  assign pg11388 = ng3654;
  assign pg17577 = ng5283;
  assign pg17674 = ng5320;
  assign pg17760 = ng6358;
  assign pg18099 = pg6745;
  assign pg20652 = ng94;
  assign pg24166 = pg72;
  assign pg24173 = pg100;
  assign pg24184 = pg135;
  assign pg29213 = ng86;
  assign pg29220 = ng128;
  assign pg34233 = pg34235;
  assign pg14597 = ng5331;
  assign pg14694 = ng5637;
  assign pg17813 = ng5673;
  assign pg21292 = ng136;
  assign pg24165 = pg64;
  assign pg24174 = pg113;
  assign pg24183 = pg134;
  assign pg29212 = ng79;
  assign pg29221 = ng136;
  assign pg32975 = pg26801;
  assign pg34234 = pg34235;
  assign pg34788 = pg33894;
  assign pg11678 = ng802;
  assign pg12923 = ng1570;
  assign pg14518 = ng4000;
  assign pg14662 = ng5290;
  assign pg14673 = ng6023;
  assign pg17607 = ng5969;
  assign pg17715 = ng6027;
  assign pg19357 = ng1399;
  assign pg24168 = pg84;
  assign pg24179 = pg124;
  assign pg25219 = ng5343;
  assign pg29215 = ng102;
  assign pg30332 = ng1242;
  assign pg16627 = ng3618;
  assign pg23612 = pg30329;
  assign pg24167 = pg73;
  assign pg29214 = ng94;
  assign pg14635 = ng5677;
  assign pg17519 = ng5276;
  assign pg17580 = ng5623;
  assign pg24177 = pg116;
  assign pg29217 = ng117;
  assign pg30330 = pg23652;
  assign pg34240 = pg34237;
  assign pg12832 = ng1;
  assign pg16722 = ng3676;
  assign pg24169 = pg90;
  assign pg24178 = pg120;
  assign pg29216 = ng106;
  assign pg7916 = ng1157;
  assign pg8919 = ng4229;
  assign pg11447 = ng4191;
  assign pg13881 = ng3672;
  assign pg16624 = ng3274;
  assign pg17711 = ng5666;
  assign pg17722 = ng6668;
  assign pg20049 = ng59;
  assign pg29219 = ng121;
  assign pg8918 = ng4226;
  assign pg11770 = ng4185;
  assign pg16874 = ng3317;
  assign pg17604 = ng5630;
  assign pg21245 = ng128;
  assign pg29218 = ng66;
  assign pg34839 = pg34956;
  assign pg8839 = ng4277;
  assign pg16603 = ng3267;
  assign pg16656 = ng3625;
  assign pg16744 = ng3661;
  assign pg17646 = ng5976;
  assign pg17743 = ng6373;
  assign pg17778 = ng6704;
  assign pg17787 = ng5327;
  assign pg18092 = pg6753;
  assign pg11418 = ng4005;
  assign pg16686 = ng3325;
  assign pg17845 = ng6365;
  assign pg21176 = ng106;
  assign pg12368 = ng637;
  assign pg13895 = ng3281;
  assign pg14779 = ng6329;
  assign pg17639 = ng5335;
  assign pg17688 = ng6661;
  assign pg18094 = pg6748;
  assign pg18881 = ng66;
  assign pg23683 = ng1242;
  assign pg10527 = ng1576;
  assign pg13865 = ng3321;
  assign pg16659 = ng3969;
  assign pg17649 = ng6315;
  assign pg17678 = ng5681;
  assign pg17685 = ng6322;
  assign pg17739 = ng6012;
  assign pg17764 = ng6719;
  assign pg18095 = pg6749;
  assign pg11349 = ng3303;
  assign pg13259 = ng1116;
  assign pg16748 = ng4027;
  assign pg16775 = ng4012;
  assign pg17316 = ng1079;
  assign pg17404 = ng1422;
  assign pg17871 = ng6711;
  assign pg18096 = pg6750;
  assign pg21270 = ng117;
  assign pg8416 = ng1239;
  assign pg9617 = ng5794;
  assign pg31863 = pg25167;
  assign pg7257 = ng4414;
  assign pg8920 = ng4232;
  assign pg9251 = ng4304;
  assign pg9817 = ng6490;
  assign pg13966 = ng3983;
  assign pg14217 = ng875;
  assign pg27831 = pg33533;
  assign pg31861 = ng5343;
  assign pg8291 = ng215;
  assign pg12238 = ng5313;
  assign pg12300 = ng5659;
  assign pg14096 = ng878;
  assign pg14201 = ng869;
  assign pg14421 = ng3298;
  assign pg16955 = ng4019;
  assign pg17400 = ng1083;
  assign pg31862 = pg25259;
  assign pg8283 = ng5002;
  assign pg8915 = ng4213;
  assign pg9019 = ng4287;
  assign pg9682 = ng6140;
  assign pg12350 = ng6005;
  assign pg12422 = ng6351;
  assign pg13049 = ng5654;
  assign pg13085 = ng6346;
  assign pg14125 = ng881;
  assign pg14147 = ng884;
  assign pg31665 = pg34437;
  assign pg8279 = ng3443;
  assign pg21698 = pg36;
  assign pg31860 = pg25114;
  assign pg8719 = ng365;
  assign pg8917 = ng4219;
  assign pg9615 = ng5452;
  assign pg9680 = ng5798;
  assign pg9743 = ng6486;
  assign pg23002 = pg30327;
  assign pg28753 = pg33959;
  assign pg31656 = pg34436;
  assign pg7946 = ng1500;
  assign pg8178 = ng4999;
  assign pg8277 = ng3096;
  assign pg8358 = ng194;
  assign pg8475 = ng1582;
  assign pg8916 = ng4216;
  assign pg9553 = ng5105;
  assign pg10306 = ng4537;
  assign pg10500 = ng1233;
  assign pg13039 = ng5308;
  assign pg23759 = pg30331;
  assign n793 = ng4005;
  assign n843 = ng1239;
  assign n868 = ng5276;
  assign n903 = ng1075;
  assign n923 = ng4449;
  assign n928 = ng1116;
  assign n953 = ng884;
  assign n968 = ng5983;
  assign n998 = ng4219;
  assign n1033 = ng4027;
  assign n1113 = pg33079;
  assign n1143 = ng4185;
  assign n1223 = ng5794;
  assign n1238 = ng6023;
  assign n1253 = ng4294;
  assign n1258 = ng1500;
  assign n1273 = ng3668;
  assign n1313 = ng3654;
  assign n1378 = ng1056;
  assign n1402 = ng5681;
  assign n1442 = ng5308;
  assign n1467 = ng194;
  assign n1482 = ng3649;
  assign n1531 = ng344;
  assign n1546 = ng4204;
  assign n1556 = ng6019;
  assign n1560 = pg33435;
  assign n1580 = ng3274;
  assign n1670 = ng5637;
  assign n1685 = ng6490;
  assign n1735 = ng6358;
  assign n1764 = ng6140;
  assign n1794 = ng5101;
  assign n1873 = ng4537;
  assign n1926 = ng3443;
  assign n1956 = ng6369;
  assign n1960 = ng3632;
  assign n1975 = ng6692;
  assign n1985 = ng4809;
  assign n2055 = ng5005;
  assign n2080 = ng5673;
  assign n2105 = ng5630;
  assign n2119 = ng5448;
  assign n2187 = ng3983;
  assign n2217 = ng4000;
  assign n2227 = ng878;
  assign n2297 = ng4194;
  assign n2327 = ng5313;
  assign n2381 = ng365;
  assign n2436 = ng6346;
  assign n2490 = ng1079;
  assign n2609 = ng6351;
  assign n2644 = ng4277;
  assign n2673 = ng4213;
  assign n2762 = ng3298;
  assign n2787 = ng4226;
  assign n2812 = ng4519;
  assign n2896 = ng4197;
  assign n2941 = ng5623;
  assign n2944 = ng6012;
  assign n2948 = ng6315;
  assign n3097 = ng5677;
  assign n3156 = ng4999;
  assign n3161 = ng1459;
  assign n3196 = ng869;
  assign n3265 = ng3672;
  assign n3538 = ng4812;
  assign n3618 = ng4210;
  assign n3652 = ng3661;
  assign n3657 = ng3794;
  assign n3700 = ng5452;
  assign n3738 = ng5654;
  assign n3762 = ng3969;
  assign n3772 = ng6000;
  assign n3825 = ng4216;
  assign n3834 = ng3281;
  assign n4009 = ng5331;
  assign n4037 = ng1570;
  assign n4042 = ng3447;
  assign n4180 = ng5105;
  assign n4190 = ng3325;
  assign n4255 = ng6668;
  assign n4338 = ng4304;
  assign n4397 = ng6697;
  assign n4407 = ng1227;
  assign n4416 = ng6365;
  assign n4424 = ng5290;
  assign n4443 = ng6322;
  assign n4451 = ng4815;
  assign n4490 = ng5659;
  assign n4524 = ng640;
  assign n4544 = ng1576;
  assign n4608 = ng3798;
  assign n4623 = ng4570;
  assign n4682 = ng5969;
  assign n4687 = ng6715;
  assign n4691 = ng1233;
  assign n4710 = ng6711;
  assign n4718 = ng5320;
  assign n4767 = ng4023;
  assign n4848 = ng875;
  assign n4891 = ng1083;
  assign n4936 = ng3303;
  assign n5015 = ng3096;
  assign n5054 = ng5976;
  assign n5077 = ng4520;
  assign n5127 = ng3321;
  assign n5181 = ng3092;
  assign n5235 = ng3676;
  assign n5312 = ng6329;
  assign n5330 = ng5327;
  assign n5353 = ng6486;
  assign n5373 = pg6752;
  assign n5477 = ng6661;
  assign n5480 = ng6675;
  assign n5509 = ng3310;
  assign n5533 = ng3267;
  assign n5566 = ng637;
  assign n5594 = ng4012;
  assign n5672 = ng5798;
  assign n5766 = ng4414;
  assign n5785 = ng4019;
  assign n5921 = ng1157;
  assign n5983 = ng1418;
  assign n6033 = ng802;
  assign n6037 = ng5666;
  assign n6045 = ng5335;
  assign n6065 = ng6005;
  assign n6088 = ng4446;
  assign n6092 = ng881;
  assign n6105 = ng4222;
  assign n6169 = ng6144;
  assign n6188 = ng5283;
  assign n6216 = ng4207;
  assign n6304 = ng6704;
  assign n6342 = ng4229;
  assign n6489 = ng1399;
  assign n6513 = ng1426;
  assign n6527 = ng1582;
  assign n6566 = ng4191;
  assign n6600 = ng859;
  assign n6614 = ng4467;
  assign n6628 = ng3976;
  assign n6810 = ng4200;
  assign n6902 = ng3618;
  assign n6916 = ng6373;
  assign n7019 = ng4188;
  assign n7027 = ng799;
  assign n7089 = ng6027;
  assign n7093 = ng4232;
  assign n7280 = ng3625;
  assign n7383 = ng4287;
  assign n7392 = ng215;
  assign n7426 = ng3317;
  assign n7537 = ng6719;
  assign n7551 = ng4571;
  assign n7584 = ng4408;
  assign n7603 = ng1422;
  assign n7641 = ng887;
  assign n7660 = ng5002;
  always @ (posedge clock) begin
    ng6215 <= n688;
    ng4332 <= n693;
    ng2837 <= n698;
    ng1135 <= n703;
    ng2485 <= n708;
    ng4375 <= n713;
    ng4304 <= n718;
    ng1171 <= n723;
    ng3235 <= n728;
    ng2852 <= n733;
    ng4135 <= n738;
    ng222 <= n743;
    ng365 <= n748;
    ng2815 <= n753;
    ng4888 <= n758;
    ng433 <= n763;
    ng3736 <= n768;
    ng246 <= n773;
    ng102 <= n778;
    ng1030 <= n783;
    ng110 <= n788;
    ng3983 <= n793;
    ng4801 <= n798;
    ng4045 <= n803;
    ng4169 <= n808;
    ng2145 <= n813;
    ng5138 <= n818;
    ng3873 <= n823;
    ng3752 <= n828;
    ng136 <= n833;
    ng1772 <= n838;
    ng990 <= n843;
    ng3171 <= n848;
    ng168 <= n853;
    ng441 <= n858;
    ng160 <= n863;
    ng5283 <= n868;
    ng1361 <= n873;
    ng6621 <= n878;
    ng5689 <= n883;
    ng6593 <= n888;
    ng55 <= n893;
    ng5827 <= n898;
    ng1079 <= n903;
    ng74 <= n908;
    ng5381 <= n913;
    ng5723 <= n918;
    ng4443 <= n923;
    ng979 <= n928;
    ng1484 <= n933;
    ng6044 <= n938;
    ng3817 <= n943;
    ng316 <= n948;
    ng887 <= n953;
    ng3080 <= n958;
    ng499 <= n963;
    ng6012 <= n968;
    ng3443 <= n973;
    ng2269 <= n978;
    ng2927 <= n983;
    ng577 <= n988;
    ng599 <= n993;
    ng4222 <= n998;
    ng781 <= n1003;
    ng6428 <= n1008;
    ng2759 <= n1013;
    ng2715 <= n1018;
    ng1870 <= n1023;
    ng1768 <= n1028;
    ng4031 <= n1033;
    ng6181 <= n1038;
    ng5731 <= n1043;
    ng2173 <= n1048;
    ng1783 <= n1053;
    ng6058 <= n1058;
    ng106 <= n1063;
    ng2711 <= n1068;
    ng2803 <= n1073;
    ng6303 <= n1078;
    ng3462 <= n1083;
    ng482 <= n1088;
    ng3085 <= n1093;
    ng1811 <= n1098;
    ng2890 <= n1103;
    ng1542 <= n1108;
    ng111 <= n1113;
    ng2161 <= n1118;
    ng947 <= n1123;
    ng546 <= n1128;
    ng3913 <= n1133;
    ng1570 <= n1138;
    ng4213 <= n1143;
    ng5599 <= n1148;
    ng3893 <= n1153;
    ng4141 <= n1158;
    ng3106 <= n1163;
    ng3841 <= n1168;
    ng2004 <= n1173;
    ng3586 <= n1178;
    ng4132 <= n1183;
    ng939 <= n1188;
    ng6195 <= n1193;
    ng925 <= n1198;
    ng6255 <= n1203;
    ng2177 <= n1208;
    ng5835 <= n1213;
    ng4543 <= n1218;
    ng5802 <= n1223;
    ng5092 <= n1228;
    ng3933 <= n1233;
    ng6027 <= n1238;
    ng911 <= n1243;
    ng3901 <= n1248;
    ng4297 <= n1253;
    ng1582 <= n1258;
    ng4049 <= n1263;
    ng3139 <= n1268;
    ng3672 <= n1273;
    ng6649 <= n1278;
    ng2599 <= n1283;
    ng4087 <= n1288;
    ng1467 <= n1293;
    ng6519 <= n1298;
    ng1700 <= n1303;
    ng1950 <= n1308;
    ng3632 <= n1313;
    ng46 <= n1318;
    ng2417 <= n1323;
    ng4741 <= n1328;
    ng475 <= n1333;
    ng3787 <= n1338;
    ng333 <= n1343;
    ng5105 <= n1348;
    ng6351 <= n1353;
    ng1779 <= n1358;
    ng2834 <= n1363;
    ng3470 <= n1368;
    ng5188 <= n1373;
    ng1116 <= n1378;
    ng504 <= n1382;
    ng3767 <= n1387;
    ng6541 <= n1392;
    ng6209 <= n1397;
    ng5685 <= n1402;
    ng1157 <= n1407;
    ng3466 <= n1412;
    ng3333 <= n1417;
    ng4922 <= n1422;
    ng6613 <= n1427;
    ng93 <= n1432;
    ng637 <= n1437;
    ng5327 <= n1442;
    ng1478 <= n1447;
    ng5413 <= n1452;
    ng63 <= n1457;
    ng2643 <= n1462;
    ng191 <= n1467;
    ng6052 <= n1472;
    ng1620 <= n1477;
    ng3668 <= n1482;
    ng2495 <= n1486;
    ng5583 <= n1491;
    ng2138 <= n1496;
    ng5244 <= n1501;
    ng936 <= n1506;
    ng429 <= n1511;
    ng4854 <= n1516;
    ng37 <= n1521;
    ng6381 <= n1526;
    ng347 <= n1531;
    ng4287 <= n1536;
    ng2767 <= n1541;
    ng4207 <= n1546;
    ng5921 <= n1551;
    ng6023 <= n1556;
    ng85 <= n1560;
    ng5069 <= n1565;
    ng1061 <= n1570;
    ng4401 <= n1575;
    ng3298 <= n1580;
    ng3431 <= n1585;
    ng3610 <= n1590;
    ng4975 <= n1595;
    ng4427 <= n1600;
    ng4145 <= n1605;
    ng1834 <= n1610;
    ng5703 <= n1615;
    ng4537 <= n1620;
    ng1141 <= n1625;
    ng6120 <= n1630;
    ng4512 <= n1635;
    ng4253 <= n1640;
    ng4570 <= n1645;
    ng1548 <= n1650;
    ng4284 <= n1655;
    ng385 <= n1660;
    ng291 <= n1665;
    ng5666 <= n1670;
    ng3111 <= n1675;
    ng718 <= n1680;
    ng6497 <= n1685;
    ng6267 <= n1690;
    ng3010 <= n1695;
    ng2399 <= n1700;
    ng2898 <= n1705;
    ng4414 <= n1710;
    ng4831 <= n1715;
    ng5889 <= n1720;
    ng822 <= n1725;
    ng43 <= n1730;
    ng6315 <= n1735;
    ng2112 <= n1740;
    ng5543 <= n1745;
    ng4449 <= n1750;
    ng142 <= n1754;
    ng5022 <= n1759;
    ng6148 <= n1764;
    ng1448 <= n1769;
    ng3961 <= n1774;
    ng1018 <= n1779;
    ng5029 <= n1784;
    ng513 <= n1789;
    ng5109 <= n1794;
    ng2016 <= n1799;
    ng5575 <= n1804;
    ng5052 <= n1809;
    ng3412 <= n1814;
    ng1992 <= n1819;
    ng2902 <= n1824;
    ng3808 <= n1829;
    ng5373 <= n1834;
    ng1608 <= n1839;
    ng5535 <= n1844;
    ng405 <= n1849;
    ng215 <= n1854;
    ng5448 <= n1859;
    ng3203 <= n1864;
    ng655 <= n1869;
    ng4423 <= n1873;
    ng4633 <= n1878;
    ng4116 <= n1883;
    ng298 <= n1888;
    ng1075 <= n1893;
    ng4501 <= n1897;
    ng6513 <= n1902;
    ng3368 <= n1907;
    ng5240 <= n1912;
    ng1002 <= n1917;
    ng896 <= n1922;
    ng3451 <= n1926;
    ng2712 <= n1931;
    ng5929 <= n1936;
    ng6486 <= n1941;
    ng837 <= n1946;
    ng2437 <= n1951;
    ng6373 <= n1956;
    ng3661 <= n1960;
    ng785 <= n1965;
    ng2575 <= n1970;
    ng6711 <= n1975;
    ng3925 <= n1980;
    ng4812 <= n1985;
    ng4765 <= n1990;
    ng1266 <= n1995;
    ng6605 <= n2000;
    ng2868 <= n2005;
    ng6573 <= n2010;
    ng5485 <= n2015;
    ng1211 <= n2020;
    ng1821 <= n2025;
    ng5124 <= n2030;
    ng5377 <= n2035;
    ng6434 <= n2040;
    ng6697 <= n2045;
    ng4932 <= n2050;
    ng5008 <= n2055;
    ng790 <= n2060;
    ng5142 <= n2065;
    ng3594 <= n2070;
    ng5953 <= n2075;
    ng5677 <= n2080;
    ng6561 <= n2085;
    ng2775 <= n2090;
    ng4366 <= n2095;
    ng5016 <= n2100;
    ng5654 <= n2105;
    ng5128 <= n2110;
    ng3763 <= n2115;
    ng5456 <= n2119;
    ng4674 <= n2124;
    ng4153 <= n2129;
    ng117 <= n2134;
    ng3239 <= n2139;
    ng1437 <= n2144;
    ng4809 <= n2149;
    ng52 <= n2153;
    ng4269 <= n2158;
    ng3343 <= n2163;
    ng2819 <= n2168;
    ng3050 <= n2173;
    ng4495 <= n2178;
    ng1070 <= n2183;
    ng4012 <= n2187;
    ng6251 <= n2192;
    ng1283 <= n2197;
    ng6537 <= n2202;
    ng2932 <= n2207;
    ng4584 <= n2212;
    ng4019 <= n2217;
    ng5798 <= n2222;
    ng881 <= n2227;
    ng2984 <= n2232;
    ng1418 <= n2237;
    ng1256 <= n2242;
    ng2841 <= n2247;
    ng2307 <= n2252;
    ng5759 <= n2257;
    ng3719 <= n2262;
    ng5452 <= n2267;
    ng31 <= n2272;
    ng3029 <= n2277;
    ng4455 <= n2282;
    ng9 <= n2287;
    ng5445 <= n2292;
    ng4197 <= n2297;
    ng4950 <= n2302;
    ng5216 <= n2307;
    ng2710 <= n2312;
    ng1936 <= n2317;
    ng1668 <= n2322;
    ng5290 <= n2327;
    ng3689 <= n2332;
    ng4146 <= n2337;
    ng4681 <= n2342;
    ng3774 <= n2347;
    ng827 <= n2352;
    ng287 <= n2357;
    ng1277 <= n2362;
    ng2799 <= n2367;
    ng1945 <= n2372;
    ng776 <= n2377;
    ng358 <= n2381;
    ng967 <= n2386;
    ng626 <= n2391;
    ng4340 <= n2396;
    ng2036 <= n2401;
    ng1249 <= n2406;
    ng2102 <= n2411;
    ng6173 <= n2416;
    ng2338 <= n2421;
    ng6741 <= n2426;
    ng65 <= n2431;
    ng6365 <= n2436;
    ng6509 <= n2441;
    ng2070 <= n2446;
    ng5563 <= n2451;
    ng4473 <= n2456;
    ng2445 <= n2461;
    ng2407 <= n2466;
    ng1677 <= n2471;
    ng86 <= n2476;
    ng2827 <= n2481;
    ng6451 <= n2486;
    ng1083 <= n2490;
    ng1306 <= n2495;
    ng1514 <= n2500;
    ng4727 <= n2505;
    ng3219 <= n2510;
    ng6597 <= n2515;
    ng5913 <= n2520;
    ng3259 <= n2525;
    ng2999 <= n2530;
    ng2472 <= n2535;
    ng3195 <= n2540;
    ng4417 <= n2545;
    ng2922 <= n2550;
    ng3401 <= n2555;
    ng3119 <= n2560;
    ng3211 <= n2565;
    ng3821 <= n2570;
    ng3191 <= n2575;
    ng2527 <= n2580;
    ng3243 <= n2585;
    ng5204 <= n2590;
    ng1862 <= n2595;
    ng6065 <= n2600;
    ng1178 <= n2605;
    ng6329 <= n2609;
    ng3530 <= n2614;
    ng4273 <= n2619;
    ng4572 <= n2624;
    ng2259 <= n2629;
    ng6191 <= n2634;
    ng6307 <= n2639;
    ng4281 <= n2644;
    ng4639 <= n2649;
    ng5037 <= n2654;
    ng6279 <= n2659;
    ng471 <= n2664;
    ng5297 <= n2669;
    ng4216 <= n2673;
    ng232 <= n2678;
    ng3759 <= n2683;
    ng3498 <= n2688;
    ng6555 <= n2693;
    ng1472 <= n2698;
    ng4760 <= n2703;
    ng2204 <= n2708;
    ng862 <= n2713;
    ng6736 <= n2718;
    ng6500 <= n2723;
    ng2724 <= n2728;
    ng2882 <= n2733;
    ng2541 <= n2738;
    ng6653 <= n2743;
    ng4894 <= n2748;
    ng2476 <= n2753;
    ng2729 <= n2758;
    ng3317 <= n2762;
    ng930 <= n2767;
    ng6682 <= n2772;
    ng2873 <= n2777;
    ng4899 <= n2782;
    ng4229 <= n2787;
    ng3484 <= n2792;
    ng604 <= n2797;
    ng1825 <= n2802;
    ng4392 <= n2807;
    ng4520 <= n2812;
    ng1395 <= n2817;
    ng714 <= n2822;
    ng79 <= n2827;
    ng6505 <= n2832;
    ng5462 <= n2837;
    ng3731 <= n2842;
    ng6423 <= n2847;
    ng5073 <= n2852;
    ng1636 <= n2857;
    ng5849 <= n2862;
    ng2197 <= n2867;
    ng4129 <= n2872;
    ng1858 <= n2877;
    ng6581 <= n2882;
    ng1902 <= n2887;
    ng2126 <= n2892;
    ng4200 <= n2896;
    ng582 <= n2901;
    ng3845 <= n2906;
    ng5747 <= n2911;
    ng2079 <= n2916;
    ng6082 <= n2921;
    ng5841 <= n2926;
    ng4239 <= n2931;
    ng5148 <= n2936;
    ng5630 <= n2941;
    ng5969 <= n2944;
    ng6322 <= n2948;
    ng128 <= n2953;
    ng2610 <= n2958;
    ng6727 <= n2963;
    ng4742 <= n2968;
    ng3143 <= n2973;
    ng4927 <= n2978;
    ng5077 <= n2983;
    ng2342 <= n2988;
    ng3574 <= n2993;
    ng4138 <= n2998;
    ng2319 <= n3003;
    ng5752 <= n3008;
    ng51 <= n3013;
    ng5791 <= n3018;
    ng1041 <= n3023;
    ng3770 <= n3028;
    ng4467 <= n3033;
    ng2279 <= n3038;
    ng859 <= n3043;
    ng2606 <= n3048;
    ng262 <= n3053;
    ng3502 <= n3058;
    ng5817 <= n3063;
    ng4944 <= n3068;
    ng3827 <= n3073;
    ng4704 <= n3078;
    ng336 <= n3083;
    ng2153 <= n3088;
    ng3480 <= n3093;
    ng5681 <= n3097;
    ng4646 <= n3101;
    ng5357 <= n3106;
    ng4907 <= n3111;
    ng3937 <= n3116;
    ng5949 <= n3121;
    ng1854 <= n3126;
    ng4064 <= n3131;
    ng6247 <= n3136;
    ng1259 <= n3141;
    ng6589 <= n3146;
    ng3004 <= n3151;
    ng5002 <= n3156;
    ng1322 <= n3161;
    ng1913 <= n3166;
    ng5489 <= n3171;
    ng182 <= n3176;
    ng1592 <= n3181;
    ng2689 <= n3186;
    ng3089 <= n3191;
    ng875 <= n3196;
    ng2509 <= n3201;
    ng3921 <= n3206;
    ng1756 <= n3211;
    ng6116 <= n3216;
    ng2950 <= n3221;
    ng446 <= n3226;
    ng4349 <= n3231;
    ng6163 <= n3236;
    ng5248 <= n3241;
    ng4446 <= n3246;
    ng4191 <= n3251;
    ng2116 <= n3256;
    ng2697 <= n3261;
    ng3676 <= n3265;
    ng49 <= n3270;
    ng2453 <= n3275;
    ng3391 <= n3280;
    ng4420 <= n3285;
    ng3606 <= n3290;
    ng843 <= n3295;
    ng3506 <= n3300;
    ng1036 <= n3305;
    ng4104 <= n3310;
    ng1706 <= n3315;
    ng6398 <= n3320;
    ng5523 <= n3325;
    ng6159 <= n3330;
    ng2960 <= n3335;
    ng5495 <= n3340;
    ng2975 <= n3345;
    ng6549 <= n3350;
    ng2315 <= n3355;
    ng2595 <= n3360;
    ng6545 <= n3365;
    ng2652 <= n3370;
    ng6235 <= n3375;
    ng3385 <= n3380;
    ng542 <= n3385;
    ng1840 <= n3390;
    ng703 <= n3395;
    ng5101 <= n3400;
    ng4072 <= n3404;
    ng3133 <= n3409;
    ng22 <= n3414;
    ng1906 <= n3419;
    ng4912 <= n3424;
    ng1959 <= n3429;
    ng3857 <= n3434;
    ng2375 <= n3439;
    ng4991 <= n3444;
    ng2946 <= n3449;
    ng2831 <= n3454;
    ng739 <= n3459;
    ng5084 <= n3464;
    ng4785 <= n3469;
    ng2791 <= n3474;
    ng6609 <= n3479;
    ng2098 <= n3484;
    ng6455 <= n3489;
    ng3546 <= n3494;
    ng2185 <= n3499;
    ng2491 <= n3504;
    ng1312 <= n3509;
    ng1129 <= n3514;
    ng1221 <= n3519;
    ng1624 <= n3524;
    ng1848 <= n3529;
    ng4859 <= n3534;
    ng4815 <= n3538;
    ng2994 <= n3543;
    ng956 <= n3548;
    ng2421 <= n3553;
    ng6533 <= n3558;
    ng370 <= n3563;
    ng1874 <= n3568;
    ng4125 <= n3573;
    ng5481 <= n3578;
    ng7 <= n3583;
    ng2361 <= n3588;
    ng2327 <= n3593;
    ng723 <= n3598;
    ng94 <= n3603;
    ng3703 <= n3608;
    ng4549 <= n3613;
    ng4180 <= n3618;
    ng1926 <= n3623;
    ng676 <= n3628;
    ng4558 <= n3633;
    ng4864 <= n3638;
    ng1532 <= n3643;
    ng1389 <= n3648;
    ng3618 <= n3652;
    ng3802 <= n3657;
    ng2255 <= n3662;
    ng5499 <= n3667;
    ng4185 <= n3672;
    ng5917 <= n3676;
    ng6167 <= n3681;
    ng3917 <= n3686;
    ng2537 <= n3691;
    ng5268 <= n3696;
    ng5459 <= n3700;
    ng3419 <= n3705;
    ng3881 <= n3710;
    ng6113 <= n3715;
    ng5256 <= n3720;
    ng5421 <= n3725;
    ng4732 <= n3730;
    ng344 <= n3735;
    ng5673 <= n3738;
    ng2878 <= n3742;
    ng933 <= n3747;
    ng4157 <= n3752;
    ng3863 <= n3757;
    ng3976 <= n3762;
    ng1657 <= n3767;
    ng6019 <= n3772;
    ng4035 <= n3776;
    ng667 <= n3781;
    ng5475 <= n3786;
    ng5603 <= n3791;
    ng2719 <= n3796;
    ng3949 <= n3801;
    ng209 <= n3806;
    ng4462 <= n3811;
    ng4249 <= n3816;
    ng5236 <= n3821;
    ng4219 <= n3825;
    ng4849 <= n3829;
    ng3310 <= n3834;
    ng2227 <= n3839;
    ng6411 <= n3844;
    ng5062 <= n3849;
    ng34 <= n3854;
    ng424 <= n3859;
    ng1280 <= n3864;
    ng650 <= n3869;
    ng2181 <= n3874;
    ng1046 <= n3879;
    ng1345 <= n3884;
    ng5694 <= n3889;
    ng2441 <= n3894;
    ng4821 <= n3899;
    ng3694 <= n3904;
    ng2779 <= n3909;
    ng376 <= n3914;
    ng907 <= n3919;
    ng699 <= n3924;
    ng3129 <= n3929;
    ng4698 <= n3934;
    ng6035 <= n3939;
    ng4507 <= n3944;
    ng4040 <= n3949;
    ng3380 <= n3954;
    ng5555 <= n3959;
    ng590 <= n3964;
    ng1752 <= n3969;
    ng4477 <= n3974;
    ng1296 <= n3979;
    ng4382 <= n3984;
    ng1052 <= n3989;
    ng1728 <= n3994;
    ng969 <= n3999;
    ng355 <= n4004;
    ng5335 <= n4009;
    ng6490 <= n4014;
    ng225 <= n4018;
    ng5869 <= n4023;
    ng153 <= n4028;
    ng2811 <= n4033;
    ng1585 <= n4037;
    ng3454 <= n4042;
    ng4108 <= n4047;
    ng5881 <= n4052;
    ng1146 <= n4057;
    ng518 <= n4062;
    ng4531 <= n4067;
    ng3045 <= n4072;
    ng468 <= n4077;
    ng5041 <= n4082;
    ng2988 <= n4087;
    ng1526 <= n4092;
    ng568 <= n4097;
    ng4294 <= n4102;
    ng3361 <= n4106;
    ng4546 <= n4111;
    ng3072 <= n4116;
    ng6098 <= n4121;
    ng6283 <= n4126;
    ng6415 <= n4131;
    ng5120 <= n4136;
    ng1399 <= n4141;
    ng4322 <= n4146;
    ng5252 <= n4151;
    ng1274 <= n4156;
    ng112 <= n4161;
    ng5033 <= n4166;
    ng4939 <= n4171;
    ng5097 <= n4176;
    ng5112 <= n4180;
    ng3408 <= n4185;
    ng3329 <= n4190;
    ng943 <= n4195;
    ng5200 <= n4200;
    ng2912 <= n4205;
    ng3352 <= n4210;
    ng3125 <= n4215;
    ng1988 <= n4220;
    ng5348 <= n4225;
    ng1 <= n4230;
    ng1878 <= n4235;
    ng2547 <= n4240;
    ng5343 <= n4245;
    ng48 <= n4250;
    ng6692 <= n4255;
    ng5567 <= n4259;
    ng1233 <= n4264;
    ng753 <= n4269;
    ng351 <= n4274;
    ng58 <= n4279;
    ng3179 <= n4284;
    ng2807 <= n4289;
    ng1682 <= n4294;
    ng5831 <= n4299;
    ng3231 <= n4304;
    ng4486 <= n4309;
    ng5579 <= n4314;
    ng6625 <= n4319;
    ng3798 <= n4324;
    ng4388 <= n4329;
    ng4564 <= n4334;
    ng4308 <= n4338;
    ng5385 <= n4343;
    ng2625 <= n4348;
    ng3897 <= n4353;
    ng2860 <= n4358;
    ng6641 <= n4363;
    ng5396 <= n4368;
    ng2151 <= n4373;
    ng3538 <= n4378;
    ng6523 <= n4383;
    ng3263 <= n4388;
    ng3562 <= n4393;
    ng6675 <= n4397;
    ng5937 <= n4402;
    ng1242 <= n4407;
    ng4771 <= n4412;
    ng6369 <= n4416;
    ng4966 <= n4420;
    ng5320 <= n4424;
    ng1199 <= n4429;
    ng5941 <= n4434;
    ng1152 <= n4439;
    ng6346 <= n4443;
    ng2856 <= n4447;
    ng4818 <= n4451;
    ng1056 <= n4456;
    ng1964 <= n4460;
    ng19 <= n4465;
    ng5401 <= n4470;
    ng5170 <= n4475;
    ng1559 <= n4480;
    ng4843 <= n4485;
    ng5637 <= n4490;
    ng6657 <= n4494;
    ng2894 <= n4499;
    ng4311 <= n4504;
    ng3223 <= n4509;
    ng3251 <= n4514;
    ng5619 <= n4519;
    ng559 <= n4524;
    ng554 <= n4529;
    ng1798 <= n4534;
    ng4871 <= n4539;
    ng1579 <= n4544;
    ng4643 <= n4549;
    ng2980 <= n4554;
    ng5901 <= n4559;
    ng479 <= n4564;
    ng4653 <= n4569;
    ng5424 <= n4574;
    ng1105 <= n4579;
    ng3889 <= n4584;
    ng4098 <= n4589;
    ng4504 <= n4594;
    ng1589 <= n4599;
    ng5990 <= n4604;
    ng3805 <= n4608;
    ng6275 <= n4613;
    ng6239 <= n4618;
    ng4571 <= n4623;
    ng5406 <= n4628;
    ng150 <= n4633;
    ng538 <= n4638;
    ng4743 <= n4643;
    ng5571 <= n4648;
    ng5196 <= n4653;
    ng2351 <= n4658;
    ng4434 <= n4663;
    ng301 <= n4668;
    ng854 <= n4673;
    ng2518 <= n4678;
    ng5976 <= n4682;
    ng6719 <= n4687;
    ng1236 <= n4691;
    ng4616 <= n4696;
    ng2523 <= n4701;
    ng2551 <= n4706;
    ng6715 <= n4710;
    ng2579 <= n4714;
    ng5276 <= n4718;
    ng3929 <= n4722;
    ng2012 <= n4727;
    ng4836 <= n4732;
    ng2108 <= n4737;
    ng2571 <= n4742;
    ng2093 <= n4747;
    ng6479 <= n4752;
    ng1554 <= n4757;
    ng3207 <= n4762;
    ng4027 <= n4767;
    ng1720 <= n4771;
    ng1193 <= n4776;
    ng3255 <= n4781;
    ng5893 <= n4786;
    ng4456 <= n4791;
    ng6140 <= n4796;
    ng1300 <= n4800;
    ng3747 <= n4805;
    ng4552 <= n4810;
    ng5417 <= n4815;
    ng3187 <= n4820;
    ng4931 <= n4825;
    ng1996 <= n4830;
    ng3654 <= n4835;
    ng3017 <= n4839;
    ng496 <= n4844;
    ng878 <= n4848;
    ng4722 <= n4852;
    ng6154 <= n4857;
    ng5264 <= n4862;
    ng3151 <= n4867;
    ng2886 <= n4872;
    ng6386 <= n4877;
    ng5736 <= n4882;
    ng4054 <= n4887;
    ng1087 <= n4891;
    ng3476 <= n4896;
    ng4575 <= n4901;
    ng5873 <= n4906;
    ng5719 <= n4911;
    ng4578 <= n4916;
    ng4459 <= n4921;
    ng6311 <= n4926;
    ng4826 <= n4931;
    ng3281 <= n4936;
    ng3338 <= n4940;
    ng1696 <= n4945;
    ng3025 <= n4950;
    ng6 <= n4955;
    ng3578 <= n4960;
    ng2380 <= n4965;
    ng2648 <= n4970;
    ng5441 <= n4975;
    ng341 <= n4980;
    ng4601 <= n4985;
    ng2567 <= n4990;
    ng890 <= n4995;
    ng2864 <= n5000;
    ng28 <= n5005;
    ng4561 <= n5010;
    ng3103 <= n5015;
    ng5156 <= n5020;
    ng2273 <= n5025;
    ng904 <= n5030;
    ng6459 <= n5035;
    ng6227 <= n5040;
    ng6203 <= n5045;
    ng66 <= n5050;
    ng6000 <= n5054;
    ng2165 <= n5058;
    ng4112 <= n5063;
    ng1982 <= n5068;
    ng4717 <= n5073;
    ng4483 <= n5077;
    ng3215 <= n5082;
    ng1367 <= n5087;
    ng2051 <= n5092;
    ng1691 <= n5097;
    ng1111 <= n5102;
    ng5821 <= n5107;
    ng411 <= n5112;
    ng4057 <= n5117;
    ng5763 <= n5122;
    ng3325 <= n5127;
    ng2661 <= n5131;
    ng3061 <= n5136;
    ng2970 <= n5141;
    ng4628 <= n5146;
    ng12 <= n5151;
    ng2771 <= n5156;
    ng3570 <= n5161;
    ng622 <= n5166;
    ng3853 <= n5171;
    ng2941 <= n5176;
    ng3100 <= n5181;
    ng4737 <= n5186;
    ng3440 <= n5191;
    ng5360 <= n5196;
    ng4754 <= n5201;
    ng4983 <= n5206;
    ng4961 <= n5211;
    ng3494 <= n5216;
    ng4749 <= n5221;
    ng2465 <= n5226;
    ng4917 <= n5231;
    ng3680 <= n5235;
    ng1748 <= n5240;
    ng3092 <= n5245;
    ng758 <= n5249;
    ng1227 <= n5254;
    ng1664 <= n5258;
    ng528 <= n5263;
    ng2848 <= n5268;
    ng1564 <= n5273;
    ng3712 <= n5278;
    ng962 <= n5283;
    ng457 <= n5288;
    ng5787 <= n5293;
    ng3831 <= n5298;
    ng4793 <= n5303;
    ng5808 <= n5308;
    ng6358 <= n5312;
    ng1890 <= n5316;
    ng799 <= n5321;
    ng5897 <= n5326;
    ng5331 <= n5330;
    ng3791 <= n5334;
    ng4093 <= n5339;
    ng2619 <= n5344;
    ng661 <= n5349;
    ng6494 <= n5353;
    ng1413 <= n5358;
    ng2311 <= n5363;
    ng5774 <= n5368;
    ng70 <= n5373;
    ng794 <= n5378;
    ng4999 <= n5383;
    ng2667 <= n5387;
    ng2555 <= n5392;
    ng4581 <= n5397;
    ng1616 <= n5402;
    ng305 <= n5407;
    ng255 <= n5412;
    ng3423 <= n5417;
    ng613 <= n5422;
    ng5390 <= n5427;
    ng3034 <= n5432;
    ng817 <= n5437;
    ng686 <= n5442;
    ng4489 <= n5447;
    ng4955 <= n5452;
    ng2675 <= n5457;
    ng25 <= n5462;
    ng391 <= n5467;
    ng329 <= n5472;
    ng6668 <= n5477;
    ng6704 <= n5480;
    ng5727 <= n5485;
    ng6439 <= n5490;
    ng2533 <= n5495;
    ng6404 <= n5500;
    ng2936 <= n5505;
    ng3267 <= n5509;
    ng6299 <= n5514;
    ng3068 <= n5519;
    ng319 <= n5524;
    ng1351 <= n5529;
    ng3274 <= n5533;
    ng728 <= n5537;
    ng2084 <= n5542;
    ng691 <= n5547;
    ng5698 <= n5552;
    ng4515 <= n5557;
    ng1882 <= n5562;
    ng640 <= n5566;
    ng6336 <= n5570;
    ng5134 <= n5575;
    ng4076 <= n5580;
    ng1495 <= n5585;
    ng3040 <= n5590;
    ng3969 <= n5594;
    ng5160 <= n5598;
    ng1189 <= n5603;
    ng3372 <= n5608;
    ng437 <= n5613;
    ng5511 <= n5618;
    ng3965 <= n5623;
    ng6483 <= n5628;
    ng6187 <= n5633;
    ng914 <= n5638;
    ng5551 <= n5643;
    ng1373 <= n5648;
    ng5712 <= n5653;
    ng632 <= n5658;
    ng1246 <= n5663;
    ng4498 <= n5668;
    ng5805 <= n5672;
    ng2241 <= n5677;
    ng2370 <= n5682;
    ng5770 <= n5687;
    ng2756 <= n5692;
    ng3436 <= n5697;
    ng2514 <= n5702;
    ng2763 <= n5707;
    ng6645 <= n5712;
    ng3869 <= n5717;
    ng2629 <= n5722;
    ng45 <= n5727;
    ng4165 <= n5732;
    ng3639 <= n5737;
    ng269 <= n5742;
    ng3957 <= n5747;
    ng1183 <= n5752;
    ng5767 <= n5757;
    ng4669 <= n5762;
    ng4411 <= n5766;
    ng3602 <= n5771;
    ng4688 <= n5776;
    ng3227 <= n5781;
    ng4023 <= n5785;
    ng2040 <= n5789;
    ng3396 <= n5794;
    ng6077 <= n5799;
    ng3021 <= n5804;
    ng5857 <= n5809;
    ng8 <= n5814;
    ng550 <= n5819;
    ng283 <= n5824;
    ng2795 <= n5829;
    ng194 <= n5834;
    ng6049 <= n5838;
    ng4082 <= n5843;
    ng1252 <= n5848;
    ng5527 <= n5853;
    ng5224 <= n5858;
    ng1287 <= n5863;
    ng1644 <= n5868;
    ng5176 <= n5873;
    ng1536 <= n5878;
    ng5228 <= n5883;
    ng3849 <= n5888;
    ng2303 <= n5893;
    ng3096 <= n5898;
    ng324 <= n5902;
    ng6527 <= n5907;
    ng5644 <= n5912;
    ng1311 <= n5917;
    ng1239 <= n5921;
    ng3953 <= n5925;
    ng164 <= n5930;
    ng1648 <= n5935;
    ng929 <= n5940;
    ng6295 <= n5945;
    ng1792 <= n5950;
    ng2583 <= n5955;
    ng3416 <= n5960;
    ng3447 <= n5965;
    ng6462 <= n5969;
    ng278 <= n5974;
    ng6395 <= n5979;
    ng1422 <= n5983;
    ng763 <= n5988;
    ng1632 <= n5993;
    ng744 <= n5998;
    ng1442 <= n6003;
    ng1454 <= n6008;
    ng2287 <= n6013;
    ng3566 <= n6018;
    ng681 <= n6023;
    ng3518 <= n6028;
    ng736 <= n6033;
    ng5623 <= n6037;
    ng3835 <= n6041;
    ng5339 <= n6045;
    ng174 <= n6050;
    ng5742 <= n6055;
    ng2783 <= n6060;
    ng5983 <= n6065;
    ng6243 <= n6069;
    ng6128 <= n6074;
    ng16 <= n6079;
    ng239 <= n6084;
    ng4452 <= n6088;
    ng884 <= n6092;
    ng2152 <= n6096;
    ng5164 <= n6101;
    ng4226 <= n6105;
    ng2461 <= n6109;
    ng4369 <= n6114;
    ng3288 <= n6119;
    ng1263 <= n6124;
    ng4664 <= n6129;
    ng2047 <= n6134;
    ng4430 <= n6139;
    ng572 <= n6144;
    ng3990 <= n6149;
    ng812 <= n6154;
    ng3684 <= n6159;
    ng401 <= n6164;
    ng6151 <= n6169;
    ng586 <= n6174;
    ng2393 <= n6179;
    ng5428 <= n6184;
    ng5308 <= n6188;
    ng2587 <= n6192;
    ng6271 <= n6197;
    ng2020 <= n6202;
    ng460 <= n6207;
    ng3247 <= n6212;
    ng4210 <= n6216;
    ng199 <= n6220;
    ng5080 <= n6225;
    ng2965 <= n6230;
    ng1404 <= n6235;
    ng617 <= n6240;
    ng3161 <= n6245;
    ng1844 <= n6250;
    ng6109 <= n6255;
    ng1955 <= n6260;
    ng6419 <= n6265;
    ng671 <= n6270;
    ng1270 <= n6275;
    ng5925 <= n6280;
    ng2787 <= n6285;
    ng6601 <= n6290;
    ng4119 <= n6295;
    ng5845 <= n6300;
    ng6661 <= n6304;
    ng3550 <= n6308;
    ng1687 <= n6313;
    ng1710 <= n6318;
    ng5152 <= n6323;
    ng2060 <= n6328;
    ng3727 <= n6333;
    ng5046 <= n6338;
    ng4232 <= n6342;
    ng4519 <= n6347;
    ng3614 <= n6352;
    ng5272 <= n6357;
    ng4358 <= n6362;
    ng3003 <= n6367;
    ng5366 <= n6372;
    ng5260 <= n6377;
    ng4300 <= n6382;
    ng71 <= n6387;
    ng2299 <= n6392;
    ng4492 <= n6397;
    ng6137 <= n6402;
    ng3794 <= n6407;
    ng3905 <= n6411;
    ng5313 <= n6416;
    ng1917 <= n6420;
    ng5965 <= n6425;
    ng5933 <= n6430;
    ng5611 <= n6435;
    ng4534 <= n6440;
    ng417 <= n6445;
    ng1604 <= n6450;
    ng2008 <= n6455;
    ng2122 <= n6460;
    ng2433 <= n6465;
    ng4164 <= n6470;
    ng6637 <= n6475;
    ng3558 <= n6480;
    ng157 <= n6485;
    ng1459 <= n6489;
    ng5961 <= n6493;
    ng6629 <= n6498;
    ng5436 <= n6503;
    ng1216 <= n6508;
    ng1430 <= n6513;
    ng3742 <= n6518;
    ng5208 <= n6523;
    ng1333 <= n6527;
    ng101 <= n6532;
    ng5706 <= n6537;
    ng1816 <= n6542;
    ng2403 <= n6547;
    ng952 <= n6552;
    ng2223 <= n6557;
    ng5957 <= n6562;
    ng4188 <= n6566;
    ng2130 <= n6571;
    ng3706 <= n6576;
    ng832 <= n6581;
    ng2823 <= n6586;
    ng6040 <= n6591;
    ng1760 <= n6596;
    ng869 <= n6600;
    ng2193 <= n6604;
    ng996 <= n6609;
    ng4474 <= n6614;
    ng4480 <= n6619;
    ng3582 <= n6624;
    ng4000 <= n6628;
    ng5467 <= n6632;
    ng4608 <= n6637;
    ng1894 <= n6642;
    ng5011 <= n6647;
    ng5863 <= n6652;
    ng6444 <= n6657;
    ng3723 <= n6662;
    ng5220 <= n6667;
    ng2384 <= n6672;
    ng4527 <= n6677;
    ng1489 <= n6682;
    ng4277 <= n6687;
    ng3347 <= n6691;
    ng2265 <= n6696;
    ng1974 <= n6701;
    ng1124 <= n6706;
    ng2429 <= n6711;
    ng1978 <= n6716;
    ng6390 <= n6721;
    ng3199 <= n6726;
    ng3065 <= n6731;
    ng1740 <= n6736;
    ng2681 <= n6741;
    ng2413 <= n6746;
    ng5352 <= n6751;
    ng6617 <= n6756;
    ng2704 <= n6761;
    ng2250 <= n6766;
    ng2357 <= n6771;
    ng5115 <= n6776;
    ng5595 <= n6781;
    ng2735 <= n6786;
    ng4659 <= n6791;
    ng1094 <= n6796;
    ng534 <= n6801;
    ng1521 <= n6806;
    ng4204 <= n6810;
    ng59 <= n6814;
    ng772 <= n6819;
    ng2563 <= n6824;
    ng3598 <= n6829;
    ng294 <= n6834;
    ng921 <= n6839;
    ng3522 <= n6844;
    ng1379 <= n6849;
    ng5587 <= n6854;
    ng1500 <= n6859;
    ng4264 <= n6863;
    ng6291 <= n6868;
    ng2955 <= n6873;
    ng3115 <= n6878;
    ng1724 <= n6883;
    ng6177 <= n6888;
    ng4593 <= n6893;
    ng1024 <= n6898;
    ng3625 <= n6902;
    ng203 <= n6907;
    ng5057 <= n6912;
    ng6377 <= n6916;
    ng4776 <= n6921;
    ng5591 <= n6926;
    ng5507 <= n6931;
    ng6088 <= n6936;
    ng452 <= n6941;
    ng807 <= n6946;
    ng1600 <= n6951;
    ng4621 <= n6956;
    ng1099 <= n6961;
    ng2024 <= n6966;
    ng901 <= n6971;
    ng4242 <= n6976;
    ng2741 <= n6981;
    ng2217 <= n6986;
    ng464 <= n6991;
    ng6219 <= n6996;
    ng1714 <= n7001;
    ng1968 <= n7006;
    ng4878 <= n7011;
    ng3303 <= n7016;
    ng4194 <= n7019;
    ng5503 <= n7023;
    ng802 <= n7027;
    ng595 <= n7031;
    ng3542 <= n7036;
    ng847 <= n7041;
    ng6005 <= n7046;
    ng1736 <= n7050;
    ng47 <= n7055;
    ng2389 <= n7060;
    ng3782 <= n7065;
    ng2638 <= n7070;
    ng2066 <= n7075;
    ng4258 <= n7080;
    ng5232 <= n7085;
    ng6031 <= n7089;
    ng4235 <= n7093;
    ng6073 <= n7098;
    ng3147 <= n7103;
    ng4438 <= n7108;
    ng5547 <= n7113;
    ng4122 <= n7118;
    ng1319 <= n7123;
    ng1612 <= n7128;
    ng5813 <= n7133;
    ng4172 <= n7138;
    ng3355 <= n7143;
    ng490 <= n7148;
    ng3457 <= n7153;
    ng2844 <= n7158;
    ng4709 <= n7163;
    ng1291 <= n7168;
    ng2449 <= n7173;
    ng5212 <= n7178;
    ng1830 <= n7183;
    ng6474 <= n7188;
    ng4408 <= n7193;
    ng3376 <= n7198;
    ng2907 <= n7203;
    ng976 <= n7208;
    ng2236 <= n7213;
    ng5659 <= n7218;
    ng6287 <= n7222;
    ng5180 <= n7227;
    ng918 <= n7232;
    ng5945 <= n7237;
    ng5517 <= n7242;
    ng4245 <= n7247;
    ng2246 <= n7252;
    ng1932 <= n7257;
    ng1576 <= n7262;
    ng3941 <= n7266;
    ng1744 <= n7271;
    ng3512 <= n7276;
    ng3649 <= n7280;
    ng2657 <= n7284;
    ng4933 <= n7289;
    ng608 <= n7294;
    ng5782 <= n7299;
    ng1886 <= n7304;
    ng1008 <= n7309;
    ng645 <= n7314;
    ng392 <= n7319;
    ng146 <= n7324;
    ng2671 <= n7329;
    ng6565 <= n7334;
    ng5909 <= n7339;
    ng4372 <= n7344;
    ng3155 <= n7349;
    ng5607 <= n7354;
    ng4521 <= n7359;
    ng562 <= n7364;
    ng6105 <= n7369;
    ng6466 <= n7374;
    ng6133 <= n7379;
    ng4291 <= n7383;
    ng3590 <= n7388;
    ng218 <= n7392;
    ng2028 <= n7397;
    ng2685 <= n7402;
    ng1802 <= n7407;
    ng3490 <= n7412;
    ng3167 <= n7417;
    ng2295 <= n7422;
    ng3321 <= n7426;
    ng3813 <= n7430;
    ng1205 <= n7435;
    ng2208 <= n7440;
    ng732 <= n7445;
    ng968 <= n7450;
    ng4176 <= n7455;
    ng6263 <= n7460;
    ng4540 <= n7465;
    ng121 <= n7470;
    ng6732 <= n7475;
    ng3554 <= n7480;
    ng749 <= n7485;
    ng5615 <= n7490;
    ng6199 <= n7495;
    ng2089 <= n7500;
    ng6144 <= n7505;
    ng3909 <= n7509;
    ng2917 <= n7514;
    ng2504 <= n7519;
    ng6093 <= n7524;
    ng4005 <= n7529;
    ng2331 <= n7533;
    ng6723 <= n7537;
    ng6585 <= n7542;
    ng6633 <= n7547;
    ng4555 <= n7551;
    ng6069 <= n7556;
    ng4567 <= n7561;
    ng1339 <= n7566;
    ng767 <= n7571;
    ng5794 <= n7576;
    ng6259 <= n7580;
    ng4405 <= n7584;
    ng3945 <= n7589;
    ng2748 <= n7594;
    ng2283 <= n7599;
    ng1426 <= n7603;
    ng3698 <= n7607;
    ng311 <= n7612;
    ng3057 <= n7617;
    ng1384 <= n7622;
    ng5853 <= n7627;
    ng5559 <= n7632;
    ng5905 <= n7637;
    ng872 <= n7641;
    ng50 <= n7646;
    ng5471 <= n7651;
    ng2169 <= n7656;
    ng5005 <= n7660;
  end
endmodule

