// Benchmark "testing" written by ABC on Thu Oct  8 22:16:31 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A74  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A74;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[209]_ ,
    \new_[210]_ , \new_[214]_ , \new_[215]_ , \new_[216]_ , \new_[220]_ ,
    \new_[221]_ , \new_[225]_ , \new_[226]_ , \new_[227]_ , \new_[228]_ ,
    \new_[232]_ , \new_[233]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ ,
    \new_[243]_ , \new_[244]_ , \new_[247]_ , \new_[250]_ , \new_[251]_ ,
    \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[258]_ , \new_[259]_ ,
    \new_[263]_ , \new_[264]_ , \new_[265]_ , \new_[269]_ , \new_[270]_ ,
    \new_[273]_ , \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ ,
    \new_[283]_ , \new_[284]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[294]_ , \new_[295]_ , \new_[298]_ , \new_[301]_ , \new_[302]_ ,
    \new_[303]_ , \new_[304]_ , \new_[305]_ , \new_[306]_ , \new_[310]_ ,
    \new_[311]_ , \new_[315]_ , \new_[316]_ , \new_[317]_ , \new_[321]_ ,
    \new_[322]_ , \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ ,
    \new_[333]_ , \new_[334]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[344]_ , \new_[345]_ , \new_[348]_ , \new_[351]_ , \new_[352]_ ,
    \new_[353]_ , \new_[354]_ , \new_[355]_ , \new_[359]_ , \new_[360]_ ,
    \new_[364]_ , \new_[365]_ , \new_[366]_ , \new_[370]_ , \new_[371]_ ,
    \new_[374]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[384]_ , \new_[385]_ , \new_[389]_ , \new_[390]_ , \new_[391]_ ,
    \new_[395]_ , \new_[396]_ , \new_[399]_ , \new_[402]_ , \new_[403]_ ,
    \new_[404]_ , \new_[405]_ , \new_[406]_ , \new_[407]_ , \new_[408]_ ,
    \new_[412]_ , \new_[413]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ ,
    \new_[423]_ , \new_[424]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[435]_ , \new_[436]_ , \new_[440]_ , \new_[441]_ ,
    \new_[442]_ , \new_[446]_ , \new_[447]_ , \new_[450]_ , \new_[453]_ ,
    \new_[454]_ , \new_[455]_ , \new_[456]_ , \new_[457]_ , \new_[461]_ ,
    \new_[462]_ , \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[472]_ ,
    \new_[473]_ , \new_[476]_ , \new_[479]_ , \new_[480]_ , \new_[481]_ ,
    \new_[482]_ , \new_[486]_ , \new_[487]_ , \new_[491]_ , \new_[492]_ ,
    \new_[493]_ , \new_[497]_ , \new_[498]_ , \new_[501]_ , \new_[504]_ ,
    \new_[505]_ , \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ ,
    \new_[513]_ , \new_[514]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[524]_ , \new_[525]_ , \new_[528]_ , \new_[531]_ , \new_[532]_ ,
    \new_[533]_ , \new_[534]_ , \new_[538]_ , \new_[539]_ , \new_[543]_ ,
    \new_[544]_ , \new_[545]_ , \new_[549]_ , \new_[550]_ , \new_[553]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[564]_ , \new_[565]_ , \new_[569]_ , \new_[570]_ , \new_[571]_ ,
    \new_[575]_ , \new_[576]_ , \new_[579]_ , \new_[582]_ , \new_[583]_ ,
    \new_[584]_ , \new_[585]_ , \new_[589]_ , \new_[590]_ , \new_[594]_ ,
    \new_[595]_ , \new_[596]_ , \new_[600]_ , \new_[601]_ , \new_[604]_ ,
    \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ , \new_[611]_ ,
    \new_[612]_ , \new_[613]_ , \new_[625]_ , \new_[629]_ , \new_[633]_ ,
    \new_[637]_ , \new_[641]_ , \new_[645]_ , \new_[649]_ , \new_[653]_ ,
    \new_[657]_ , \new_[661]_ , \new_[664]_ , \new_[667]_ , \new_[670]_ ,
    \new_[673]_ , \new_[676]_ , \new_[679]_ , \new_[682]_ , \new_[685]_ ,
    \new_[688]_ , \new_[691]_ , \new_[694]_ , \new_[697]_ , \new_[700]_ ,
    \new_[703]_ , \new_[706]_ , \new_[709]_ , \new_[712]_ , \new_[715]_ ,
    \new_[718]_ , \new_[721]_ , \new_[724]_ , \new_[727]_ , \new_[730]_ ,
    \new_[733]_ , \new_[736]_ , \new_[739]_ , \new_[742]_ , \new_[745]_ ,
    \new_[748]_ , \new_[751]_ , \new_[754]_ , \new_[757]_ , \new_[760]_ ,
    \new_[764]_ , \new_[765]_ , \new_[768]_ , \new_[772]_ , \new_[773]_ ,
    \new_[776]_ , \new_[780]_ , \new_[781]_ , \new_[784]_ , \new_[788]_ ,
    \new_[789]_ , \new_[792]_ , \new_[796]_ , \new_[797]_ , \new_[800]_ ,
    \new_[804]_ , \new_[805]_ , \new_[808]_ , \new_[812]_ , \new_[813]_ ,
    \new_[816]_ , \new_[820]_ , \new_[821]_ , \new_[824]_ , \new_[828]_ ,
    \new_[829]_ , \new_[832]_ , \new_[836]_ , \new_[837]_ , \new_[840]_ ,
    \new_[844]_ , \new_[845]_ , \new_[848]_ , \new_[852]_ , \new_[853]_ ,
    \new_[856]_ , \new_[860]_ , \new_[861]_ , \new_[864]_ , \new_[868]_ ,
    \new_[869]_ , \new_[872]_ , \new_[876]_ , \new_[877]_ , \new_[880]_ ,
    \new_[884]_ , \new_[885]_ , \new_[888]_ , \new_[892]_ , \new_[893]_ ,
    \new_[896]_ , \new_[900]_ , \new_[901]_ , \new_[904]_ , \new_[908]_ ,
    \new_[909]_ , \new_[912]_ , \new_[916]_ , \new_[917]_ , \new_[921]_ ,
    \new_[922]_ , \new_[926]_ , \new_[927]_ , \new_[931]_ , \new_[932]_ ,
    \new_[936]_ , \new_[937]_ , \new_[941]_ , \new_[942]_ , \new_[946]_ ,
    \new_[947]_ , \new_[951]_ , \new_[952]_ , \new_[956]_ , \new_[957]_ ,
    \new_[961]_ , \new_[962]_ , \new_[966]_ , \new_[967]_ , \new_[971]_ ,
    \new_[972]_ , \new_[976]_ , \new_[977]_ , \new_[981]_ , \new_[982]_ ,
    \new_[986]_ , \new_[987]_ , \new_[991]_ , \new_[992]_ , \new_[996]_ ,
    \new_[997]_ , \new_[1001]_ , \new_[1002]_ , \new_[1006]_ ,
    \new_[1007]_ , \new_[1011]_ , \new_[1012]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1021]_ , \new_[1022]_ , \new_[1026]_ ,
    \new_[1027]_ , \new_[1031]_ , \new_[1032]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1041]_ , \new_[1042]_ , \new_[1046]_ ,
    \new_[1047]_ , \new_[1051]_ , \new_[1052]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1061]_ , \new_[1062]_ , \new_[1066]_ ,
    \new_[1067]_ , \new_[1071]_ , \new_[1072]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1081]_ , \new_[1082]_ , \new_[1086]_ ,
    \new_[1087]_ , \new_[1091]_ , \new_[1092]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1101]_ , \new_[1102]_ , \new_[1106]_ ,
    \new_[1107]_ , \new_[1111]_ , \new_[1112]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1121]_ , \new_[1122]_ , \new_[1126]_ ,
    \new_[1127]_ , \new_[1131]_ , \new_[1132]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1141]_ , \new_[1142]_ , \new_[1146]_ ,
    \new_[1147]_ , \new_[1151]_ , \new_[1152]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1161]_ , \new_[1162]_ , \new_[1166]_ ,
    \new_[1167]_ , \new_[1171]_ , \new_[1172]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1181]_ , \new_[1182]_ , \new_[1185]_ ,
    \new_[1188]_ , \new_[1189]_ , \new_[1193]_ , \new_[1194]_ ,
    \new_[1197]_ , \new_[1200]_ , \new_[1201]_ , \new_[1205]_ ,
    \new_[1206]_ , \new_[1209]_ , \new_[1212]_ , \new_[1213]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1221]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1229]_ , \new_[1230]_ , \new_[1233]_ ,
    \new_[1236]_ , \new_[1237]_ , \new_[1241]_ , \new_[1242]_ ,
    \new_[1245]_ , \new_[1248]_ , \new_[1249]_ , \new_[1253]_ ,
    \new_[1254]_ , \new_[1257]_ , \new_[1260]_ , \new_[1261]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1269]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1277]_ , \new_[1278]_ , \new_[1281]_ ,
    \new_[1284]_ , \new_[1285]_ , \new_[1289]_ , \new_[1290]_ ,
    \new_[1293]_ , \new_[1296]_ , \new_[1297]_ , \new_[1301]_ ,
    \new_[1302]_ , \new_[1305]_ , \new_[1308]_ , \new_[1309]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1317]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1325]_ , \new_[1326]_ , \new_[1329]_ ,
    \new_[1332]_ , \new_[1333]_ , \new_[1337]_ , \new_[1338]_ ,
    \new_[1341]_ , \new_[1344]_ , \new_[1345]_ , \new_[1349]_ ,
    \new_[1350]_ , \new_[1353]_ , \new_[1356]_ , \new_[1357]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1365]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1373]_ , \new_[1374]_ , \new_[1377]_ ,
    \new_[1380]_ , \new_[1381]_ , \new_[1385]_ , \new_[1386]_ ,
    \new_[1389]_ , \new_[1392]_ , \new_[1393]_ , \new_[1397]_ ,
    \new_[1398]_ , \new_[1401]_ , \new_[1404]_ , \new_[1405]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1413]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1421]_ , \new_[1422]_ , \new_[1425]_ ,
    \new_[1428]_ , \new_[1429]_ , \new_[1433]_ , \new_[1434]_ ,
    \new_[1437]_ , \new_[1440]_ , \new_[1441]_ , \new_[1445]_ ,
    \new_[1446]_ , \new_[1449]_ , \new_[1452]_ , \new_[1453]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1461]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1469]_ , \new_[1470]_ , \new_[1473]_ ,
    \new_[1476]_ , \new_[1477]_ , \new_[1481]_ , \new_[1482]_ ,
    \new_[1485]_ , \new_[1488]_ , \new_[1489]_ , \new_[1493]_ ,
    \new_[1494]_ , \new_[1497]_ , \new_[1500]_ , \new_[1501]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1509]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1517]_ , \new_[1518]_ , \new_[1521]_ ,
    \new_[1524]_ , \new_[1525]_ , \new_[1529]_ , \new_[1530]_ ,
    \new_[1533]_ , \new_[1536]_ , \new_[1537]_ , \new_[1541]_ ,
    \new_[1542]_ , \new_[1545]_ , \new_[1548]_ , \new_[1549]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1557]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1565]_ , \new_[1566]_ , \new_[1569]_ ,
    \new_[1572]_ , \new_[1573]_ , \new_[1577]_ , \new_[1578]_ ,
    \new_[1581]_ , \new_[1584]_ , \new_[1585]_ , \new_[1589]_ ,
    \new_[1590]_ , \new_[1593]_ , \new_[1596]_ , \new_[1597]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1605]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1613]_ , \new_[1614]_ , \new_[1617]_ ,
    \new_[1620]_ , \new_[1621]_ , \new_[1625]_ , \new_[1626]_ ,
    \new_[1629]_ , \new_[1632]_ , \new_[1633]_ , \new_[1637]_ ,
    \new_[1638]_ , \new_[1641]_ , \new_[1644]_ , \new_[1645]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1653]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1660]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1667]_ , \new_[1670]_ , \new_[1671]_ , \new_[1674]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1681]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1688]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1695]_ , \new_[1698]_ , \new_[1699]_ , \new_[1702]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1709]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1716]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1723]_ , \new_[1726]_ , \new_[1727]_ , \new_[1730]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1737]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1744]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1751]_ , \new_[1754]_ , \new_[1755]_ , \new_[1758]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1765]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1772]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1779]_ , \new_[1782]_ , \new_[1783]_ , \new_[1786]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1793]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1800]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1807]_ , \new_[1810]_ , \new_[1811]_ , \new_[1814]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1821]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1828]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1835]_ , \new_[1838]_ , \new_[1839]_ , \new_[1842]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1849]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1856]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1863]_ , \new_[1866]_ , \new_[1867]_ , \new_[1870]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1877]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1884]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1891]_ , \new_[1894]_ , \new_[1895]_ , \new_[1898]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1905]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1912]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1919]_ , \new_[1922]_ , \new_[1923]_ , \new_[1926]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1933]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1940]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1947]_ , \new_[1950]_ , \new_[1951]_ , \new_[1954]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1961]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1968]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1975]_ , \new_[1978]_ , \new_[1979]_ , \new_[1982]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1989]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1996]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2003]_ , \new_[2006]_ , \new_[2007]_ , \new_[2010]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2017]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2024]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2031]_ , \new_[2034]_ , \new_[2035]_ , \new_[2038]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2045]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2052]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2059]_ , \new_[2062]_ , \new_[2063]_ , \new_[2066]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2073]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2080]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2087]_ , \new_[2090]_ , \new_[2091]_ , \new_[2094]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2101]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2108]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2115]_ , \new_[2118]_ , \new_[2119]_ , \new_[2122]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2129]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2136]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2143]_ , \new_[2146]_ , \new_[2147]_ , \new_[2150]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2157]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2164]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2171]_ , \new_[2174]_ , \new_[2175]_ , \new_[2178]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2185]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2192]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2199]_ , \new_[2202]_ , \new_[2203]_ , \new_[2206]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2213]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2220]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2227]_ , \new_[2230]_ , \new_[2231]_ , \new_[2234]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2241]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2248]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2255]_ , \new_[2258]_ , \new_[2259]_ , \new_[2262]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2269]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2276]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2283]_ , \new_[2286]_ , \new_[2287]_ , \new_[2290]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2297]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2304]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2311]_ , \new_[2314]_ , \new_[2315]_ , \new_[2318]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2325]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2332]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2339]_ , \new_[2343]_ , \new_[2344]_ , \new_[2345]_ ,
    \new_[2348]_ , \new_[2351]_ , \new_[2352]_ , \new_[2355]_ ,
    \new_[2359]_ , \new_[2360]_ , \new_[2361]_ , \new_[2364]_ ,
    \new_[2367]_ , \new_[2368]_ , \new_[2371]_ , \new_[2375]_ ,
    \new_[2376]_ , \new_[2377]_ , \new_[2380]_ , \new_[2383]_ ,
    \new_[2384]_ , \new_[2387]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2396]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2403]_ , \new_[2407]_ , \new_[2408]_ , \new_[2409]_ ,
    \new_[2412]_ , \new_[2415]_ , \new_[2416]_ , \new_[2419]_ ,
    \new_[2423]_ , \new_[2424]_ , \new_[2425]_ , \new_[2428]_ ,
    \new_[2431]_ , \new_[2432]_ , \new_[2435]_ , \new_[2439]_ ,
    \new_[2440]_ , \new_[2441]_ , \new_[2444]_ , \new_[2447]_ ,
    \new_[2448]_ , \new_[2451]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2460]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2467]_ , \new_[2471]_ , \new_[2472]_ , \new_[2473]_ ,
    \new_[2476]_ , \new_[2479]_ , \new_[2480]_ , \new_[2483]_ ,
    \new_[2487]_ , \new_[2488]_ , \new_[2489]_ , \new_[2492]_ ,
    \new_[2495]_ , \new_[2496]_ , \new_[2499]_ , \new_[2503]_ ,
    \new_[2504]_ , \new_[2505]_ , \new_[2508]_ , \new_[2511]_ ,
    \new_[2512]_ , \new_[2515]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2524]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2531]_ , \new_[2535]_ , \new_[2536]_ , \new_[2537]_ ,
    \new_[2540]_ , \new_[2543]_ , \new_[2544]_ , \new_[2547]_ ,
    \new_[2551]_ , \new_[2552]_ , \new_[2553]_ , \new_[2556]_ ,
    \new_[2559]_ , \new_[2560]_ , \new_[2563]_ , \new_[2567]_ ,
    \new_[2568]_ , \new_[2569]_ , \new_[2572]_ , \new_[2575]_ ,
    \new_[2576]_ , \new_[2579]_ , \new_[2583]_ , \new_[2584]_ ,
    \new_[2585]_ , \new_[2588]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2595]_ , \new_[2599]_ , \new_[2600]_ , \new_[2601]_ ,
    \new_[2604]_ , \new_[2607]_ , \new_[2608]_ , \new_[2611]_ ,
    \new_[2615]_ , \new_[2616]_ , \new_[2617]_ , \new_[2620]_ ,
    \new_[2623]_ , \new_[2624]_ , \new_[2627]_ , \new_[2631]_ ,
    \new_[2632]_ , \new_[2633]_ , \new_[2636]_ , \new_[2639]_ ,
    \new_[2640]_ , \new_[2643]_ , \new_[2647]_ , \new_[2648]_ ,
    \new_[2649]_ , \new_[2652]_ , \new_[2655]_ , \new_[2656]_ ,
    \new_[2659]_ , \new_[2663]_ , \new_[2664]_ , \new_[2665]_ ,
    \new_[2668]_ , \new_[2671]_ , \new_[2672]_ , \new_[2675]_ ,
    \new_[2679]_ , \new_[2680]_ , \new_[2681]_ , \new_[2684]_ ,
    \new_[2687]_ , \new_[2688]_ , \new_[2691]_ , \new_[2695]_ ,
    \new_[2696]_ , \new_[2697]_ , \new_[2700]_ , \new_[2703]_ ,
    \new_[2704]_ , \new_[2707]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2716]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2723]_ , \new_[2727]_ , \new_[2728]_ , \new_[2729]_ ,
    \new_[2732]_ , \new_[2735]_ , \new_[2736]_ , \new_[2739]_ ,
    \new_[2743]_ , \new_[2744]_ , \new_[2745]_ , \new_[2748]_ ,
    \new_[2751]_ , \new_[2752]_ , \new_[2755]_ , \new_[2759]_ ,
    \new_[2760]_ , \new_[2761]_ , \new_[2764]_ , \new_[2767]_ ,
    \new_[2768]_ , \new_[2771]_ , \new_[2775]_ , \new_[2776]_ ,
    \new_[2777]_ , \new_[2780]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2787]_ , \new_[2791]_ , \new_[2792]_ , \new_[2793]_ ,
    \new_[2796]_ , \new_[2799]_ , \new_[2800]_ , \new_[2803]_ ,
    \new_[2807]_ , \new_[2808]_ , \new_[2809]_ , \new_[2812]_ ,
    \new_[2815]_ , \new_[2816]_ , \new_[2819]_ , \new_[2823]_ ,
    \new_[2824]_ , \new_[2825]_ , \new_[2828]_ , \new_[2831]_ ,
    \new_[2832]_ , \new_[2835]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2844]_ , \new_[2848]_ , \new_[2849]_ ,
    \new_[2850]_ , \new_[2853]_ , \new_[2857]_ , \new_[2858]_ ,
    \new_[2859]_ , \new_[2862]_ , \new_[2866]_ , \new_[2867]_ ,
    \new_[2868]_ , \new_[2871]_ , \new_[2875]_ , \new_[2876]_ ,
    \new_[2877]_ , \new_[2880]_ , \new_[2884]_ , \new_[2885]_ ,
    \new_[2886]_ , \new_[2889]_ , \new_[2893]_ , \new_[2894]_ ,
    \new_[2895]_ , \new_[2898]_ , \new_[2902]_ , \new_[2903]_ ,
    \new_[2904]_ , \new_[2907]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2916]_ , \new_[2920]_ , \new_[2921]_ ,
    \new_[2922]_ , \new_[2925]_ , \new_[2929]_ , \new_[2930]_ ,
    \new_[2931]_ , \new_[2934]_ , \new_[2938]_ , \new_[2939]_ ,
    \new_[2940]_ , \new_[2943]_ , \new_[2947]_ , \new_[2948]_ ,
    \new_[2949]_ , \new_[2952]_ , \new_[2956]_ , \new_[2957]_ ,
    \new_[2958]_ , \new_[2961]_ , \new_[2965]_ , \new_[2966]_ ,
    \new_[2967]_ , \new_[2970]_ , \new_[2974]_ , \new_[2975]_ ,
    \new_[2976]_ , \new_[2979]_ , \new_[2983]_ , \new_[2984]_ ,
    \new_[2985]_ ;
  assign A74 = \new_[613]_  | \new_[408]_ ;
  assign \new_[1]_  = \new_[2985]_  & \new_[2976]_ ;
  assign \new_[2]_  = \new_[2967]_  & \new_[2958]_ ;
  assign \new_[3]_  = \new_[2949]_  & \new_[2940]_ ;
  assign \new_[4]_  = \new_[2931]_  & \new_[2922]_ ;
  assign \new_[5]_  = \new_[2913]_  & \new_[2904]_ ;
  assign \new_[6]_  = \new_[2895]_  & \new_[2886]_ ;
  assign \new_[7]_  = \new_[2877]_  & \new_[2868]_ ;
  assign \new_[8]_  = \new_[2859]_  & \new_[2850]_ ;
  assign \new_[9]_  = \new_[2841]_  & \new_[2832]_ ;
  assign \new_[10]_  = \new_[2825]_  & \new_[2816]_ ;
  assign \new_[11]_  = \new_[2809]_  & \new_[2800]_ ;
  assign \new_[12]_  = \new_[2793]_  & \new_[2784]_ ;
  assign \new_[13]_  = \new_[2777]_  & \new_[2768]_ ;
  assign \new_[14]_  = \new_[2761]_  & \new_[2752]_ ;
  assign \new_[15]_  = \new_[2745]_  & \new_[2736]_ ;
  assign \new_[16]_  = \new_[2729]_  & \new_[2720]_ ;
  assign \new_[17]_  = \new_[2713]_  & \new_[2704]_ ;
  assign \new_[18]_  = \new_[2697]_  & \new_[2688]_ ;
  assign \new_[19]_  = \new_[2681]_  & \new_[2672]_ ;
  assign \new_[20]_  = \new_[2665]_  & \new_[2656]_ ;
  assign \new_[21]_  = \new_[2649]_  & \new_[2640]_ ;
  assign \new_[22]_  = \new_[2633]_  & \new_[2624]_ ;
  assign \new_[23]_  = \new_[2617]_  & \new_[2608]_ ;
  assign \new_[24]_  = \new_[2601]_  & \new_[2592]_ ;
  assign \new_[25]_  = \new_[2585]_  & \new_[2576]_ ;
  assign \new_[26]_  = \new_[2569]_  & \new_[2560]_ ;
  assign \new_[27]_  = \new_[2553]_  & \new_[2544]_ ;
  assign \new_[28]_  = \new_[2537]_  & \new_[2528]_ ;
  assign \new_[29]_  = \new_[2521]_  & \new_[2512]_ ;
  assign \new_[30]_  = \new_[2505]_  & \new_[2496]_ ;
  assign \new_[31]_  = \new_[2489]_  & \new_[2480]_ ;
  assign \new_[32]_  = \new_[2473]_  & \new_[2464]_ ;
  assign \new_[33]_  = \new_[2457]_  & \new_[2448]_ ;
  assign \new_[34]_  = \new_[2441]_  & \new_[2432]_ ;
  assign \new_[35]_  = \new_[2425]_  & \new_[2416]_ ;
  assign \new_[36]_  = \new_[2409]_  & \new_[2400]_ ;
  assign \new_[37]_  = \new_[2393]_  & \new_[2384]_ ;
  assign \new_[38]_  = \new_[2377]_  & \new_[2368]_ ;
  assign \new_[39]_  = \new_[2361]_  & \new_[2352]_ ;
  assign \new_[40]_  = \new_[2345]_  & \new_[2336]_ ;
  assign \new_[41]_  = \new_[2329]_  & \new_[2322]_ ;
  assign \new_[42]_  = \new_[2315]_  & \new_[2308]_ ;
  assign \new_[43]_  = \new_[2301]_  & \new_[2294]_ ;
  assign \new_[44]_  = \new_[2287]_  & \new_[2280]_ ;
  assign \new_[45]_  = \new_[2273]_  & \new_[2266]_ ;
  assign \new_[46]_  = \new_[2259]_  & \new_[2252]_ ;
  assign \new_[47]_  = \new_[2245]_  & \new_[2238]_ ;
  assign \new_[48]_  = \new_[2231]_  & \new_[2224]_ ;
  assign \new_[49]_  = \new_[2217]_  & \new_[2210]_ ;
  assign \new_[50]_  = \new_[2203]_  & \new_[2196]_ ;
  assign \new_[51]_  = \new_[2189]_  & \new_[2182]_ ;
  assign \new_[52]_  = \new_[2175]_  & \new_[2168]_ ;
  assign \new_[53]_  = \new_[2161]_  & \new_[2154]_ ;
  assign \new_[54]_  = \new_[2147]_  & \new_[2140]_ ;
  assign \new_[55]_  = \new_[2133]_  & \new_[2126]_ ;
  assign \new_[56]_  = \new_[2119]_  & \new_[2112]_ ;
  assign \new_[57]_  = \new_[2105]_  & \new_[2098]_ ;
  assign \new_[58]_  = \new_[2091]_  & \new_[2084]_ ;
  assign \new_[59]_  = \new_[2077]_  & \new_[2070]_ ;
  assign \new_[60]_  = \new_[2063]_  & \new_[2056]_ ;
  assign \new_[61]_  = \new_[2049]_  & \new_[2042]_ ;
  assign \new_[62]_  = \new_[2035]_  & \new_[2028]_ ;
  assign \new_[63]_  = \new_[2021]_  & \new_[2014]_ ;
  assign \new_[64]_  = \new_[2007]_  & \new_[2000]_ ;
  assign \new_[65]_  = \new_[1993]_  & \new_[1986]_ ;
  assign \new_[66]_  = \new_[1979]_  & \new_[1972]_ ;
  assign \new_[67]_  = \new_[1965]_  & \new_[1958]_ ;
  assign \new_[68]_  = \new_[1951]_  & \new_[1944]_ ;
  assign \new_[69]_  = \new_[1937]_  & \new_[1930]_ ;
  assign \new_[70]_  = \new_[1923]_  & \new_[1916]_ ;
  assign \new_[71]_  = \new_[1909]_  & \new_[1902]_ ;
  assign \new_[72]_  = \new_[1895]_  & \new_[1888]_ ;
  assign \new_[73]_  = \new_[1881]_  & \new_[1874]_ ;
  assign \new_[74]_  = \new_[1867]_  & \new_[1860]_ ;
  assign \new_[75]_  = \new_[1853]_  & \new_[1846]_ ;
  assign \new_[76]_  = \new_[1839]_  & \new_[1832]_ ;
  assign \new_[77]_  = \new_[1825]_  & \new_[1818]_ ;
  assign \new_[78]_  = \new_[1811]_  & \new_[1804]_ ;
  assign \new_[79]_  = \new_[1797]_  & \new_[1790]_ ;
  assign \new_[80]_  = \new_[1783]_  & \new_[1776]_ ;
  assign \new_[81]_  = \new_[1769]_  & \new_[1762]_ ;
  assign \new_[82]_  = \new_[1755]_  & \new_[1748]_ ;
  assign \new_[83]_  = \new_[1741]_  & \new_[1734]_ ;
  assign \new_[84]_  = \new_[1727]_  & \new_[1720]_ ;
  assign \new_[85]_  = \new_[1713]_  & \new_[1706]_ ;
  assign \new_[86]_  = \new_[1699]_  & \new_[1692]_ ;
  assign \new_[87]_  = \new_[1685]_  & \new_[1678]_ ;
  assign \new_[88]_  = \new_[1671]_  & \new_[1664]_ ;
  assign \new_[89]_  = \new_[1657]_  & \new_[1650]_ ;
  assign \new_[90]_  = \new_[1645]_  & \new_[1638]_ ;
  assign \new_[91]_  = \new_[1633]_  & \new_[1626]_ ;
  assign \new_[92]_  = \new_[1621]_  & \new_[1614]_ ;
  assign \new_[93]_  = \new_[1609]_  & \new_[1602]_ ;
  assign \new_[94]_  = \new_[1597]_  & \new_[1590]_ ;
  assign \new_[95]_  = \new_[1585]_  & \new_[1578]_ ;
  assign \new_[96]_  = \new_[1573]_  & \new_[1566]_ ;
  assign \new_[97]_  = \new_[1561]_  & \new_[1554]_ ;
  assign \new_[98]_  = \new_[1549]_  & \new_[1542]_ ;
  assign \new_[99]_  = \new_[1537]_  & \new_[1530]_ ;
  assign \new_[100]_  = \new_[1525]_  & \new_[1518]_ ;
  assign \new_[101]_  = \new_[1513]_  & \new_[1506]_ ;
  assign \new_[102]_  = \new_[1501]_  & \new_[1494]_ ;
  assign \new_[103]_  = \new_[1489]_  & \new_[1482]_ ;
  assign \new_[104]_  = \new_[1477]_  & \new_[1470]_ ;
  assign \new_[105]_  = \new_[1465]_  & \new_[1458]_ ;
  assign \new_[106]_  = \new_[1453]_  & \new_[1446]_ ;
  assign \new_[107]_  = \new_[1441]_  & \new_[1434]_ ;
  assign \new_[108]_  = \new_[1429]_  & \new_[1422]_ ;
  assign \new_[109]_  = \new_[1417]_  & \new_[1410]_ ;
  assign \new_[110]_  = \new_[1405]_  & \new_[1398]_ ;
  assign \new_[111]_  = \new_[1393]_  & \new_[1386]_ ;
  assign \new_[112]_  = \new_[1381]_  & \new_[1374]_ ;
  assign \new_[113]_  = \new_[1369]_  & \new_[1362]_ ;
  assign \new_[114]_  = \new_[1357]_  & \new_[1350]_ ;
  assign \new_[115]_  = \new_[1345]_  & \new_[1338]_ ;
  assign \new_[116]_  = \new_[1333]_  & \new_[1326]_ ;
  assign \new_[117]_  = \new_[1321]_  & \new_[1314]_ ;
  assign \new_[118]_  = \new_[1309]_  & \new_[1302]_ ;
  assign \new_[119]_  = \new_[1297]_  & \new_[1290]_ ;
  assign \new_[120]_  = \new_[1285]_  & \new_[1278]_ ;
  assign \new_[121]_  = \new_[1273]_  & \new_[1266]_ ;
  assign \new_[122]_  = \new_[1261]_  & \new_[1254]_ ;
  assign \new_[123]_  = \new_[1249]_  & \new_[1242]_ ;
  assign \new_[124]_  = \new_[1237]_  & \new_[1230]_ ;
  assign \new_[125]_  = \new_[1225]_  & \new_[1218]_ ;
  assign \new_[126]_  = \new_[1213]_  & \new_[1206]_ ;
  assign \new_[127]_  = \new_[1201]_  & \new_[1194]_ ;
  assign \new_[128]_  = \new_[1189]_  & \new_[1182]_ ;
  assign \new_[129]_  = \new_[1177]_  & \new_[1172]_ ;
  assign \new_[130]_  = \new_[1167]_  & \new_[1162]_ ;
  assign \new_[131]_  = \new_[1157]_  & \new_[1152]_ ;
  assign \new_[132]_  = \new_[1147]_  & \new_[1142]_ ;
  assign \new_[133]_  = \new_[1137]_  & \new_[1132]_ ;
  assign \new_[134]_  = \new_[1127]_  & \new_[1122]_ ;
  assign \new_[135]_  = \new_[1117]_  & \new_[1112]_ ;
  assign \new_[136]_  = \new_[1107]_  & \new_[1102]_ ;
  assign \new_[137]_  = \new_[1097]_  & \new_[1092]_ ;
  assign \new_[138]_  = \new_[1087]_  & \new_[1082]_ ;
  assign \new_[139]_  = \new_[1077]_  & \new_[1072]_ ;
  assign \new_[140]_  = \new_[1067]_  & \new_[1062]_ ;
  assign \new_[141]_  = \new_[1057]_  & \new_[1052]_ ;
  assign \new_[142]_  = \new_[1047]_  & \new_[1042]_ ;
  assign \new_[143]_  = \new_[1037]_  & \new_[1032]_ ;
  assign \new_[144]_  = \new_[1027]_  & \new_[1022]_ ;
  assign \new_[145]_  = \new_[1017]_  & \new_[1012]_ ;
  assign \new_[146]_  = \new_[1007]_  & \new_[1002]_ ;
  assign \new_[147]_  = \new_[997]_  & \new_[992]_ ;
  assign \new_[148]_  = \new_[987]_  & \new_[982]_ ;
  assign \new_[149]_  = \new_[977]_  & \new_[972]_ ;
  assign \new_[150]_  = \new_[967]_  & \new_[962]_ ;
  assign \new_[151]_  = \new_[957]_  & \new_[952]_ ;
  assign \new_[152]_  = \new_[947]_  & \new_[942]_ ;
  assign \new_[153]_  = \new_[937]_  & \new_[932]_ ;
  assign \new_[154]_  = \new_[927]_  & \new_[922]_ ;
  assign \new_[155]_  = \new_[917]_  & \new_[912]_ ;
  assign \new_[156]_  = \new_[909]_  & \new_[904]_ ;
  assign \new_[157]_  = \new_[901]_  & \new_[896]_ ;
  assign \new_[158]_  = \new_[893]_  & \new_[888]_ ;
  assign \new_[159]_  = \new_[885]_  & \new_[880]_ ;
  assign \new_[160]_  = \new_[877]_  & \new_[872]_ ;
  assign \new_[161]_  = \new_[869]_  & \new_[864]_ ;
  assign \new_[162]_  = \new_[861]_  & \new_[856]_ ;
  assign \new_[163]_  = \new_[853]_  & \new_[848]_ ;
  assign \new_[164]_  = \new_[845]_  & \new_[840]_ ;
  assign \new_[165]_  = \new_[837]_  & \new_[832]_ ;
  assign \new_[166]_  = \new_[829]_  & \new_[824]_ ;
  assign \new_[167]_  = \new_[821]_  & \new_[816]_ ;
  assign \new_[168]_  = \new_[813]_  & \new_[808]_ ;
  assign \new_[169]_  = \new_[805]_  & \new_[800]_ ;
  assign \new_[170]_  = \new_[797]_  & \new_[792]_ ;
  assign \new_[171]_  = \new_[789]_  & \new_[784]_ ;
  assign \new_[172]_  = \new_[781]_  & \new_[776]_ ;
  assign \new_[173]_  = \new_[773]_  & \new_[768]_ ;
  assign \new_[174]_  = \new_[765]_  & \new_[760]_ ;
  assign \new_[175]_  = \new_[757]_  & \new_[754]_ ;
  assign \new_[176]_  = \new_[751]_  & \new_[748]_ ;
  assign \new_[177]_  = \new_[745]_  & \new_[742]_ ;
  assign \new_[178]_  = \new_[739]_  & \new_[736]_ ;
  assign \new_[179]_  = \new_[733]_  & \new_[730]_ ;
  assign \new_[180]_  = \new_[727]_  & \new_[724]_ ;
  assign \new_[181]_  = \new_[721]_  & \new_[718]_ ;
  assign \new_[182]_  = \new_[715]_  & \new_[712]_ ;
  assign \new_[183]_  = \new_[709]_  & \new_[706]_ ;
  assign \new_[184]_  = \new_[703]_  & \new_[700]_ ;
  assign \new_[185]_  = \new_[697]_  & \new_[694]_ ;
  assign \new_[186]_  = \new_[691]_  & \new_[688]_ ;
  assign \new_[187]_  = \new_[685]_  & \new_[682]_ ;
  assign \new_[188]_  = \new_[679]_  & \new_[676]_ ;
  assign \new_[189]_  = \new_[673]_  & \new_[670]_ ;
  assign \new_[190]_  = \new_[667]_  & \new_[664]_ ;
  assign \new_[191]_  = A169 & \new_[661]_ ;
  assign \new_[192]_  = A169 & \new_[657]_ ;
  assign \new_[193]_  = A168 & \new_[653]_ ;
  assign \new_[194]_  = A168 & \new_[649]_ ;
  assign \new_[195]_  = A200 & \new_[645]_ ;
  assign \new_[196]_  = A199 & \new_[641]_ ;
  assign \new_[197]_  = A202 & \new_[637]_ ;
  assign \new_[198]_  = A202 & \new_[633]_ ;
  assign \new_[199]_  = A265 & \new_[629]_ ;
  assign \new_[200]_  = ~A265 & \new_[625]_ ;
  assign \new_[201]_  = A235 & A169;
  assign \new_[202]_  = A235 & A202;
  assign \new_[203]_  = A267 & A266;
  assign \new_[204]_  = A267 & A265;
  assign \new_[209]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[210]_  = A268 | \new_[209]_ ;
  assign \new_[214]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[215]_  = \new_[202]_  | \new_[214]_ ;
  assign \new_[216]_  = \new_[215]_  | \new_[210]_ ;
  assign \new_[220]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[221]_  = \new_[199]_  | \new_[220]_ ;
  assign \new_[225]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[226]_  = \new_[196]_  | \new_[225]_ ;
  assign \new_[227]_  = \new_[226]_  | \new_[221]_ ;
  assign \new_[228]_  = \new_[227]_  | \new_[216]_ ;
  assign \new_[232]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[233]_  = \new_[193]_  | \new_[232]_ ;
  assign \new_[237]_  = \new_[188]_  | \new_[189]_ ;
  assign \new_[238]_  = \new_[190]_  | \new_[237]_ ;
  assign \new_[239]_  = \new_[238]_  | \new_[233]_ ;
  assign \new_[243]_  = \new_[185]_  | \new_[186]_ ;
  assign \new_[244]_  = \new_[187]_  | \new_[243]_ ;
  assign \new_[247]_  = \new_[183]_  | \new_[184]_ ;
  assign \new_[250]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[251]_  = \new_[250]_  | \new_[247]_ ;
  assign \new_[252]_  = \new_[251]_  | \new_[244]_ ;
  assign \new_[253]_  = \new_[252]_  | \new_[239]_ ;
  assign \new_[254]_  = \new_[253]_  | \new_[228]_ ;
  assign \new_[258]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[259]_  = \new_[180]_  | \new_[258]_ ;
  assign \new_[263]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[264]_  = \new_[177]_  | \new_[263]_ ;
  assign \new_[265]_  = \new_[264]_  | \new_[259]_ ;
  assign \new_[269]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[270]_  = \new_[174]_  | \new_[269]_ ;
  assign \new_[273]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[276]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[277]_  = \new_[276]_  | \new_[273]_ ;
  assign \new_[278]_  = \new_[277]_  | \new_[270]_ ;
  assign \new_[279]_  = \new_[278]_  | \new_[265]_ ;
  assign \new_[283]_  = \new_[165]_  | \new_[166]_ ;
  assign \new_[284]_  = \new_[167]_  | \new_[283]_ ;
  assign \new_[288]_  = \new_[162]_  | \new_[163]_ ;
  assign \new_[289]_  = \new_[164]_  | \new_[288]_ ;
  assign \new_[290]_  = \new_[289]_  | \new_[284]_ ;
  assign \new_[294]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[295]_  = \new_[161]_  | \new_[294]_ ;
  assign \new_[298]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[301]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[302]_  = \new_[301]_  | \new_[298]_ ;
  assign \new_[303]_  = \new_[302]_  | \new_[295]_ ;
  assign \new_[304]_  = \new_[303]_  | \new_[290]_ ;
  assign \new_[305]_  = \new_[304]_  | \new_[279]_ ;
  assign \new_[306]_  = \new_[305]_  | \new_[254]_ ;
  assign \new_[310]_  = \new_[152]_  | \new_[153]_ ;
  assign \new_[311]_  = \new_[154]_  | \new_[310]_ ;
  assign \new_[315]_  = \new_[149]_  | \new_[150]_ ;
  assign \new_[316]_  = \new_[151]_  | \new_[315]_ ;
  assign \new_[317]_  = \new_[316]_  | \new_[311]_ ;
  assign \new_[321]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[322]_  = \new_[148]_  | \new_[321]_ ;
  assign \new_[326]_  = \new_[143]_  | \new_[144]_ ;
  assign \new_[327]_  = \new_[145]_  | \new_[326]_ ;
  assign \new_[328]_  = \new_[327]_  | \new_[322]_ ;
  assign \new_[329]_  = \new_[328]_  | \new_[317]_ ;
  assign \new_[333]_  = \new_[140]_  | \new_[141]_ ;
  assign \new_[334]_  = \new_[142]_  | \new_[333]_ ;
  assign \new_[338]_  = \new_[137]_  | \new_[138]_ ;
  assign \new_[339]_  = \new_[139]_  | \new_[338]_ ;
  assign \new_[340]_  = \new_[339]_  | \new_[334]_ ;
  assign \new_[344]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[345]_  = \new_[136]_  | \new_[344]_ ;
  assign \new_[348]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[351]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[352]_  = \new_[351]_  | \new_[348]_ ;
  assign \new_[353]_  = \new_[352]_  | \new_[345]_ ;
  assign \new_[354]_  = \new_[353]_  | \new_[340]_ ;
  assign \new_[355]_  = \new_[354]_  | \new_[329]_ ;
  assign \new_[359]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[360]_  = \new_[129]_  | \new_[359]_ ;
  assign \new_[364]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[365]_  = \new_[126]_  | \new_[364]_ ;
  assign \new_[366]_  = \new_[365]_  | \new_[360]_ ;
  assign \new_[370]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[371]_  = \new_[123]_  | \new_[370]_ ;
  assign \new_[374]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[377]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[378]_  = \new_[377]_  | \new_[374]_ ;
  assign \new_[379]_  = \new_[378]_  | \new_[371]_ ;
  assign \new_[380]_  = \new_[379]_  | \new_[366]_ ;
  assign \new_[384]_  = \new_[114]_  | \new_[115]_ ;
  assign \new_[385]_  = \new_[116]_  | \new_[384]_ ;
  assign \new_[389]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[390]_  = \new_[113]_  | \new_[389]_ ;
  assign \new_[391]_  = \new_[390]_  | \new_[385]_ ;
  assign \new_[395]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[396]_  = \new_[110]_  | \new_[395]_ ;
  assign \new_[399]_  = \new_[106]_  | \new_[107]_ ;
  assign \new_[402]_  = \new_[104]_  | \new_[105]_ ;
  assign \new_[403]_  = \new_[402]_  | \new_[399]_ ;
  assign \new_[404]_  = \new_[403]_  | \new_[396]_ ;
  assign \new_[405]_  = \new_[404]_  | \new_[391]_ ;
  assign \new_[406]_  = \new_[405]_  | \new_[380]_ ;
  assign \new_[407]_  = \new_[406]_  | \new_[355]_ ;
  assign \new_[408]_  = \new_[407]_  | \new_[306]_ ;
  assign \new_[412]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[413]_  = \new_[103]_  | \new_[412]_ ;
  assign \new_[417]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[418]_  = \new_[100]_  | \new_[417]_ ;
  assign \new_[419]_  = \new_[418]_  | \new_[413]_ ;
  assign \new_[423]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[424]_  = \new_[97]_  | \new_[423]_ ;
  assign \new_[428]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[429]_  = \new_[94]_  | \new_[428]_ ;
  assign \new_[430]_  = \new_[429]_  | \new_[424]_ ;
  assign \new_[431]_  = \new_[430]_  | \new_[419]_ ;
  assign \new_[435]_  = \new_[89]_  | \new_[90]_ ;
  assign \new_[436]_  = \new_[91]_  | \new_[435]_ ;
  assign \new_[440]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[441]_  = \new_[88]_  | \new_[440]_ ;
  assign \new_[442]_  = \new_[441]_  | \new_[436]_ ;
  assign \new_[446]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[447]_  = \new_[85]_  | \new_[446]_ ;
  assign \new_[450]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[453]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[454]_  = \new_[453]_  | \new_[450]_ ;
  assign \new_[455]_  = \new_[454]_  | \new_[447]_ ;
  assign \new_[456]_  = \new_[455]_  | \new_[442]_ ;
  assign \new_[457]_  = \new_[456]_  | \new_[431]_ ;
  assign \new_[461]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[462]_  = \new_[78]_  | \new_[461]_ ;
  assign \new_[466]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[467]_  = \new_[75]_  | \new_[466]_ ;
  assign \new_[468]_  = \new_[467]_  | \new_[462]_ ;
  assign \new_[472]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[473]_  = \new_[72]_  | \new_[472]_ ;
  assign \new_[476]_  = \new_[68]_  | \new_[69]_ ;
  assign \new_[479]_  = \new_[66]_  | \new_[67]_ ;
  assign \new_[480]_  = \new_[479]_  | \new_[476]_ ;
  assign \new_[481]_  = \new_[480]_  | \new_[473]_ ;
  assign \new_[482]_  = \new_[481]_  | \new_[468]_ ;
  assign \new_[486]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[487]_  = \new_[65]_  | \new_[486]_ ;
  assign \new_[491]_  = \new_[60]_  | \new_[61]_ ;
  assign \new_[492]_  = \new_[62]_  | \new_[491]_ ;
  assign \new_[493]_  = \new_[492]_  | \new_[487]_ ;
  assign \new_[497]_  = \new_[57]_  | \new_[58]_ ;
  assign \new_[498]_  = \new_[59]_  | \new_[497]_ ;
  assign \new_[501]_  = \new_[55]_  | \new_[56]_ ;
  assign \new_[504]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[505]_  = \new_[504]_  | \new_[501]_ ;
  assign \new_[506]_  = \new_[505]_  | \new_[498]_ ;
  assign \new_[507]_  = \new_[506]_  | \new_[493]_ ;
  assign \new_[508]_  = \new_[507]_  | \new_[482]_ ;
  assign \new_[509]_  = \new_[508]_  | \new_[457]_ ;
  assign \new_[513]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[514]_  = \new_[52]_  | \new_[513]_ ;
  assign \new_[518]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[519]_  = \new_[49]_  | \new_[518]_ ;
  assign \new_[520]_  = \new_[519]_  | \new_[514]_ ;
  assign \new_[524]_  = \new_[44]_  | \new_[45]_ ;
  assign \new_[525]_  = \new_[46]_  | \new_[524]_ ;
  assign \new_[528]_  = \new_[42]_  | \new_[43]_ ;
  assign \new_[531]_  = \new_[40]_  | \new_[41]_ ;
  assign \new_[532]_  = \new_[531]_  | \new_[528]_ ;
  assign \new_[533]_  = \new_[532]_  | \new_[525]_ ;
  assign \new_[534]_  = \new_[533]_  | \new_[520]_ ;
  assign \new_[538]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[539]_  = \new_[39]_  | \new_[538]_ ;
  assign \new_[543]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[544]_  = \new_[36]_  | \new_[543]_ ;
  assign \new_[545]_  = \new_[544]_  | \new_[539]_ ;
  assign \new_[549]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[550]_  = \new_[33]_  | \new_[549]_ ;
  assign \new_[553]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[556]_  = \new_[27]_  | \new_[28]_ ;
  assign \new_[557]_  = \new_[556]_  | \new_[553]_ ;
  assign \new_[558]_  = \new_[557]_  | \new_[550]_ ;
  assign \new_[559]_  = \new_[558]_  | \new_[545]_ ;
  assign \new_[560]_  = \new_[559]_  | \new_[534]_ ;
  assign \new_[564]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[565]_  = \new_[26]_  | \new_[564]_ ;
  assign \new_[569]_  = \new_[21]_  | \new_[22]_ ;
  assign \new_[570]_  = \new_[23]_  | \new_[569]_ ;
  assign \new_[571]_  = \new_[570]_  | \new_[565]_ ;
  assign \new_[575]_  = \new_[18]_  | \new_[19]_ ;
  assign \new_[576]_  = \new_[20]_  | \new_[575]_ ;
  assign \new_[579]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[582]_  = \new_[14]_  | \new_[15]_ ;
  assign \new_[583]_  = \new_[582]_  | \new_[579]_ ;
  assign \new_[584]_  = \new_[583]_  | \new_[576]_ ;
  assign \new_[585]_  = \new_[584]_  | \new_[571]_ ;
  assign \new_[589]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[590]_  = \new_[13]_  | \new_[589]_ ;
  assign \new_[594]_  = \new_[8]_  | \new_[9]_ ;
  assign \new_[595]_  = \new_[10]_  | \new_[594]_ ;
  assign \new_[596]_  = \new_[595]_  | \new_[590]_ ;
  assign \new_[600]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[601]_  = \new_[7]_  | \new_[600]_ ;
  assign \new_[604]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[607]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[608]_  = \new_[607]_  | \new_[604]_ ;
  assign \new_[609]_  = \new_[608]_  | \new_[601]_ ;
  assign \new_[610]_  = \new_[609]_  | \new_[596]_ ;
  assign \new_[611]_  = \new_[610]_  | \new_[585]_ ;
  assign \new_[612]_  = \new_[611]_  | \new_[560]_ ;
  assign \new_[613]_  = \new_[612]_  | \new_[509]_ ;
  assign \new_[625]_  = A269 & A266;
  assign \new_[629]_  = A269 & ~A266;
  assign \new_[633]_  = A234 & A232;
  assign \new_[637]_  = A234 & A233;
  assign \new_[641]_  = A235 & A201;
  assign \new_[645]_  = A235 & A201;
  assign \new_[649]_  = A235 & A166;
  assign \new_[653]_  = A235 & A167;
  assign \new_[657]_  = A234 & A232;
  assign \new_[661]_  = A234 & A233;
  assign \new_[664]_  = ~A232 & A202;
  assign \new_[667]_  = A236 & A233;
  assign \new_[670]_  = A232 & A202;
  assign \new_[673]_  = A236 & ~A233;
  assign \new_[676]_  = A201 & A199;
  assign \new_[679]_  = A234 & A232;
  assign \new_[682]_  = A201 & A199;
  assign \new_[685]_  = A234 & A233;
  assign \new_[688]_  = A201 & A200;
  assign \new_[691]_  = A234 & A232;
  assign \new_[694]_  = A201 & A200;
  assign \new_[697]_  = A234 & A233;
  assign \new_[700]_  = A200 & ~A199;
  assign \new_[703]_  = A235 & A203;
  assign \new_[706]_  = ~A200 & A199;
  assign \new_[709]_  = A235 & A203;
  assign \new_[712]_  = A166 & A168;
  assign \new_[715]_  = A234 & A232;
  assign \new_[718]_  = A166 & A168;
  assign \new_[721]_  = A234 & A233;
  assign \new_[724]_  = A167 & A168;
  assign \new_[727]_  = A234 & A232;
  assign \new_[730]_  = A167 & A168;
  assign \new_[733]_  = A234 & A233;
  assign \new_[736]_  = A167 & A170;
  assign \new_[739]_  = A235 & ~A166;
  assign \new_[742]_  = ~A167 & A170;
  assign \new_[745]_  = A235 & A166;
  assign \new_[748]_  = ~A232 & A169;
  assign \new_[751]_  = A236 & A233;
  assign \new_[754]_  = A232 & A169;
  assign \new_[757]_  = A236 & ~A233;
  assign \new_[760]_  = A201 & A199;
  assign \new_[764]_  = A236 & A233;
  assign \new_[765]_  = ~A232 & \new_[764]_ ;
  assign \new_[768]_  = A201 & A199;
  assign \new_[772]_  = A236 & ~A233;
  assign \new_[773]_  = A232 & \new_[772]_ ;
  assign \new_[776]_  = A201 & A200;
  assign \new_[780]_  = A236 & A233;
  assign \new_[781]_  = ~A232 & \new_[780]_ ;
  assign \new_[784]_  = A201 & A200;
  assign \new_[788]_  = A236 & ~A233;
  assign \new_[789]_  = A232 & \new_[788]_ ;
  assign \new_[792]_  = A200 & ~A199;
  assign \new_[796]_  = A234 & A232;
  assign \new_[797]_  = A203 & \new_[796]_ ;
  assign \new_[800]_  = A200 & ~A199;
  assign \new_[804]_  = A234 & A233;
  assign \new_[805]_  = A203 & \new_[804]_ ;
  assign \new_[808]_  = ~A200 & A199;
  assign \new_[812]_  = A234 & A232;
  assign \new_[813]_  = A203 & \new_[812]_ ;
  assign \new_[816]_  = ~A200 & A199;
  assign \new_[820]_  = A234 & A233;
  assign \new_[821]_  = A203 & \new_[820]_ ;
  assign \new_[824]_  = A166 & A168;
  assign \new_[828]_  = A236 & A233;
  assign \new_[829]_  = ~A232 & \new_[828]_ ;
  assign \new_[832]_  = A166 & A168;
  assign \new_[836]_  = A236 & ~A233;
  assign \new_[837]_  = A232 & \new_[836]_ ;
  assign \new_[840]_  = A167 & A168;
  assign \new_[844]_  = A236 & A233;
  assign \new_[845]_  = ~A232 & \new_[844]_ ;
  assign \new_[848]_  = A167 & A168;
  assign \new_[852]_  = A236 & ~A233;
  assign \new_[853]_  = A232 & \new_[852]_ ;
  assign \new_[856]_  = A167 & A170;
  assign \new_[860]_  = A234 & A232;
  assign \new_[861]_  = ~A166 & \new_[860]_ ;
  assign \new_[864]_  = A167 & A170;
  assign \new_[868]_  = A234 & A233;
  assign \new_[869]_  = ~A166 & \new_[868]_ ;
  assign \new_[872]_  = ~A167 & A170;
  assign \new_[876]_  = A234 & A232;
  assign \new_[877]_  = A166 & \new_[876]_ ;
  assign \new_[880]_  = ~A167 & A170;
  assign \new_[884]_  = A234 & A233;
  assign \new_[885]_  = A166 & \new_[884]_ ;
  assign \new_[888]_  = ~A201 & A169;
  assign \new_[892]_  = A301 & ~A203;
  assign \new_[893]_  = ~A202 & \new_[892]_ ;
  assign \new_[896]_  = ~A199 & A169;
  assign \new_[900]_  = A301 & ~A202;
  assign \new_[901]_  = ~A200 & \new_[900]_ ;
  assign \new_[904]_  = ~A167 & ~A169;
  assign \new_[908]_  = A301 & A202;
  assign \new_[909]_  = ~A166 & \new_[908]_ ;
  assign \new_[912]_  = ~A169 & ~A170;
  assign \new_[916]_  = A301 & A202;
  assign \new_[917]_  = ~A168 & \new_[916]_ ;
  assign \new_[921]_  = A203 & A200;
  assign \new_[922]_  = ~A199 & \new_[921]_ ;
  assign \new_[926]_  = A236 & A233;
  assign \new_[927]_  = ~A232 & \new_[926]_ ;
  assign \new_[931]_  = A203 & A200;
  assign \new_[932]_  = ~A199 & \new_[931]_ ;
  assign \new_[936]_  = A236 & ~A233;
  assign \new_[937]_  = A232 & \new_[936]_ ;
  assign \new_[941]_  = A203 & ~A200;
  assign \new_[942]_  = A199 & \new_[941]_ ;
  assign \new_[946]_  = A236 & A233;
  assign \new_[947]_  = ~A232 & \new_[946]_ ;
  assign \new_[951]_  = A203 & ~A200;
  assign \new_[952]_  = A199 & \new_[951]_ ;
  assign \new_[956]_  = A236 & ~A233;
  assign \new_[957]_  = A232 & \new_[956]_ ;
  assign \new_[961]_  = ~A201 & A166;
  assign \new_[962]_  = A168 & \new_[961]_ ;
  assign \new_[966]_  = A301 & ~A203;
  assign \new_[967]_  = ~A202 & \new_[966]_ ;
  assign \new_[971]_  = ~A199 & A166;
  assign \new_[972]_  = A168 & \new_[971]_ ;
  assign \new_[976]_  = A301 & ~A202;
  assign \new_[977]_  = ~A200 & \new_[976]_ ;
  assign \new_[981]_  = ~A201 & A167;
  assign \new_[982]_  = A168 & \new_[981]_ ;
  assign \new_[986]_  = A301 & ~A203;
  assign \new_[987]_  = ~A202 & \new_[986]_ ;
  assign \new_[991]_  = ~A199 & A167;
  assign \new_[992]_  = A168 & \new_[991]_ ;
  assign \new_[996]_  = A301 & ~A202;
  assign \new_[997]_  = ~A200 & \new_[996]_ ;
  assign \new_[1001]_  = ~A166 & A167;
  assign \new_[1002]_  = A170 & \new_[1001]_ ;
  assign \new_[1006]_  = A236 & A233;
  assign \new_[1007]_  = ~A232 & \new_[1006]_ ;
  assign \new_[1011]_  = ~A166 & A167;
  assign \new_[1012]_  = A170 & \new_[1011]_ ;
  assign \new_[1016]_  = A236 & ~A233;
  assign \new_[1017]_  = A232 & \new_[1016]_ ;
  assign \new_[1021]_  = A166 & ~A167;
  assign \new_[1022]_  = A170 & \new_[1021]_ ;
  assign \new_[1026]_  = A236 & A233;
  assign \new_[1027]_  = ~A232 & \new_[1026]_ ;
  assign \new_[1031]_  = A166 & ~A167;
  assign \new_[1032]_  = A170 & \new_[1031]_ ;
  assign \new_[1036]_  = A236 & ~A233;
  assign \new_[1037]_  = A232 & \new_[1036]_ ;
  assign \new_[1041]_  = ~A202 & ~A201;
  assign \new_[1042]_  = A169 & \new_[1041]_ ;
  assign \new_[1046]_  = A300 & A299;
  assign \new_[1047]_  = ~A203 & \new_[1046]_ ;
  assign \new_[1051]_  = ~A202 & ~A201;
  assign \new_[1052]_  = A169 & \new_[1051]_ ;
  assign \new_[1056]_  = A300 & A298;
  assign \new_[1057]_  = ~A203 & \new_[1056]_ ;
  assign \new_[1061]_  = A200 & A199;
  assign \new_[1062]_  = A169 & \new_[1061]_ ;
  assign \new_[1066]_  = A301 & ~A202;
  assign \new_[1067]_  = ~A201 & \new_[1066]_ ;
  assign \new_[1071]_  = ~A200 & ~A199;
  assign \new_[1072]_  = A169 & \new_[1071]_ ;
  assign \new_[1076]_  = A300 & A299;
  assign \new_[1077]_  = ~A202 & \new_[1076]_ ;
  assign \new_[1081]_  = ~A200 & ~A199;
  assign \new_[1082]_  = A169 & \new_[1081]_ ;
  assign \new_[1086]_  = A300 & A298;
  assign \new_[1087]_  = ~A202 & \new_[1086]_ ;
  assign \new_[1091]_  = ~A166 & ~A167;
  assign \new_[1092]_  = ~A169 & \new_[1091]_ ;
  assign \new_[1096]_  = A300 & A299;
  assign \new_[1097]_  = A202 & \new_[1096]_ ;
  assign \new_[1101]_  = ~A166 & ~A167;
  assign \new_[1102]_  = ~A169 & \new_[1101]_ ;
  assign \new_[1106]_  = A300 & A298;
  assign \new_[1107]_  = A202 & \new_[1106]_ ;
  assign \new_[1111]_  = ~A166 & ~A167;
  assign \new_[1112]_  = ~A169 & \new_[1111]_ ;
  assign \new_[1116]_  = A301 & A201;
  assign \new_[1117]_  = A199 & \new_[1116]_ ;
  assign \new_[1121]_  = ~A166 & ~A167;
  assign \new_[1122]_  = ~A169 & \new_[1121]_ ;
  assign \new_[1126]_  = A301 & A201;
  assign \new_[1127]_  = A200 & \new_[1126]_ ;
  assign \new_[1131]_  = A167 & ~A168;
  assign \new_[1132]_  = ~A169 & \new_[1131]_ ;
  assign \new_[1136]_  = A301 & A202;
  assign \new_[1137]_  = A166 & \new_[1136]_ ;
  assign \new_[1141]_  = ~A168 & ~A169;
  assign \new_[1142]_  = ~A170 & \new_[1141]_ ;
  assign \new_[1146]_  = A300 & A299;
  assign \new_[1147]_  = A202 & \new_[1146]_ ;
  assign \new_[1151]_  = ~A168 & ~A169;
  assign \new_[1152]_  = ~A170 & \new_[1151]_ ;
  assign \new_[1156]_  = A300 & A298;
  assign \new_[1157]_  = A202 & \new_[1156]_ ;
  assign \new_[1161]_  = ~A168 & ~A169;
  assign \new_[1162]_  = ~A170 & \new_[1161]_ ;
  assign \new_[1166]_  = A301 & A201;
  assign \new_[1167]_  = A199 & \new_[1166]_ ;
  assign \new_[1171]_  = ~A168 & ~A169;
  assign \new_[1172]_  = ~A170 & \new_[1171]_ ;
  assign \new_[1176]_  = A301 & A201;
  assign \new_[1177]_  = A200 & \new_[1176]_ ;
  assign \new_[1181]_  = ~A201 & A166;
  assign \new_[1182]_  = A168 & \new_[1181]_ ;
  assign \new_[1185]_  = ~A203 & ~A202;
  assign \new_[1188]_  = A300 & A299;
  assign \new_[1189]_  = \new_[1188]_  & \new_[1185]_ ;
  assign \new_[1193]_  = ~A201 & A166;
  assign \new_[1194]_  = A168 & \new_[1193]_ ;
  assign \new_[1197]_  = ~A203 & ~A202;
  assign \new_[1200]_  = A300 & A298;
  assign \new_[1201]_  = \new_[1200]_  & \new_[1197]_ ;
  assign \new_[1205]_  = A199 & A166;
  assign \new_[1206]_  = A168 & \new_[1205]_ ;
  assign \new_[1209]_  = ~A201 & A200;
  assign \new_[1212]_  = A301 & ~A202;
  assign \new_[1213]_  = \new_[1212]_  & \new_[1209]_ ;
  assign \new_[1217]_  = ~A199 & A166;
  assign \new_[1218]_  = A168 & \new_[1217]_ ;
  assign \new_[1221]_  = ~A202 & ~A200;
  assign \new_[1224]_  = A300 & A299;
  assign \new_[1225]_  = \new_[1224]_  & \new_[1221]_ ;
  assign \new_[1229]_  = ~A199 & A166;
  assign \new_[1230]_  = A168 & \new_[1229]_ ;
  assign \new_[1233]_  = ~A202 & ~A200;
  assign \new_[1236]_  = A300 & A298;
  assign \new_[1237]_  = \new_[1236]_  & \new_[1233]_ ;
  assign \new_[1241]_  = ~A201 & A167;
  assign \new_[1242]_  = A168 & \new_[1241]_ ;
  assign \new_[1245]_  = ~A203 & ~A202;
  assign \new_[1248]_  = A300 & A299;
  assign \new_[1249]_  = \new_[1248]_  & \new_[1245]_ ;
  assign \new_[1253]_  = ~A201 & A167;
  assign \new_[1254]_  = A168 & \new_[1253]_ ;
  assign \new_[1257]_  = ~A203 & ~A202;
  assign \new_[1260]_  = A300 & A298;
  assign \new_[1261]_  = \new_[1260]_  & \new_[1257]_ ;
  assign \new_[1265]_  = A199 & A167;
  assign \new_[1266]_  = A168 & \new_[1265]_ ;
  assign \new_[1269]_  = ~A201 & A200;
  assign \new_[1272]_  = A301 & ~A202;
  assign \new_[1273]_  = \new_[1272]_  & \new_[1269]_ ;
  assign \new_[1277]_  = ~A199 & A167;
  assign \new_[1278]_  = A168 & \new_[1277]_ ;
  assign \new_[1281]_  = ~A202 & ~A200;
  assign \new_[1284]_  = A300 & A299;
  assign \new_[1285]_  = \new_[1284]_  & \new_[1281]_ ;
  assign \new_[1289]_  = ~A199 & A167;
  assign \new_[1290]_  = A168 & \new_[1289]_ ;
  assign \new_[1293]_  = ~A202 & ~A200;
  assign \new_[1296]_  = A300 & A298;
  assign \new_[1297]_  = \new_[1296]_  & \new_[1293]_ ;
  assign \new_[1301]_  = ~A166 & A167;
  assign \new_[1302]_  = A170 & \new_[1301]_ ;
  assign \new_[1305]_  = ~A202 & ~A201;
  assign \new_[1308]_  = A301 & ~A203;
  assign \new_[1309]_  = \new_[1308]_  & \new_[1305]_ ;
  assign \new_[1313]_  = ~A166 & A167;
  assign \new_[1314]_  = A170 & \new_[1313]_ ;
  assign \new_[1317]_  = ~A200 & ~A199;
  assign \new_[1320]_  = A301 & ~A202;
  assign \new_[1321]_  = \new_[1320]_  & \new_[1317]_ ;
  assign \new_[1325]_  = A166 & ~A167;
  assign \new_[1326]_  = A170 & \new_[1325]_ ;
  assign \new_[1329]_  = ~A202 & ~A201;
  assign \new_[1332]_  = A301 & ~A203;
  assign \new_[1333]_  = \new_[1332]_  & \new_[1329]_ ;
  assign \new_[1337]_  = A166 & ~A167;
  assign \new_[1338]_  = A170 & \new_[1337]_ ;
  assign \new_[1341]_  = ~A200 & ~A199;
  assign \new_[1344]_  = A301 & ~A202;
  assign \new_[1345]_  = \new_[1344]_  & \new_[1341]_ ;
  assign \new_[1349]_  = ~A202 & ~A201;
  assign \new_[1350]_  = A169 & \new_[1349]_ ;
  assign \new_[1353]_  = A298 & ~A203;
  assign \new_[1356]_  = A302 & ~A299;
  assign \new_[1357]_  = \new_[1356]_  & \new_[1353]_ ;
  assign \new_[1361]_  = ~A202 & ~A201;
  assign \new_[1362]_  = A169 & \new_[1361]_ ;
  assign \new_[1365]_  = ~A298 & ~A203;
  assign \new_[1368]_  = A302 & A299;
  assign \new_[1369]_  = \new_[1368]_  & \new_[1365]_ ;
  assign \new_[1373]_  = A200 & A199;
  assign \new_[1374]_  = A169 & \new_[1373]_ ;
  assign \new_[1377]_  = ~A202 & ~A201;
  assign \new_[1380]_  = A300 & A299;
  assign \new_[1381]_  = \new_[1380]_  & \new_[1377]_ ;
  assign \new_[1385]_  = A200 & A199;
  assign \new_[1386]_  = A169 & \new_[1385]_ ;
  assign \new_[1389]_  = ~A202 & ~A201;
  assign \new_[1392]_  = A300 & A298;
  assign \new_[1393]_  = \new_[1392]_  & \new_[1389]_ ;
  assign \new_[1397]_  = ~A200 & ~A199;
  assign \new_[1398]_  = A169 & \new_[1397]_ ;
  assign \new_[1401]_  = A298 & ~A202;
  assign \new_[1404]_  = A302 & ~A299;
  assign \new_[1405]_  = \new_[1404]_  & \new_[1401]_ ;
  assign \new_[1409]_  = ~A200 & ~A199;
  assign \new_[1410]_  = A169 & \new_[1409]_ ;
  assign \new_[1413]_  = ~A298 & ~A202;
  assign \new_[1416]_  = A302 & A299;
  assign \new_[1417]_  = \new_[1416]_  & \new_[1413]_ ;
  assign \new_[1421]_  = ~A166 & ~A167;
  assign \new_[1422]_  = ~A169 & \new_[1421]_ ;
  assign \new_[1425]_  = A298 & A202;
  assign \new_[1428]_  = A302 & ~A299;
  assign \new_[1429]_  = \new_[1428]_  & \new_[1425]_ ;
  assign \new_[1433]_  = ~A166 & ~A167;
  assign \new_[1434]_  = ~A169 & \new_[1433]_ ;
  assign \new_[1437]_  = ~A298 & A202;
  assign \new_[1440]_  = A302 & A299;
  assign \new_[1441]_  = \new_[1440]_  & \new_[1437]_ ;
  assign \new_[1445]_  = ~A166 & ~A167;
  assign \new_[1446]_  = ~A169 & \new_[1445]_ ;
  assign \new_[1449]_  = A201 & A199;
  assign \new_[1452]_  = A300 & A299;
  assign \new_[1453]_  = \new_[1452]_  & \new_[1449]_ ;
  assign \new_[1457]_  = ~A166 & ~A167;
  assign \new_[1458]_  = ~A169 & \new_[1457]_ ;
  assign \new_[1461]_  = A201 & A199;
  assign \new_[1464]_  = A300 & A298;
  assign \new_[1465]_  = \new_[1464]_  & \new_[1461]_ ;
  assign \new_[1469]_  = ~A166 & ~A167;
  assign \new_[1470]_  = ~A169 & \new_[1469]_ ;
  assign \new_[1473]_  = A201 & A200;
  assign \new_[1476]_  = A300 & A299;
  assign \new_[1477]_  = \new_[1476]_  & \new_[1473]_ ;
  assign \new_[1481]_  = ~A166 & ~A167;
  assign \new_[1482]_  = ~A169 & \new_[1481]_ ;
  assign \new_[1485]_  = A201 & A200;
  assign \new_[1488]_  = A300 & A298;
  assign \new_[1489]_  = \new_[1488]_  & \new_[1485]_ ;
  assign \new_[1493]_  = ~A166 & ~A167;
  assign \new_[1494]_  = ~A169 & \new_[1493]_ ;
  assign \new_[1497]_  = A200 & ~A199;
  assign \new_[1500]_  = A301 & A203;
  assign \new_[1501]_  = \new_[1500]_  & \new_[1497]_ ;
  assign \new_[1505]_  = ~A166 & ~A167;
  assign \new_[1506]_  = ~A169 & \new_[1505]_ ;
  assign \new_[1509]_  = ~A200 & A199;
  assign \new_[1512]_  = A301 & A203;
  assign \new_[1513]_  = \new_[1512]_  & \new_[1509]_ ;
  assign \new_[1517]_  = A167 & ~A168;
  assign \new_[1518]_  = ~A169 & \new_[1517]_ ;
  assign \new_[1521]_  = A202 & A166;
  assign \new_[1524]_  = A300 & A299;
  assign \new_[1525]_  = \new_[1524]_  & \new_[1521]_ ;
  assign \new_[1529]_  = A167 & ~A168;
  assign \new_[1530]_  = ~A169 & \new_[1529]_ ;
  assign \new_[1533]_  = A202 & A166;
  assign \new_[1536]_  = A300 & A298;
  assign \new_[1537]_  = \new_[1536]_  & \new_[1533]_ ;
  assign \new_[1541]_  = A167 & ~A168;
  assign \new_[1542]_  = ~A169 & \new_[1541]_ ;
  assign \new_[1545]_  = A199 & A166;
  assign \new_[1548]_  = A301 & A201;
  assign \new_[1549]_  = \new_[1548]_  & \new_[1545]_ ;
  assign \new_[1553]_  = A167 & ~A168;
  assign \new_[1554]_  = ~A169 & \new_[1553]_ ;
  assign \new_[1557]_  = A200 & A166;
  assign \new_[1560]_  = A301 & A201;
  assign \new_[1561]_  = \new_[1560]_  & \new_[1557]_ ;
  assign \new_[1565]_  = ~A168 & ~A169;
  assign \new_[1566]_  = ~A170 & \new_[1565]_ ;
  assign \new_[1569]_  = A298 & A202;
  assign \new_[1572]_  = A302 & ~A299;
  assign \new_[1573]_  = \new_[1572]_  & \new_[1569]_ ;
  assign \new_[1577]_  = ~A168 & ~A169;
  assign \new_[1578]_  = ~A170 & \new_[1577]_ ;
  assign \new_[1581]_  = ~A298 & A202;
  assign \new_[1584]_  = A302 & A299;
  assign \new_[1585]_  = \new_[1584]_  & \new_[1581]_ ;
  assign \new_[1589]_  = ~A168 & ~A169;
  assign \new_[1590]_  = ~A170 & \new_[1589]_ ;
  assign \new_[1593]_  = A201 & A199;
  assign \new_[1596]_  = A300 & A299;
  assign \new_[1597]_  = \new_[1596]_  & \new_[1593]_ ;
  assign \new_[1601]_  = ~A168 & ~A169;
  assign \new_[1602]_  = ~A170 & \new_[1601]_ ;
  assign \new_[1605]_  = A201 & A199;
  assign \new_[1608]_  = A300 & A298;
  assign \new_[1609]_  = \new_[1608]_  & \new_[1605]_ ;
  assign \new_[1613]_  = ~A168 & ~A169;
  assign \new_[1614]_  = ~A170 & \new_[1613]_ ;
  assign \new_[1617]_  = A201 & A200;
  assign \new_[1620]_  = A300 & A299;
  assign \new_[1621]_  = \new_[1620]_  & \new_[1617]_ ;
  assign \new_[1625]_  = ~A168 & ~A169;
  assign \new_[1626]_  = ~A170 & \new_[1625]_ ;
  assign \new_[1629]_  = A201 & A200;
  assign \new_[1632]_  = A300 & A298;
  assign \new_[1633]_  = \new_[1632]_  & \new_[1629]_ ;
  assign \new_[1637]_  = ~A168 & ~A169;
  assign \new_[1638]_  = ~A170 & \new_[1637]_ ;
  assign \new_[1641]_  = A200 & ~A199;
  assign \new_[1644]_  = A301 & A203;
  assign \new_[1645]_  = \new_[1644]_  & \new_[1641]_ ;
  assign \new_[1649]_  = ~A168 & ~A169;
  assign \new_[1650]_  = ~A170 & \new_[1649]_ ;
  assign \new_[1653]_  = ~A200 & A199;
  assign \new_[1656]_  = A301 & A203;
  assign \new_[1657]_  = \new_[1656]_  & \new_[1653]_ ;
  assign \new_[1660]_  = A166 & A168;
  assign \new_[1663]_  = ~A202 & ~A201;
  assign \new_[1664]_  = \new_[1663]_  & \new_[1660]_ ;
  assign \new_[1667]_  = A298 & ~A203;
  assign \new_[1670]_  = A302 & ~A299;
  assign \new_[1671]_  = \new_[1670]_  & \new_[1667]_ ;
  assign \new_[1674]_  = A166 & A168;
  assign \new_[1677]_  = ~A202 & ~A201;
  assign \new_[1678]_  = \new_[1677]_  & \new_[1674]_ ;
  assign \new_[1681]_  = ~A298 & ~A203;
  assign \new_[1684]_  = A302 & A299;
  assign \new_[1685]_  = \new_[1684]_  & \new_[1681]_ ;
  assign \new_[1688]_  = A166 & A168;
  assign \new_[1691]_  = A200 & A199;
  assign \new_[1692]_  = \new_[1691]_  & \new_[1688]_ ;
  assign \new_[1695]_  = ~A202 & ~A201;
  assign \new_[1698]_  = A300 & A299;
  assign \new_[1699]_  = \new_[1698]_  & \new_[1695]_ ;
  assign \new_[1702]_  = A166 & A168;
  assign \new_[1705]_  = A200 & A199;
  assign \new_[1706]_  = \new_[1705]_  & \new_[1702]_ ;
  assign \new_[1709]_  = ~A202 & ~A201;
  assign \new_[1712]_  = A300 & A298;
  assign \new_[1713]_  = \new_[1712]_  & \new_[1709]_ ;
  assign \new_[1716]_  = A166 & A168;
  assign \new_[1719]_  = ~A200 & ~A199;
  assign \new_[1720]_  = \new_[1719]_  & \new_[1716]_ ;
  assign \new_[1723]_  = A298 & ~A202;
  assign \new_[1726]_  = A302 & ~A299;
  assign \new_[1727]_  = \new_[1726]_  & \new_[1723]_ ;
  assign \new_[1730]_  = A166 & A168;
  assign \new_[1733]_  = ~A200 & ~A199;
  assign \new_[1734]_  = \new_[1733]_  & \new_[1730]_ ;
  assign \new_[1737]_  = ~A298 & ~A202;
  assign \new_[1740]_  = A302 & A299;
  assign \new_[1741]_  = \new_[1740]_  & \new_[1737]_ ;
  assign \new_[1744]_  = A167 & A168;
  assign \new_[1747]_  = ~A202 & ~A201;
  assign \new_[1748]_  = \new_[1747]_  & \new_[1744]_ ;
  assign \new_[1751]_  = A298 & ~A203;
  assign \new_[1754]_  = A302 & ~A299;
  assign \new_[1755]_  = \new_[1754]_  & \new_[1751]_ ;
  assign \new_[1758]_  = A167 & A168;
  assign \new_[1761]_  = ~A202 & ~A201;
  assign \new_[1762]_  = \new_[1761]_  & \new_[1758]_ ;
  assign \new_[1765]_  = ~A298 & ~A203;
  assign \new_[1768]_  = A302 & A299;
  assign \new_[1769]_  = \new_[1768]_  & \new_[1765]_ ;
  assign \new_[1772]_  = A167 & A168;
  assign \new_[1775]_  = A200 & A199;
  assign \new_[1776]_  = \new_[1775]_  & \new_[1772]_ ;
  assign \new_[1779]_  = ~A202 & ~A201;
  assign \new_[1782]_  = A300 & A299;
  assign \new_[1783]_  = \new_[1782]_  & \new_[1779]_ ;
  assign \new_[1786]_  = A167 & A168;
  assign \new_[1789]_  = A200 & A199;
  assign \new_[1790]_  = \new_[1789]_  & \new_[1786]_ ;
  assign \new_[1793]_  = ~A202 & ~A201;
  assign \new_[1796]_  = A300 & A298;
  assign \new_[1797]_  = \new_[1796]_  & \new_[1793]_ ;
  assign \new_[1800]_  = A167 & A168;
  assign \new_[1803]_  = ~A200 & ~A199;
  assign \new_[1804]_  = \new_[1803]_  & \new_[1800]_ ;
  assign \new_[1807]_  = A298 & ~A202;
  assign \new_[1810]_  = A302 & ~A299;
  assign \new_[1811]_  = \new_[1810]_  & \new_[1807]_ ;
  assign \new_[1814]_  = A167 & A168;
  assign \new_[1817]_  = ~A200 & ~A199;
  assign \new_[1818]_  = \new_[1817]_  & \new_[1814]_ ;
  assign \new_[1821]_  = ~A298 & ~A202;
  assign \new_[1824]_  = A302 & A299;
  assign \new_[1825]_  = \new_[1824]_  & \new_[1821]_ ;
  assign \new_[1828]_  = A167 & A170;
  assign \new_[1831]_  = ~A201 & ~A166;
  assign \new_[1832]_  = \new_[1831]_  & \new_[1828]_ ;
  assign \new_[1835]_  = ~A203 & ~A202;
  assign \new_[1838]_  = A300 & A299;
  assign \new_[1839]_  = \new_[1838]_  & \new_[1835]_ ;
  assign \new_[1842]_  = A167 & A170;
  assign \new_[1845]_  = ~A201 & ~A166;
  assign \new_[1846]_  = \new_[1845]_  & \new_[1842]_ ;
  assign \new_[1849]_  = ~A203 & ~A202;
  assign \new_[1852]_  = A300 & A298;
  assign \new_[1853]_  = \new_[1852]_  & \new_[1849]_ ;
  assign \new_[1856]_  = A167 & A170;
  assign \new_[1859]_  = A199 & ~A166;
  assign \new_[1860]_  = \new_[1859]_  & \new_[1856]_ ;
  assign \new_[1863]_  = ~A201 & A200;
  assign \new_[1866]_  = A301 & ~A202;
  assign \new_[1867]_  = \new_[1866]_  & \new_[1863]_ ;
  assign \new_[1870]_  = A167 & A170;
  assign \new_[1873]_  = ~A199 & ~A166;
  assign \new_[1874]_  = \new_[1873]_  & \new_[1870]_ ;
  assign \new_[1877]_  = ~A202 & ~A200;
  assign \new_[1880]_  = A300 & A299;
  assign \new_[1881]_  = \new_[1880]_  & \new_[1877]_ ;
  assign \new_[1884]_  = A167 & A170;
  assign \new_[1887]_  = ~A199 & ~A166;
  assign \new_[1888]_  = \new_[1887]_  & \new_[1884]_ ;
  assign \new_[1891]_  = ~A202 & ~A200;
  assign \new_[1894]_  = A300 & A298;
  assign \new_[1895]_  = \new_[1894]_  & \new_[1891]_ ;
  assign \new_[1898]_  = ~A167 & A170;
  assign \new_[1901]_  = ~A201 & A166;
  assign \new_[1902]_  = \new_[1901]_  & \new_[1898]_ ;
  assign \new_[1905]_  = ~A203 & ~A202;
  assign \new_[1908]_  = A300 & A299;
  assign \new_[1909]_  = \new_[1908]_  & \new_[1905]_ ;
  assign \new_[1912]_  = ~A167 & A170;
  assign \new_[1915]_  = ~A201 & A166;
  assign \new_[1916]_  = \new_[1915]_  & \new_[1912]_ ;
  assign \new_[1919]_  = ~A203 & ~A202;
  assign \new_[1922]_  = A300 & A298;
  assign \new_[1923]_  = \new_[1922]_  & \new_[1919]_ ;
  assign \new_[1926]_  = ~A167 & A170;
  assign \new_[1929]_  = A199 & A166;
  assign \new_[1930]_  = \new_[1929]_  & \new_[1926]_ ;
  assign \new_[1933]_  = ~A201 & A200;
  assign \new_[1936]_  = A301 & ~A202;
  assign \new_[1937]_  = \new_[1936]_  & \new_[1933]_ ;
  assign \new_[1940]_  = ~A167 & A170;
  assign \new_[1943]_  = ~A199 & A166;
  assign \new_[1944]_  = \new_[1943]_  & \new_[1940]_ ;
  assign \new_[1947]_  = ~A202 & ~A200;
  assign \new_[1950]_  = A300 & A299;
  assign \new_[1951]_  = \new_[1950]_  & \new_[1947]_ ;
  assign \new_[1954]_  = ~A167 & A170;
  assign \new_[1957]_  = ~A199 & A166;
  assign \new_[1958]_  = \new_[1957]_  & \new_[1954]_ ;
  assign \new_[1961]_  = ~A202 & ~A200;
  assign \new_[1964]_  = A300 & A298;
  assign \new_[1965]_  = \new_[1964]_  & \new_[1961]_ ;
  assign \new_[1968]_  = A199 & A169;
  assign \new_[1971]_  = ~A201 & A200;
  assign \new_[1972]_  = \new_[1971]_  & \new_[1968]_ ;
  assign \new_[1975]_  = A298 & ~A202;
  assign \new_[1978]_  = A302 & ~A299;
  assign \new_[1979]_  = \new_[1978]_  & \new_[1975]_ ;
  assign \new_[1982]_  = A199 & A169;
  assign \new_[1985]_  = ~A201 & A200;
  assign \new_[1986]_  = \new_[1985]_  & \new_[1982]_ ;
  assign \new_[1989]_  = ~A298 & ~A202;
  assign \new_[1992]_  = A302 & A299;
  assign \new_[1993]_  = \new_[1992]_  & \new_[1989]_ ;
  assign \new_[1996]_  = ~A167 & ~A169;
  assign \new_[1999]_  = A199 & ~A166;
  assign \new_[2000]_  = \new_[1999]_  & \new_[1996]_ ;
  assign \new_[2003]_  = A298 & A201;
  assign \new_[2006]_  = A302 & ~A299;
  assign \new_[2007]_  = \new_[2006]_  & \new_[2003]_ ;
  assign \new_[2010]_  = ~A167 & ~A169;
  assign \new_[2013]_  = A199 & ~A166;
  assign \new_[2014]_  = \new_[2013]_  & \new_[2010]_ ;
  assign \new_[2017]_  = ~A298 & A201;
  assign \new_[2020]_  = A302 & A299;
  assign \new_[2021]_  = \new_[2020]_  & \new_[2017]_ ;
  assign \new_[2024]_  = ~A167 & ~A169;
  assign \new_[2027]_  = A200 & ~A166;
  assign \new_[2028]_  = \new_[2027]_  & \new_[2024]_ ;
  assign \new_[2031]_  = A298 & A201;
  assign \new_[2034]_  = A302 & ~A299;
  assign \new_[2035]_  = \new_[2034]_  & \new_[2031]_ ;
  assign \new_[2038]_  = ~A167 & ~A169;
  assign \new_[2041]_  = A200 & ~A166;
  assign \new_[2042]_  = \new_[2041]_  & \new_[2038]_ ;
  assign \new_[2045]_  = ~A298 & A201;
  assign \new_[2048]_  = A302 & A299;
  assign \new_[2049]_  = \new_[2048]_  & \new_[2045]_ ;
  assign \new_[2052]_  = ~A167 & ~A169;
  assign \new_[2055]_  = ~A199 & ~A166;
  assign \new_[2056]_  = \new_[2055]_  & \new_[2052]_ ;
  assign \new_[2059]_  = A203 & A200;
  assign \new_[2062]_  = A300 & A299;
  assign \new_[2063]_  = \new_[2062]_  & \new_[2059]_ ;
  assign \new_[2066]_  = ~A167 & ~A169;
  assign \new_[2069]_  = ~A199 & ~A166;
  assign \new_[2070]_  = \new_[2069]_  & \new_[2066]_ ;
  assign \new_[2073]_  = A203 & A200;
  assign \new_[2076]_  = A300 & A298;
  assign \new_[2077]_  = \new_[2076]_  & \new_[2073]_ ;
  assign \new_[2080]_  = ~A167 & ~A169;
  assign \new_[2083]_  = A199 & ~A166;
  assign \new_[2084]_  = \new_[2083]_  & \new_[2080]_ ;
  assign \new_[2087]_  = A203 & ~A200;
  assign \new_[2090]_  = A300 & A299;
  assign \new_[2091]_  = \new_[2090]_  & \new_[2087]_ ;
  assign \new_[2094]_  = ~A167 & ~A169;
  assign \new_[2097]_  = A199 & ~A166;
  assign \new_[2098]_  = \new_[2097]_  & \new_[2094]_ ;
  assign \new_[2101]_  = A203 & ~A200;
  assign \new_[2104]_  = A300 & A298;
  assign \new_[2105]_  = \new_[2104]_  & \new_[2101]_ ;
  assign \new_[2108]_  = ~A168 & ~A169;
  assign \new_[2111]_  = A166 & A167;
  assign \new_[2112]_  = \new_[2111]_  & \new_[2108]_ ;
  assign \new_[2115]_  = A298 & A202;
  assign \new_[2118]_  = A302 & ~A299;
  assign \new_[2119]_  = \new_[2118]_  & \new_[2115]_ ;
  assign \new_[2122]_  = ~A168 & ~A169;
  assign \new_[2125]_  = A166 & A167;
  assign \new_[2126]_  = \new_[2125]_  & \new_[2122]_ ;
  assign \new_[2129]_  = ~A298 & A202;
  assign \new_[2132]_  = A302 & A299;
  assign \new_[2133]_  = \new_[2132]_  & \new_[2129]_ ;
  assign \new_[2136]_  = ~A168 & ~A169;
  assign \new_[2139]_  = A166 & A167;
  assign \new_[2140]_  = \new_[2139]_  & \new_[2136]_ ;
  assign \new_[2143]_  = A201 & A199;
  assign \new_[2146]_  = A300 & A299;
  assign \new_[2147]_  = \new_[2146]_  & \new_[2143]_ ;
  assign \new_[2150]_  = ~A168 & ~A169;
  assign \new_[2153]_  = A166 & A167;
  assign \new_[2154]_  = \new_[2153]_  & \new_[2150]_ ;
  assign \new_[2157]_  = A201 & A199;
  assign \new_[2160]_  = A300 & A298;
  assign \new_[2161]_  = \new_[2160]_  & \new_[2157]_ ;
  assign \new_[2164]_  = ~A168 & ~A169;
  assign \new_[2167]_  = A166 & A167;
  assign \new_[2168]_  = \new_[2167]_  & \new_[2164]_ ;
  assign \new_[2171]_  = A201 & A200;
  assign \new_[2174]_  = A300 & A299;
  assign \new_[2175]_  = \new_[2174]_  & \new_[2171]_ ;
  assign \new_[2178]_  = ~A168 & ~A169;
  assign \new_[2181]_  = A166 & A167;
  assign \new_[2182]_  = \new_[2181]_  & \new_[2178]_ ;
  assign \new_[2185]_  = A201 & A200;
  assign \new_[2188]_  = A300 & A298;
  assign \new_[2189]_  = \new_[2188]_  & \new_[2185]_ ;
  assign \new_[2192]_  = ~A168 & ~A169;
  assign \new_[2195]_  = A166 & A167;
  assign \new_[2196]_  = \new_[2195]_  & \new_[2192]_ ;
  assign \new_[2199]_  = A200 & ~A199;
  assign \new_[2202]_  = A301 & A203;
  assign \new_[2203]_  = \new_[2202]_  & \new_[2199]_ ;
  assign \new_[2206]_  = ~A168 & ~A169;
  assign \new_[2209]_  = A166 & A167;
  assign \new_[2210]_  = \new_[2209]_  & \new_[2206]_ ;
  assign \new_[2213]_  = ~A200 & A199;
  assign \new_[2216]_  = A301 & A203;
  assign \new_[2217]_  = \new_[2216]_  & \new_[2213]_ ;
  assign \new_[2220]_  = ~A169 & ~A170;
  assign \new_[2223]_  = A199 & ~A168;
  assign \new_[2224]_  = \new_[2223]_  & \new_[2220]_ ;
  assign \new_[2227]_  = A298 & A201;
  assign \new_[2230]_  = A302 & ~A299;
  assign \new_[2231]_  = \new_[2230]_  & \new_[2227]_ ;
  assign \new_[2234]_  = ~A169 & ~A170;
  assign \new_[2237]_  = A199 & ~A168;
  assign \new_[2238]_  = \new_[2237]_  & \new_[2234]_ ;
  assign \new_[2241]_  = ~A298 & A201;
  assign \new_[2244]_  = A302 & A299;
  assign \new_[2245]_  = \new_[2244]_  & \new_[2241]_ ;
  assign \new_[2248]_  = ~A169 & ~A170;
  assign \new_[2251]_  = A200 & ~A168;
  assign \new_[2252]_  = \new_[2251]_  & \new_[2248]_ ;
  assign \new_[2255]_  = A298 & A201;
  assign \new_[2258]_  = A302 & ~A299;
  assign \new_[2259]_  = \new_[2258]_  & \new_[2255]_ ;
  assign \new_[2262]_  = ~A169 & ~A170;
  assign \new_[2265]_  = A200 & ~A168;
  assign \new_[2266]_  = \new_[2265]_  & \new_[2262]_ ;
  assign \new_[2269]_  = ~A298 & A201;
  assign \new_[2272]_  = A302 & A299;
  assign \new_[2273]_  = \new_[2272]_  & \new_[2269]_ ;
  assign \new_[2276]_  = ~A169 & ~A170;
  assign \new_[2279]_  = ~A199 & ~A168;
  assign \new_[2280]_  = \new_[2279]_  & \new_[2276]_ ;
  assign \new_[2283]_  = A203 & A200;
  assign \new_[2286]_  = A300 & A299;
  assign \new_[2287]_  = \new_[2286]_  & \new_[2283]_ ;
  assign \new_[2290]_  = ~A169 & ~A170;
  assign \new_[2293]_  = ~A199 & ~A168;
  assign \new_[2294]_  = \new_[2293]_  & \new_[2290]_ ;
  assign \new_[2297]_  = A203 & A200;
  assign \new_[2300]_  = A300 & A298;
  assign \new_[2301]_  = \new_[2300]_  & \new_[2297]_ ;
  assign \new_[2304]_  = ~A169 & ~A170;
  assign \new_[2307]_  = A199 & ~A168;
  assign \new_[2308]_  = \new_[2307]_  & \new_[2304]_ ;
  assign \new_[2311]_  = A203 & ~A200;
  assign \new_[2314]_  = A300 & A299;
  assign \new_[2315]_  = \new_[2314]_  & \new_[2311]_ ;
  assign \new_[2318]_  = ~A169 & ~A170;
  assign \new_[2321]_  = A199 & ~A168;
  assign \new_[2322]_  = \new_[2321]_  & \new_[2318]_ ;
  assign \new_[2325]_  = A203 & ~A200;
  assign \new_[2328]_  = A300 & A298;
  assign \new_[2329]_  = \new_[2328]_  & \new_[2325]_ ;
  assign \new_[2332]_  = A166 & A168;
  assign \new_[2335]_  = A200 & A199;
  assign \new_[2336]_  = \new_[2335]_  & \new_[2332]_ ;
  assign \new_[2339]_  = ~A202 & ~A201;
  assign \new_[2343]_  = A302 & ~A299;
  assign \new_[2344]_  = A298 & \new_[2343]_ ;
  assign \new_[2345]_  = \new_[2344]_  & \new_[2339]_ ;
  assign \new_[2348]_  = A166 & A168;
  assign \new_[2351]_  = A200 & A199;
  assign \new_[2352]_  = \new_[2351]_  & \new_[2348]_ ;
  assign \new_[2355]_  = ~A202 & ~A201;
  assign \new_[2359]_  = A302 & A299;
  assign \new_[2360]_  = ~A298 & \new_[2359]_ ;
  assign \new_[2361]_  = \new_[2360]_  & \new_[2355]_ ;
  assign \new_[2364]_  = A167 & A168;
  assign \new_[2367]_  = A200 & A199;
  assign \new_[2368]_  = \new_[2367]_  & \new_[2364]_ ;
  assign \new_[2371]_  = ~A202 & ~A201;
  assign \new_[2375]_  = A302 & ~A299;
  assign \new_[2376]_  = A298 & \new_[2375]_ ;
  assign \new_[2377]_  = \new_[2376]_  & \new_[2371]_ ;
  assign \new_[2380]_  = A167 & A168;
  assign \new_[2383]_  = A200 & A199;
  assign \new_[2384]_  = \new_[2383]_  & \new_[2380]_ ;
  assign \new_[2387]_  = ~A202 & ~A201;
  assign \new_[2391]_  = A302 & A299;
  assign \new_[2392]_  = ~A298 & \new_[2391]_ ;
  assign \new_[2393]_  = \new_[2392]_  & \new_[2387]_ ;
  assign \new_[2396]_  = A167 & A170;
  assign \new_[2399]_  = ~A201 & ~A166;
  assign \new_[2400]_  = \new_[2399]_  & \new_[2396]_ ;
  assign \new_[2403]_  = ~A203 & ~A202;
  assign \new_[2407]_  = A302 & ~A299;
  assign \new_[2408]_  = A298 & \new_[2407]_ ;
  assign \new_[2409]_  = \new_[2408]_  & \new_[2403]_ ;
  assign \new_[2412]_  = A167 & A170;
  assign \new_[2415]_  = ~A201 & ~A166;
  assign \new_[2416]_  = \new_[2415]_  & \new_[2412]_ ;
  assign \new_[2419]_  = ~A203 & ~A202;
  assign \new_[2423]_  = A302 & A299;
  assign \new_[2424]_  = ~A298 & \new_[2423]_ ;
  assign \new_[2425]_  = \new_[2424]_  & \new_[2419]_ ;
  assign \new_[2428]_  = A167 & A170;
  assign \new_[2431]_  = A199 & ~A166;
  assign \new_[2432]_  = \new_[2431]_  & \new_[2428]_ ;
  assign \new_[2435]_  = ~A201 & A200;
  assign \new_[2439]_  = A300 & A299;
  assign \new_[2440]_  = ~A202 & \new_[2439]_ ;
  assign \new_[2441]_  = \new_[2440]_  & \new_[2435]_ ;
  assign \new_[2444]_  = A167 & A170;
  assign \new_[2447]_  = A199 & ~A166;
  assign \new_[2448]_  = \new_[2447]_  & \new_[2444]_ ;
  assign \new_[2451]_  = ~A201 & A200;
  assign \new_[2455]_  = A300 & A298;
  assign \new_[2456]_  = ~A202 & \new_[2455]_ ;
  assign \new_[2457]_  = \new_[2456]_  & \new_[2451]_ ;
  assign \new_[2460]_  = A167 & A170;
  assign \new_[2463]_  = ~A199 & ~A166;
  assign \new_[2464]_  = \new_[2463]_  & \new_[2460]_ ;
  assign \new_[2467]_  = ~A202 & ~A200;
  assign \new_[2471]_  = A302 & ~A299;
  assign \new_[2472]_  = A298 & \new_[2471]_ ;
  assign \new_[2473]_  = \new_[2472]_  & \new_[2467]_ ;
  assign \new_[2476]_  = A167 & A170;
  assign \new_[2479]_  = ~A199 & ~A166;
  assign \new_[2480]_  = \new_[2479]_  & \new_[2476]_ ;
  assign \new_[2483]_  = ~A202 & ~A200;
  assign \new_[2487]_  = A302 & A299;
  assign \new_[2488]_  = ~A298 & \new_[2487]_ ;
  assign \new_[2489]_  = \new_[2488]_  & \new_[2483]_ ;
  assign \new_[2492]_  = ~A167 & A170;
  assign \new_[2495]_  = ~A201 & A166;
  assign \new_[2496]_  = \new_[2495]_  & \new_[2492]_ ;
  assign \new_[2499]_  = ~A203 & ~A202;
  assign \new_[2503]_  = A302 & ~A299;
  assign \new_[2504]_  = A298 & \new_[2503]_ ;
  assign \new_[2505]_  = \new_[2504]_  & \new_[2499]_ ;
  assign \new_[2508]_  = ~A167 & A170;
  assign \new_[2511]_  = ~A201 & A166;
  assign \new_[2512]_  = \new_[2511]_  & \new_[2508]_ ;
  assign \new_[2515]_  = ~A203 & ~A202;
  assign \new_[2519]_  = A302 & A299;
  assign \new_[2520]_  = ~A298 & \new_[2519]_ ;
  assign \new_[2521]_  = \new_[2520]_  & \new_[2515]_ ;
  assign \new_[2524]_  = ~A167 & A170;
  assign \new_[2527]_  = A199 & A166;
  assign \new_[2528]_  = \new_[2527]_  & \new_[2524]_ ;
  assign \new_[2531]_  = ~A201 & A200;
  assign \new_[2535]_  = A300 & A299;
  assign \new_[2536]_  = ~A202 & \new_[2535]_ ;
  assign \new_[2537]_  = \new_[2536]_  & \new_[2531]_ ;
  assign \new_[2540]_  = ~A167 & A170;
  assign \new_[2543]_  = A199 & A166;
  assign \new_[2544]_  = \new_[2543]_  & \new_[2540]_ ;
  assign \new_[2547]_  = ~A201 & A200;
  assign \new_[2551]_  = A300 & A298;
  assign \new_[2552]_  = ~A202 & \new_[2551]_ ;
  assign \new_[2553]_  = \new_[2552]_  & \new_[2547]_ ;
  assign \new_[2556]_  = ~A167 & A170;
  assign \new_[2559]_  = ~A199 & A166;
  assign \new_[2560]_  = \new_[2559]_  & \new_[2556]_ ;
  assign \new_[2563]_  = ~A202 & ~A200;
  assign \new_[2567]_  = A302 & ~A299;
  assign \new_[2568]_  = A298 & \new_[2567]_ ;
  assign \new_[2569]_  = \new_[2568]_  & \new_[2563]_ ;
  assign \new_[2572]_  = ~A167 & A170;
  assign \new_[2575]_  = ~A199 & A166;
  assign \new_[2576]_  = \new_[2575]_  & \new_[2572]_ ;
  assign \new_[2579]_  = ~A202 & ~A200;
  assign \new_[2583]_  = A302 & A299;
  assign \new_[2584]_  = ~A298 & \new_[2583]_ ;
  assign \new_[2585]_  = \new_[2584]_  & \new_[2579]_ ;
  assign \new_[2588]_  = ~A167 & ~A169;
  assign \new_[2591]_  = ~A199 & ~A166;
  assign \new_[2592]_  = \new_[2591]_  & \new_[2588]_ ;
  assign \new_[2595]_  = A203 & A200;
  assign \new_[2599]_  = A302 & ~A299;
  assign \new_[2600]_  = A298 & \new_[2599]_ ;
  assign \new_[2601]_  = \new_[2600]_  & \new_[2595]_ ;
  assign \new_[2604]_  = ~A167 & ~A169;
  assign \new_[2607]_  = ~A199 & ~A166;
  assign \new_[2608]_  = \new_[2607]_  & \new_[2604]_ ;
  assign \new_[2611]_  = A203 & A200;
  assign \new_[2615]_  = A302 & A299;
  assign \new_[2616]_  = ~A298 & \new_[2615]_ ;
  assign \new_[2617]_  = \new_[2616]_  & \new_[2611]_ ;
  assign \new_[2620]_  = ~A167 & ~A169;
  assign \new_[2623]_  = A199 & ~A166;
  assign \new_[2624]_  = \new_[2623]_  & \new_[2620]_ ;
  assign \new_[2627]_  = A203 & ~A200;
  assign \new_[2631]_  = A302 & ~A299;
  assign \new_[2632]_  = A298 & \new_[2631]_ ;
  assign \new_[2633]_  = \new_[2632]_  & \new_[2627]_ ;
  assign \new_[2636]_  = ~A167 & ~A169;
  assign \new_[2639]_  = A199 & ~A166;
  assign \new_[2640]_  = \new_[2639]_  & \new_[2636]_ ;
  assign \new_[2643]_  = A203 & ~A200;
  assign \new_[2647]_  = A302 & A299;
  assign \new_[2648]_  = ~A298 & \new_[2647]_ ;
  assign \new_[2649]_  = \new_[2648]_  & \new_[2643]_ ;
  assign \new_[2652]_  = ~A168 & ~A169;
  assign \new_[2655]_  = A166 & A167;
  assign \new_[2656]_  = \new_[2655]_  & \new_[2652]_ ;
  assign \new_[2659]_  = A201 & A199;
  assign \new_[2663]_  = A302 & ~A299;
  assign \new_[2664]_  = A298 & \new_[2663]_ ;
  assign \new_[2665]_  = \new_[2664]_  & \new_[2659]_ ;
  assign \new_[2668]_  = ~A168 & ~A169;
  assign \new_[2671]_  = A166 & A167;
  assign \new_[2672]_  = \new_[2671]_  & \new_[2668]_ ;
  assign \new_[2675]_  = A201 & A199;
  assign \new_[2679]_  = A302 & A299;
  assign \new_[2680]_  = ~A298 & \new_[2679]_ ;
  assign \new_[2681]_  = \new_[2680]_  & \new_[2675]_ ;
  assign \new_[2684]_  = ~A168 & ~A169;
  assign \new_[2687]_  = A166 & A167;
  assign \new_[2688]_  = \new_[2687]_  & \new_[2684]_ ;
  assign \new_[2691]_  = A201 & A200;
  assign \new_[2695]_  = A302 & ~A299;
  assign \new_[2696]_  = A298 & \new_[2695]_ ;
  assign \new_[2697]_  = \new_[2696]_  & \new_[2691]_ ;
  assign \new_[2700]_  = ~A168 & ~A169;
  assign \new_[2703]_  = A166 & A167;
  assign \new_[2704]_  = \new_[2703]_  & \new_[2700]_ ;
  assign \new_[2707]_  = A201 & A200;
  assign \new_[2711]_  = A302 & A299;
  assign \new_[2712]_  = ~A298 & \new_[2711]_ ;
  assign \new_[2713]_  = \new_[2712]_  & \new_[2707]_ ;
  assign \new_[2716]_  = ~A168 & ~A169;
  assign \new_[2719]_  = A166 & A167;
  assign \new_[2720]_  = \new_[2719]_  & \new_[2716]_ ;
  assign \new_[2723]_  = A200 & ~A199;
  assign \new_[2727]_  = A300 & A299;
  assign \new_[2728]_  = A203 & \new_[2727]_ ;
  assign \new_[2729]_  = \new_[2728]_  & \new_[2723]_ ;
  assign \new_[2732]_  = ~A168 & ~A169;
  assign \new_[2735]_  = A166 & A167;
  assign \new_[2736]_  = \new_[2735]_  & \new_[2732]_ ;
  assign \new_[2739]_  = A200 & ~A199;
  assign \new_[2743]_  = A300 & A298;
  assign \new_[2744]_  = A203 & \new_[2743]_ ;
  assign \new_[2745]_  = \new_[2744]_  & \new_[2739]_ ;
  assign \new_[2748]_  = ~A168 & ~A169;
  assign \new_[2751]_  = A166 & A167;
  assign \new_[2752]_  = \new_[2751]_  & \new_[2748]_ ;
  assign \new_[2755]_  = ~A200 & A199;
  assign \new_[2759]_  = A300 & A299;
  assign \new_[2760]_  = A203 & \new_[2759]_ ;
  assign \new_[2761]_  = \new_[2760]_  & \new_[2755]_ ;
  assign \new_[2764]_  = ~A168 & ~A169;
  assign \new_[2767]_  = A166 & A167;
  assign \new_[2768]_  = \new_[2767]_  & \new_[2764]_ ;
  assign \new_[2771]_  = ~A200 & A199;
  assign \new_[2775]_  = A300 & A298;
  assign \new_[2776]_  = A203 & \new_[2775]_ ;
  assign \new_[2777]_  = \new_[2776]_  & \new_[2771]_ ;
  assign \new_[2780]_  = ~A169 & ~A170;
  assign \new_[2783]_  = ~A199 & ~A168;
  assign \new_[2784]_  = \new_[2783]_  & \new_[2780]_ ;
  assign \new_[2787]_  = A203 & A200;
  assign \new_[2791]_  = A302 & ~A299;
  assign \new_[2792]_  = A298 & \new_[2791]_ ;
  assign \new_[2793]_  = \new_[2792]_  & \new_[2787]_ ;
  assign \new_[2796]_  = ~A169 & ~A170;
  assign \new_[2799]_  = ~A199 & ~A168;
  assign \new_[2800]_  = \new_[2799]_  & \new_[2796]_ ;
  assign \new_[2803]_  = A203 & A200;
  assign \new_[2807]_  = A302 & A299;
  assign \new_[2808]_  = ~A298 & \new_[2807]_ ;
  assign \new_[2809]_  = \new_[2808]_  & \new_[2803]_ ;
  assign \new_[2812]_  = ~A169 & ~A170;
  assign \new_[2815]_  = A199 & ~A168;
  assign \new_[2816]_  = \new_[2815]_  & \new_[2812]_ ;
  assign \new_[2819]_  = A203 & ~A200;
  assign \new_[2823]_  = A302 & ~A299;
  assign \new_[2824]_  = A298 & \new_[2823]_ ;
  assign \new_[2825]_  = \new_[2824]_  & \new_[2819]_ ;
  assign \new_[2828]_  = ~A169 & ~A170;
  assign \new_[2831]_  = A199 & ~A168;
  assign \new_[2832]_  = \new_[2831]_  & \new_[2828]_ ;
  assign \new_[2835]_  = A203 & ~A200;
  assign \new_[2839]_  = A302 & A299;
  assign \new_[2840]_  = ~A298 & \new_[2839]_ ;
  assign \new_[2841]_  = \new_[2840]_  & \new_[2835]_ ;
  assign \new_[2844]_  = A167 & A170;
  assign \new_[2848]_  = A200 & A199;
  assign \new_[2849]_  = ~A166 & \new_[2848]_ ;
  assign \new_[2850]_  = \new_[2849]_  & \new_[2844]_ ;
  assign \new_[2853]_  = ~A202 & ~A201;
  assign \new_[2857]_  = A302 & ~A299;
  assign \new_[2858]_  = A298 & \new_[2857]_ ;
  assign \new_[2859]_  = \new_[2858]_  & \new_[2853]_ ;
  assign \new_[2862]_  = A167 & A170;
  assign \new_[2866]_  = A200 & A199;
  assign \new_[2867]_  = ~A166 & \new_[2866]_ ;
  assign \new_[2868]_  = \new_[2867]_  & \new_[2862]_ ;
  assign \new_[2871]_  = ~A202 & ~A201;
  assign \new_[2875]_  = A302 & A299;
  assign \new_[2876]_  = ~A298 & \new_[2875]_ ;
  assign \new_[2877]_  = \new_[2876]_  & \new_[2871]_ ;
  assign \new_[2880]_  = ~A167 & A170;
  assign \new_[2884]_  = A200 & A199;
  assign \new_[2885]_  = A166 & \new_[2884]_ ;
  assign \new_[2886]_  = \new_[2885]_  & \new_[2880]_ ;
  assign \new_[2889]_  = ~A202 & ~A201;
  assign \new_[2893]_  = A302 & ~A299;
  assign \new_[2894]_  = A298 & \new_[2893]_ ;
  assign \new_[2895]_  = \new_[2894]_  & \new_[2889]_ ;
  assign \new_[2898]_  = ~A167 & A170;
  assign \new_[2902]_  = A200 & A199;
  assign \new_[2903]_  = A166 & \new_[2902]_ ;
  assign \new_[2904]_  = \new_[2903]_  & \new_[2898]_ ;
  assign \new_[2907]_  = ~A202 & ~A201;
  assign \new_[2911]_  = A302 & A299;
  assign \new_[2912]_  = ~A298 & \new_[2911]_ ;
  assign \new_[2913]_  = \new_[2912]_  & \new_[2907]_ ;
  assign \new_[2916]_  = ~A168 & ~A169;
  assign \new_[2920]_  = ~A199 & A166;
  assign \new_[2921]_  = A167 & \new_[2920]_ ;
  assign \new_[2922]_  = \new_[2921]_  & \new_[2916]_ ;
  assign \new_[2925]_  = A203 & A200;
  assign \new_[2929]_  = A302 & ~A299;
  assign \new_[2930]_  = A298 & \new_[2929]_ ;
  assign \new_[2931]_  = \new_[2930]_  & \new_[2925]_ ;
  assign \new_[2934]_  = ~A168 & ~A169;
  assign \new_[2938]_  = ~A199 & A166;
  assign \new_[2939]_  = A167 & \new_[2938]_ ;
  assign \new_[2940]_  = \new_[2939]_  & \new_[2934]_ ;
  assign \new_[2943]_  = A203 & A200;
  assign \new_[2947]_  = A302 & A299;
  assign \new_[2948]_  = ~A298 & \new_[2947]_ ;
  assign \new_[2949]_  = \new_[2948]_  & \new_[2943]_ ;
  assign \new_[2952]_  = ~A168 & ~A169;
  assign \new_[2956]_  = A199 & A166;
  assign \new_[2957]_  = A167 & \new_[2956]_ ;
  assign \new_[2958]_  = \new_[2957]_  & \new_[2952]_ ;
  assign \new_[2961]_  = A203 & ~A200;
  assign \new_[2965]_  = A302 & ~A299;
  assign \new_[2966]_  = A298 & \new_[2965]_ ;
  assign \new_[2967]_  = \new_[2966]_  & \new_[2961]_ ;
  assign \new_[2970]_  = ~A168 & ~A169;
  assign \new_[2974]_  = A199 & A166;
  assign \new_[2975]_  = A167 & \new_[2974]_ ;
  assign \new_[2976]_  = \new_[2975]_  & \new_[2970]_ ;
  assign \new_[2979]_  = A203 & ~A200;
  assign \new_[2983]_  = A302 & A299;
  assign \new_[2984]_  = ~A298 & \new_[2983]_ ;
  assign \new_[2985]_  = \new_[2984]_  & \new_[2979]_ ;
endmodule


