// Benchmark "testing" written by ABC on Thu Oct  8 22:16:31 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A75  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A75;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[768]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[778]_ ,
    \new_[779]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ , \new_[786]_ ,
    \new_[790]_ , \new_[791]_ , \new_[795]_ , \new_[796]_ , \new_[797]_ ,
    \new_[801]_ , \new_[802]_ , \new_[806]_ , \new_[807]_ , \new_[808]_ ,
    \new_[809]_ , \new_[810]_ , \new_[814]_ , \new_[815]_ , \new_[819]_ ,
    \new_[820]_ , \new_[821]_ , \new_[825]_ , \new_[826]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[837]_ , \new_[838]_ ,
    \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[848]_ , \new_[849]_ ,
    \new_[853]_ , \new_[854]_ , \new_[855]_ , \new_[856]_ , \new_[857]_ ,
    \new_[858]_ , \new_[862]_ , \new_[863]_ , \new_[867]_ , \new_[868]_ ,
    \new_[869]_ , \new_[873]_ , \new_[874]_ , \new_[878]_ , \new_[879]_ ,
    \new_[880]_ , \new_[881]_ , \new_[885]_ , \new_[886]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[896]_ , \new_[897]_ , \new_[901]_ ,
    \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ , \new_[909]_ ,
    \new_[910]_ , \new_[914]_ , \new_[915]_ , \new_[916]_ , \new_[920]_ ,
    \new_[921]_ , \new_[925]_ , \new_[926]_ , \new_[927]_ , \new_[928]_ ,
    \new_[932]_ , \new_[933]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ ,
    \new_[943]_ , \new_[944]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[958]_ ,
    \new_[959]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ , \new_[969]_ ,
    \new_[970]_ , \new_[974]_ , \new_[975]_ , \new_[976]_ , \new_[977]_ ,
    \new_[981]_ , \new_[982]_ , \new_[986]_ , \new_[987]_ , \new_[988]_ ,
    \new_[992]_ , \new_[993]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ ,
    \new_[1000]_ , \new_[1001]_ , \new_[1005]_ , \new_[1006]_ ,
    \new_[1010]_ , \new_[1011]_ , \new_[1012]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1021]_ , \new_[1022]_ , \new_[1023]_ ,
    \new_[1024]_ , \new_[1028]_ , \new_[1029]_ , \new_[1033]_ ,
    \new_[1034]_ , \new_[1035]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1044]_ , \new_[1045]_ , \new_[1046]_ , \new_[1047]_ ,
    \new_[1048]_ , \new_[1049]_ , \new_[1053]_ , \new_[1054]_ ,
    \new_[1058]_ , \new_[1059]_ , \new_[1060]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1069]_ , \new_[1070]_ , \new_[1071]_ ,
    \new_[1072]_ , \new_[1076]_ , \new_[1077]_ , \new_[1081]_ ,
    \new_[1082]_ , \new_[1083]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1092]_ , \new_[1093]_ , \new_[1094]_ , \new_[1095]_ ,
    \new_[1096]_ , \new_[1100]_ , \new_[1101]_ , \new_[1105]_ ,
    \new_[1106]_ , \new_[1107]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1116]_ , \new_[1117]_ , \new_[1118]_ , \new_[1119]_ ,
    \new_[1123]_ , \new_[1124]_ , \new_[1128]_ , \new_[1129]_ ,
    \new_[1130]_ , \new_[1134]_ , \new_[1135]_ , \new_[1139]_ ,
    \new_[1140]_ , \new_[1141]_ , \new_[1142]_ , \new_[1143]_ ,
    \new_[1144]_ , \new_[1145]_ , \new_[1146]_ , \new_[1149]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1159]_ ,
    \new_[1160]_ , \new_[1164]_ , \new_[1165]_ , \new_[1166]_ ,
    \new_[1167]_ , \new_[1171]_ , \new_[1172]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1182]_ , \new_[1183]_ ,
    \new_[1187]_ , \new_[1188]_ , \new_[1189]_ , \new_[1190]_ ,
    \new_[1191]_ , \new_[1195]_ , \new_[1196]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1206]_ , \new_[1207]_ ,
    \new_[1211]_ , \new_[1212]_ , \new_[1213]_ , \new_[1214]_ ,
    \new_[1218]_ , \new_[1219]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1229]_ , \new_[1230]_ , \new_[1234]_ ,
    \new_[1235]_ , \new_[1236]_ , \new_[1237]_ , \new_[1238]_ ,
    \new_[1239]_ , \new_[1243]_ , \new_[1244]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1254]_ , \new_[1255]_ ,
    \new_[1259]_ , \new_[1260]_ , \new_[1261]_ , \new_[1262]_ ,
    \new_[1266]_ , \new_[1267]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1277]_ , \new_[1278]_ , \new_[1282]_ ,
    \new_[1283]_ , \new_[1284]_ , \new_[1285]_ , \new_[1286]_ ,
    \new_[1290]_ , \new_[1291]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1301]_ , \new_[1302]_ , \new_[1306]_ ,
    \new_[1307]_ , \new_[1308]_ , \new_[1309]_ , \new_[1313]_ ,
    \new_[1314]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1324]_ , \new_[1325]_ , \new_[1329]_ , \new_[1330]_ ,
    \new_[1331]_ , \new_[1332]_ , \new_[1333]_ , \new_[1334]_ ,
    \new_[1335]_ , \new_[1339]_ , \new_[1340]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1350]_ , \new_[1351]_ ,
    \new_[1355]_ , \new_[1356]_ , \new_[1357]_ , \new_[1358]_ ,
    \new_[1362]_ , \new_[1363]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1373]_ , \new_[1374]_ , \new_[1378]_ ,
    \new_[1379]_ , \new_[1380]_ , \new_[1381]_ , \new_[1382]_ ,
    \new_[1386]_ , \new_[1387]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1397]_ , \new_[1398]_ , \new_[1402]_ ,
    \new_[1403]_ , \new_[1404]_ , \new_[1405]_ , \new_[1409]_ ,
    \new_[1410]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1420]_ , \new_[1421]_ , \new_[1425]_ , \new_[1426]_ ,
    \new_[1427]_ , \new_[1428]_ , \new_[1429]_ , \new_[1430]_ ,
    \new_[1434]_ , \new_[1435]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1445]_ , \new_[1446]_ , \new_[1450]_ ,
    \new_[1451]_ , \new_[1452]_ , \new_[1453]_ , \new_[1457]_ ,
    \new_[1458]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1468]_ , \new_[1469]_ , \new_[1473]_ , \new_[1474]_ ,
    \new_[1475]_ , \new_[1476]_ , \new_[1477]_ , \new_[1481]_ ,
    \new_[1482]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1492]_ , \new_[1493]_ , \new_[1497]_ , \new_[1498]_ ,
    \new_[1499]_ , \new_[1500]_ , \new_[1504]_ , \new_[1505]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1515]_ ,
    \new_[1516]_ , \new_[1520]_ , \new_[1521]_ , \new_[1522]_ ,
    \new_[1523]_ , \new_[1524]_ , \new_[1525]_ , \new_[1526]_ ,
    \new_[1527]_ , \new_[1528]_ , \new_[1531]_ , \new_[1535]_ ,
    \new_[1536]_ , \new_[1537]_ , \new_[1541]_ , \new_[1542]_ ,
    \new_[1546]_ , \new_[1547]_ , \new_[1548]_ , \new_[1549]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1558]_ , \new_[1559]_ ,
    \new_[1560]_ , \new_[1564]_ , \new_[1565]_ , \new_[1569]_ ,
    \new_[1570]_ , \new_[1571]_ , \new_[1572]_ , \new_[1573]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1582]_ , \new_[1583]_ ,
    \new_[1584]_ , \new_[1588]_ , \new_[1589]_ , \new_[1593]_ ,
    \new_[1594]_ , \new_[1595]_ , \new_[1596]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1605]_ , \new_[1606]_ , \new_[1607]_ ,
    \new_[1611]_ , \new_[1612]_ , \new_[1616]_ , \new_[1617]_ ,
    \new_[1618]_ , \new_[1619]_ , \new_[1620]_ , \new_[1621]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1630]_ , \new_[1631]_ ,
    \new_[1632]_ , \new_[1636]_ , \new_[1637]_ , \new_[1641]_ ,
    \new_[1642]_ , \new_[1643]_ , \new_[1644]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1653]_ , \new_[1654]_ , \new_[1655]_ ,
    \new_[1659]_ , \new_[1660]_ , \new_[1664]_ , \new_[1665]_ ,
    \new_[1666]_ , \new_[1667]_ , \new_[1668]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1677]_ , \new_[1678]_ , \new_[1679]_ ,
    \new_[1683]_ , \new_[1684]_ , \new_[1688]_ , \new_[1689]_ ,
    \new_[1690]_ , \new_[1691]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1700]_ , \new_[1701]_ , \new_[1702]_ , \new_[1706]_ ,
    \new_[1707]_ , \new_[1711]_ , \new_[1712]_ , \new_[1713]_ ,
    \new_[1714]_ , \new_[1715]_ , \new_[1716]_ , \new_[1717]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1726]_ , \new_[1727]_ ,
    \new_[1728]_ , \new_[1732]_ , \new_[1733]_ , \new_[1737]_ ,
    \new_[1738]_ , \new_[1739]_ , \new_[1740]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1749]_ , \new_[1750]_ , \new_[1751]_ ,
    \new_[1755]_ , \new_[1756]_ , \new_[1760]_ , \new_[1761]_ ,
    \new_[1762]_ , \new_[1763]_ , \new_[1764]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1773]_ , \new_[1774]_ , \new_[1775]_ ,
    \new_[1779]_ , \new_[1780]_ , \new_[1784]_ , \new_[1785]_ ,
    \new_[1786]_ , \new_[1787]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1796]_ , \new_[1797]_ , \new_[1798]_ , \new_[1802]_ ,
    \new_[1803]_ , \new_[1807]_ , \new_[1808]_ , \new_[1809]_ ,
    \new_[1810]_ , \new_[1811]_ , \new_[1812]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1821]_ , \new_[1822]_ , \new_[1823]_ ,
    \new_[1827]_ , \new_[1828]_ , \new_[1832]_ , \new_[1833]_ ,
    \new_[1834]_ , \new_[1835]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1844]_ , \new_[1845]_ , \new_[1846]_ , \new_[1850]_ ,
    \new_[1851]_ , \new_[1855]_ , \new_[1856]_ , \new_[1857]_ ,
    \new_[1858]_ , \new_[1859]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1868]_ , \new_[1869]_ , \new_[1870]_ , \new_[1874]_ ,
    \new_[1875]_ , \new_[1879]_ , \new_[1880]_ , \new_[1881]_ ,
    \new_[1882]_ , \new_[1886]_ , \new_[1887]_ , \new_[1891]_ ,
    \new_[1892]_ , \new_[1893]_ , \new_[1897]_ , \new_[1898]_ ,
    \new_[1902]_ , \new_[1903]_ , \new_[1904]_ , \new_[1905]_ ,
    \new_[1906]_ , \new_[1907]_ , \new_[1908]_ , \new_[1909]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1918]_ , \new_[1919]_ ,
    \new_[1920]_ , \new_[1924]_ , \new_[1925]_ , \new_[1929]_ ,
    \new_[1930]_ , \new_[1931]_ , \new_[1932]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1941]_ , \new_[1942]_ , \new_[1943]_ ,
    \new_[1947]_ , \new_[1948]_ , \new_[1952]_ , \new_[1953]_ ,
    \new_[1954]_ , \new_[1955]_ , \new_[1956]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1965]_ , \new_[1966]_ , \new_[1967]_ ,
    \new_[1971]_ , \new_[1972]_ , \new_[1976]_ , \new_[1977]_ ,
    \new_[1978]_ , \new_[1979]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1988]_ , \new_[1989]_ , \new_[1990]_ , \new_[1994]_ ,
    \new_[1995]_ , \new_[1999]_ , \new_[2000]_ , \new_[2001]_ ,
    \new_[2002]_ , \new_[2003]_ , \new_[2004]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2013]_ , \new_[2014]_ , \new_[2015]_ ,
    \new_[2019]_ , \new_[2020]_ , \new_[2024]_ , \new_[2025]_ ,
    \new_[2026]_ , \new_[2027]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2036]_ , \new_[2037]_ , \new_[2038]_ , \new_[2042]_ ,
    \new_[2043]_ , \new_[2047]_ , \new_[2048]_ , \new_[2049]_ ,
    \new_[2050]_ , \new_[2051]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2060]_ , \new_[2061]_ , \new_[2062]_ , \new_[2066]_ ,
    \new_[2067]_ , \new_[2071]_ , \new_[2072]_ , \new_[2073]_ ,
    \new_[2074]_ , \new_[2078]_ , \new_[2079]_ , \new_[2083]_ ,
    \new_[2084]_ , \new_[2085]_ , \new_[2089]_ , \new_[2090]_ ,
    \new_[2094]_ , \new_[2095]_ , \new_[2096]_ , \new_[2097]_ ,
    \new_[2098]_ , \new_[2099]_ , \new_[2100]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2109]_ , \new_[2110]_ , \new_[2111]_ ,
    \new_[2115]_ , \new_[2116]_ , \new_[2120]_ , \new_[2121]_ ,
    \new_[2122]_ , \new_[2123]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2132]_ , \new_[2133]_ , \new_[2134]_ , \new_[2138]_ ,
    \new_[2139]_ , \new_[2143]_ , \new_[2144]_ , \new_[2145]_ ,
    \new_[2146]_ , \new_[2147]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2156]_ , \new_[2157]_ , \new_[2158]_ , \new_[2162]_ ,
    \new_[2163]_ , \new_[2167]_ , \new_[2168]_ , \new_[2169]_ ,
    \new_[2170]_ , \new_[2174]_ , \new_[2175]_ , \new_[2179]_ ,
    \new_[2180]_ , \new_[2181]_ , \new_[2185]_ , \new_[2186]_ ,
    \new_[2190]_ , \new_[2191]_ , \new_[2192]_ , \new_[2193]_ ,
    \new_[2194]_ , \new_[2195]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2204]_ , \new_[2205]_ , \new_[2206]_ , \new_[2210]_ ,
    \new_[2211]_ , \new_[2215]_ , \new_[2216]_ , \new_[2217]_ ,
    \new_[2218]_ , \new_[2222]_ , \new_[2223]_ , \new_[2227]_ ,
    \new_[2228]_ , \new_[2229]_ , \new_[2233]_ , \new_[2234]_ ,
    \new_[2238]_ , \new_[2239]_ , \new_[2240]_ , \new_[2241]_ ,
    \new_[2242]_ , \new_[2246]_ , \new_[2247]_ , \new_[2251]_ ,
    \new_[2252]_ , \new_[2253]_ , \new_[2257]_ , \new_[2258]_ ,
    \new_[2262]_ , \new_[2263]_ , \new_[2264]_ , \new_[2265]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2274]_ , \new_[2275]_ ,
    \new_[2276]_ , \new_[2280]_ , \new_[2281]_ , \new_[2285]_ ,
    \new_[2286]_ , \new_[2287]_ , \new_[2288]_ , \new_[2289]_ ,
    \new_[2290]_ , \new_[2291]_ , \new_[2292]_ , \new_[2293]_ ,
    \new_[2296]_ , \new_[2299]_ , \new_[2302]_ , \new_[2305]_ ,
    \new_[2308]_ , \new_[2312]_ , \new_[2313]_ , \new_[2316]_ ,
    \new_[2320]_ , \new_[2321]_ , \new_[2324]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2332]_ , \new_[2336]_ , \new_[2337]_ ,
    \new_[2340]_ , \new_[2344]_ , \new_[2345]_ , \new_[2349]_ ,
    \new_[2350]_ , \new_[2354]_ , \new_[2355]_ , \new_[2359]_ ,
    \new_[2360]_ , \new_[2364]_ , \new_[2365]_ , \new_[2369]_ ,
    \new_[2370]_ , \new_[2374]_ , \new_[2375]_ , \new_[2379]_ ,
    \new_[2380]_ , \new_[2384]_ , \new_[2385]_ , \new_[2389]_ ,
    \new_[2390]_ , \new_[2394]_ , \new_[2395]_ , \new_[2399]_ ,
    \new_[2400]_ , \new_[2404]_ , \new_[2405]_ , \new_[2409]_ ,
    \new_[2410]_ , \new_[2414]_ , \new_[2415]_ , \new_[2419]_ ,
    \new_[2420]_ , \new_[2424]_ , \new_[2425]_ , \new_[2429]_ ,
    \new_[2430]_ , \new_[2434]_ , \new_[2435]_ , \new_[2439]_ ,
    \new_[2440]_ , \new_[2444]_ , \new_[2445]_ , \new_[2449]_ ,
    \new_[2450]_ , \new_[2453]_ , \new_[2456]_ , \new_[2457]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2465]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2473]_ , \new_[2474]_ , \new_[2477]_ ,
    \new_[2480]_ , \new_[2481]_ , \new_[2485]_ , \new_[2486]_ ,
    \new_[2489]_ , \new_[2492]_ , \new_[2493]_ , \new_[2497]_ ,
    \new_[2498]_ , \new_[2501]_ , \new_[2504]_ , \new_[2505]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2513]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2521]_ , \new_[2522]_ , \new_[2525]_ ,
    \new_[2528]_ , \new_[2529]_ , \new_[2533]_ , \new_[2534]_ ,
    \new_[2537]_ , \new_[2540]_ , \new_[2541]_ , \new_[2545]_ ,
    \new_[2546]_ , \new_[2549]_ , \new_[2552]_ , \new_[2553]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2561]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2569]_ , \new_[2570]_ , \new_[2573]_ ,
    \new_[2576]_ , \new_[2577]_ , \new_[2581]_ , \new_[2582]_ ,
    \new_[2585]_ , \new_[2588]_ , \new_[2589]_ , \new_[2593]_ ,
    \new_[2594]_ , \new_[2597]_ , \new_[2600]_ , \new_[2601]_ ,
    \new_[2605]_ , \new_[2606]_ , \new_[2609]_ , \new_[2612]_ ,
    \new_[2613]_ , \new_[2617]_ , \new_[2618]_ , \new_[2621]_ ,
    \new_[2624]_ , \new_[2625]_ , \new_[2629]_ , \new_[2630]_ ,
    \new_[2633]_ , \new_[2636]_ , \new_[2637]_ , \new_[2641]_ ,
    \new_[2642]_ , \new_[2645]_ , \new_[2648]_ , \new_[2649]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2657]_ , \new_[2660]_ ,
    \new_[2661]_ , \new_[2665]_ , \new_[2666]_ , \new_[2669]_ ,
    \new_[2672]_ , \new_[2673]_ , \new_[2677]_ , \new_[2678]_ ,
    \new_[2681]_ , \new_[2684]_ , \new_[2685]_ , \new_[2689]_ ,
    \new_[2690]_ , \new_[2693]_ , \new_[2696]_ , \new_[2697]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2705]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2713]_ , \new_[2714]_ , \new_[2717]_ ,
    \new_[2720]_ , \new_[2721]_ , \new_[2725]_ , \new_[2726]_ ,
    \new_[2729]_ , \new_[2732]_ , \new_[2733]_ , \new_[2737]_ ,
    \new_[2738]_ , \new_[2741]_ , \new_[2744]_ , \new_[2745]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2753]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2761]_ , \new_[2762]_ , \new_[2765]_ ,
    \new_[2768]_ , \new_[2769]_ , \new_[2773]_ , \new_[2774]_ ,
    \new_[2777]_ , \new_[2780]_ , \new_[2781]_ , \new_[2784]_ ,
    \new_[2787]_ , \new_[2788]_ , \new_[2791]_ , \new_[2794]_ ,
    \new_[2795]_ , \new_[2798]_ , \new_[2801]_ , \new_[2802]_ ,
    \new_[2805]_ , \new_[2808]_ , \new_[2809]_ , \new_[2812]_ ,
    \new_[2815]_ , \new_[2816]_ , \new_[2819]_ , \new_[2822]_ ,
    \new_[2823]_ , \new_[2826]_ , \new_[2829]_ , \new_[2830]_ ,
    \new_[2833]_ , \new_[2836]_ , \new_[2837]_ , \new_[2840]_ ,
    \new_[2843]_ , \new_[2844]_ , \new_[2847]_ , \new_[2850]_ ,
    \new_[2851]_ , \new_[2854]_ , \new_[2857]_ , \new_[2858]_ ,
    \new_[2861]_ , \new_[2864]_ , \new_[2865]_ , \new_[2868]_ ,
    \new_[2871]_ , \new_[2872]_ , \new_[2875]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2882]_ , \new_[2885]_ , \new_[2886]_ ,
    \new_[2889]_ , \new_[2892]_ , \new_[2893]_ , \new_[2896]_ ,
    \new_[2899]_ , \new_[2900]_ , \new_[2903]_ , \new_[2906]_ ,
    \new_[2907]_ , \new_[2910]_ , \new_[2913]_ , \new_[2914]_ ,
    \new_[2917]_ , \new_[2920]_ , \new_[2921]_ , \new_[2924]_ ,
    \new_[2927]_ , \new_[2928]_ , \new_[2931]_ , \new_[2934]_ ,
    \new_[2935]_ , \new_[2938]_ , \new_[2941]_ , \new_[2942]_ ,
    \new_[2945]_ , \new_[2948]_ , \new_[2949]_ , \new_[2952]_ ,
    \new_[2955]_ , \new_[2956]_ , \new_[2959]_ , \new_[2962]_ ,
    \new_[2963]_ , \new_[2966]_ , \new_[2969]_ , \new_[2970]_ ,
    \new_[2973]_ , \new_[2976]_ , \new_[2977]_ , \new_[2980]_ ,
    \new_[2983]_ , \new_[2984]_ , \new_[2987]_ , \new_[2990]_ ,
    \new_[2991]_ , \new_[2994]_ , \new_[2997]_ , \new_[2998]_ ,
    \new_[3001]_ , \new_[3004]_ , \new_[3005]_ , \new_[3008]_ ,
    \new_[3011]_ , \new_[3012]_ , \new_[3015]_ , \new_[3018]_ ,
    \new_[3019]_ , \new_[3022]_ , \new_[3025]_ , \new_[3026]_ ,
    \new_[3029]_ , \new_[3032]_ , \new_[3033]_ , \new_[3036]_ ,
    \new_[3039]_ , \new_[3040]_ , \new_[3043]_ , \new_[3046]_ ,
    \new_[3047]_ , \new_[3050]_ , \new_[3053]_ , \new_[3054]_ ,
    \new_[3057]_ , \new_[3060]_ , \new_[3061]_ , \new_[3064]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3071]_ , \new_[3074]_ ,
    \new_[3075]_ , \new_[3078]_ , \new_[3081]_ , \new_[3082]_ ,
    \new_[3085]_ , \new_[3088]_ , \new_[3089]_ , \new_[3092]_ ,
    \new_[3095]_ , \new_[3096]_ , \new_[3099]_ , \new_[3102]_ ,
    \new_[3103]_ , \new_[3106]_ , \new_[3109]_ , \new_[3110]_ ,
    \new_[3113]_ , \new_[3116]_ , \new_[3117]_ , \new_[3120]_ ,
    \new_[3123]_ , \new_[3124]_ , \new_[3127]_ , \new_[3130]_ ,
    \new_[3131]_ , \new_[3134]_ , \new_[3137]_ , \new_[3138]_ ,
    \new_[3141]_ , \new_[3144]_ , \new_[3145]_ , \new_[3148]_ ,
    \new_[3151]_ , \new_[3152]_ , \new_[3155]_ , \new_[3158]_ ,
    \new_[3159]_ , \new_[3162]_ , \new_[3165]_ , \new_[3166]_ ,
    \new_[3169]_ , \new_[3172]_ , \new_[3173]_ , \new_[3176]_ ,
    \new_[3179]_ , \new_[3180]_ , \new_[3183]_ , \new_[3186]_ ,
    \new_[3187]_ , \new_[3190]_ , \new_[3193]_ , \new_[3194]_ ,
    \new_[3197]_ , \new_[3200]_ , \new_[3201]_ , \new_[3204]_ ,
    \new_[3207]_ , \new_[3208]_ , \new_[3211]_ , \new_[3214]_ ,
    \new_[3215]_ , \new_[3218]_ , \new_[3221]_ , \new_[3222]_ ,
    \new_[3225]_ , \new_[3228]_ , \new_[3229]_ , \new_[3232]_ ,
    \new_[3235]_ , \new_[3236]_ , \new_[3239]_ , \new_[3242]_ ,
    \new_[3243]_ , \new_[3246]_ , \new_[3249]_ , \new_[3250]_ ,
    \new_[3253]_ , \new_[3256]_ , \new_[3257]_ , \new_[3260]_ ,
    \new_[3263]_ , \new_[3264]_ , \new_[3267]_ , \new_[3270]_ ,
    \new_[3271]_ , \new_[3274]_ , \new_[3277]_ , \new_[3278]_ ,
    \new_[3281]_ , \new_[3284]_ , \new_[3285]_ , \new_[3288]_ ,
    \new_[3291]_ , \new_[3292]_ , \new_[3295]_ , \new_[3298]_ ,
    \new_[3299]_ , \new_[3302]_ , \new_[3305]_ , \new_[3306]_ ,
    \new_[3309]_ , \new_[3312]_ , \new_[3313]_ , \new_[3316]_ ,
    \new_[3319]_ , \new_[3320]_ , \new_[3323]_ , \new_[3326]_ ,
    \new_[3327]_ , \new_[3330]_ , \new_[3333]_ , \new_[3334]_ ,
    \new_[3337]_ , \new_[3340]_ , \new_[3341]_ , \new_[3344]_ ,
    \new_[3347]_ , \new_[3348]_ , \new_[3351]_ , \new_[3354]_ ,
    \new_[3355]_ , \new_[3358]_ , \new_[3361]_ , \new_[3362]_ ,
    \new_[3365]_ , \new_[3368]_ , \new_[3369]_ , \new_[3372]_ ,
    \new_[3375]_ , \new_[3376]_ , \new_[3379]_ , \new_[3382]_ ,
    \new_[3383]_ , \new_[3386]_ , \new_[3389]_ , \new_[3390]_ ,
    \new_[3393]_ , \new_[3396]_ , \new_[3397]_ , \new_[3400]_ ,
    \new_[3403]_ , \new_[3404]_ , \new_[3407]_ , \new_[3410]_ ,
    \new_[3411]_ , \new_[3414]_ , \new_[3417]_ , \new_[3418]_ ,
    \new_[3421]_ , \new_[3424]_ , \new_[3425]_ , \new_[3428]_ ,
    \new_[3431]_ , \new_[3432]_ , \new_[3435]_ , \new_[3438]_ ,
    \new_[3439]_ , \new_[3442]_ , \new_[3445]_ , \new_[3446]_ ,
    \new_[3449]_ , \new_[3452]_ , \new_[3453]_ , \new_[3456]_ ,
    \new_[3459]_ , \new_[3460]_ , \new_[3463]_ , \new_[3466]_ ,
    \new_[3467]_ , \new_[3470]_ , \new_[3473]_ , \new_[3474]_ ,
    \new_[3477]_ , \new_[3480]_ , \new_[3481]_ , \new_[3484]_ ,
    \new_[3487]_ , \new_[3488]_ , \new_[3491]_ , \new_[3494]_ ,
    \new_[3495]_ , \new_[3498]_ , \new_[3501]_ , \new_[3502]_ ,
    \new_[3505]_ , \new_[3508]_ , \new_[3509]_ , \new_[3512]_ ,
    \new_[3515]_ , \new_[3516]_ , \new_[3519]_ , \new_[3522]_ ,
    \new_[3523]_ , \new_[3526]_ , \new_[3529]_ , \new_[3530]_ ,
    \new_[3533]_ , \new_[3536]_ , \new_[3537]_ , \new_[3540]_ ,
    \new_[3543]_ , \new_[3544]_ , \new_[3547]_ , \new_[3550]_ ,
    \new_[3551]_ , \new_[3554]_ , \new_[3557]_ , \new_[3558]_ ,
    \new_[3561]_ , \new_[3564]_ , \new_[3565]_ , \new_[3568]_ ,
    \new_[3571]_ , \new_[3572]_ , \new_[3575]_ , \new_[3578]_ ,
    \new_[3579]_ , \new_[3582]_ , \new_[3585]_ , \new_[3586]_ ,
    \new_[3589]_ , \new_[3592]_ , \new_[3593]_ , \new_[3596]_ ,
    \new_[3599]_ , \new_[3600]_ , \new_[3603]_ , \new_[3606]_ ,
    \new_[3607]_ , \new_[3610]_ , \new_[3613]_ , \new_[3614]_ ,
    \new_[3617]_ , \new_[3620]_ , \new_[3621]_ , \new_[3624]_ ,
    \new_[3627]_ , \new_[3628]_ , \new_[3631]_ , \new_[3634]_ ,
    \new_[3635]_ , \new_[3638]_ , \new_[3641]_ , \new_[3642]_ ,
    \new_[3645]_ , \new_[3648]_ , \new_[3649]_ , \new_[3652]_ ,
    \new_[3655]_ , \new_[3656]_ , \new_[3659]_ , \new_[3662]_ ,
    \new_[3663]_ , \new_[3666]_ , \new_[3669]_ , \new_[3670]_ ,
    \new_[3673]_ , \new_[3676]_ , \new_[3677]_ , \new_[3680]_ ,
    \new_[3683]_ , \new_[3684]_ , \new_[3687]_ , \new_[3690]_ ,
    \new_[3691]_ , \new_[3694]_ , \new_[3697]_ , \new_[3698]_ ,
    \new_[3701]_ , \new_[3704]_ , \new_[3705]_ , \new_[3708]_ ,
    \new_[3711]_ , \new_[3712]_ , \new_[3715]_ , \new_[3718]_ ,
    \new_[3719]_ , \new_[3722]_ , \new_[3725]_ , \new_[3726]_ ,
    \new_[3729]_ , \new_[3732]_ , \new_[3733]_ , \new_[3736]_ ,
    \new_[3739]_ , \new_[3740]_ , \new_[3743]_ , \new_[3746]_ ,
    \new_[3747]_ , \new_[3750]_ , \new_[3753]_ , \new_[3754]_ ,
    \new_[3757]_ , \new_[3760]_ , \new_[3761]_ , \new_[3764]_ ,
    \new_[3767]_ , \new_[3768]_ , \new_[3771]_ , \new_[3774]_ ,
    \new_[3775]_ , \new_[3778]_ , \new_[3781]_ , \new_[3782]_ ,
    \new_[3785]_ , \new_[3788]_ , \new_[3789]_ , \new_[3792]_ ,
    \new_[3795]_ , \new_[3796]_ , \new_[3799]_ , \new_[3802]_ ,
    \new_[3803]_ , \new_[3806]_ , \new_[3809]_ , \new_[3810]_ ,
    \new_[3813]_ , \new_[3816]_ , \new_[3817]_ , \new_[3820]_ ,
    \new_[3823]_ , \new_[3824]_ , \new_[3827]_ , \new_[3830]_ ,
    \new_[3831]_ , \new_[3834]_ , \new_[3837]_ , \new_[3838]_ ,
    \new_[3841]_ , \new_[3844]_ , \new_[3845]_ , \new_[3848]_ ,
    \new_[3851]_ , \new_[3852]_ , \new_[3855]_ , \new_[3858]_ ,
    \new_[3859]_ , \new_[3862]_ , \new_[3865]_ , \new_[3866]_ ,
    \new_[3869]_ , \new_[3872]_ , \new_[3873]_ , \new_[3876]_ ,
    \new_[3879]_ , \new_[3880]_ , \new_[3883]_ , \new_[3886]_ ,
    \new_[3887]_ , \new_[3890]_ , \new_[3893]_ , \new_[3894]_ ,
    \new_[3897]_ , \new_[3900]_ , \new_[3901]_ , \new_[3904]_ ,
    \new_[3907]_ , \new_[3908]_ , \new_[3911]_ , \new_[3914]_ ,
    \new_[3915]_ , \new_[3918]_ , \new_[3921]_ , \new_[3922]_ ,
    \new_[3925]_ , \new_[3928]_ , \new_[3929]_ , \new_[3932]_ ,
    \new_[3935]_ , \new_[3936]_ , \new_[3939]_ , \new_[3942]_ ,
    \new_[3943]_ , \new_[3946]_ , \new_[3949]_ , \new_[3950]_ ,
    \new_[3953]_ , \new_[3956]_ , \new_[3957]_ , \new_[3960]_ ,
    \new_[3963]_ , \new_[3964]_ , \new_[3967]_ , \new_[3971]_ ,
    \new_[3972]_ , \new_[3973]_ , \new_[3976]_ , \new_[3979]_ ,
    \new_[3980]_ , \new_[3983]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3989]_ , \new_[3992]_ , \new_[3995]_ , \new_[3996]_ ,
    \new_[3999]_ , \new_[4003]_ , \new_[4004]_ , \new_[4005]_ ,
    \new_[4008]_ , \new_[4011]_ , \new_[4012]_ , \new_[4015]_ ,
    \new_[4019]_ , \new_[4020]_ , \new_[4021]_ , \new_[4024]_ ,
    \new_[4027]_ , \new_[4028]_ , \new_[4031]_ , \new_[4035]_ ,
    \new_[4036]_ , \new_[4037]_ , \new_[4040]_ , \new_[4043]_ ,
    \new_[4044]_ , \new_[4047]_ , \new_[4051]_ , \new_[4052]_ ,
    \new_[4053]_ , \new_[4056]_ , \new_[4059]_ , \new_[4060]_ ,
    \new_[4063]_ , \new_[4067]_ , \new_[4068]_ , \new_[4069]_ ,
    \new_[4072]_ , \new_[4075]_ , \new_[4076]_ , \new_[4079]_ ,
    \new_[4083]_ , \new_[4084]_ , \new_[4085]_ , \new_[4088]_ ,
    \new_[4091]_ , \new_[4092]_ , \new_[4095]_ , \new_[4099]_ ,
    \new_[4100]_ , \new_[4101]_ , \new_[4104]_ , \new_[4107]_ ,
    \new_[4108]_ , \new_[4111]_ , \new_[4115]_ , \new_[4116]_ ,
    \new_[4117]_ , \new_[4120]_ , \new_[4123]_ , \new_[4124]_ ,
    \new_[4127]_ , \new_[4131]_ , \new_[4132]_ , \new_[4133]_ ,
    \new_[4136]_ , \new_[4139]_ , \new_[4140]_ , \new_[4143]_ ,
    \new_[4147]_ , \new_[4148]_ , \new_[4149]_ , \new_[4152]_ ,
    \new_[4155]_ , \new_[4156]_ , \new_[4159]_ , \new_[4163]_ ,
    \new_[4164]_ , \new_[4165]_ , \new_[4168]_ , \new_[4171]_ ,
    \new_[4172]_ , \new_[4175]_ , \new_[4179]_ , \new_[4180]_ ,
    \new_[4181]_ , \new_[4184]_ , \new_[4187]_ , \new_[4188]_ ,
    \new_[4191]_ , \new_[4195]_ , \new_[4196]_ , \new_[4197]_ ,
    \new_[4200]_ , \new_[4203]_ , \new_[4204]_ , \new_[4207]_ ,
    \new_[4211]_ , \new_[4212]_ , \new_[4213]_ , \new_[4216]_ ,
    \new_[4219]_ , \new_[4220]_ , \new_[4223]_ , \new_[4227]_ ,
    \new_[4228]_ , \new_[4229]_ , \new_[4232]_ , \new_[4235]_ ,
    \new_[4236]_ , \new_[4239]_ , \new_[4243]_ , \new_[4244]_ ,
    \new_[4245]_ , \new_[4248]_ , \new_[4251]_ , \new_[4252]_ ,
    \new_[4255]_ , \new_[4259]_ , \new_[4260]_ , \new_[4261]_ ,
    \new_[4264]_ , \new_[4267]_ , \new_[4268]_ , \new_[4271]_ ,
    \new_[4275]_ , \new_[4276]_ , \new_[4277]_ , \new_[4280]_ ,
    \new_[4283]_ , \new_[4284]_ , \new_[4287]_ , \new_[4291]_ ,
    \new_[4292]_ , \new_[4293]_ , \new_[4296]_ , \new_[4299]_ ,
    \new_[4300]_ , \new_[4303]_ , \new_[4307]_ , \new_[4308]_ ,
    \new_[4309]_ , \new_[4312]_ , \new_[4315]_ , \new_[4316]_ ,
    \new_[4319]_ , \new_[4323]_ , \new_[4324]_ , \new_[4325]_ ,
    \new_[4328]_ , \new_[4331]_ , \new_[4332]_ , \new_[4335]_ ,
    \new_[4339]_ , \new_[4340]_ , \new_[4341]_ , \new_[4344]_ ,
    \new_[4347]_ , \new_[4348]_ , \new_[4351]_ , \new_[4355]_ ,
    \new_[4356]_ , \new_[4357]_ , \new_[4360]_ , \new_[4363]_ ,
    \new_[4364]_ , \new_[4367]_ , \new_[4371]_ , \new_[4372]_ ,
    \new_[4373]_ , \new_[4376]_ , \new_[4379]_ , \new_[4380]_ ,
    \new_[4383]_ , \new_[4387]_ , \new_[4388]_ , \new_[4389]_ ,
    \new_[4392]_ , \new_[4395]_ , \new_[4396]_ , \new_[4399]_ ,
    \new_[4403]_ , \new_[4404]_ , \new_[4405]_ , \new_[4408]_ ,
    \new_[4411]_ , \new_[4412]_ , \new_[4415]_ , \new_[4419]_ ,
    \new_[4420]_ , \new_[4421]_ , \new_[4424]_ , \new_[4427]_ ,
    \new_[4428]_ , \new_[4431]_ , \new_[4435]_ , \new_[4436]_ ,
    \new_[4437]_ , \new_[4440]_ , \new_[4443]_ , \new_[4444]_ ,
    \new_[4447]_ , \new_[4451]_ , \new_[4452]_ , \new_[4453]_ ,
    \new_[4456]_ , \new_[4459]_ , \new_[4460]_ , \new_[4463]_ ,
    \new_[4467]_ , \new_[4468]_ , \new_[4469]_ , \new_[4472]_ ,
    \new_[4475]_ , \new_[4476]_ , \new_[4479]_ , \new_[4483]_ ,
    \new_[4484]_ , \new_[4485]_ , \new_[4488]_ , \new_[4491]_ ,
    \new_[4492]_ , \new_[4495]_ , \new_[4499]_ , \new_[4500]_ ,
    \new_[4501]_ , \new_[4504]_ , \new_[4507]_ , \new_[4508]_ ,
    \new_[4511]_ , \new_[4515]_ , \new_[4516]_ , \new_[4517]_ ,
    \new_[4520]_ , \new_[4523]_ , \new_[4524]_ , \new_[4527]_ ,
    \new_[4531]_ , \new_[4532]_ , \new_[4533]_ , \new_[4536]_ ,
    \new_[4539]_ , \new_[4540]_ , \new_[4543]_ , \new_[4547]_ ,
    \new_[4548]_ , \new_[4549]_ , \new_[4552]_ , \new_[4555]_ ,
    \new_[4556]_ , \new_[4559]_ , \new_[4563]_ , \new_[4564]_ ,
    \new_[4565]_ , \new_[4568]_ , \new_[4571]_ , \new_[4572]_ ,
    \new_[4575]_ , \new_[4579]_ , \new_[4580]_ , \new_[4581]_ ,
    \new_[4584]_ , \new_[4587]_ , \new_[4588]_ , \new_[4591]_ ,
    \new_[4595]_ , \new_[4596]_ , \new_[4597]_ , \new_[4600]_ ,
    \new_[4603]_ , \new_[4604]_ , \new_[4607]_ , \new_[4611]_ ,
    \new_[4612]_ , \new_[4613]_ , \new_[4616]_ , \new_[4619]_ ,
    \new_[4620]_ , \new_[4623]_ , \new_[4627]_ , \new_[4628]_ ,
    \new_[4629]_ , \new_[4632]_ , \new_[4635]_ , \new_[4636]_ ,
    \new_[4639]_ , \new_[4643]_ , \new_[4644]_ , \new_[4645]_ ,
    \new_[4648]_ , \new_[4651]_ , \new_[4652]_ , \new_[4655]_ ,
    \new_[4659]_ , \new_[4660]_ , \new_[4661]_ , \new_[4664]_ ,
    \new_[4667]_ , \new_[4668]_ , \new_[4671]_ , \new_[4675]_ ,
    \new_[4676]_ , \new_[4677]_ , \new_[4680]_ , \new_[4683]_ ,
    \new_[4684]_ , \new_[4687]_ , \new_[4691]_ , \new_[4692]_ ,
    \new_[4693]_ , \new_[4696]_ , \new_[4699]_ , \new_[4700]_ ,
    \new_[4703]_ , \new_[4707]_ , \new_[4708]_ , \new_[4709]_ ,
    \new_[4712]_ , \new_[4715]_ , \new_[4716]_ , \new_[4719]_ ,
    \new_[4723]_ , \new_[4724]_ , \new_[4725]_ , \new_[4728]_ ,
    \new_[4731]_ , \new_[4732]_ , \new_[4735]_ , \new_[4739]_ ,
    \new_[4740]_ , \new_[4741]_ , \new_[4744]_ , \new_[4747]_ ,
    \new_[4748]_ , \new_[4751]_ , \new_[4755]_ , \new_[4756]_ ,
    \new_[4757]_ , \new_[4760]_ , \new_[4763]_ , \new_[4764]_ ,
    \new_[4767]_ , \new_[4771]_ , \new_[4772]_ , \new_[4773]_ ,
    \new_[4776]_ , \new_[4779]_ , \new_[4780]_ , \new_[4783]_ ,
    \new_[4787]_ , \new_[4788]_ , \new_[4789]_ , \new_[4792]_ ,
    \new_[4795]_ , \new_[4796]_ , \new_[4799]_ , \new_[4803]_ ,
    \new_[4804]_ , \new_[4805]_ , \new_[4808]_ , \new_[4811]_ ,
    \new_[4812]_ , \new_[4815]_ , \new_[4819]_ , \new_[4820]_ ,
    \new_[4821]_ , \new_[4824]_ , \new_[4827]_ , \new_[4828]_ ,
    \new_[4831]_ , \new_[4835]_ , \new_[4836]_ , \new_[4837]_ ,
    \new_[4840]_ , \new_[4843]_ , \new_[4844]_ , \new_[4847]_ ,
    \new_[4851]_ , \new_[4852]_ , \new_[4853]_ , \new_[4856]_ ,
    \new_[4859]_ , \new_[4860]_ , \new_[4863]_ , \new_[4867]_ ,
    \new_[4868]_ , \new_[4869]_ , \new_[4872]_ , \new_[4875]_ ,
    \new_[4876]_ , \new_[4879]_ , \new_[4883]_ , \new_[4884]_ ,
    \new_[4885]_ , \new_[4888]_ , \new_[4891]_ , \new_[4892]_ ,
    \new_[4895]_ , \new_[4899]_ , \new_[4900]_ , \new_[4901]_ ,
    \new_[4904]_ , \new_[4907]_ , \new_[4908]_ , \new_[4911]_ ,
    \new_[4915]_ , \new_[4916]_ , \new_[4917]_ , \new_[4920]_ ,
    \new_[4923]_ , \new_[4924]_ , \new_[4927]_ , \new_[4931]_ ,
    \new_[4932]_ , \new_[4933]_ , \new_[4936]_ , \new_[4939]_ ,
    \new_[4940]_ , \new_[4943]_ , \new_[4947]_ , \new_[4948]_ ,
    \new_[4949]_ , \new_[4952]_ , \new_[4955]_ , \new_[4956]_ ,
    \new_[4959]_ , \new_[4963]_ , \new_[4964]_ , \new_[4965]_ ,
    \new_[4968]_ , \new_[4971]_ , \new_[4972]_ , \new_[4975]_ ,
    \new_[4979]_ , \new_[4980]_ , \new_[4981]_ , \new_[4984]_ ,
    \new_[4987]_ , \new_[4988]_ , \new_[4991]_ , \new_[4995]_ ,
    \new_[4996]_ , \new_[4997]_ , \new_[5000]_ , \new_[5003]_ ,
    \new_[5004]_ , \new_[5007]_ , \new_[5011]_ , \new_[5012]_ ,
    \new_[5013]_ , \new_[5016]_ , \new_[5019]_ , \new_[5020]_ ,
    \new_[5023]_ , \new_[5027]_ , \new_[5028]_ , \new_[5029]_ ,
    \new_[5032]_ , \new_[5035]_ , \new_[5036]_ , \new_[5039]_ ,
    \new_[5043]_ , \new_[5044]_ , \new_[5045]_ , \new_[5048]_ ,
    \new_[5051]_ , \new_[5052]_ , \new_[5055]_ , \new_[5059]_ ,
    \new_[5060]_ , \new_[5061]_ , \new_[5064]_ , \new_[5067]_ ,
    \new_[5068]_ , \new_[5071]_ , \new_[5075]_ , \new_[5076]_ ,
    \new_[5077]_ , \new_[5080]_ , \new_[5083]_ , \new_[5084]_ ,
    \new_[5087]_ , \new_[5091]_ , \new_[5092]_ , \new_[5093]_ ,
    \new_[5096]_ , \new_[5099]_ , \new_[5100]_ , \new_[5103]_ ,
    \new_[5107]_ , \new_[5108]_ , \new_[5109]_ , \new_[5112]_ ,
    \new_[5115]_ , \new_[5116]_ , \new_[5119]_ , \new_[5123]_ ,
    \new_[5124]_ , \new_[5125]_ , \new_[5128]_ , \new_[5131]_ ,
    \new_[5132]_ , \new_[5135]_ , \new_[5139]_ , \new_[5140]_ ,
    \new_[5141]_ , \new_[5144]_ , \new_[5147]_ , \new_[5148]_ ,
    \new_[5151]_ , \new_[5155]_ , \new_[5156]_ , \new_[5157]_ ,
    \new_[5160]_ , \new_[5163]_ , \new_[5164]_ , \new_[5167]_ ,
    \new_[5171]_ , \new_[5172]_ , \new_[5173]_ , \new_[5176]_ ,
    \new_[5179]_ , \new_[5180]_ , \new_[5183]_ , \new_[5187]_ ,
    \new_[5188]_ , \new_[5189]_ , \new_[5192]_ , \new_[5195]_ ,
    \new_[5196]_ , \new_[5199]_ , \new_[5203]_ , \new_[5204]_ ,
    \new_[5205]_ , \new_[5208]_ , \new_[5211]_ , \new_[5212]_ ,
    \new_[5215]_ , \new_[5219]_ , \new_[5220]_ , \new_[5221]_ ,
    \new_[5224]_ , \new_[5227]_ , \new_[5228]_ , \new_[5231]_ ,
    \new_[5235]_ , \new_[5236]_ , \new_[5237]_ , \new_[5240]_ ,
    \new_[5243]_ , \new_[5244]_ , \new_[5247]_ , \new_[5251]_ ,
    \new_[5252]_ , \new_[5253]_ , \new_[5256]_ , \new_[5259]_ ,
    \new_[5260]_ , \new_[5263]_ , \new_[5267]_ , \new_[5268]_ ,
    \new_[5269]_ , \new_[5272]_ , \new_[5275]_ , \new_[5276]_ ,
    \new_[5279]_ , \new_[5283]_ , \new_[5284]_ , \new_[5285]_ ,
    \new_[5288]_ , \new_[5291]_ , \new_[5292]_ , \new_[5295]_ ,
    \new_[5299]_ , \new_[5300]_ , \new_[5301]_ , \new_[5304]_ ,
    \new_[5307]_ , \new_[5308]_ , \new_[5311]_ , \new_[5315]_ ,
    \new_[5316]_ , \new_[5317]_ , \new_[5320]_ , \new_[5323]_ ,
    \new_[5324]_ , \new_[5327]_ , \new_[5331]_ , \new_[5332]_ ,
    \new_[5333]_ , \new_[5336]_ , \new_[5339]_ , \new_[5340]_ ,
    \new_[5343]_ , \new_[5347]_ , \new_[5348]_ , \new_[5349]_ ,
    \new_[5352]_ , \new_[5355]_ , \new_[5356]_ , \new_[5359]_ ,
    \new_[5363]_ , \new_[5364]_ , \new_[5365]_ , \new_[5368]_ ,
    \new_[5371]_ , \new_[5372]_ , \new_[5375]_ , \new_[5379]_ ,
    \new_[5380]_ , \new_[5381]_ , \new_[5384]_ , \new_[5387]_ ,
    \new_[5388]_ , \new_[5391]_ , \new_[5395]_ , \new_[5396]_ ,
    \new_[5397]_ , \new_[5400]_ , \new_[5403]_ , \new_[5404]_ ,
    \new_[5407]_ , \new_[5411]_ , \new_[5412]_ , \new_[5413]_ ,
    \new_[5416]_ , \new_[5419]_ , \new_[5420]_ , \new_[5423]_ ,
    \new_[5427]_ , \new_[5428]_ , \new_[5429]_ , \new_[5432]_ ,
    \new_[5435]_ , \new_[5436]_ , \new_[5439]_ , \new_[5443]_ ,
    \new_[5444]_ , \new_[5445]_ , \new_[5448]_ , \new_[5451]_ ,
    \new_[5452]_ , \new_[5455]_ , \new_[5459]_ , \new_[5460]_ ,
    \new_[5461]_ , \new_[5464]_ , \new_[5467]_ , \new_[5468]_ ,
    \new_[5471]_ , \new_[5475]_ , \new_[5476]_ , \new_[5477]_ ,
    \new_[5480]_ , \new_[5483]_ , \new_[5484]_ , \new_[5487]_ ,
    \new_[5491]_ , \new_[5492]_ , \new_[5493]_ , \new_[5496]_ ,
    \new_[5499]_ , \new_[5500]_ , \new_[5503]_ , \new_[5507]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5512]_ , \new_[5515]_ ,
    \new_[5516]_ , \new_[5519]_ , \new_[5523]_ , \new_[5524]_ ,
    \new_[5525]_ , \new_[5528]_ , \new_[5531]_ , \new_[5532]_ ,
    \new_[5535]_ , \new_[5539]_ , \new_[5540]_ , \new_[5541]_ ,
    \new_[5544]_ , \new_[5547]_ , \new_[5548]_ , \new_[5551]_ ,
    \new_[5555]_ , \new_[5556]_ , \new_[5557]_ , \new_[5560]_ ,
    \new_[5563]_ , \new_[5564]_ , \new_[5567]_ , \new_[5571]_ ,
    \new_[5572]_ , \new_[5573]_ , \new_[5576]_ , \new_[5579]_ ,
    \new_[5580]_ , \new_[5583]_ , \new_[5587]_ , \new_[5588]_ ,
    \new_[5589]_ , \new_[5592]_ , \new_[5595]_ , \new_[5596]_ ,
    \new_[5599]_ , \new_[5603]_ , \new_[5604]_ , \new_[5605]_ ,
    \new_[5608]_ , \new_[5611]_ , \new_[5612]_ , \new_[5615]_ ,
    \new_[5619]_ , \new_[5620]_ , \new_[5621]_ , \new_[5624]_ ,
    \new_[5627]_ , \new_[5628]_ , \new_[5631]_ , \new_[5635]_ ,
    \new_[5636]_ , \new_[5637]_ , \new_[5640]_ , \new_[5643]_ ,
    \new_[5644]_ , \new_[5647]_ , \new_[5651]_ , \new_[5652]_ ,
    \new_[5653]_ , \new_[5656]_ , \new_[5659]_ , \new_[5660]_ ,
    \new_[5663]_ , \new_[5667]_ , \new_[5668]_ , \new_[5669]_ ,
    \new_[5672]_ , \new_[5675]_ , \new_[5676]_ , \new_[5679]_ ,
    \new_[5683]_ , \new_[5684]_ , \new_[5685]_ , \new_[5688]_ ,
    \new_[5691]_ , \new_[5692]_ , \new_[5695]_ , \new_[5699]_ ,
    \new_[5700]_ , \new_[5701]_ , \new_[5704]_ , \new_[5707]_ ,
    \new_[5708]_ , \new_[5711]_ , \new_[5715]_ , \new_[5716]_ ,
    \new_[5717]_ , \new_[5720]_ , \new_[5723]_ , \new_[5724]_ ,
    \new_[5727]_ , \new_[5731]_ , \new_[5732]_ , \new_[5733]_ ,
    \new_[5736]_ , \new_[5739]_ , \new_[5740]_ , \new_[5743]_ ,
    \new_[5747]_ , \new_[5748]_ , \new_[5749]_ , \new_[5752]_ ,
    \new_[5755]_ , \new_[5756]_ , \new_[5759]_ , \new_[5763]_ ,
    \new_[5764]_ , \new_[5765]_ , \new_[5768]_ , \new_[5771]_ ,
    \new_[5772]_ , \new_[5775]_ , \new_[5779]_ , \new_[5780]_ ,
    \new_[5781]_ , \new_[5784]_ , \new_[5787]_ , \new_[5788]_ ,
    \new_[5791]_ , \new_[5795]_ , \new_[5796]_ , \new_[5797]_ ,
    \new_[5800]_ , \new_[5803]_ , \new_[5804]_ , \new_[5807]_ ,
    \new_[5811]_ , \new_[5812]_ , \new_[5813]_ , \new_[5816]_ ,
    \new_[5819]_ , \new_[5820]_ , \new_[5823]_ , \new_[5827]_ ,
    \new_[5828]_ , \new_[5829]_ , \new_[5832]_ , \new_[5835]_ ,
    \new_[5836]_ , \new_[5839]_ , \new_[5843]_ , \new_[5844]_ ,
    \new_[5845]_ , \new_[5848]_ , \new_[5851]_ , \new_[5852]_ ,
    \new_[5855]_ , \new_[5859]_ , \new_[5860]_ , \new_[5861]_ ,
    \new_[5864]_ , \new_[5867]_ , \new_[5868]_ , \new_[5871]_ ,
    \new_[5875]_ , \new_[5876]_ , \new_[5877]_ , \new_[5880]_ ,
    \new_[5883]_ , \new_[5884]_ , \new_[5887]_ , \new_[5891]_ ,
    \new_[5892]_ , \new_[5893]_ , \new_[5896]_ , \new_[5899]_ ,
    \new_[5900]_ , \new_[5903]_ , \new_[5907]_ , \new_[5908]_ ,
    \new_[5909]_ , \new_[5912]_ , \new_[5915]_ , \new_[5916]_ ,
    \new_[5919]_ , \new_[5923]_ , \new_[5924]_ , \new_[5925]_ ,
    \new_[5928]_ , \new_[5931]_ , \new_[5932]_ , \new_[5935]_ ,
    \new_[5939]_ , \new_[5940]_ , \new_[5941]_ , \new_[5944]_ ,
    \new_[5947]_ , \new_[5948]_ , \new_[5951]_ , \new_[5955]_ ,
    \new_[5956]_ , \new_[5957]_ , \new_[5960]_ , \new_[5963]_ ,
    \new_[5964]_ , \new_[5967]_ , \new_[5971]_ , \new_[5972]_ ,
    \new_[5973]_ , \new_[5976]_ , \new_[5979]_ , \new_[5980]_ ,
    \new_[5983]_ , \new_[5987]_ , \new_[5988]_ , \new_[5989]_ ,
    \new_[5992]_ , \new_[5995]_ , \new_[5996]_ , \new_[5999]_ ,
    \new_[6003]_ , \new_[6004]_ , \new_[6005]_ , \new_[6008]_ ,
    \new_[6011]_ , \new_[6012]_ , \new_[6015]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6021]_ , \new_[6024]_ , \new_[6027]_ ,
    \new_[6028]_ , \new_[6031]_ , \new_[6035]_ , \new_[6036]_ ,
    \new_[6037]_ , \new_[6040]_ , \new_[6043]_ , \new_[6044]_ ,
    \new_[6047]_ , \new_[6051]_ , \new_[6052]_ , \new_[6053]_ ,
    \new_[6056]_ , \new_[6059]_ , \new_[6060]_ , \new_[6063]_ ,
    \new_[6067]_ , \new_[6068]_ , \new_[6069]_ , \new_[6072]_ ,
    \new_[6075]_ , \new_[6076]_ , \new_[6079]_ , \new_[6083]_ ,
    \new_[6084]_ , \new_[6085]_ , \new_[6088]_ , \new_[6091]_ ,
    \new_[6092]_ , \new_[6095]_ , \new_[6099]_ , \new_[6100]_ ,
    \new_[6101]_ , \new_[6104]_ , \new_[6107]_ , \new_[6108]_ ,
    \new_[6111]_ , \new_[6115]_ , \new_[6116]_ , \new_[6117]_ ,
    \new_[6120]_ , \new_[6123]_ , \new_[6124]_ , \new_[6127]_ ,
    \new_[6131]_ , \new_[6132]_ , \new_[6133]_ , \new_[6136]_ ,
    \new_[6139]_ , \new_[6140]_ , \new_[6143]_ , \new_[6147]_ ,
    \new_[6148]_ , \new_[6149]_ , \new_[6152]_ , \new_[6155]_ ,
    \new_[6156]_ , \new_[6159]_ , \new_[6163]_ , \new_[6164]_ ,
    \new_[6165]_ , \new_[6168]_ , \new_[6171]_ , \new_[6172]_ ,
    \new_[6175]_ , \new_[6179]_ , \new_[6180]_ , \new_[6181]_ ,
    \new_[6184]_ , \new_[6187]_ , \new_[6188]_ , \new_[6191]_ ,
    \new_[6195]_ , \new_[6196]_ , \new_[6197]_ , \new_[6200]_ ,
    \new_[6203]_ , \new_[6204]_ , \new_[6207]_ , \new_[6211]_ ,
    \new_[6212]_ , \new_[6213]_ , \new_[6216]_ , \new_[6219]_ ,
    \new_[6220]_ , \new_[6223]_ , \new_[6227]_ , \new_[6228]_ ,
    \new_[6229]_ , \new_[6232]_ , \new_[6235]_ , \new_[6236]_ ,
    \new_[6239]_ , \new_[6243]_ , \new_[6244]_ , \new_[6245]_ ,
    \new_[6248]_ , \new_[6251]_ , \new_[6252]_ , \new_[6255]_ ,
    \new_[6259]_ , \new_[6260]_ , \new_[6261]_ , \new_[6264]_ ,
    \new_[6267]_ , \new_[6268]_ , \new_[6271]_ , \new_[6275]_ ,
    \new_[6276]_ , \new_[6277]_ , \new_[6280]_ , \new_[6283]_ ,
    \new_[6284]_ , \new_[6287]_ , \new_[6291]_ , \new_[6292]_ ,
    \new_[6293]_ , \new_[6296]_ , \new_[6299]_ , \new_[6300]_ ,
    \new_[6303]_ , \new_[6307]_ , \new_[6308]_ , \new_[6309]_ ,
    \new_[6312]_ , \new_[6315]_ , \new_[6316]_ , \new_[6319]_ ,
    \new_[6323]_ , \new_[6324]_ , \new_[6325]_ , \new_[6328]_ ,
    \new_[6331]_ , \new_[6332]_ , \new_[6335]_ , \new_[6339]_ ,
    \new_[6340]_ , \new_[6341]_ , \new_[6344]_ , \new_[6347]_ ,
    \new_[6348]_ , \new_[6351]_ , \new_[6355]_ , \new_[6356]_ ,
    \new_[6357]_ , \new_[6360]_ , \new_[6363]_ , \new_[6364]_ ,
    \new_[6367]_ , \new_[6371]_ , \new_[6372]_ , \new_[6373]_ ,
    \new_[6376]_ , \new_[6379]_ , \new_[6380]_ , \new_[6383]_ ,
    \new_[6387]_ , \new_[6388]_ , \new_[6389]_ , \new_[6392]_ ,
    \new_[6395]_ , \new_[6396]_ , \new_[6399]_ , \new_[6403]_ ,
    \new_[6404]_ , \new_[6405]_ , \new_[6408]_ , \new_[6411]_ ,
    \new_[6412]_ , \new_[6415]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6421]_ , \new_[6424]_ , \new_[6427]_ , \new_[6428]_ ,
    \new_[6431]_ , \new_[6435]_ , \new_[6436]_ , \new_[6437]_ ,
    \new_[6440]_ , \new_[6443]_ , \new_[6444]_ , \new_[6447]_ ,
    \new_[6451]_ , \new_[6452]_ , \new_[6453]_ , \new_[6456]_ ,
    \new_[6459]_ , \new_[6460]_ , \new_[6463]_ , \new_[6467]_ ,
    \new_[6468]_ , \new_[6469]_ , \new_[6472]_ , \new_[6475]_ ,
    \new_[6476]_ , \new_[6479]_ , \new_[6483]_ , \new_[6484]_ ,
    \new_[6485]_ , \new_[6488]_ , \new_[6491]_ , \new_[6492]_ ,
    \new_[6495]_ , \new_[6499]_ , \new_[6500]_ , \new_[6501]_ ,
    \new_[6504]_ , \new_[6507]_ , \new_[6508]_ , \new_[6511]_ ,
    \new_[6515]_ , \new_[6516]_ , \new_[6517]_ , \new_[6520]_ ,
    \new_[6523]_ , \new_[6524]_ , \new_[6527]_ , \new_[6531]_ ,
    \new_[6532]_ , \new_[6533]_ , \new_[6536]_ , \new_[6539]_ ,
    \new_[6540]_ , \new_[6543]_ , \new_[6547]_ , \new_[6548]_ ,
    \new_[6549]_ , \new_[6552]_ , \new_[6555]_ , \new_[6556]_ ,
    \new_[6559]_ , \new_[6563]_ , \new_[6564]_ , \new_[6565]_ ,
    \new_[6568]_ , \new_[6571]_ , \new_[6572]_ , \new_[6575]_ ,
    \new_[6579]_ , \new_[6580]_ , \new_[6581]_ , \new_[6584]_ ,
    \new_[6588]_ , \new_[6589]_ , \new_[6590]_ , \new_[6593]_ ,
    \new_[6597]_ , \new_[6598]_ , \new_[6599]_ , \new_[6602]_ ,
    \new_[6606]_ , \new_[6607]_ , \new_[6608]_ , \new_[6611]_ ,
    \new_[6615]_ , \new_[6616]_ , \new_[6617]_ , \new_[6620]_ ,
    \new_[6624]_ , \new_[6625]_ , \new_[6626]_ , \new_[6629]_ ,
    \new_[6633]_ , \new_[6634]_ , \new_[6635]_ , \new_[6638]_ ,
    \new_[6642]_ , \new_[6643]_ , \new_[6644]_ , \new_[6647]_ ,
    \new_[6651]_ , \new_[6652]_ , \new_[6653]_ , \new_[6656]_ ,
    \new_[6660]_ , \new_[6661]_ , \new_[6662]_ , \new_[6665]_ ,
    \new_[6669]_ , \new_[6670]_ , \new_[6671]_ , \new_[6674]_ ,
    \new_[6678]_ , \new_[6679]_ , \new_[6680]_ , \new_[6683]_ ,
    \new_[6687]_ , \new_[6688]_ , \new_[6689]_ , \new_[6692]_ ,
    \new_[6696]_ , \new_[6697]_ , \new_[6698]_ , \new_[6701]_ ,
    \new_[6705]_ , \new_[6706]_ , \new_[6707]_ , \new_[6710]_ ,
    \new_[6714]_ , \new_[6715]_ , \new_[6716]_ , \new_[6719]_ ,
    \new_[6723]_ , \new_[6724]_ , \new_[6725]_ , \new_[6728]_ ,
    \new_[6732]_ , \new_[6733]_ , \new_[6734]_ , \new_[6737]_ ,
    \new_[6741]_ , \new_[6742]_ , \new_[6743]_ , \new_[6746]_ ,
    \new_[6750]_ , \new_[6751]_ , \new_[6752]_ , \new_[6755]_ ,
    \new_[6759]_ , \new_[6760]_ , \new_[6761]_ , \new_[6764]_ ,
    \new_[6768]_ , \new_[6769]_ , \new_[6770]_ , \new_[6773]_ ,
    \new_[6777]_ , \new_[6778]_ , \new_[6779]_ , \new_[6782]_ ,
    \new_[6786]_ , \new_[6787]_ , \new_[6788]_ , \new_[6791]_ ,
    \new_[6795]_ , \new_[6796]_ , \new_[6797]_ , \new_[6800]_ ,
    \new_[6804]_ , \new_[6805]_ , \new_[6806]_ , \new_[6809]_ ,
    \new_[6813]_ , \new_[6814]_ , \new_[6815]_ , \new_[6818]_ ,
    \new_[6822]_ , \new_[6823]_ , \new_[6824]_ , \new_[6827]_ ,
    \new_[6831]_ , \new_[6832]_ , \new_[6833]_ , \new_[6836]_ ,
    \new_[6840]_ , \new_[6841]_ , \new_[6842]_ , \new_[6845]_ ,
    \new_[6849]_ , \new_[6850]_ , \new_[6851]_ , \new_[6854]_ ,
    \new_[6858]_ , \new_[6859]_ , \new_[6860]_ , \new_[6863]_ ,
    \new_[6867]_ , \new_[6868]_ , \new_[6869]_ , \new_[6872]_ ,
    \new_[6876]_ , \new_[6877]_ , \new_[6878]_ , \new_[6881]_ ,
    \new_[6885]_ , \new_[6886]_ , \new_[6887]_ , \new_[6890]_ ,
    \new_[6894]_ , \new_[6895]_ , \new_[6896]_ , \new_[6899]_ ,
    \new_[6903]_ , \new_[6904]_ , \new_[6905]_ , \new_[6908]_ ,
    \new_[6912]_ , \new_[6913]_ , \new_[6914]_ , \new_[6917]_ ,
    \new_[6921]_ , \new_[6922]_ , \new_[6923]_ , \new_[6926]_ ,
    \new_[6930]_ , \new_[6931]_ , \new_[6932]_ , \new_[6935]_ ,
    \new_[6939]_ , \new_[6940]_ , \new_[6941]_ , \new_[6944]_ ,
    \new_[6948]_ , \new_[6949]_ , \new_[6950]_ , \new_[6953]_ ,
    \new_[6957]_ , \new_[6958]_ , \new_[6959]_ , \new_[6962]_ ,
    \new_[6966]_ , \new_[6967]_ , \new_[6968]_ , \new_[6971]_ ,
    \new_[6975]_ , \new_[6976]_ , \new_[6977]_ , \new_[6980]_ ,
    \new_[6984]_ , \new_[6985]_ , \new_[6986]_ , \new_[6989]_ ,
    \new_[6993]_ , \new_[6994]_ , \new_[6995]_ , \new_[6998]_ ,
    \new_[7002]_ , \new_[7003]_ , \new_[7004]_ , \new_[7007]_ ,
    \new_[7011]_ , \new_[7012]_ , \new_[7013]_ , \new_[7016]_ ,
    \new_[7020]_ , \new_[7021]_ , \new_[7022]_ , \new_[7025]_ ,
    \new_[7029]_ , \new_[7030]_ , \new_[7031]_ , \new_[7034]_ ,
    \new_[7038]_ , \new_[7039]_ , \new_[7040]_ , \new_[7043]_ ,
    \new_[7047]_ , \new_[7048]_ , \new_[7049]_ , \new_[7052]_ ,
    \new_[7056]_ , \new_[7057]_ , \new_[7058]_ , \new_[7061]_ ,
    \new_[7065]_ , \new_[7066]_ , \new_[7067]_ , \new_[7070]_ ,
    \new_[7074]_ , \new_[7075]_ , \new_[7076]_ , \new_[7079]_ ,
    \new_[7083]_ , \new_[7084]_ , \new_[7085]_ , \new_[7088]_ ,
    \new_[7092]_ , \new_[7093]_ , \new_[7094]_ , \new_[7097]_ ,
    \new_[7101]_ , \new_[7102]_ , \new_[7103]_ , \new_[7106]_ ,
    \new_[7110]_ , \new_[7111]_ , \new_[7112]_ , \new_[7115]_ ,
    \new_[7119]_ , \new_[7120]_ , \new_[7121]_ , \new_[7124]_ ,
    \new_[7128]_ , \new_[7129]_ , \new_[7130]_ , \new_[7133]_ ,
    \new_[7137]_ , \new_[7138]_ , \new_[7139]_ , \new_[7142]_ ,
    \new_[7146]_ , \new_[7147]_ , \new_[7148]_ , \new_[7151]_ ,
    \new_[7155]_ , \new_[7156]_ , \new_[7157]_ , \new_[7160]_ ,
    \new_[7164]_ , \new_[7165]_ , \new_[7166]_ , \new_[7169]_ ,
    \new_[7173]_ , \new_[7174]_ , \new_[7175]_ , \new_[7178]_ ,
    \new_[7182]_ , \new_[7183]_ , \new_[7184]_ , \new_[7187]_ ,
    \new_[7191]_ , \new_[7192]_ , \new_[7193]_ , \new_[7196]_ ,
    \new_[7200]_ , \new_[7201]_ , \new_[7202]_ , \new_[7205]_ ,
    \new_[7209]_ , \new_[7210]_ , \new_[7211]_ , \new_[7214]_ ,
    \new_[7218]_ , \new_[7219]_ , \new_[7220]_ , \new_[7223]_ ,
    \new_[7227]_ , \new_[7228]_ , \new_[7229]_ , \new_[7232]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7241]_ ,
    \new_[7245]_ , \new_[7246]_ , \new_[7247]_ , \new_[7250]_ ,
    \new_[7254]_ , \new_[7255]_ , \new_[7256]_ , \new_[7259]_ ,
    \new_[7263]_ , \new_[7264]_ , \new_[7265]_ , \new_[7268]_ ,
    \new_[7272]_ , \new_[7273]_ , \new_[7274]_ , \new_[7277]_ ,
    \new_[7281]_ , \new_[7282]_ , \new_[7283]_ , \new_[7286]_ ,
    \new_[7290]_ , \new_[7291]_ , \new_[7292]_ , \new_[7295]_ ,
    \new_[7299]_ , \new_[7300]_ , \new_[7301]_ , \new_[7304]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7310]_ , \new_[7313]_ ,
    \new_[7317]_ , \new_[7318]_ , \new_[7319]_ , \new_[7322]_ ,
    \new_[7326]_ , \new_[7327]_ , \new_[7328]_ , \new_[7331]_ ,
    \new_[7335]_ , \new_[7336]_ , \new_[7337]_ , \new_[7340]_ ,
    \new_[7344]_ , \new_[7345]_ , \new_[7346]_ , \new_[7349]_ ,
    \new_[7353]_ , \new_[7354]_ , \new_[7355]_ , \new_[7358]_ ,
    \new_[7362]_ , \new_[7363]_ , \new_[7364]_ , \new_[7367]_ ,
    \new_[7371]_ , \new_[7372]_ , \new_[7373]_ , \new_[7376]_ ,
    \new_[7380]_ , \new_[7381]_ , \new_[7382]_ , \new_[7385]_ ,
    \new_[7389]_ , \new_[7390]_ , \new_[7391]_ , \new_[7394]_ ,
    \new_[7398]_ , \new_[7399]_ , \new_[7400]_ , \new_[7403]_ ,
    \new_[7407]_ , \new_[7408]_ , \new_[7409]_ , \new_[7412]_ ,
    \new_[7416]_ , \new_[7417]_ , \new_[7418]_ , \new_[7421]_ ,
    \new_[7425]_ , \new_[7426]_ , \new_[7427]_ , \new_[7430]_ ,
    \new_[7434]_ , \new_[7435]_ , \new_[7436]_ , \new_[7439]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7445]_ , \new_[7448]_ ,
    \new_[7452]_ , \new_[7453]_ , \new_[7454]_ , \new_[7457]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7466]_ ,
    \new_[7470]_ , \new_[7471]_ , \new_[7472]_ , \new_[7475]_ ,
    \new_[7479]_ , \new_[7480]_ , \new_[7481]_ , \new_[7484]_ ,
    \new_[7488]_ , \new_[7489]_ , \new_[7490]_ , \new_[7493]_ ,
    \new_[7497]_ , \new_[7498]_ , \new_[7499]_ , \new_[7502]_ ,
    \new_[7506]_ , \new_[7507]_ , \new_[7508]_ , \new_[7511]_ ,
    \new_[7515]_ , \new_[7516]_ , \new_[7517]_ , \new_[7520]_ ,
    \new_[7524]_ , \new_[7525]_ , \new_[7526]_ , \new_[7529]_ ,
    \new_[7533]_ , \new_[7534]_ , \new_[7535]_ , \new_[7538]_ ,
    \new_[7542]_ , \new_[7543]_ , \new_[7544]_ , \new_[7547]_ ,
    \new_[7551]_ , \new_[7552]_ , \new_[7553]_ , \new_[7556]_ ,
    \new_[7560]_ , \new_[7561]_ , \new_[7562]_ , \new_[7565]_ ,
    \new_[7569]_ , \new_[7570]_ , \new_[7571]_ , \new_[7574]_ ,
    \new_[7578]_ , \new_[7579]_ , \new_[7580]_ , \new_[7583]_ ,
    \new_[7587]_ , \new_[7588]_ , \new_[7589]_ , \new_[7592]_ ,
    \new_[7596]_ , \new_[7597]_ , \new_[7598]_ , \new_[7601]_ ,
    \new_[7605]_ , \new_[7606]_ , \new_[7607]_ , \new_[7610]_ ,
    \new_[7614]_ , \new_[7615]_ , \new_[7616]_ , \new_[7619]_ ,
    \new_[7623]_ , \new_[7624]_ , \new_[7625]_ , \new_[7628]_ ,
    \new_[7632]_ , \new_[7633]_ , \new_[7634]_ , \new_[7637]_ ,
    \new_[7641]_ , \new_[7642]_ , \new_[7643]_ , \new_[7646]_ ,
    \new_[7650]_ , \new_[7651]_ , \new_[7652]_ , \new_[7655]_ ,
    \new_[7659]_ , \new_[7660]_ , \new_[7661]_ , \new_[7664]_ ,
    \new_[7668]_ , \new_[7669]_ , \new_[7670]_ , \new_[7673]_ ,
    \new_[7677]_ , \new_[7678]_ , \new_[7679]_ , \new_[7682]_ ,
    \new_[7686]_ , \new_[7687]_ , \new_[7688]_ , \new_[7691]_ ,
    \new_[7695]_ , \new_[7696]_ , \new_[7697]_ , \new_[7700]_ ,
    \new_[7704]_ , \new_[7705]_ , \new_[7706]_ , \new_[7709]_ ,
    \new_[7713]_ , \new_[7714]_ , \new_[7715]_ , \new_[7718]_ ,
    \new_[7722]_ , \new_[7723]_ , \new_[7724]_ , \new_[7727]_ ,
    \new_[7731]_ , \new_[7732]_ , \new_[7733]_ , \new_[7736]_ ,
    \new_[7740]_ , \new_[7741]_ , \new_[7742]_ , \new_[7745]_ ,
    \new_[7749]_ , \new_[7750]_ , \new_[7751]_ , \new_[7754]_ ,
    \new_[7758]_ , \new_[7759]_ , \new_[7760]_ , \new_[7763]_ ,
    \new_[7767]_ , \new_[7768]_ , \new_[7769]_ , \new_[7772]_ ,
    \new_[7776]_ , \new_[7777]_ , \new_[7778]_ , \new_[7781]_ ,
    \new_[7785]_ , \new_[7786]_ , \new_[7787]_ , \new_[7790]_ ,
    \new_[7794]_ , \new_[7795]_ , \new_[7796]_ , \new_[7799]_ ,
    \new_[7803]_ , \new_[7804]_ , \new_[7805]_ , \new_[7808]_ ,
    \new_[7812]_ , \new_[7813]_ , \new_[7814]_ , \new_[7817]_ ,
    \new_[7821]_ , \new_[7822]_ , \new_[7823]_ , \new_[7826]_ ,
    \new_[7830]_ , \new_[7831]_ , \new_[7832]_ , \new_[7835]_ ,
    \new_[7839]_ , \new_[7840]_ , \new_[7841]_ , \new_[7844]_ ,
    \new_[7848]_ , \new_[7849]_ , \new_[7850]_ , \new_[7853]_ ,
    \new_[7857]_ , \new_[7858]_ , \new_[7859]_ , \new_[7862]_ ,
    \new_[7866]_ , \new_[7867]_ , \new_[7868]_ , \new_[7871]_ ,
    \new_[7875]_ , \new_[7876]_ , \new_[7877]_ , \new_[7880]_ ,
    \new_[7884]_ , \new_[7885]_ , \new_[7886]_ , \new_[7889]_ ,
    \new_[7893]_ , \new_[7894]_ , \new_[7895]_ , \new_[7898]_ ,
    \new_[7902]_ , \new_[7903]_ , \new_[7904]_ , \new_[7907]_ ,
    \new_[7911]_ , \new_[7912]_ , \new_[7913]_ , \new_[7916]_ ,
    \new_[7920]_ , \new_[7921]_ , \new_[7922]_ , \new_[7925]_ ,
    \new_[7929]_ , \new_[7930]_ , \new_[7931]_ , \new_[7934]_ ,
    \new_[7938]_ , \new_[7939]_ , \new_[7940]_ , \new_[7943]_ ,
    \new_[7947]_ , \new_[7948]_ , \new_[7949]_ , \new_[7952]_ ,
    \new_[7956]_ , \new_[7957]_ , \new_[7958]_ , \new_[7961]_ ,
    \new_[7965]_ , \new_[7966]_ , \new_[7967]_ , \new_[7970]_ ,
    \new_[7974]_ , \new_[7975]_ , \new_[7976]_ , \new_[7979]_ ,
    \new_[7983]_ , \new_[7984]_ , \new_[7985]_ , \new_[7988]_ ,
    \new_[7992]_ , \new_[7993]_ , \new_[7994]_ , \new_[7997]_ ,
    \new_[8001]_ , \new_[8002]_ , \new_[8003]_ , \new_[8006]_ ,
    \new_[8010]_ , \new_[8011]_ , \new_[8012]_ , \new_[8015]_ ,
    \new_[8019]_ , \new_[8020]_ , \new_[8021]_ , \new_[8024]_ ,
    \new_[8028]_ , \new_[8029]_ , \new_[8030]_ , \new_[8033]_ ,
    \new_[8037]_ , \new_[8038]_ , \new_[8039]_ , \new_[8042]_ ,
    \new_[8046]_ , \new_[8047]_ , \new_[8048]_ , \new_[8051]_ ,
    \new_[8055]_ , \new_[8056]_ , \new_[8057]_ , \new_[8060]_ ,
    \new_[8064]_ , \new_[8065]_ , \new_[8066]_ , \new_[8069]_ ,
    \new_[8073]_ , \new_[8074]_ , \new_[8075]_ , \new_[8078]_ ,
    \new_[8082]_ , \new_[8083]_ , \new_[8084]_ , \new_[8087]_ ,
    \new_[8091]_ , \new_[8092]_ , \new_[8093]_ , \new_[8096]_ ,
    \new_[8100]_ , \new_[8101]_ , \new_[8102]_ , \new_[8105]_ ,
    \new_[8109]_ , \new_[8110]_ , \new_[8111]_ , \new_[8114]_ ,
    \new_[8118]_ , \new_[8119]_ , \new_[8120]_ , \new_[8123]_ ,
    \new_[8127]_ , \new_[8128]_ , \new_[8129]_ , \new_[8132]_ ,
    \new_[8136]_ , \new_[8137]_ , \new_[8138]_ , \new_[8141]_ ,
    \new_[8145]_ , \new_[8146]_ , \new_[8147]_ , \new_[8150]_ ,
    \new_[8154]_ , \new_[8155]_ , \new_[8156]_ , \new_[8159]_ ,
    \new_[8163]_ , \new_[8164]_ , \new_[8165]_ , \new_[8168]_ ,
    \new_[8172]_ , \new_[8173]_ , \new_[8174]_ , \new_[8177]_ ,
    \new_[8181]_ , \new_[8182]_ , \new_[8183]_ , \new_[8186]_ ,
    \new_[8190]_ , \new_[8191]_ , \new_[8192]_ , \new_[8195]_ ,
    \new_[8199]_ , \new_[8200]_ , \new_[8201]_ , \new_[8204]_ ,
    \new_[8208]_ , \new_[8209]_ , \new_[8210]_ , \new_[8213]_ ,
    \new_[8217]_ , \new_[8218]_ , \new_[8219]_ , \new_[8222]_ ,
    \new_[8226]_ , \new_[8227]_ , \new_[8228]_ , \new_[8231]_ ,
    \new_[8235]_ , \new_[8236]_ , \new_[8237]_ , \new_[8240]_ ,
    \new_[8244]_ , \new_[8245]_ , \new_[8246]_ , \new_[8249]_ ,
    \new_[8253]_ , \new_[8254]_ , \new_[8255]_ , \new_[8258]_ ,
    \new_[8262]_ , \new_[8263]_ , \new_[8264]_ , \new_[8267]_ ,
    \new_[8271]_ , \new_[8272]_ , \new_[8273]_ , \new_[8276]_ ,
    \new_[8280]_ , \new_[8281]_ , \new_[8282]_ , \new_[8285]_ ,
    \new_[8289]_ , \new_[8290]_ , \new_[8291]_ , \new_[8294]_ ,
    \new_[8298]_ , \new_[8299]_ , \new_[8300]_ , \new_[8303]_ ,
    \new_[8307]_ , \new_[8308]_ , \new_[8309]_ , \new_[8312]_ ,
    \new_[8316]_ , \new_[8317]_ , \new_[8318]_ , \new_[8321]_ ,
    \new_[8325]_ , \new_[8326]_ , \new_[8327]_ , \new_[8330]_ ,
    \new_[8334]_ , \new_[8335]_ , \new_[8336]_ , \new_[8339]_ ,
    \new_[8343]_ , \new_[8344]_ , \new_[8345]_ , \new_[8348]_ ,
    \new_[8352]_ , \new_[8353]_ , \new_[8354]_ , \new_[8357]_ ,
    \new_[8361]_ , \new_[8362]_ , \new_[8363]_ , \new_[8366]_ ,
    \new_[8370]_ , \new_[8371]_ , \new_[8372]_ , \new_[8375]_ ,
    \new_[8379]_ , \new_[8380]_ , \new_[8381]_ , \new_[8384]_ ,
    \new_[8388]_ , \new_[8389]_ , \new_[8390]_ , \new_[8393]_ ,
    \new_[8397]_ , \new_[8398]_ , \new_[8399]_ , \new_[8402]_ ,
    \new_[8406]_ , \new_[8407]_ , \new_[8408]_ , \new_[8411]_ ,
    \new_[8415]_ , \new_[8416]_ , \new_[8417]_ , \new_[8420]_ ,
    \new_[8424]_ , \new_[8425]_ , \new_[8426]_ , \new_[8429]_ ,
    \new_[8433]_ , \new_[8434]_ , \new_[8435]_ , \new_[8438]_ ,
    \new_[8442]_ , \new_[8443]_ , \new_[8444]_ , \new_[8447]_ ,
    \new_[8451]_ , \new_[8452]_ , \new_[8453]_ , \new_[8456]_ ,
    \new_[8460]_ , \new_[8461]_ , \new_[8462]_ , \new_[8465]_ ,
    \new_[8469]_ , \new_[8470]_ , \new_[8471]_ , \new_[8474]_ ,
    \new_[8478]_ , \new_[8479]_ , \new_[8480]_ , \new_[8483]_ ,
    \new_[8487]_ , \new_[8488]_ , \new_[8489]_ , \new_[8492]_ ,
    \new_[8496]_ , \new_[8497]_ , \new_[8498]_ , \new_[8501]_ ,
    \new_[8505]_ , \new_[8506]_ , \new_[8507]_ , \new_[8510]_ ,
    \new_[8514]_ , \new_[8515]_ , \new_[8516]_ , \new_[8519]_ ,
    \new_[8523]_ , \new_[8524]_ , \new_[8525]_ , \new_[8528]_ ,
    \new_[8532]_ , \new_[8533]_ , \new_[8534]_ , \new_[8537]_ ,
    \new_[8541]_ , \new_[8542]_ , \new_[8543]_ , \new_[8546]_ ,
    \new_[8550]_ , \new_[8551]_ , \new_[8552]_ , \new_[8555]_ ,
    \new_[8559]_ , \new_[8560]_ , \new_[8561]_ , \new_[8564]_ ,
    \new_[8568]_ , \new_[8569]_ , \new_[8570]_ , \new_[8573]_ ,
    \new_[8577]_ , \new_[8578]_ , \new_[8579]_ , \new_[8582]_ ,
    \new_[8586]_ , \new_[8587]_ , \new_[8588]_ , \new_[8591]_ ,
    \new_[8595]_ , \new_[8596]_ , \new_[8597]_ , \new_[8600]_ ,
    \new_[8604]_ , \new_[8605]_ , \new_[8606]_ , \new_[8609]_ ,
    \new_[8613]_ , \new_[8614]_ , \new_[8615]_ , \new_[8618]_ ,
    \new_[8622]_ , \new_[8623]_ , \new_[8624]_ , \new_[8627]_ ,
    \new_[8631]_ , \new_[8632]_ , \new_[8633]_ , \new_[8636]_ ,
    \new_[8640]_ , \new_[8641]_ , \new_[8642]_ , \new_[8645]_ ,
    \new_[8649]_ , \new_[8650]_ , \new_[8651]_ , \new_[8654]_ ,
    \new_[8658]_ , \new_[8659]_ , \new_[8660]_ , \new_[8663]_ ,
    \new_[8667]_ , \new_[8668]_ , \new_[8669]_ , \new_[8672]_ ,
    \new_[8676]_ , \new_[8677]_ , \new_[8678]_ , \new_[8681]_ ,
    \new_[8685]_ , \new_[8686]_ , \new_[8687]_ , \new_[8690]_ ,
    \new_[8694]_ , \new_[8695]_ , \new_[8696]_ , \new_[8699]_ ,
    \new_[8703]_ , \new_[8704]_ , \new_[8705]_ , \new_[8708]_ ,
    \new_[8712]_ , \new_[8713]_ , \new_[8714]_ , \new_[8717]_ ,
    \new_[8721]_ , \new_[8722]_ , \new_[8723]_ , \new_[8726]_ ,
    \new_[8730]_ , \new_[8731]_ , \new_[8732]_ , \new_[8735]_ ,
    \new_[8739]_ , \new_[8740]_ , \new_[8741]_ , \new_[8744]_ ,
    \new_[8748]_ , \new_[8749]_ , \new_[8750]_ , \new_[8753]_ ,
    \new_[8757]_ , \new_[8758]_ , \new_[8759]_ , \new_[8762]_ ,
    \new_[8766]_ , \new_[8767]_ , \new_[8768]_ , \new_[8771]_ ,
    \new_[8775]_ , \new_[8776]_ , \new_[8777]_ , \new_[8780]_ ,
    \new_[8784]_ , \new_[8785]_ , \new_[8786]_ , \new_[8789]_ ,
    \new_[8793]_ , \new_[8794]_ , \new_[8795]_ , \new_[8798]_ ,
    \new_[8802]_ , \new_[8803]_ , \new_[8804]_ , \new_[8807]_ ,
    \new_[8811]_ , \new_[8812]_ , \new_[8813]_ , \new_[8816]_ ,
    \new_[8820]_ , \new_[8821]_ , \new_[8822]_ , \new_[8825]_ ,
    \new_[8829]_ , \new_[8830]_ , \new_[8831]_ , \new_[8834]_ ,
    \new_[8838]_ , \new_[8839]_ , \new_[8840]_ , \new_[8843]_ ,
    \new_[8847]_ , \new_[8848]_ , \new_[8849]_ , \new_[8852]_ ,
    \new_[8856]_ , \new_[8857]_ , \new_[8858]_ , \new_[8861]_ ,
    \new_[8865]_ , \new_[8866]_ , \new_[8867]_ , \new_[8870]_ ,
    \new_[8874]_ , \new_[8875]_ , \new_[8876]_ , \new_[8879]_ ,
    \new_[8883]_ , \new_[8884]_ , \new_[8885]_ , \new_[8888]_ ,
    \new_[8892]_ , \new_[8893]_ , \new_[8894]_ , \new_[8897]_ ,
    \new_[8901]_ , \new_[8902]_ , \new_[8903]_ , \new_[8906]_ ,
    \new_[8910]_ , \new_[8911]_ , \new_[8912]_ , \new_[8915]_ ,
    \new_[8919]_ , \new_[8920]_ , \new_[8921]_ , \new_[8924]_ ,
    \new_[8928]_ , \new_[8929]_ , \new_[8930]_ , \new_[8933]_ ,
    \new_[8937]_ , \new_[8938]_ , \new_[8939]_ , \new_[8942]_ ,
    \new_[8946]_ , \new_[8947]_ , \new_[8948]_ , \new_[8951]_ ,
    \new_[8955]_ , \new_[8956]_ , \new_[8957]_ , \new_[8960]_ ,
    \new_[8964]_ , \new_[8965]_ , \new_[8966]_ , \new_[8969]_ ,
    \new_[8973]_ , \new_[8974]_ , \new_[8975]_ , \new_[8978]_ ,
    \new_[8982]_ , \new_[8983]_ , \new_[8984]_ , \new_[8987]_ ,
    \new_[8991]_ , \new_[8992]_ , \new_[8993]_ , \new_[8996]_ ,
    \new_[9000]_ , \new_[9001]_ , \new_[9002]_ , \new_[9005]_ ,
    \new_[9009]_ , \new_[9010]_ , \new_[9011]_ , \new_[9014]_ ,
    \new_[9018]_ , \new_[9019]_ , \new_[9020]_ , \new_[9023]_ ,
    \new_[9027]_ , \new_[9028]_ , \new_[9029]_ , \new_[9032]_ ,
    \new_[9036]_ , \new_[9037]_ , \new_[9038]_ , \new_[9041]_ ,
    \new_[9045]_ , \new_[9046]_ , \new_[9047]_ , \new_[9050]_ ,
    \new_[9054]_ , \new_[9055]_ , \new_[9056]_ , \new_[9059]_ ,
    \new_[9063]_ , \new_[9064]_ , \new_[9065]_ , \new_[9068]_ ,
    \new_[9072]_ , \new_[9073]_ , \new_[9074]_ , \new_[9077]_ ,
    \new_[9081]_ , \new_[9082]_ , \new_[9083]_ , \new_[9086]_ ,
    \new_[9090]_ , \new_[9091]_ , \new_[9092]_ , \new_[9095]_ ,
    \new_[9099]_ , \new_[9100]_ , \new_[9101]_ , \new_[9104]_ ,
    \new_[9108]_ , \new_[9109]_ , \new_[9110]_ , \new_[9113]_ ,
    \new_[9117]_ , \new_[9118]_ , \new_[9119]_ , \new_[9122]_ ,
    \new_[9126]_ , \new_[9127]_ , \new_[9128]_ , \new_[9131]_ ,
    \new_[9135]_ , \new_[9136]_ , \new_[9137]_ , \new_[9140]_ ,
    \new_[9144]_ , \new_[9145]_ , \new_[9146]_ , \new_[9149]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9155]_ , \new_[9158]_ ,
    \new_[9162]_ , \new_[9163]_ , \new_[9164]_ , \new_[9167]_ ,
    \new_[9171]_ , \new_[9172]_ , \new_[9173]_ , \new_[9176]_ ,
    \new_[9180]_ , \new_[9181]_ , \new_[9182]_ , \new_[9185]_ ,
    \new_[9189]_ , \new_[9190]_ , \new_[9191]_ , \new_[9194]_ ,
    \new_[9198]_ , \new_[9199]_ , \new_[9200]_ , \new_[9203]_ ,
    \new_[9207]_ , \new_[9208]_ , \new_[9209]_ , \new_[9212]_ ,
    \new_[9216]_ , \new_[9217]_ , \new_[9218]_ , \new_[9221]_ ,
    \new_[9225]_ , \new_[9226]_ , \new_[9227]_ , \new_[9230]_ ,
    \new_[9234]_ , \new_[9235]_ , \new_[9236]_ , \new_[9239]_ ,
    \new_[9243]_ , \new_[9244]_ , \new_[9245]_ , \new_[9248]_ ,
    \new_[9252]_ , \new_[9253]_ , \new_[9254]_ , \new_[9257]_ ,
    \new_[9261]_ , \new_[9262]_ , \new_[9263]_ , \new_[9266]_ ,
    \new_[9270]_ , \new_[9271]_ , \new_[9272]_ , \new_[9275]_ ,
    \new_[9279]_ , \new_[9280]_ , \new_[9281]_ , \new_[9284]_ ,
    \new_[9288]_ , \new_[9289]_ , \new_[9290]_ , \new_[9293]_ ,
    \new_[9297]_ , \new_[9298]_ , \new_[9299]_ , \new_[9302]_ ,
    \new_[9306]_ , \new_[9307]_ , \new_[9308]_ , \new_[9311]_ ,
    \new_[9315]_ , \new_[9316]_ , \new_[9317]_ , \new_[9320]_ ,
    \new_[9324]_ , \new_[9325]_ , \new_[9326]_ , \new_[9329]_ ,
    \new_[9333]_ , \new_[9334]_ , \new_[9335]_ , \new_[9338]_ ,
    \new_[9342]_ , \new_[9343]_ , \new_[9344]_ , \new_[9347]_ ,
    \new_[9351]_ , \new_[9352]_ , \new_[9353]_ , \new_[9356]_ ,
    \new_[9360]_ , \new_[9361]_ , \new_[9362]_ , \new_[9365]_ ,
    \new_[9369]_ , \new_[9370]_ , \new_[9371]_ , \new_[9374]_ ,
    \new_[9378]_ , \new_[9379]_ , \new_[9380]_ , \new_[9383]_ ,
    \new_[9387]_ , \new_[9388]_ , \new_[9389]_ , \new_[9392]_ ,
    \new_[9396]_ , \new_[9397]_ , \new_[9398]_ , \new_[9401]_ ,
    \new_[9405]_ , \new_[9406]_ , \new_[9407]_ , \new_[9410]_ ,
    \new_[9414]_ , \new_[9415]_ , \new_[9416]_ , \new_[9419]_ ,
    \new_[9423]_ , \new_[9424]_ , \new_[9425]_ , \new_[9428]_ ,
    \new_[9432]_ , \new_[9433]_ , \new_[9434]_ , \new_[9437]_ ,
    \new_[9441]_ , \new_[9442]_ , \new_[9443]_ , \new_[9446]_ ,
    \new_[9450]_ , \new_[9451]_ , \new_[9452]_ , \new_[9455]_ ,
    \new_[9459]_ , \new_[9460]_ , \new_[9461]_ , \new_[9464]_ ,
    \new_[9468]_ , \new_[9469]_ , \new_[9470]_ , \new_[9473]_ ,
    \new_[9477]_ , \new_[9478]_ , \new_[9479]_ , \new_[9482]_ ,
    \new_[9486]_ , \new_[9487]_ , \new_[9488]_ , \new_[9491]_ ,
    \new_[9495]_ , \new_[9496]_ , \new_[9497]_ , \new_[9500]_ ,
    \new_[9504]_ , \new_[9505]_ , \new_[9506]_ , \new_[9509]_ ,
    \new_[9513]_ , \new_[9514]_ , \new_[9515]_ , \new_[9518]_ ,
    \new_[9522]_ , \new_[9523]_ , \new_[9524]_ , \new_[9527]_ ,
    \new_[9531]_ , \new_[9532]_ , \new_[9533]_ , \new_[9536]_ ,
    \new_[9540]_ , \new_[9541]_ , \new_[9542]_ , \new_[9545]_ ,
    \new_[9549]_ , \new_[9550]_ , \new_[9551]_ , \new_[9554]_ ,
    \new_[9558]_ , \new_[9559]_ , \new_[9560]_ , \new_[9563]_ ,
    \new_[9567]_ , \new_[9568]_ , \new_[9569]_ , \new_[9572]_ ,
    \new_[9576]_ , \new_[9577]_ , \new_[9578]_ , \new_[9581]_ ,
    \new_[9585]_ , \new_[9586]_ , \new_[9587]_ , \new_[9590]_ ,
    \new_[9594]_ , \new_[9595]_ , \new_[9596]_ , \new_[9599]_ ,
    \new_[9603]_ , \new_[9604]_ , \new_[9605]_ , \new_[9608]_ ,
    \new_[9612]_ , \new_[9613]_ , \new_[9614]_ , \new_[9617]_ ,
    \new_[9621]_ , \new_[9622]_ , \new_[9623]_ , \new_[9626]_ ,
    \new_[9630]_ , \new_[9631]_ , \new_[9632]_ , \new_[9635]_ ,
    \new_[9639]_ , \new_[9640]_ , \new_[9641]_ , \new_[9644]_ ,
    \new_[9648]_ , \new_[9649]_ , \new_[9650]_ , \new_[9653]_ ,
    \new_[9657]_ , \new_[9658]_ , \new_[9659]_ , \new_[9662]_ ,
    \new_[9666]_ , \new_[9667]_ , \new_[9668]_ , \new_[9671]_ ,
    \new_[9675]_ , \new_[9676]_ , \new_[9677]_ , \new_[9680]_ ,
    \new_[9684]_ , \new_[9685]_ , \new_[9686]_ , \new_[9689]_ ,
    \new_[9693]_ , \new_[9694]_ , \new_[9695]_ , \new_[9698]_ ,
    \new_[9702]_ , \new_[9703]_ , \new_[9704]_ , \new_[9707]_ ,
    \new_[9711]_ , \new_[9712]_ , \new_[9713]_ , \new_[9716]_ ,
    \new_[9720]_ , \new_[9721]_ , \new_[9722]_ , \new_[9725]_ ,
    \new_[9729]_ , \new_[9730]_ , \new_[9731]_ , \new_[9734]_ ,
    \new_[9738]_ , \new_[9739]_ , \new_[9740]_ , \new_[9743]_ ,
    \new_[9747]_ , \new_[9748]_ , \new_[9749]_ , \new_[9752]_ ,
    \new_[9756]_ , \new_[9757]_ , \new_[9758]_ , \new_[9761]_ ,
    \new_[9765]_ , \new_[9766]_ , \new_[9767]_ , \new_[9770]_ ,
    \new_[9774]_ , \new_[9775]_ , \new_[9776]_ , \new_[9779]_ ,
    \new_[9783]_ , \new_[9784]_ , \new_[9785]_ , \new_[9788]_ ,
    \new_[9792]_ , \new_[9793]_ , \new_[9794]_ , \new_[9797]_ ,
    \new_[9801]_ , \new_[9802]_ , \new_[9803]_ , \new_[9806]_ ,
    \new_[9810]_ , \new_[9811]_ , \new_[9812]_ , \new_[9815]_ ,
    \new_[9819]_ , \new_[9820]_ , \new_[9821]_ , \new_[9824]_ ,
    \new_[9828]_ , \new_[9829]_ , \new_[9830]_ , \new_[9833]_ ,
    \new_[9837]_ , \new_[9838]_ , \new_[9839]_ , \new_[9842]_ ,
    \new_[9846]_ , \new_[9847]_ , \new_[9848]_ , \new_[9851]_ ,
    \new_[9855]_ , \new_[9856]_ , \new_[9857]_ , \new_[9860]_ ,
    \new_[9864]_ , \new_[9865]_ , \new_[9866]_ , \new_[9869]_ ,
    \new_[9873]_ , \new_[9874]_ , \new_[9875]_ , \new_[9878]_ ,
    \new_[9882]_ , \new_[9883]_ , \new_[9884]_ , \new_[9887]_ ,
    \new_[9891]_ , \new_[9892]_ , \new_[9893]_ , \new_[9896]_ ,
    \new_[9900]_ , \new_[9901]_ , \new_[9902]_ , \new_[9905]_ ,
    \new_[9909]_ , \new_[9910]_ , \new_[9911]_ , \new_[9914]_ ,
    \new_[9918]_ , \new_[9919]_ , \new_[9920]_ , \new_[9923]_ ,
    \new_[9927]_ , \new_[9928]_ , \new_[9929]_ , \new_[9932]_ ,
    \new_[9936]_ , \new_[9937]_ , \new_[9938]_ , \new_[9941]_ ,
    \new_[9945]_ , \new_[9946]_ , \new_[9947]_ , \new_[9950]_ ,
    \new_[9954]_ , \new_[9955]_ , \new_[9956]_ , \new_[9959]_ ,
    \new_[9963]_ , \new_[9964]_ , \new_[9965]_ , \new_[9968]_ ,
    \new_[9972]_ , \new_[9973]_ , \new_[9974]_ , \new_[9977]_ ,
    \new_[9981]_ , \new_[9982]_ , \new_[9983]_ , \new_[9986]_ ,
    \new_[9990]_ , \new_[9991]_ , \new_[9992]_ , \new_[9995]_ ,
    \new_[9999]_ , \new_[10000]_ , \new_[10001]_ , \new_[10004]_ ,
    \new_[10008]_ , \new_[10009]_ , \new_[10010]_ , \new_[10013]_ ,
    \new_[10017]_ , \new_[10018]_ , \new_[10019]_ , \new_[10022]_ ,
    \new_[10026]_ , \new_[10027]_ , \new_[10028]_ , \new_[10031]_ ,
    \new_[10035]_ , \new_[10036]_ , \new_[10037]_ , \new_[10040]_ ,
    \new_[10044]_ , \new_[10045]_ , \new_[10046]_ , \new_[10049]_ ,
    \new_[10053]_ , \new_[10054]_ , \new_[10055]_ , \new_[10058]_ ,
    \new_[10062]_ , \new_[10063]_ , \new_[10064]_ , \new_[10067]_ ,
    \new_[10071]_ , \new_[10072]_ , \new_[10073]_ , \new_[10076]_ ,
    \new_[10080]_ , \new_[10081]_ , \new_[10082]_ , \new_[10085]_ ,
    \new_[10089]_ , \new_[10090]_ , \new_[10091]_ , \new_[10094]_ ,
    \new_[10098]_ , \new_[10099]_ , \new_[10100]_ , \new_[10103]_ ,
    \new_[10107]_ , \new_[10108]_ , \new_[10109]_ , \new_[10112]_ ,
    \new_[10116]_ , \new_[10117]_ , \new_[10118]_ , \new_[10121]_ ,
    \new_[10125]_ , \new_[10126]_ , \new_[10127]_ , \new_[10130]_ ,
    \new_[10134]_ , \new_[10135]_ , \new_[10136]_ , \new_[10139]_ ,
    \new_[10143]_ , \new_[10144]_ , \new_[10145]_ , \new_[10148]_ ,
    \new_[10152]_ , \new_[10153]_ , \new_[10154]_ , \new_[10157]_ ,
    \new_[10161]_ , \new_[10162]_ , \new_[10163]_ , \new_[10166]_ ,
    \new_[10170]_ , \new_[10171]_ , \new_[10172]_ , \new_[10175]_ ,
    \new_[10179]_ , \new_[10180]_ , \new_[10181]_ , \new_[10184]_ ,
    \new_[10188]_ , \new_[10189]_ , \new_[10190]_ , \new_[10193]_ ,
    \new_[10197]_ , \new_[10198]_ , \new_[10199]_ , \new_[10202]_ ,
    \new_[10206]_ , \new_[10207]_ , \new_[10208]_ , \new_[10211]_ ,
    \new_[10215]_ , \new_[10216]_ , \new_[10217]_ , \new_[10220]_ ,
    \new_[10224]_ , \new_[10225]_ , \new_[10226]_ , \new_[10229]_ ,
    \new_[10233]_ , \new_[10234]_ , \new_[10235]_ , \new_[10238]_ ,
    \new_[10242]_ , \new_[10243]_ , \new_[10244]_ , \new_[10247]_ ,
    \new_[10251]_ , \new_[10252]_ , \new_[10253]_ , \new_[10256]_ ,
    \new_[10260]_ , \new_[10261]_ , \new_[10262]_ , \new_[10265]_ ,
    \new_[10269]_ , \new_[10270]_ , \new_[10271]_ , \new_[10274]_ ,
    \new_[10278]_ , \new_[10279]_ , \new_[10280]_ , \new_[10283]_ ,
    \new_[10287]_ , \new_[10288]_ , \new_[10289]_ , \new_[10292]_ ,
    \new_[10296]_ , \new_[10297]_ , \new_[10298]_ , \new_[10301]_ ,
    \new_[10305]_ , \new_[10306]_ , \new_[10307]_ , \new_[10310]_ ,
    \new_[10314]_ , \new_[10315]_ , \new_[10316]_ , \new_[10319]_ ,
    \new_[10323]_ , \new_[10324]_ , \new_[10325]_ , \new_[10328]_ ,
    \new_[10332]_ , \new_[10333]_ , \new_[10334]_ , \new_[10338]_ ,
    \new_[10339]_ , \new_[10343]_ , \new_[10344]_ , \new_[10345]_ ,
    \new_[10348]_ , \new_[10352]_ , \new_[10353]_ , \new_[10354]_ ,
    \new_[10358]_ , \new_[10359]_ , \new_[10363]_ , \new_[10364]_ ,
    \new_[10365]_ , \new_[10368]_ , \new_[10372]_ , \new_[10373]_ ,
    \new_[10374]_ , \new_[10378]_ , \new_[10379]_ , \new_[10383]_ ,
    \new_[10384]_ , \new_[10385]_ , \new_[10388]_ , \new_[10392]_ ,
    \new_[10393]_ , \new_[10394]_ , \new_[10398]_ , \new_[10399]_ ,
    \new_[10403]_ , \new_[10404]_ , \new_[10405]_ , \new_[10408]_ ,
    \new_[10412]_ , \new_[10413]_ , \new_[10414]_ , \new_[10418]_ ,
    \new_[10419]_ , \new_[10423]_ , \new_[10424]_ , \new_[10425]_ ,
    \new_[10428]_ , \new_[10432]_ , \new_[10433]_ , \new_[10434]_ ,
    \new_[10438]_ , \new_[10439]_ , \new_[10443]_ , \new_[10444]_ ,
    \new_[10445]_ , \new_[10448]_ , \new_[10452]_ , \new_[10453]_ ,
    \new_[10454]_ , \new_[10458]_ , \new_[10459]_ , \new_[10463]_ ,
    \new_[10464]_ , \new_[10465]_ , \new_[10468]_ , \new_[10472]_ ,
    \new_[10473]_ , \new_[10474]_ , \new_[10478]_ , \new_[10479]_ ,
    \new_[10483]_ , \new_[10484]_ , \new_[10485]_ , \new_[10488]_ ,
    \new_[10492]_ , \new_[10493]_ , \new_[10494]_ , \new_[10498]_ ,
    \new_[10499]_ , \new_[10503]_ , \new_[10504]_ , \new_[10505]_ ,
    \new_[10508]_ , \new_[10512]_ , \new_[10513]_ , \new_[10514]_ ,
    \new_[10518]_ , \new_[10519]_ , \new_[10523]_ , \new_[10524]_ ,
    \new_[10525]_ , \new_[10528]_ , \new_[10532]_ , \new_[10533]_ ,
    \new_[10534]_ , \new_[10538]_ , \new_[10539]_ , \new_[10543]_ ,
    \new_[10544]_ , \new_[10545]_ , \new_[10548]_ , \new_[10552]_ ,
    \new_[10553]_ , \new_[10554]_ , \new_[10558]_ , \new_[10559]_ ,
    \new_[10563]_ , \new_[10564]_ , \new_[10565]_ , \new_[10568]_ ,
    \new_[10572]_ , \new_[10573]_ , \new_[10574]_ , \new_[10578]_ ,
    \new_[10579]_ , \new_[10583]_ , \new_[10584]_ , \new_[10585]_ ,
    \new_[10588]_ , \new_[10592]_ , \new_[10593]_ , \new_[10594]_ ,
    \new_[10598]_ , \new_[10599]_ , \new_[10603]_ , \new_[10604]_ ,
    \new_[10605]_ , \new_[10608]_ , \new_[10612]_ , \new_[10613]_ ,
    \new_[10614]_ , \new_[10618]_ , \new_[10619]_ , \new_[10623]_ ,
    \new_[10624]_ , \new_[10625]_ , \new_[10628]_ , \new_[10632]_ ,
    \new_[10633]_ , \new_[10634]_ , \new_[10638]_ , \new_[10639]_ ,
    \new_[10643]_ , \new_[10644]_ , \new_[10645]_ , \new_[10648]_ ,
    \new_[10652]_ , \new_[10653]_ , \new_[10654]_ , \new_[10658]_ ,
    \new_[10659]_ , \new_[10663]_ , \new_[10664]_ , \new_[10665]_ ,
    \new_[10668]_ , \new_[10672]_ , \new_[10673]_ , \new_[10674]_ ,
    \new_[10678]_ , \new_[10679]_ , \new_[10683]_ , \new_[10684]_ ,
    \new_[10685]_ , \new_[10688]_ , \new_[10692]_ , \new_[10693]_ ,
    \new_[10694]_ , \new_[10698]_ , \new_[10699]_ , \new_[10703]_ ,
    \new_[10704]_ , \new_[10705]_ , \new_[10708]_ , \new_[10712]_ ,
    \new_[10713]_ , \new_[10714]_ , \new_[10718]_ , \new_[10719]_ ,
    \new_[10723]_ , \new_[10724]_ , \new_[10725]_ , \new_[10728]_ ,
    \new_[10732]_ , \new_[10733]_ , \new_[10734]_ , \new_[10738]_ ,
    \new_[10739]_ , \new_[10743]_ , \new_[10744]_ , \new_[10745]_ ,
    \new_[10748]_ , \new_[10752]_ , \new_[10753]_ , \new_[10754]_ ,
    \new_[10758]_ , \new_[10759]_ , \new_[10763]_ , \new_[10764]_ ,
    \new_[10765]_ , \new_[10768]_ , \new_[10772]_ , \new_[10773]_ ,
    \new_[10774]_ , \new_[10778]_ , \new_[10779]_ , \new_[10783]_ ,
    \new_[10784]_ , \new_[10785]_ , \new_[10788]_ , \new_[10792]_ ,
    \new_[10793]_ , \new_[10794]_ , \new_[10798]_ , \new_[10799]_ ,
    \new_[10803]_ , \new_[10804]_ , \new_[10805]_ , \new_[10808]_ ,
    \new_[10812]_ , \new_[10813]_ , \new_[10814]_ , \new_[10818]_ ,
    \new_[10819]_ , \new_[10823]_ , \new_[10824]_ , \new_[10825]_ ,
    \new_[10828]_ , \new_[10832]_ , \new_[10833]_ , \new_[10834]_ ,
    \new_[10838]_ , \new_[10839]_ , \new_[10843]_ , \new_[10844]_ ,
    \new_[10845]_ , \new_[10848]_ , \new_[10852]_ , \new_[10853]_ ,
    \new_[10854]_ , \new_[10858]_ , \new_[10859]_ , \new_[10863]_ ,
    \new_[10864]_ , \new_[10865]_ , \new_[10868]_ , \new_[10872]_ ,
    \new_[10873]_ , \new_[10874]_ , \new_[10878]_ , \new_[10879]_ ,
    \new_[10883]_ , \new_[10884]_ , \new_[10885]_ , \new_[10888]_ ,
    \new_[10892]_ , \new_[10893]_ , \new_[10894]_ , \new_[10898]_ ,
    \new_[10899]_ , \new_[10903]_ , \new_[10904]_ , \new_[10905]_ ,
    \new_[10908]_ , \new_[10912]_ , \new_[10913]_ , \new_[10914]_ ,
    \new_[10918]_ , \new_[10919]_ , \new_[10923]_ , \new_[10924]_ ,
    \new_[10925]_ , \new_[10928]_ , \new_[10932]_ , \new_[10933]_ ,
    \new_[10934]_ , \new_[10938]_ , \new_[10939]_ , \new_[10943]_ ,
    \new_[10944]_ , \new_[10945]_ , \new_[10948]_ , \new_[10952]_ ,
    \new_[10953]_ , \new_[10954]_ , \new_[10958]_ , \new_[10959]_ ,
    \new_[10963]_ , \new_[10964]_ , \new_[10965]_ , \new_[10968]_ ,
    \new_[10972]_ , \new_[10973]_ , \new_[10974]_ , \new_[10978]_ ,
    \new_[10979]_ , \new_[10983]_ , \new_[10984]_ , \new_[10985]_ ,
    \new_[10988]_ , \new_[10992]_ , \new_[10993]_ , \new_[10994]_ ,
    \new_[10998]_ , \new_[10999]_ , \new_[11003]_ , \new_[11004]_ ,
    \new_[11005]_ , \new_[11008]_ , \new_[11012]_ , \new_[11013]_ ,
    \new_[11014]_ , \new_[11018]_ , \new_[11019]_ , \new_[11023]_ ,
    \new_[11024]_ , \new_[11025]_ , \new_[11028]_ , \new_[11032]_ ,
    \new_[11033]_ , \new_[11034]_ , \new_[11038]_ , \new_[11039]_ ,
    \new_[11043]_ , \new_[11044]_ , \new_[11045]_ , \new_[11048]_ ,
    \new_[11052]_ , \new_[11053]_ , \new_[11054]_ , \new_[11058]_ ,
    \new_[11059]_ , \new_[11063]_ , \new_[11064]_ , \new_[11065]_ ,
    \new_[11068]_ , \new_[11072]_ , \new_[11073]_ , \new_[11074]_ ,
    \new_[11078]_ , \new_[11079]_ , \new_[11083]_ , \new_[11084]_ ,
    \new_[11085]_ , \new_[11088]_ , \new_[11092]_ , \new_[11093]_ ,
    \new_[11094]_ , \new_[11098]_ , \new_[11099]_ , \new_[11103]_ ,
    \new_[11104]_ , \new_[11105]_ , \new_[11108]_ , \new_[11112]_ ,
    \new_[11113]_ , \new_[11114]_ , \new_[11118]_ , \new_[11119]_ ,
    \new_[11123]_ , \new_[11124]_ , \new_[11125]_ , \new_[11128]_ ,
    \new_[11132]_ , \new_[11133]_ , \new_[11134]_ , \new_[11138]_ ,
    \new_[11139]_ , \new_[11143]_ , \new_[11144]_ , \new_[11145]_ ,
    \new_[11148]_ , \new_[11152]_ , \new_[11153]_ , \new_[11154]_ ,
    \new_[11158]_ , \new_[11159]_ , \new_[11163]_ , \new_[11164]_ ,
    \new_[11165]_ , \new_[11168]_ , \new_[11172]_ , \new_[11173]_ ,
    \new_[11174]_ , \new_[11178]_ , \new_[11179]_ , \new_[11183]_ ,
    \new_[11184]_ , \new_[11185]_ , \new_[11188]_ , \new_[11192]_ ,
    \new_[11193]_ , \new_[11194]_ , \new_[11198]_ , \new_[11199]_ ,
    \new_[11203]_ , \new_[11204]_ , \new_[11205]_ , \new_[11208]_ ,
    \new_[11212]_ , \new_[11213]_ , \new_[11214]_ , \new_[11218]_ ,
    \new_[11219]_ , \new_[11223]_ , \new_[11224]_ , \new_[11225]_ ,
    \new_[11228]_ , \new_[11232]_ , \new_[11233]_ , \new_[11234]_ ,
    \new_[11238]_ , \new_[11239]_ , \new_[11243]_ , \new_[11244]_ ,
    \new_[11245]_ , \new_[11248]_ , \new_[11252]_ , \new_[11253]_ ,
    \new_[11254]_ , \new_[11258]_ , \new_[11259]_ , \new_[11263]_ ,
    \new_[11264]_ , \new_[11265]_ , \new_[11268]_ , \new_[11272]_ ,
    \new_[11273]_ , \new_[11274]_ , \new_[11278]_ , \new_[11279]_ ,
    \new_[11283]_ , \new_[11284]_ , \new_[11285]_ , \new_[11288]_ ,
    \new_[11292]_ , \new_[11293]_ , \new_[11294]_ , \new_[11298]_ ,
    \new_[11299]_ , \new_[11303]_ , \new_[11304]_ , \new_[11305]_ ,
    \new_[11308]_ , \new_[11312]_ , \new_[11313]_ , \new_[11314]_ ,
    \new_[11318]_ , \new_[11319]_ , \new_[11323]_ , \new_[11324]_ ,
    \new_[11325]_ , \new_[11328]_ , \new_[11332]_ , \new_[11333]_ ,
    \new_[11334]_ , \new_[11338]_ , \new_[11339]_ , \new_[11343]_ ,
    \new_[11344]_ , \new_[11345]_ , \new_[11348]_ , \new_[11352]_ ,
    \new_[11353]_ , \new_[11354]_ , \new_[11358]_ , \new_[11359]_ ,
    \new_[11363]_ , \new_[11364]_ , \new_[11365]_ , \new_[11368]_ ,
    \new_[11372]_ , \new_[11373]_ , \new_[11374]_ , \new_[11378]_ ,
    \new_[11379]_ , \new_[11383]_ , \new_[11384]_ , \new_[11385]_ ,
    \new_[11388]_ , \new_[11392]_ , \new_[11393]_ , \new_[11394]_ ,
    \new_[11398]_ , \new_[11399]_ , \new_[11403]_ , \new_[11404]_ ,
    \new_[11405]_ , \new_[11408]_ , \new_[11412]_ , \new_[11413]_ ,
    \new_[11414]_ , \new_[11418]_ , \new_[11419]_ , \new_[11423]_ ,
    \new_[11424]_ , \new_[11425]_ , \new_[11428]_ , \new_[11432]_ ,
    \new_[11433]_ , \new_[11434]_ , \new_[11438]_ , \new_[11439]_ ,
    \new_[11443]_ , \new_[11444]_ , \new_[11445]_ , \new_[11448]_ ,
    \new_[11452]_ , \new_[11453]_ , \new_[11454]_ , \new_[11458]_ ,
    \new_[11459]_ , \new_[11463]_ , \new_[11464]_ , \new_[11465]_ ,
    \new_[11468]_ , \new_[11472]_ , \new_[11473]_ , \new_[11474]_ ,
    \new_[11478]_ , \new_[11479]_ , \new_[11483]_ , \new_[11484]_ ,
    \new_[11485]_ , \new_[11488]_ , \new_[11492]_ , \new_[11493]_ ,
    \new_[11494]_ , \new_[11498]_ , \new_[11499]_ , \new_[11503]_ ,
    \new_[11504]_ , \new_[11505]_ , \new_[11508]_ , \new_[11512]_ ,
    \new_[11513]_ , \new_[11514]_ , \new_[11518]_ , \new_[11519]_ ,
    \new_[11523]_ , \new_[11524]_ , \new_[11525]_ , \new_[11528]_ ,
    \new_[11532]_ , \new_[11533]_ , \new_[11534]_ , \new_[11538]_ ,
    \new_[11539]_ , \new_[11543]_ , \new_[11544]_ , \new_[11545]_ ,
    \new_[11548]_ , \new_[11552]_ , \new_[11553]_ , \new_[11554]_ ,
    \new_[11558]_ , \new_[11559]_ , \new_[11563]_ , \new_[11564]_ ,
    \new_[11565]_ , \new_[11568]_ , \new_[11572]_ , \new_[11573]_ ,
    \new_[11574]_ , \new_[11578]_ , \new_[11579]_ , \new_[11583]_ ,
    \new_[11584]_ , \new_[11585]_ , \new_[11588]_ , \new_[11592]_ ,
    \new_[11593]_ , \new_[11594]_ , \new_[11598]_ , \new_[11599]_ ,
    \new_[11603]_ , \new_[11604]_ , \new_[11605]_ , \new_[11608]_ ,
    \new_[11612]_ , \new_[11613]_ , \new_[11614]_ , \new_[11618]_ ,
    \new_[11619]_ , \new_[11623]_ , \new_[11624]_ , \new_[11625]_ ,
    \new_[11628]_ , \new_[11632]_ , \new_[11633]_ , \new_[11634]_ ,
    \new_[11638]_ , \new_[11639]_ , \new_[11643]_ , \new_[11644]_ ,
    \new_[11645]_ , \new_[11648]_ , \new_[11652]_ , \new_[11653]_ ,
    \new_[11654]_ , \new_[11658]_ , \new_[11659]_ , \new_[11663]_ ,
    \new_[11664]_ , \new_[11665]_ , \new_[11668]_ , \new_[11672]_ ,
    \new_[11673]_ , \new_[11674]_ , \new_[11678]_ , \new_[11679]_ ,
    \new_[11683]_ , \new_[11684]_ , \new_[11685]_ , \new_[11688]_ ,
    \new_[11692]_ , \new_[11693]_ , \new_[11694]_ , \new_[11698]_ ,
    \new_[11699]_ , \new_[11703]_ , \new_[11704]_ , \new_[11705]_ ,
    \new_[11708]_ , \new_[11712]_ , \new_[11713]_ , \new_[11714]_ ,
    \new_[11718]_ , \new_[11719]_ , \new_[11723]_ , \new_[11724]_ ,
    \new_[11725]_ , \new_[11728]_ , \new_[11732]_ , \new_[11733]_ ,
    \new_[11734]_ , \new_[11738]_ , \new_[11739]_ , \new_[11743]_ ,
    \new_[11744]_ , \new_[11745]_ , \new_[11748]_ , \new_[11752]_ ,
    \new_[11753]_ , \new_[11754]_ , \new_[11758]_ , \new_[11759]_ ,
    \new_[11763]_ , \new_[11764]_ , \new_[11765]_ , \new_[11768]_ ,
    \new_[11772]_ , \new_[11773]_ , \new_[11774]_ , \new_[11778]_ ,
    \new_[11779]_ , \new_[11783]_ , \new_[11784]_ , \new_[11785]_ ,
    \new_[11788]_ , \new_[11792]_ , \new_[11793]_ , \new_[11794]_ ,
    \new_[11798]_ , \new_[11799]_ , \new_[11803]_ , \new_[11804]_ ,
    \new_[11805]_ , \new_[11808]_ , \new_[11812]_ , \new_[11813]_ ,
    \new_[11814]_ , \new_[11818]_ , \new_[11819]_ , \new_[11823]_ ,
    \new_[11824]_ , \new_[11825]_ , \new_[11828]_ , \new_[11832]_ ,
    \new_[11833]_ , \new_[11834]_ , \new_[11838]_ , \new_[11839]_ ,
    \new_[11843]_ , \new_[11844]_ , \new_[11845]_ , \new_[11848]_ ,
    \new_[11852]_ , \new_[11853]_ , \new_[11854]_ , \new_[11858]_ ,
    \new_[11859]_ , \new_[11863]_ , \new_[11864]_ , \new_[11865]_ ,
    \new_[11868]_ , \new_[11872]_ , \new_[11873]_ , \new_[11874]_ ,
    \new_[11878]_ , \new_[11879]_ , \new_[11883]_ , \new_[11884]_ ,
    \new_[11885]_ , \new_[11888]_ , \new_[11892]_ , \new_[11893]_ ,
    \new_[11894]_ , \new_[11898]_ , \new_[11899]_ , \new_[11903]_ ,
    \new_[11904]_ , \new_[11905]_ , \new_[11908]_ , \new_[11912]_ ,
    \new_[11913]_ , \new_[11914]_ , \new_[11918]_ , \new_[11919]_ ,
    \new_[11923]_ , \new_[11924]_ , \new_[11925]_ , \new_[11928]_ ,
    \new_[11932]_ , \new_[11933]_ , \new_[11934]_ , \new_[11938]_ ,
    \new_[11939]_ , \new_[11943]_ , \new_[11944]_ , \new_[11945]_ ,
    \new_[11948]_ , \new_[11952]_ , \new_[11953]_ , \new_[11954]_ ,
    \new_[11958]_ , \new_[11959]_ , \new_[11963]_ , \new_[11964]_ ,
    \new_[11965]_ , \new_[11968]_ , \new_[11972]_ , \new_[11973]_ ,
    \new_[11974]_ , \new_[11978]_ , \new_[11979]_ , \new_[11983]_ ,
    \new_[11984]_ , \new_[11985]_ , \new_[11988]_ , \new_[11992]_ ,
    \new_[11993]_ , \new_[11994]_ , \new_[11998]_ , \new_[11999]_ ,
    \new_[12003]_ , \new_[12004]_ , \new_[12005]_ , \new_[12008]_ ,
    \new_[12012]_ , \new_[12013]_ , \new_[12014]_ , \new_[12018]_ ,
    \new_[12019]_ , \new_[12023]_ , \new_[12024]_ , \new_[12025]_ ,
    \new_[12028]_ , \new_[12032]_ , \new_[12033]_ , \new_[12034]_ ,
    \new_[12038]_ , \new_[12039]_ , \new_[12043]_ , \new_[12044]_ ,
    \new_[12045]_ , \new_[12048]_ , \new_[12052]_ , \new_[12053]_ ,
    \new_[12054]_ , \new_[12058]_ , \new_[12059]_ , \new_[12063]_ ,
    \new_[12064]_ , \new_[12065]_ , \new_[12068]_ , \new_[12072]_ ,
    \new_[12073]_ , \new_[12074]_ , \new_[12078]_ , \new_[12079]_ ,
    \new_[12083]_ , \new_[12084]_ , \new_[12085]_ , \new_[12088]_ ,
    \new_[12092]_ , \new_[12093]_ , \new_[12094]_ , \new_[12098]_ ,
    \new_[12099]_ , \new_[12103]_ , \new_[12104]_ , \new_[12105]_ ,
    \new_[12108]_ , \new_[12112]_ , \new_[12113]_ , \new_[12114]_ ,
    \new_[12118]_ , \new_[12119]_ , \new_[12123]_ , \new_[12124]_ ,
    \new_[12125]_ , \new_[12128]_ , \new_[12132]_ , \new_[12133]_ ,
    \new_[12134]_ , \new_[12138]_ , \new_[12139]_ , \new_[12143]_ ,
    \new_[12144]_ , \new_[12145]_ , \new_[12148]_ , \new_[12152]_ ,
    \new_[12153]_ , \new_[12154]_ , \new_[12158]_ , \new_[12159]_ ,
    \new_[12163]_ , \new_[12164]_ , \new_[12165]_ , \new_[12168]_ ,
    \new_[12172]_ , \new_[12173]_ , \new_[12174]_ , \new_[12178]_ ,
    \new_[12179]_ , \new_[12183]_ , \new_[12184]_ , \new_[12185]_ ,
    \new_[12188]_ , \new_[12192]_ , \new_[12193]_ , \new_[12194]_ ,
    \new_[12198]_ , \new_[12199]_ , \new_[12203]_ , \new_[12204]_ ,
    \new_[12205]_ , \new_[12208]_ , \new_[12212]_ , \new_[12213]_ ,
    \new_[12214]_ , \new_[12218]_ , \new_[12219]_ , \new_[12223]_ ,
    \new_[12224]_ , \new_[12225]_ , \new_[12228]_ , \new_[12232]_ ,
    \new_[12233]_ , \new_[12234]_ , \new_[12238]_ , \new_[12239]_ ,
    \new_[12243]_ , \new_[12244]_ , \new_[12245]_ , \new_[12248]_ ,
    \new_[12252]_ , \new_[12253]_ , \new_[12254]_ , \new_[12258]_ ,
    \new_[12259]_ , \new_[12263]_ , \new_[12264]_ , \new_[12265]_ ,
    \new_[12268]_ , \new_[12272]_ , \new_[12273]_ , \new_[12274]_ ,
    \new_[12278]_ , \new_[12279]_ , \new_[12283]_ , \new_[12284]_ ,
    \new_[12285]_ , \new_[12288]_ , \new_[12292]_ , \new_[12293]_ ,
    \new_[12294]_ , \new_[12298]_ , \new_[12299]_ , \new_[12303]_ ,
    \new_[12304]_ , \new_[12305]_ , \new_[12308]_ , \new_[12312]_ ,
    \new_[12313]_ , \new_[12314]_ , \new_[12318]_ , \new_[12319]_ ,
    \new_[12323]_ , \new_[12324]_ , \new_[12325]_ , \new_[12328]_ ,
    \new_[12332]_ , \new_[12333]_ , \new_[12334]_ , \new_[12338]_ ,
    \new_[12339]_ , \new_[12343]_ , \new_[12344]_ , \new_[12345]_ ,
    \new_[12348]_ , \new_[12352]_ , \new_[12353]_ , \new_[12354]_ ,
    \new_[12358]_ , \new_[12359]_ , \new_[12363]_ , \new_[12364]_ ,
    \new_[12365]_ , \new_[12368]_ , \new_[12372]_ , \new_[12373]_ ,
    \new_[12374]_ , \new_[12378]_ , \new_[12379]_ , \new_[12383]_ ,
    \new_[12384]_ , \new_[12385]_ , \new_[12388]_ , \new_[12392]_ ,
    \new_[12393]_ , \new_[12394]_ , \new_[12398]_ , \new_[12399]_ ,
    \new_[12403]_ , \new_[12404]_ , \new_[12405]_ , \new_[12408]_ ,
    \new_[12412]_ , \new_[12413]_ , \new_[12414]_ , \new_[12418]_ ,
    \new_[12419]_ , \new_[12423]_ , \new_[12424]_ , \new_[12425]_ ,
    \new_[12428]_ , \new_[12432]_ , \new_[12433]_ , \new_[12434]_ ,
    \new_[12438]_ , \new_[12439]_ , \new_[12443]_ , \new_[12444]_ ,
    \new_[12445]_ , \new_[12448]_ , \new_[12452]_ , \new_[12453]_ ,
    \new_[12454]_ , \new_[12458]_ , \new_[12459]_ , \new_[12463]_ ,
    \new_[12464]_ , \new_[12465]_ , \new_[12468]_ , \new_[12472]_ ,
    \new_[12473]_ , \new_[12474]_ , \new_[12478]_ , \new_[12479]_ ,
    \new_[12483]_ , \new_[12484]_ , \new_[12485]_ , \new_[12488]_ ,
    \new_[12492]_ , \new_[12493]_ , \new_[12494]_ , \new_[12498]_ ,
    \new_[12499]_ , \new_[12503]_ , \new_[12504]_ , \new_[12505]_ ,
    \new_[12508]_ , \new_[12512]_ , \new_[12513]_ , \new_[12514]_ ,
    \new_[12518]_ , \new_[12519]_ , \new_[12523]_ , \new_[12524]_ ,
    \new_[12525]_ , \new_[12528]_ , \new_[12532]_ , \new_[12533]_ ,
    \new_[12534]_ , \new_[12538]_ , \new_[12539]_ , \new_[12543]_ ,
    \new_[12544]_ , \new_[12545]_ , \new_[12548]_ , \new_[12552]_ ,
    \new_[12553]_ , \new_[12554]_ , \new_[12558]_ , \new_[12559]_ ,
    \new_[12563]_ , \new_[12564]_ , \new_[12565]_ , \new_[12568]_ ,
    \new_[12572]_ , \new_[12573]_ , \new_[12574]_ , \new_[12578]_ ,
    \new_[12579]_ , \new_[12583]_ , \new_[12584]_ , \new_[12585]_ ,
    \new_[12588]_ , \new_[12592]_ , \new_[12593]_ , \new_[12594]_ ,
    \new_[12598]_ , \new_[12599]_ , \new_[12603]_ , \new_[12604]_ ,
    \new_[12605]_ , \new_[12608]_ , \new_[12612]_ , \new_[12613]_ ,
    \new_[12614]_ , \new_[12618]_ , \new_[12619]_ , \new_[12623]_ ,
    \new_[12624]_ , \new_[12625]_ , \new_[12628]_ , \new_[12632]_ ,
    \new_[12633]_ , \new_[12634]_ , \new_[12638]_ , \new_[12639]_ ,
    \new_[12643]_ , \new_[12644]_ , \new_[12645]_ , \new_[12648]_ ,
    \new_[12652]_ , \new_[12653]_ , \new_[12654]_ , \new_[12658]_ ,
    \new_[12659]_ , \new_[12663]_ , \new_[12664]_ , \new_[12665]_ ,
    \new_[12668]_ , \new_[12672]_ , \new_[12673]_ , \new_[12674]_ ,
    \new_[12678]_ , \new_[12679]_ , \new_[12683]_ , \new_[12684]_ ,
    \new_[12685]_ , \new_[12688]_ , \new_[12692]_ , \new_[12693]_ ,
    \new_[12694]_ , \new_[12698]_ , \new_[12699]_ , \new_[12703]_ ,
    \new_[12704]_ , \new_[12705]_ , \new_[12708]_ , \new_[12712]_ ,
    \new_[12713]_ , \new_[12714]_ , \new_[12718]_ , \new_[12719]_ ,
    \new_[12723]_ , \new_[12724]_ , \new_[12725]_ , \new_[12728]_ ,
    \new_[12732]_ , \new_[12733]_ , \new_[12734]_ , \new_[12738]_ ,
    \new_[12739]_ , \new_[12743]_ , \new_[12744]_ , \new_[12745]_ ,
    \new_[12748]_ , \new_[12752]_ , \new_[12753]_ , \new_[12754]_ ,
    \new_[12758]_ , \new_[12759]_ , \new_[12763]_ , \new_[12764]_ ,
    \new_[12765]_ , \new_[12768]_ , \new_[12772]_ , \new_[12773]_ ,
    \new_[12774]_ , \new_[12778]_ , \new_[12779]_ , \new_[12783]_ ,
    \new_[12784]_ , \new_[12785]_ , \new_[12788]_ , \new_[12792]_ ,
    \new_[12793]_ , \new_[12794]_ , \new_[12798]_ , \new_[12799]_ ,
    \new_[12803]_ , \new_[12804]_ , \new_[12805]_ , \new_[12808]_ ,
    \new_[12812]_ , \new_[12813]_ , \new_[12814]_ , \new_[12818]_ ,
    \new_[12819]_ , \new_[12823]_ , \new_[12824]_ , \new_[12825]_ ,
    \new_[12828]_ , \new_[12832]_ , \new_[12833]_ , \new_[12834]_ ,
    \new_[12838]_ , \new_[12839]_ , \new_[12843]_ , \new_[12844]_ ,
    \new_[12845]_ , \new_[12848]_ , \new_[12852]_ , \new_[12853]_ ,
    \new_[12854]_ , \new_[12858]_ , \new_[12859]_ , \new_[12863]_ ,
    \new_[12864]_ , \new_[12865]_ , \new_[12868]_ , \new_[12872]_ ,
    \new_[12873]_ , \new_[12874]_ , \new_[12878]_ , \new_[12879]_ ,
    \new_[12883]_ , \new_[12884]_ , \new_[12885]_ , \new_[12888]_ ,
    \new_[12892]_ , \new_[12893]_ , \new_[12894]_ , \new_[12898]_ ,
    \new_[12899]_ , \new_[12903]_ , \new_[12904]_ , \new_[12905]_ ,
    \new_[12908]_ , \new_[12912]_ , \new_[12913]_ , \new_[12914]_ ,
    \new_[12918]_ , \new_[12919]_ , \new_[12923]_ , \new_[12924]_ ,
    \new_[12925]_ , \new_[12928]_ , \new_[12932]_ , \new_[12933]_ ,
    \new_[12934]_ , \new_[12938]_ , \new_[12939]_ , \new_[12943]_ ,
    \new_[12944]_ , \new_[12945]_ , \new_[12948]_ , \new_[12952]_ ,
    \new_[12953]_ , \new_[12954]_ , \new_[12958]_ , \new_[12959]_ ,
    \new_[12963]_ , \new_[12964]_ , \new_[12965]_ , \new_[12968]_ ,
    \new_[12972]_ , \new_[12973]_ , \new_[12974]_ , \new_[12978]_ ,
    \new_[12979]_ , \new_[12983]_ , \new_[12984]_ , \new_[12985]_ ,
    \new_[12988]_ , \new_[12992]_ , \new_[12993]_ , \new_[12994]_ ,
    \new_[12998]_ , \new_[12999]_ , \new_[13003]_ , \new_[13004]_ ,
    \new_[13005]_ , \new_[13008]_ , \new_[13012]_ , \new_[13013]_ ,
    \new_[13014]_ , \new_[13018]_ , \new_[13019]_ , \new_[13023]_ ,
    \new_[13024]_ , \new_[13025]_ , \new_[13028]_ , \new_[13032]_ ,
    \new_[13033]_ , \new_[13034]_ , \new_[13038]_ , \new_[13039]_ ,
    \new_[13043]_ , \new_[13044]_ , \new_[13045]_ , \new_[13048]_ ,
    \new_[13052]_ , \new_[13053]_ , \new_[13054]_ , \new_[13058]_ ,
    \new_[13059]_ , \new_[13063]_ , \new_[13064]_ , \new_[13065]_ ,
    \new_[13068]_ , \new_[13072]_ , \new_[13073]_ , \new_[13074]_ ,
    \new_[13078]_ , \new_[13079]_ , \new_[13083]_ , \new_[13084]_ ,
    \new_[13085]_ , \new_[13088]_ , \new_[13092]_ , \new_[13093]_ ,
    \new_[13094]_ , \new_[13098]_ , \new_[13099]_ , \new_[13103]_ ,
    \new_[13104]_ , \new_[13105]_ , \new_[13108]_ , \new_[13112]_ ,
    \new_[13113]_ , \new_[13114]_ , \new_[13118]_ , \new_[13119]_ ,
    \new_[13123]_ , \new_[13124]_ , \new_[13125]_ , \new_[13128]_ ,
    \new_[13132]_ , \new_[13133]_ , \new_[13134]_ , \new_[13138]_ ,
    \new_[13139]_ , \new_[13143]_ , \new_[13144]_ , \new_[13145]_ ,
    \new_[13148]_ , \new_[13152]_ , \new_[13153]_ , \new_[13154]_ ,
    \new_[13158]_ , \new_[13159]_ , \new_[13163]_ , \new_[13164]_ ,
    \new_[13165]_ , \new_[13168]_ , \new_[13172]_ , \new_[13173]_ ,
    \new_[13174]_ , \new_[13178]_ , \new_[13179]_ , \new_[13183]_ ,
    \new_[13184]_ , \new_[13185]_ , \new_[13188]_ , \new_[13192]_ ,
    \new_[13193]_ , \new_[13194]_ , \new_[13198]_ , \new_[13199]_ ,
    \new_[13203]_ , \new_[13204]_ , \new_[13205]_ , \new_[13208]_ ,
    \new_[13212]_ , \new_[13213]_ , \new_[13214]_ , \new_[13218]_ ,
    \new_[13219]_ , \new_[13223]_ , \new_[13224]_ , \new_[13225]_ ,
    \new_[13228]_ , \new_[13232]_ , \new_[13233]_ , \new_[13234]_ ,
    \new_[13238]_ , \new_[13239]_ , \new_[13243]_ , \new_[13244]_ ,
    \new_[13245]_ , \new_[13248]_ , \new_[13252]_ , \new_[13253]_ ,
    \new_[13254]_ , \new_[13258]_ , \new_[13259]_ , \new_[13263]_ ,
    \new_[13264]_ , \new_[13265]_ , \new_[13268]_ , \new_[13272]_ ,
    \new_[13273]_ , \new_[13274]_ , \new_[13278]_ , \new_[13279]_ ,
    \new_[13283]_ , \new_[13284]_ , \new_[13285]_ , \new_[13288]_ ,
    \new_[13292]_ , \new_[13293]_ , \new_[13294]_ , \new_[13298]_ ,
    \new_[13299]_ , \new_[13303]_ , \new_[13304]_ , \new_[13305]_ ,
    \new_[13308]_ , \new_[13312]_ , \new_[13313]_ , \new_[13314]_ ,
    \new_[13318]_ , \new_[13319]_ , \new_[13323]_ , \new_[13324]_ ,
    \new_[13325]_ , \new_[13328]_ , \new_[13332]_ , \new_[13333]_ ,
    \new_[13334]_ , \new_[13338]_ , \new_[13339]_ , \new_[13343]_ ,
    \new_[13344]_ , \new_[13345]_ , \new_[13348]_ , \new_[13352]_ ,
    \new_[13353]_ , \new_[13354]_ , \new_[13358]_ , \new_[13359]_ ,
    \new_[13363]_ , \new_[13364]_ , \new_[13365]_ , \new_[13368]_ ,
    \new_[13372]_ , \new_[13373]_ , \new_[13374]_ , \new_[13378]_ ,
    \new_[13379]_ , \new_[13383]_ , \new_[13384]_ , \new_[13385]_ ,
    \new_[13388]_ , \new_[13392]_ , \new_[13393]_ , \new_[13394]_ ,
    \new_[13398]_ , \new_[13399]_ , \new_[13403]_ , \new_[13404]_ ,
    \new_[13405]_ , \new_[13408]_ , \new_[13412]_ , \new_[13413]_ ,
    \new_[13414]_ , \new_[13418]_ , \new_[13419]_ , \new_[13423]_ ,
    \new_[13424]_ , \new_[13425]_ , \new_[13428]_ , \new_[13432]_ ,
    \new_[13433]_ , \new_[13434]_ , \new_[13438]_ , \new_[13439]_ ,
    \new_[13443]_ , \new_[13444]_ , \new_[13445]_ , \new_[13448]_ ,
    \new_[13452]_ , \new_[13453]_ , \new_[13454]_ , \new_[13458]_ ,
    \new_[13459]_ , \new_[13463]_ , \new_[13464]_ , \new_[13465]_ ,
    \new_[13468]_ , \new_[13472]_ , \new_[13473]_ , \new_[13474]_ ,
    \new_[13478]_ , \new_[13479]_ , \new_[13483]_ , \new_[13484]_ ,
    \new_[13485]_ , \new_[13488]_ , \new_[13492]_ , \new_[13493]_ ,
    \new_[13494]_ , \new_[13498]_ , \new_[13499]_ , \new_[13503]_ ,
    \new_[13504]_ , \new_[13505]_ , \new_[13508]_ , \new_[13512]_ ,
    \new_[13513]_ , \new_[13514]_ , \new_[13518]_ , \new_[13519]_ ,
    \new_[13523]_ , \new_[13524]_ , \new_[13525]_ , \new_[13528]_ ,
    \new_[13532]_ , \new_[13533]_ , \new_[13534]_ , \new_[13538]_ ,
    \new_[13539]_ , \new_[13543]_ , \new_[13544]_ , \new_[13545]_ ,
    \new_[13548]_ , \new_[13552]_ , \new_[13553]_ , \new_[13554]_ ,
    \new_[13558]_ , \new_[13559]_ , \new_[13563]_ , \new_[13564]_ ,
    \new_[13565]_ , \new_[13568]_ , \new_[13572]_ , \new_[13573]_ ,
    \new_[13574]_ , \new_[13578]_ , \new_[13579]_ , \new_[13583]_ ,
    \new_[13584]_ , \new_[13585]_ , \new_[13588]_ , \new_[13592]_ ,
    \new_[13593]_ , \new_[13594]_ , \new_[13598]_ , \new_[13599]_ ,
    \new_[13603]_ , \new_[13604]_ , \new_[13605]_ , \new_[13608]_ ,
    \new_[13612]_ , \new_[13613]_ , \new_[13614]_ , \new_[13618]_ ,
    \new_[13619]_ , \new_[13623]_ , \new_[13624]_ , \new_[13625]_ ,
    \new_[13628]_ , \new_[13632]_ , \new_[13633]_ , \new_[13634]_ ,
    \new_[13638]_ , \new_[13639]_ , \new_[13643]_ , \new_[13644]_ ,
    \new_[13645]_ , \new_[13648]_ , \new_[13652]_ , \new_[13653]_ ,
    \new_[13654]_ , \new_[13658]_ , \new_[13659]_ , \new_[13663]_ ,
    \new_[13664]_ , \new_[13665]_ , \new_[13668]_ , \new_[13672]_ ,
    \new_[13673]_ , \new_[13674]_ , \new_[13678]_ , \new_[13679]_ ,
    \new_[13683]_ , \new_[13684]_ , \new_[13685]_ , \new_[13689]_ ,
    \new_[13690]_ , \new_[13694]_ , \new_[13695]_ , \new_[13696]_ ,
    \new_[13700]_ , \new_[13701]_ , \new_[13705]_ , \new_[13706]_ ,
    \new_[13707]_ , \new_[13711]_ , \new_[13712]_ , \new_[13716]_ ,
    \new_[13717]_ , \new_[13718]_ , \new_[13722]_ , \new_[13723]_ ,
    \new_[13727]_ , \new_[13728]_ , \new_[13729]_ , \new_[13733]_ ,
    \new_[13734]_ , \new_[13738]_ , \new_[13739]_ , \new_[13740]_ ,
    \new_[13744]_ , \new_[13745]_ , \new_[13749]_ , \new_[13750]_ ,
    \new_[13751]_ , \new_[13755]_ , \new_[13756]_ , \new_[13760]_ ,
    \new_[13761]_ , \new_[13762]_ , \new_[13766]_ , \new_[13767]_ ,
    \new_[13771]_ , \new_[13772]_ , \new_[13773]_ , \new_[13777]_ ,
    \new_[13778]_ , \new_[13782]_ , \new_[13783]_ , \new_[13784]_ ,
    \new_[13788]_ , \new_[13789]_ , \new_[13793]_ , \new_[13794]_ ,
    \new_[13795]_ , \new_[13799]_ , \new_[13800]_ , \new_[13804]_ ,
    \new_[13805]_ , \new_[13806]_ , \new_[13810]_ , \new_[13811]_ ,
    \new_[13815]_ , \new_[13816]_ , \new_[13817]_ , \new_[13821]_ ,
    \new_[13822]_ , \new_[13826]_ , \new_[13827]_ , \new_[13828]_ ,
    \new_[13832]_ , \new_[13833]_ , \new_[13837]_ , \new_[13838]_ ,
    \new_[13839]_ , \new_[13843]_ , \new_[13844]_ , \new_[13848]_ ,
    \new_[13849]_ , \new_[13850]_ , \new_[13854]_ , \new_[13855]_ ,
    \new_[13859]_ , \new_[13860]_ , \new_[13861]_ , \new_[13865]_ ,
    \new_[13866]_ , \new_[13870]_ , \new_[13871]_ , \new_[13872]_ ,
    \new_[13876]_ , \new_[13877]_ , \new_[13881]_ , \new_[13882]_ ,
    \new_[13883]_ , \new_[13887]_ , \new_[13888]_ , \new_[13892]_ ,
    \new_[13893]_ , \new_[13894]_ , \new_[13898]_ , \new_[13899]_ ,
    \new_[13903]_ , \new_[13904]_ , \new_[13905]_ , \new_[13909]_ ,
    \new_[13910]_ , \new_[13914]_ , \new_[13915]_ , \new_[13916]_ ,
    \new_[13920]_ , \new_[13921]_ , \new_[13925]_ , \new_[13926]_ ,
    \new_[13927]_ , \new_[13931]_ , \new_[13932]_ , \new_[13936]_ ,
    \new_[13937]_ , \new_[13938]_ , \new_[13942]_ , \new_[13943]_ ,
    \new_[13947]_ , \new_[13948]_ , \new_[13949]_ , \new_[13953]_ ,
    \new_[13954]_ , \new_[13958]_ , \new_[13959]_ , \new_[13960]_ ,
    \new_[13964]_ , \new_[13965]_ , \new_[13969]_ , \new_[13970]_ ,
    \new_[13971]_ , \new_[13975]_ , \new_[13976]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13982]_ , \new_[13986]_ , \new_[13987]_ ,
    \new_[13991]_ , \new_[13992]_ , \new_[13993]_ , \new_[13997]_ ,
    \new_[13998]_ , \new_[14002]_ , \new_[14003]_ , \new_[14004]_ ,
    \new_[14008]_ , \new_[14009]_ , \new_[14013]_ , \new_[14014]_ ,
    \new_[14015]_ , \new_[14019]_ , \new_[14020]_ , \new_[14024]_ ,
    \new_[14025]_ , \new_[14026]_ , \new_[14030]_ , \new_[14031]_ ,
    \new_[14035]_ , \new_[14036]_ , \new_[14037]_ , \new_[14041]_ ,
    \new_[14042]_ , \new_[14046]_ , \new_[14047]_ , \new_[14048]_ ,
    \new_[14052]_ , \new_[14053]_ , \new_[14057]_ , \new_[14058]_ ,
    \new_[14059]_ , \new_[14063]_ , \new_[14064]_ , \new_[14068]_ ,
    \new_[14069]_ , \new_[14070]_ , \new_[14074]_ , \new_[14075]_ ,
    \new_[14079]_ , \new_[14080]_ , \new_[14081]_ , \new_[14085]_ ,
    \new_[14086]_ , \new_[14090]_ , \new_[14091]_ , \new_[14092]_ ,
    \new_[14096]_ , \new_[14097]_ , \new_[14101]_ , \new_[14102]_ ,
    \new_[14103]_ , \new_[14107]_ , \new_[14108]_ , \new_[14112]_ ,
    \new_[14113]_ , \new_[14114]_ , \new_[14118]_ , \new_[14119]_ ,
    \new_[14123]_ , \new_[14124]_ , \new_[14125]_ , \new_[14129]_ ,
    \new_[14130]_ , \new_[14134]_ , \new_[14135]_ , \new_[14136]_ ,
    \new_[14140]_ , \new_[14141]_ , \new_[14145]_ , \new_[14146]_ ,
    \new_[14147]_ , \new_[14151]_ , \new_[14152]_ , \new_[14156]_ ,
    \new_[14157]_ , \new_[14158]_ , \new_[14162]_ , \new_[14163]_ ,
    \new_[14167]_ , \new_[14168]_ , \new_[14169]_ , \new_[14173]_ ,
    \new_[14174]_ , \new_[14178]_ , \new_[14179]_ , \new_[14180]_ ,
    \new_[14184]_ , \new_[14185]_ , \new_[14189]_ , \new_[14190]_ ,
    \new_[14191]_ , \new_[14195]_ , \new_[14196]_ , \new_[14200]_ ,
    \new_[14201]_ , \new_[14202]_ , \new_[14206]_ , \new_[14207]_ ,
    \new_[14211]_ , \new_[14212]_ , \new_[14213]_ , \new_[14217]_ ,
    \new_[14218]_ , \new_[14222]_ , \new_[14223]_ , \new_[14224]_ ,
    \new_[14228]_ , \new_[14229]_ , \new_[14233]_ , \new_[14234]_ ,
    \new_[14235]_ , \new_[14239]_ , \new_[14240]_ , \new_[14244]_ ,
    \new_[14245]_ , \new_[14246]_ , \new_[14250]_ , \new_[14251]_ ,
    \new_[14255]_ , \new_[14256]_ , \new_[14257]_ , \new_[14261]_ ,
    \new_[14262]_ , \new_[14266]_ , \new_[14267]_ , \new_[14268]_ ,
    \new_[14272]_ , \new_[14273]_ , \new_[14277]_ , \new_[14278]_ ,
    \new_[14279]_ , \new_[14283]_ , \new_[14284]_ , \new_[14288]_ ,
    \new_[14289]_ , \new_[14290]_ , \new_[14294]_ , \new_[14295]_ ,
    \new_[14299]_ , \new_[14300]_ , \new_[14301]_ , \new_[14305]_ ,
    \new_[14306]_ , \new_[14310]_ , \new_[14311]_ , \new_[14312]_ ,
    \new_[14316]_ , \new_[14317]_ , \new_[14321]_ , \new_[14322]_ ,
    \new_[14323]_ , \new_[14327]_ , \new_[14328]_ , \new_[14332]_ ,
    \new_[14333]_ , \new_[14334]_ , \new_[14338]_ , \new_[14339]_ ,
    \new_[14343]_ , \new_[14344]_ , \new_[14345]_ , \new_[14349]_ ,
    \new_[14350]_ , \new_[14354]_ , \new_[14355]_ , \new_[14356]_ ,
    \new_[14360]_ , \new_[14361]_ , \new_[14365]_ , \new_[14366]_ ,
    \new_[14367]_ , \new_[14371]_ , \new_[14372]_ , \new_[14376]_ ,
    \new_[14377]_ , \new_[14378]_ , \new_[14382]_ , \new_[14383]_ ,
    \new_[14387]_ , \new_[14388]_ , \new_[14389]_ , \new_[14393]_ ,
    \new_[14394]_ , \new_[14398]_ , \new_[14399]_ , \new_[14400]_ ,
    \new_[14404]_ , \new_[14405]_ , \new_[14409]_ , \new_[14410]_ ,
    \new_[14411]_ , \new_[14415]_ , \new_[14416]_ , \new_[14420]_ ,
    \new_[14421]_ , \new_[14422]_ , \new_[14426]_ , \new_[14427]_ ,
    \new_[14431]_ , \new_[14432]_ , \new_[14433]_ , \new_[14437]_ ,
    \new_[14438]_ , \new_[14442]_ , \new_[14443]_ , \new_[14444]_ ,
    \new_[14448]_ , \new_[14449]_ , \new_[14453]_ , \new_[14454]_ ,
    \new_[14455]_ , \new_[14459]_ , \new_[14460]_ , \new_[14464]_ ,
    \new_[14465]_ , \new_[14466]_ , \new_[14470]_ , \new_[14471]_ ,
    \new_[14475]_ , \new_[14476]_ , \new_[14477]_ , \new_[14481]_ ,
    \new_[14482]_ , \new_[14486]_ , \new_[14487]_ , \new_[14488]_ ,
    \new_[14492]_ , \new_[14493]_ , \new_[14497]_ , \new_[14498]_ ,
    \new_[14499]_ , \new_[14503]_ , \new_[14504]_ , \new_[14508]_ ,
    \new_[14509]_ , \new_[14510]_ , \new_[14514]_ , \new_[14515]_ ,
    \new_[14519]_ , \new_[14520]_ , \new_[14521]_ , \new_[14525]_ ,
    \new_[14526]_ , \new_[14530]_ , \new_[14531]_ , \new_[14532]_ ,
    \new_[14536]_ , \new_[14537]_ , \new_[14541]_ , \new_[14542]_ ,
    \new_[14543]_ , \new_[14547]_ , \new_[14548]_ , \new_[14552]_ ,
    \new_[14553]_ , \new_[14554]_ , \new_[14558]_ , \new_[14559]_ ,
    \new_[14563]_ , \new_[14564]_ , \new_[14565]_ , \new_[14569]_ ,
    \new_[14570]_ , \new_[14574]_ , \new_[14575]_ , \new_[14576]_ ,
    \new_[14580]_ , \new_[14581]_ , \new_[14585]_ , \new_[14586]_ ,
    \new_[14587]_ , \new_[14591]_ , \new_[14592]_ , \new_[14596]_ ,
    \new_[14597]_ , \new_[14598]_ , \new_[14602]_ , \new_[14603]_ ,
    \new_[14607]_ , \new_[14608]_ , \new_[14609]_ , \new_[14613]_ ,
    \new_[14614]_ , \new_[14618]_ , \new_[14619]_ , \new_[14620]_ ,
    \new_[14624]_ , \new_[14625]_ , \new_[14629]_ , \new_[14630]_ ,
    \new_[14631]_ , \new_[14635]_ , \new_[14636]_ , \new_[14640]_ ,
    \new_[14641]_ , \new_[14642]_ , \new_[14646]_ , \new_[14647]_ ,
    \new_[14651]_ , \new_[14652]_ , \new_[14653]_ , \new_[14657]_ ,
    \new_[14658]_ , \new_[14662]_ , \new_[14663]_ , \new_[14664]_ ,
    \new_[14668]_ , \new_[14669]_ , \new_[14673]_ , \new_[14674]_ ,
    \new_[14675]_ , \new_[14679]_ , \new_[14680]_ , \new_[14684]_ ,
    \new_[14685]_ , \new_[14686]_ , \new_[14690]_ , \new_[14691]_ ,
    \new_[14695]_ , \new_[14696]_ , \new_[14697]_ , \new_[14701]_ ,
    \new_[14702]_ , \new_[14706]_ , \new_[14707]_ , \new_[14708]_ ,
    \new_[14712]_ , \new_[14713]_ , \new_[14717]_ , \new_[14718]_ ,
    \new_[14719]_ , \new_[14723]_ , \new_[14724]_ , \new_[14728]_ ,
    \new_[14729]_ , \new_[14730]_ , \new_[14734]_ , \new_[14735]_ ,
    \new_[14739]_ , \new_[14740]_ , \new_[14741]_ , \new_[14745]_ ,
    \new_[14746]_ , \new_[14750]_ , \new_[14751]_ , \new_[14752]_ ,
    \new_[14756]_ , \new_[14757]_ , \new_[14761]_ , \new_[14762]_ ,
    \new_[14763]_ , \new_[14767]_ , \new_[14768]_ , \new_[14772]_ ,
    \new_[14773]_ , \new_[14774]_ , \new_[14778]_ , \new_[14779]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14785]_ , \new_[14789]_ ,
    \new_[14790]_ , \new_[14794]_ , \new_[14795]_ , \new_[14796]_ ,
    \new_[14800]_ , \new_[14801]_ , \new_[14805]_ , \new_[14806]_ ,
    \new_[14807]_ , \new_[14811]_ , \new_[14812]_ , \new_[14816]_ ,
    \new_[14817]_ , \new_[14818]_ , \new_[14822]_ , \new_[14823]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14829]_ , \new_[14833]_ ,
    \new_[14834]_ , \new_[14838]_ , \new_[14839]_ , \new_[14840]_ ,
    \new_[14844]_ , \new_[14845]_ , \new_[14849]_ , \new_[14850]_ ,
    \new_[14851]_ , \new_[14855]_ , \new_[14856]_ , \new_[14860]_ ,
    \new_[14861]_ , \new_[14862]_ , \new_[14866]_ , \new_[14867]_ ,
    \new_[14871]_ , \new_[14872]_ , \new_[14873]_ , \new_[14877]_ ,
    \new_[14878]_ , \new_[14882]_ , \new_[14883]_ , \new_[14884]_ ,
    \new_[14888]_ , \new_[14889]_ , \new_[14893]_ , \new_[14894]_ ,
    \new_[14895]_ , \new_[14899]_ , \new_[14900]_ , \new_[14904]_ ,
    \new_[14905]_ , \new_[14906]_ , \new_[14910]_ , \new_[14911]_ ,
    \new_[14915]_ , \new_[14916]_ , \new_[14917]_ , \new_[14921]_ ,
    \new_[14922]_ , \new_[14926]_ , \new_[14927]_ , \new_[14928]_ ,
    \new_[14932]_ , \new_[14933]_ , \new_[14937]_ , \new_[14938]_ ,
    \new_[14939]_ , \new_[14943]_ , \new_[14944]_ , \new_[14948]_ ,
    \new_[14949]_ , \new_[14950]_ , \new_[14954]_ , \new_[14955]_ ,
    \new_[14959]_ , \new_[14960]_ , \new_[14961]_ , \new_[14965]_ ,
    \new_[14966]_ , \new_[14970]_ , \new_[14971]_ , \new_[14972]_ ,
    \new_[14976]_ , \new_[14977]_ , \new_[14981]_ , \new_[14982]_ ,
    \new_[14983]_ , \new_[14987]_ , \new_[14988]_ , \new_[14992]_ ,
    \new_[14993]_ , \new_[14994]_ , \new_[14998]_ , \new_[14999]_ ,
    \new_[15003]_ , \new_[15004]_ , \new_[15005]_ , \new_[15009]_ ,
    \new_[15010]_ , \new_[15014]_ , \new_[15015]_ , \new_[15016]_ ,
    \new_[15020]_ , \new_[15021]_ , \new_[15025]_ , \new_[15026]_ ,
    \new_[15027]_ , \new_[15031]_ , \new_[15032]_ , \new_[15036]_ ,
    \new_[15037]_ , \new_[15038]_ , \new_[15042]_ , \new_[15043]_ ,
    \new_[15047]_ , \new_[15048]_ , \new_[15049]_ , \new_[15053]_ ,
    \new_[15054]_ , \new_[15058]_ , \new_[15059]_ , \new_[15060]_ ,
    \new_[15064]_ , \new_[15065]_ , \new_[15069]_ , \new_[15070]_ ,
    \new_[15071]_ , \new_[15075]_ , \new_[15076]_ , \new_[15080]_ ,
    \new_[15081]_ , \new_[15082]_ , \new_[15086]_ , \new_[15087]_ ,
    \new_[15091]_ , \new_[15092]_ , \new_[15093]_ , \new_[15097]_ ,
    \new_[15098]_ , \new_[15102]_ , \new_[15103]_ , \new_[15104]_ ,
    \new_[15108]_ , \new_[15109]_ , \new_[15113]_ , \new_[15114]_ ,
    \new_[15115]_ , \new_[15119]_ , \new_[15120]_ , \new_[15124]_ ,
    \new_[15125]_ , \new_[15126]_ , \new_[15130]_ , \new_[15131]_ ,
    \new_[15135]_ , \new_[15136]_ , \new_[15137]_ , \new_[15141]_ ,
    \new_[15142]_ , \new_[15146]_ , \new_[15147]_ , \new_[15148]_ ,
    \new_[15152]_ , \new_[15153]_ , \new_[15157]_ , \new_[15158]_ ,
    \new_[15159]_ , \new_[15163]_ , \new_[15164]_ , \new_[15168]_ ,
    \new_[15169]_ , \new_[15170]_ , \new_[15174]_ , \new_[15175]_ ,
    \new_[15179]_ , \new_[15180]_ , \new_[15181]_ , \new_[15185]_ ,
    \new_[15186]_ , \new_[15190]_ , \new_[15191]_ , \new_[15192]_ ,
    \new_[15196]_ , \new_[15197]_ , \new_[15201]_ , \new_[15202]_ ,
    \new_[15203]_ , \new_[15207]_ , \new_[15208]_ , \new_[15212]_ ,
    \new_[15213]_ , \new_[15214]_ , \new_[15218]_ , \new_[15219]_ ,
    \new_[15223]_ , \new_[15224]_ , \new_[15225]_ , \new_[15229]_ ,
    \new_[15230]_ , \new_[15234]_ , \new_[15235]_ , \new_[15236]_ ,
    \new_[15240]_ , \new_[15241]_ , \new_[15245]_ , \new_[15246]_ ,
    \new_[15247]_ , \new_[15251]_ , \new_[15252]_ , \new_[15256]_ ,
    \new_[15257]_ , \new_[15258]_ , \new_[15262]_ , \new_[15263]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15269]_ , \new_[15273]_ ,
    \new_[15274]_ , \new_[15278]_ , \new_[15279]_ , \new_[15280]_ ,
    \new_[15284]_ , \new_[15285]_ , \new_[15289]_ , \new_[15290]_ ,
    \new_[15291]_ , \new_[15295]_ , \new_[15296]_ , \new_[15300]_ ,
    \new_[15301]_ , \new_[15302]_ , \new_[15306]_ , \new_[15307]_ ,
    \new_[15311]_ , \new_[15312]_ , \new_[15313]_ , \new_[15317]_ ,
    \new_[15318]_ , \new_[15322]_ , \new_[15323]_ , \new_[15324]_ ,
    \new_[15328]_ , \new_[15329]_ , \new_[15333]_ , \new_[15334]_ ,
    \new_[15335]_ , \new_[15339]_ , \new_[15340]_ , \new_[15344]_ ,
    \new_[15345]_ , \new_[15346]_ , \new_[15350]_ , \new_[15351]_ ,
    \new_[15355]_ , \new_[15356]_ , \new_[15357]_ , \new_[15361]_ ,
    \new_[15362]_ , \new_[15366]_ , \new_[15367]_ , \new_[15368]_ ,
    \new_[15372]_ , \new_[15373]_ , \new_[15377]_ , \new_[15378]_ ,
    \new_[15379]_ , \new_[15383]_ , \new_[15384]_ , \new_[15388]_ ,
    \new_[15389]_ , \new_[15390]_ , \new_[15394]_ , \new_[15395]_ ,
    \new_[15399]_ , \new_[15400]_ , \new_[15401]_ , \new_[15405]_ ,
    \new_[15406]_ , \new_[15410]_ , \new_[15411]_ , \new_[15412]_ ,
    \new_[15416]_ , \new_[15417]_ , \new_[15421]_ , \new_[15422]_ ,
    \new_[15423]_ , \new_[15427]_ , \new_[15428]_ , \new_[15432]_ ,
    \new_[15433]_ , \new_[15434]_ , \new_[15438]_ , \new_[15439]_ ,
    \new_[15443]_ , \new_[15444]_ , \new_[15445]_ , \new_[15449]_ ,
    \new_[15450]_ , \new_[15454]_ , \new_[15455]_ , \new_[15456]_ ,
    \new_[15460]_ , \new_[15461]_ , \new_[15464]_ , \new_[15467]_ ,
    \new_[15468]_ , \new_[15469]_ , \new_[15473]_ , \new_[15474]_ ,
    \new_[15478]_ , \new_[15479]_ , \new_[15480]_ , \new_[15484]_ ,
    \new_[15485]_ , \new_[15488]_ , \new_[15491]_ , \new_[15492]_ ,
    \new_[15493]_ , \new_[15497]_ , \new_[15498]_ , \new_[15502]_ ,
    \new_[15503]_ , \new_[15504]_ , \new_[15508]_ , \new_[15509]_ ,
    \new_[15512]_ , \new_[15515]_ , \new_[15516]_ , \new_[15517]_ ,
    \new_[15521]_ , \new_[15522]_ , \new_[15526]_ , \new_[15527]_ ,
    \new_[15528]_ , \new_[15532]_ , \new_[15533]_ , \new_[15536]_ ,
    \new_[15539]_ , \new_[15540]_ , \new_[15541]_ , \new_[15545]_ ,
    \new_[15546]_ , \new_[15550]_ , \new_[15551]_ , \new_[15552]_ ,
    \new_[15556]_ , \new_[15557]_ , \new_[15560]_ , \new_[15563]_ ,
    \new_[15564]_ , \new_[15565]_ , \new_[15569]_ , \new_[15570]_ ,
    \new_[15574]_ , \new_[15575]_ , \new_[15576]_ , \new_[15580]_ ,
    \new_[15581]_ , \new_[15584]_ , \new_[15587]_ , \new_[15588]_ ,
    \new_[15589]_ , \new_[15593]_ , \new_[15594]_ , \new_[15598]_ ,
    \new_[15599]_ , \new_[15600]_ , \new_[15604]_ , \new_[15605]_ ,
    \new_[15608]_ , \new_[15611]_ , \new_[15612]_ , \new_[15613]_ ,
    \new_[15617]_ , \new_[15618]_ , \new_[15622]_ , \new_[15623]_ ,
    \new_[15624]_ , \new_[15628]_ , \new_[15629]_ , \new_[15632]_ ,
    \new_[15635]_ , \new_[15636]_ , \new_[15637]_ , \new_[15641]_ ,
    \new_[15642]_ , \new_[15646]_ , \new_[15647]_ , \new_[15648]_ ,
    \new_[15652]_ , \new_[15653]_ , \new_[15656]_ , \new_[15659]_ ,
    \new_[15660]_ , \new_[15661]_ , \new_[15665]_ , \new_[15666]_ ,
    \new_[15670]_ , \new_[15671]_ , \new_[15672]_ , \new_[15676]_ ,
    \new_[15677]_ , \new_[15680]_ , \new_[15683]_ , \new_[15684]_ ,
    \new_[15685]_ , \new_[15689]_ , \new_[15690]_ , \new_[15694]_ ,
    \new_[15695]_ , \new_[15696]_ , \new_[15700]_ , \new_[15701]_ ,
    \new_[15704]_ , \new_[15707]_ , \new_[15708]_ , \new_[15709]_ ,
    \new_[15713]_ , \new_[15714]_ , \new_[15718]_ , \new_[15719]_ ,
    \new_[15720]_ , \new_[15724]_ , \new_[15725]_ , \new_[15728]_ ,
    \new_[15731]_ , \new_[15732]_ , \new_[15733]_ , \new_[15737]_ ,
    \new_[15738]_ , \new_[15742]_ , \new_[15743]_ , \new_[15744]_ ,
    \new_[15748]_ , \new_[15749]_ , \new_[15752]_ , \new_[15755]_ ,
    \new_[15756]_ , \new_[15757]_ , \new_[15761]_ , \new_[15762]_ ,
    \new_[15766]_ , \new_[15767]_ , \new_[15768]_ , \new_[15772]_ ,
    \new_[15773]_ , \new_[15776]_ , \new_[15779]_ , \new_[15780]_ ,
    \new_[15781]_ , \new_[15785]_ , \new_[15786]_ , \new_[15790]_ ,
    \new_[15791]_ , \new_[15792]_ , \new_[15796]_ , \new_[15797]_ ,
    \new_[15800]_ , \new_[15803]_ , \new_[15804]_ , \new_[15805]_ ,
    \new_[15809]_ , \new_[15810]_ , \new_[15814]_ , \new_[15815]_ ,
    \new_[15816]_ , \new_[15820]_ , \new_[15821]_ , \new_[15824]_ ,
    \new_[15827]_ , \new_[15828]_ , \new_[15829]_ ;
  assign A75 = \new_[2293]_  | \new_[1528]_ ;
  assign \new_[1]_  = \new_[15829]_  & \new_[15816]_ ;
  assign \new_[2]_  = \new_[15805]_  & \new_[15792]_ ;
  assign \new_[3]_  = \new_[15781]_  & \new_[15768]_ ;
  assign \new_[4]_  = \new_[15757]_  & \new_[15744]_ ;
  assign \new_[5]_  = \new_[15733]_  & \new_[15720]_ ;
  assign \new_[6]_  = \new_[15709]_  & \new_[15696]_ ;
  assign \new_[7]_  = \new_[15685]_  & \new_[15672]_ ;
  assign \new_[8]_  = \new_[15661]_  & \new_[15648]_ ;
  assign \new_[9]_  = \new_[15637]_  & \new_[15624]_ ;
  assign \new_[10]_  = \new_[15613]_  & \new_[15600]_ ;
  assign \new_[11]_  = \new_[15589]_  & \new_[15576]_ ;
  assign \new_[12]_  = \new_[15565]_  & \new_[15552]_ ;
  assign \new_[13]_  = \new_[15541]_  & \new_[15528]_ ;
  assign \new_[14]_  = \new_[15517]_  & \new_[15504]_ ;
  assign \new_[15]_  = \new_[15493]_  & \new_[15480]_ ;
  assign \new_[16]_  = \new_[15469]_  & \new_[15456]_ ;
  assign \new_[17]_  = \new_[15445]_  & \new_[15434]_ ;
  assign \new_[18]_  = \new_[15423]_  & \new_[15412]_ ;
  assign \new_[19]_  = \new_[15401]_  & \new_[15390]_ ;
  assign \new_[20]_  = \new_[15379]_  & \new_[15368]_ ;
  assign \new_[21]_  = \new_[15357]_  & \new_[15346]_ ;
  assign \new_[22]_  = \new_[15335]_  & \new_[15324]_ ;
  assign \new_[23]_  = \new_[15313]_  & \new_[15302]_ ;
  assign \new_[24]_  = \new_[15291]_  & \new_[15280]_ ;
  assign \new_[25]_  = \new_[15269]_  & \new_[15258]_ ;
  assign \new_[26]_  = \new_[15247]_  & \new_[15236]_ ;
  assign \new_[27]_  = \new_[15225]_  & \new_[15214]_ ;
  assign \new_[28]_  = \new_[15203]_  & \new_[15192]_ ;
  assign \new_[29]_  = \new_[15181]_  & \new_[15170]_ ;
  assign \new_[30]_  = \new_[15159]_  & \new_[15148]_ ;
  assign \new_[31]_  = \new_[15137]_  & \new_[15126]_ ;
  assign \new_[32]_  = \new_[15115]_  & \new_[15104]_ ;
  assign \new_[33]_  = \new_[15093]_  & \new_[15082]_ ;
  assign \new_[34]_  = \new_[15071]_  & \new_[15060]_ ;
  assign \new_[35]_  = \new_[15049]_  & \new_[15038]_ ;
  assign \new_[36]_  = \new_[15027]_  & \new_[15016]_ ;
  assign \new_[37]_  = \new_[15005]_  & \new_[14994]_ ;
  assign \new_[38]_  = \new_[14983]_  & \new_[14972]_ ;
  assign \new_[39]_  = \new_[14961]_  & \new_[14950]_ ;
  assign \new_[40]_  = \new_[14939]_  & \new_[14928]_ ;
  assign \new_[41]_  = \new_[14917]_  & \new_[14906]_ ;
  assign \new_[42]_  = \new_[14895]_  & \new_[14884]_ ;
  assign \new_[43]_  = \new_[14873]_  & \new_[14862]_ ;
  assign \new_[44]_  = \new_[14851]_  & \new_[14840]_ ;
  assign \new_[45]_  = \new_[14829]_  & \new_[14818]_ ;
  assign \new_[46]_  = \new_[14807]_  & \new_[14796]_ ;
  assign \new_[47]_  = \new_[14785]_  & \new_[14774]_ ;
  assign \new_[48]_  = \new_[14763]_  & \new_[14752]_ ;
  assign \new_[49]_  = \new_[14741]_  & \new_[14730]_ ;
  assign \new_[50]_  = \new_[14719]_  & \new_[14708]_ ;
  assign \new_[51]_  = \new_[14697]_  & \new_[14686]_ ;
  assign \new_[52]_  = \new_[14675]_  & \new_[14664]_ ;
  assign \new_[53]_  = \new_[14653]_  & \new_[14642]_ ;
  assign \new_[54]_  = \new_[14631]_  & \new_[14620]_ ;
  assign \new_[55]_  = \new_[14609]_  & \new_[14598]_ ;
  assign \new_[56]_  = \new_[14587]_  & \new_[14576]_ ;
  assign \new_[57]_  = \new_[14565]_  & \new_[14554]_ ;
  assign \new_[58]_  = \new_[14543]_  & \new_[14532]_ ;
  assign \new_[59]_  = \new_[14521]_  & \new_[14510]_ ;
  assign \new_[60]_  = \new_[14499]_  & \new_[14488]_ ;
  assign \new_[61]_  = \new_[14477]_  & \new_[14466]_ ;
  assign \new_[62]_  = \new_[14455]_  & \new_[14444]_ ;
  assign \new_[63]_  = \new_[14433]_  & \new_[14422]_ ;
  assign \new_[64]_  = \new_[14411]_  & \new_[14400]_ ;
  assign \new_[65]_  = \new_[14389]_  & \new_[14378]_ ;
  assign \new_[66]_  = \new_[14367]_  & \new_[14356]_ ;
  assign \new_[67]_  = \new_[14345]_  & \new_[14334]_ ;
  assign \new_[68]_  = \new_[14323]_  & \new_[14312]_ ;
  assign \new_[69]_  = \new_[14301]_  & \new_[14290]_ ;
  assign \new_[70]_  = \new_[14279]_  & \new_[14268]_ ;
  assign \new_[71]_  = \new_[14257]_  & \new_[14246]_ ;
  assign \new_[72]_  = \new_[14235]_  & \new_[14224]_ ;
  assign \new_[73]_  = \new_[14213]_  & \new_[14202]_ ;
  assign \new_[74]_  = \new_[14191]_  & \new_[14180]_ ;
  assign \new_[75]_  = \new_[14169]_  & \new_[14158]_ ;
  assign \new_[76]_  = \new_[14147]_  & \new_[14136]_ ;
  assign \new_[77]_  = \new_[14125]_  & \new_[14114]_ ;
  assign \new_[78]_  = \new_[14103]_  & \new_[14092]_ ;
  assign \new_[79]_  = \new_[14081]_  & \new_[14070]_ ;
  assign \new_[80]_  = \new_[14059]_  & \new_[14048]_ ;
  assign \new_[81]_  = \new_[14037]_  & \new_[14026]_ ;
  assign \new_[82]_  = \new_[14015]_  & \new_[14004]_ ;
  assign \new_[83]_  = \new_[13993]_  & \new_[13982]_ ;
  assign \new_[84]_  = \new_[13971]_  & \new_[13960]_ ;
  assign \new_[85]_  = \new_[13949]_  & \new_[13938]_ ;
  assign \new_[86]_  = \new_[13927]_  & \new_[13916]_ ;
  assign \new_[87]_  = \new_[13905]_  & \new_[13894]_ ;
  assign \new_[88]_  = \new_[13883]_  & \new_[13872]_ ;
  assign \new_[89]_  = \new_[13861]_  & \new_[13850]_ ;
  assign \new_[90]_  = \new_[13839]_  & \new_[13828]_ ;
  assign \new_[91]_  = \new_[13817]_  & \new_[13806]_ ;
  assign \new_[92]_  = \new_[13795]_  & \new_[13784]_ ;
  assign \new_[93]_  = \new_[13773]_  & \new_[13762]_ ;
  assign \new_[94]_  = \new_[13751]_  & \new_[13740]_ ;
  assign \new_[95]_  = \new_[13729]_  & \new_[13718]_ ;
  assign \new_[96]_  = \new_[13707]_  & \new_[13696]_ ;
  assign \new_[97]_  = \new_[13685]_  & \new_[13674]_ ;
  assign \new_[98]_  = \new_[13665]_  & \new_[13654]_ ;
  assign \new_[99]_  = \new_[13645]_  & \new_[13634]_ ;
  assign \new_[100]_  = \new_[13625]_  & \new_[13614]_ ;
  assign \new_[101]_  = \new_[13605]_  & \new_[13594]_ ;
  assign \new_[102]_  = \new_[13585]_  & \new_[13574]_ ;
  assign \new_[103]_  = \new_[13565]_  & \new_[13554]_ ;
  assign \new_[104]_  = \new_[13545]_  & \new_[13534]_ ;
  assign \new_[105]_  = \new_[13525]_  & \new_[13514]_ ;
  assign \new_[106]_  = \new_[13505]_  & \new_[13494]_ ;
  assign \new_[107]_  = \new_[13485]_  & \new_[13474]_ ;
  assign \new_[108]_  = \new_[13465]_  & \new_[13454]_ ;
  assign \new_[109]_  = \new_[13445]_  & \new_[13434]_ ;
  assign \new_[110]_  = \new_[13425]_  & \new_[13414]_ ;
  assign \new_[111]_  = \new_[13405]_  & \new_[13394]_ ;
  assign \new_[112]_  = \new_[13385]_  & \new_[13374]_ ;
  assign \new_[113]_  = \new_[13365]_  & \new_[13354]_ ;
  assign \new_[114]_  = \new_[13345]_  & \new_[13334]_ ;
  assign \new_[115]_  = \new_[13325]_  & \new_[13314]_ ;
  assign \new_[116]_  = \new_[13305]_  & \new_[13294]_ ;
  assign \new_[117]_  = \new_[13285]_  & \new_[13274]_ ;
  assign \new_[118]_  = \new_[13265]_  & \new_[13254]_ ;
  assign \new_[119]_  = \new_[13245]_  & \new_[13234]_ ;
  assign \new_[120]_  = \new_[13225]_  & \new_[13214]_ ;
  assign \new_[121]_  = \new_[13205]_  & \new_[13194]_ ;
  assign \new_[122]_  = \new_[13185]_  & \new_[13174]_ ;
  assign \new_[123]_  = \new_[13165]_  & \new_[13154]_ ;
  assign \new_[124]_  = \new_[13145]_  & \new_[13134]_ ;
  assign \new_[125]_  = \new_[13125]_  & \new_[13114]_ ;
  assign \new_[126]_  = \new_[13105]_  & \new_[13094]_ ;
  assign \new_[127]_  = \new_[13085]_  & \new_[13074]_ ;
  assign \new_[128]_  = \new_[13065]_  & \new_[13054]_ ;
  assign \new_[129]_  = \new_[13045]_  & \new_[13034]_ ;
  assign \new_[130]_  = \new_[13025]_  & \new_[13014]_ ;
  assign \new_[131]_  = \new_[13005]_  & \new_[12994]_ ;
  assign \new_[132]_  = \new_[12985]_  & \new_[12974]_ ;
  assign \new_[133]_  = \new_[12965]_  & \new_[12954]_ ;
  assign \new_[134]_  = \new_[12945]_  & \new_[12934]_ ;
  assign \new_[135]_  = \new_[12925]_  & \new_[12914]_ ;
  assign \new_[136]_  = \new_[12905]_  & \new_[12894]_ ;
  assign \new_[137]_  = \new_[12885]_  & \new_[12874]_ ;
  assign \new_[138]_  = \new_[12865]_  & \new_[12854]_ ;
  assign \new_[139]_  = \new_[12845]_  & \new_[12834]_ ;
  assign \new_[140]_  = \new_[12825]_  & \new_[12814]_ ;
  assign \new_[141]_  = \new_[12805]_  & \new_[12794]_ ;
  assign \new_[142]_  = \new_[12785]_  & \new_[12774]_ ;
  assign \new_[143]_  = \new_[12765]_  & \new_[12754]_ ;
  assign \new_[144]_  = \new_[12745]_  & \new_[12734]_ ;
  assign \new_[145]_  = \new_[12725]_  & \new_[12714]_ ;
  assign \new_[146]_  = \new_[12705]_  & \new_[12694]_ ;
  assign \new_[147]_  = \new_[12685]_  & \new_[12674]_ ;
  assign \new_[148]_  = \new_[12665]_  & \new_[12654]_ ;
  assign \new_[149]_  = \new_[12645]_  & \new_[12634]_ ;
  assign \new_[150]_  = \new_[12625]_  & \new_[12614]_ ;
  assign \new_[151]_  = \new_[12605]_  & \new_[12594]_ ;
  assign \new_[152]_  = \new_[12585]_  & \new_[12574]_ ;
  assign \new_[153]_  = \new_[12565]_  & \new_[12554]_ ;
  assign \new_[154]_  = \new_[12545]_  & \new_[12534]_ ;
  assign \new_[155]_  = \new_[12525]_  & \new_[12514]_ ;
  assign \new_[156]_  = \new_[12505]_  & \new_[12494]_ ;
  assign \new_[157]_  = \new_[12485]_  & \new_[12474]_ ;
  assign \new_[158]_  = \new_[12465]_  & \new_[12454]_ ;
  assign \new_[159]_  = \new_[12445]_  & \new_[12434]_ ;
  assign \new_[160]_  = \new_[12425]_  & \new_[12414]_ ;
  assign \new_[161]_  = \new_[12405]_  & \new_[12394]_ ;
  assign \new_[162]_  = \new_[12385]_  & \new_[12374]_ ;
  assign \new_[163]_  = \new_[12365]_  & \new_[12354]_ ;
  assign \new_[164]_  = \new_[12345]_  & \new_[12334]_ ;
  assign \new_[165]_  = \new_[12325]_  & \new_[12314]_ ;
  assign \new_[166]_  = \new_[12305]_  & \new_[12294]_ ;
  assign \new_[167]_  = \new_[12285]_  & \new_[12274]_ ;
  assign \new_[168]_  = \new_[12265]_  & \new_[12254]_ ;
  assign \new_[169]_  = \new_[12245]_  & \new_[12234]_ ;
  assign \new_[170]_  = \new_[12225]_  & \new_[12214]_ ;
  assign \new_[171]_  = \new_[12205]_  & \new_[12194]_ ;
  assign \new_[172]_  = \new_[12185]_  & \new_[12174]_ ;
  assign \new_[173]_  = \new_[12165]_  & \new_[12154]_ ;
  assign \new_[174]_  = \new_[12145]_  & \new_[12134]_ ;
  assign \new_[175]_  = \new_[12125]_  & \new_[12114]_ ;
  assign \new_[176]_  = \new_[12105]_  & \new_[12094]_ ;
  assign \new_[177]_  = \new_[12085]_  & \new_[12074]_ ;
  assign \new_[178]_  = \new_[12065]_  & \new_[12054]_ ;
  assign \new_[179]_  = \new_[12045]_  & \new_[12034]_ ;
  assign \new_[180]_  = \new_[12025]_  & \new_[12014]_ ;
  assign \new_[181]_  = \new_[12005]_  & \new_[11994]_ ;
  assign \new_[182]_  = \new_[11985]_  & \new_[11974]_ ;
  assign \new_[183]_  = \new_[11965]_  & \new_[11954]_ ;
  assign \new_[184]_  = \new_[11945]_  & \new_[11934]_ ;
  assign \new_[185]_  = \new_[11925]_  & \new_[11914]_ ;
  assign \new_[186]_  = \new_[11905]_  & \new_[11894]_ ;
  assign \new_[187]_  = \new_[11885]_  & \new_[11874]_ ;
  assign \new_[188]_  = \new_[11865]_  & \new_[11854]_ ;
  assign \new_[189]_  = \new_[11845]_  & \new_[11834]_ ;
  assign \new_[190]_  = \new_[11825]_  & \new_[11814]_ ;
  assign \new_[191]_  = \new_[11805]_  & \new_[11794]_ ;
  assign \new_[192]_  = \new_[11785]_  & \new_[11774]_ ;
  assign \new_[193]_  = \new_[11765]_  & \new_[11754]_ ;
  assign \new_[194]_  = \new_[11745]_  & \new_[11734]_ ;
  assign \new_[195]_  = \new_[11725]_  & \new_[11714]_ ;
  assign \new_[196]_  = \new_[11705]_  & \new_[11694]_ ;
  assign \new_[197]_  = \new_[11685]_  & \new_[11674]_ ;
  assign \new_[198]_  = \new_[11665]_  & \new_[11654]_ ;
  assign \new_[199]_  = \new_[11645]_  & \new_[11634]_ ;
  assign \new_[200]_  = \new_[11625]_  & \new_[11614]_ ;
  assign \new_[201]_  = \new_[11605]_  & \new_[11594]_ ;
  assign \new_[202]_  = \new_[11585]_  & \new_[11574]_ ;
  assign \new_[203]_  = \new_[11565]_  & \new_[11554]_ ;
  assign \new_[204]_  = \new_[11545]_  & \new_[11534]_ ;
  assign \new_[205]_  = \new_[11525]_  & \new_[11514]_ ;
  assign \new_[206]_  = \new_[11505]_  & \new_[11494]_ ;
  assign \new_[207]_  = \new_[11485]_  & \new_[11474]_ ;
  assign \new_[208]_  = \new_[11465]_  & \new_[11454]_ ;
  assign \new_[209]_  = \new_[11445]_  & \new_[11434]_ ;
  assign \new_[210]_  = \new_[11425]_  & \new_[11414]_ ;
  assign \new_[211]_  = \new_[11405]_  & \new_[11394]_ ;
  assign \new_[212]_  = \new_[11385]_  & \new_[11374]_ ;
  assign \new_[213]_  = \new_[11365]_  & \new_[11354]_ ;
  assign \new_[214]_  = \new_[11345]_  & \new_[11334]_ ;
  assign \new_[215]_  = \new_[11325]_  & \new_[11314]_ ;
  assign \new_[216]_  = \new_[11305]_  & \new_[11294]_ ;
  assign \new_[217]_  = \new_[11285]_  & \new_[11274]_ ;
  assign \new_[218]_  = \new_[11265]_  & \new_[11254]_ ;
  assign \new_[219]_  = \new_[11245]_  & \new_[11234]_ ;
  assign \new_[220]_  = \new_[11225]_  & \new_[11214]_ ;
  assign \new_[221]_  = \new_[11205]_  & \new_[11194]_ ;
  assign \new_[222]_  = \new_[11185]_  & \new_[11174]_ ;
  assign \new_[223]_  = \new_[11165]_  & \new_[11154]_ ;
  assign \new_[224]_  = \new_[11145]_  & \new_[11134]_ ;
  assign \new_[225]_  = \new_[11125]_  & \new_[11114]_ ;
  assign \new_[226]_  = \new_[11105]_  & \new_[11094]_ ;
  assign \new_[227]_  = \new_[11085]_  & \new_[11074]_ ;
  assign \new_[228]_  = \new_[11065]_  & \new_[11054]_ ;
  assign \new_[229]_  = \new_[11045]_  & \new_[11034]_ ;
  assign \new_[230]_  = \new_[11025]_  & \new_[11014]_ ;
  assign \new_[231]_  = \new_[11005]_  & \new_[10994]_ ;
  assign \new_[232]_  = \new_[10985]_  & \new_[10974]_ ;
  assign \new_[233]_  = \new_[10965]_  & \new_[10954]_ ;
  assign \new_[234]_  = \new_[10945]_  & \new_[10934]_ ;
  assign \new_[235]_  = \new_[10925]_  & \new_[10914]_ ;
  assign \new_[236]_  = \new_[10905]_  & \new_[10894]_ ;
  assign \new_[237]_  = \new_[10885]_  & \new_[10874]_ ;
  assign \new_[238]_  = \new_[10865]_  & \new_[10854]_ ;
  assign \new_[239]_  = \new_[10845]_  & \new_[10834]_ ;
  assign \new_[240]_  = \new_[10825]_  & \new_[10814]_ ;
  assign \new_[241]_  = \new_[10805]_  & \new_[10794]_ ;
  assign \new_[242]_  = \new_[10785]_  & \new_[10774]_ ;
  assign \new_[243]_  = \new_[10765]_  & \new_[10754]_ ;
  assign \new_[244]_  = \new_[10745]_  & \new_[10734]_ ;
  assign \new_[245]_  = \new_[10725]_  & \new_[10714]_ ;
  assign \new_[246]_  = \new_[10705]_  & \new_[10694]_ ;
  assign \new_[247]_  = \new_[10685]_  & \new_[10674]_ ;
  assign \new_[248]_  = \new_[10665]_  & \new_[10654]_ ;
  assign \new_[249]_  = \new_[10645]_  & \new_[10634]_ ;
  assign \new_[250]_  = \new_[10625]_  & \new_[10614]_ ;
  assign \new_[251]_  = \new_[10605]_  & \new_[10594]_ ;
  assign \new_[252]_  = \new_[10585]_  & \new_[10574]_ ;
  assign \new_[253]_  = \new_[10565]_  & \new_[10554]_ ;
  assign \new_[254]_  = \new_[10545]_  & \new_[10534]_ ;
  assign \new_[255]_  = \new_[10525]_  & \new_[10514]_ ;
  assign \new_[256]_  = \new_[10505]_  & \new_[10494]_ ;
  assign \new_[257]_  = \new_[10485]_  & \new_[10474]_ ;
  assign \new_[258]_  = \new_[10465]_  & \new_[10454]_ ;
  assign \new_[259]_  = \new_[10445]_  & \new_[10434]_ ;
  assign \new_[260]_  = \new_[10425]_  & \new_[10414]_ ;
  assign \new_[261]_  = \new_[10405]_  & \new_[10394]_ ;
  assign \new_[262]_  = \new_[10385]_  & \new_[10374]_ ;
  assign \new_[263]_  = \new_[10365]_  & \new_[10354]_ ;
  assign \new_[264]_  = \new_[10345]_  & \new_[10334]_ ;
  assign \new_[265]_  = \new_[10325]_  & \new_[10316]_ ;
  assign \new_[266]_  = \new_[10307]_  & \new_[10298]_ ;
  assign \new_[267]_  = \new_[10289]_  & \new_[10280]_ ;
  assign \new_[268]_  = \new_[10271]_  & \new_[10262]_ ;
  assign \new_[269]_  = \new_[10253]_  & \new_[10244]_ ;
  assign \new_[270]_  = \new_[10235]_  & \new_[10226]_ ;
  assign \new_[271]_  = \new_[10217]_  & \new_[10208]_ ;
  assign \new_[272]_  = \new_[10199]_  & \new_[10190]_ ;
  assign \new_[273]_  = \new_[10181]_  & \new_[10172]_ ;
  assign \new_[274]_  = \new_[10163]_  & \new_[10154]_ ;
  assign \new_[275]_  = \new_[10145]_  & \new_[10136]_ ;
  assign \new_[276]_  = \new_[10127]_  & \new_[10118]_ ;
  assign \new_[277]_  = \new_[10109]_  & \new_[10100]_ ;
  assign \new_[278]_  = \new_[10091]_  & \new_[10082]_ ;
  assign \new_[279]_  = \new_[10073]_  & \new_[10064]_ ;
  assign \new_[280]_  = \new_[10055]_  & \new_[10046]_ ;
  assign \new_[281]_  = \new_[10037]_  & \new_[10028]_ ;
  assign \new_[282]_  = \new_[10019]_  & \new_[10010]_ ;
  assign \new_[283]_  = \new_[10001]_  & \new_[9992]_ ;
  assign \new_[284]_  = \new_[9983]_  & \new_[9974]_ ;
  assign \new_[285]_  = \new_[9965]_  & \new_[9956]_ ;
  assign \new_[286]_  = \new_[9947]_  & \new_[9938]_ ;
  assign \new_[287]_  = \new_[9929]_  & \new_[9920]_ ;
  assign \new_[288]_  = \new_[9911]_  & \new_[9902]_ ;
  assign \new_[289]_  = \new_[9893]_  & \new_[9884]_ ;
  assign \new_[290]_  = \new_[9875]_  & \new_[9866]_ ;
  assign \new_[291]_  = \new_[9857]_  & \new_[9848]_ ;
  assign \new_[292]_  = \new_[9839]_  & \new_[9830]_ ;
  assign \new_[293]_  = \new_[9821]_  & \new_[9812]_ ;
  assign \new_[294]_  = \new_[9803]_  & \new_[9794]_ ;
  assign \new_[295]_  = \new_[9785]_  & \new_[9776]_ ;
  assign \new_[296]_  = \new_[9767]_  & \new_[9758]_ ;
  assign \new_[297]_  = \new_[9749]_  & \new_[9740]_ ;
  assign \new_[298]_  = \new_[9731]_  & \new_[9722]_ ;
  assign \new_[299]_  = \new_[9713]_  & \new_[9704]_ ;
  assign \new_[300]_  = \new_[9695]_  & \new_[9686]_ ;
  assign \new_[301]_  = \new_[9677]_  & \new_[9668]_ ;
  assign \new_[302]_  = \new_[9659]_  & \new_[9650]_ ;
  assign \new_[303]_  = \new_[9641]_  & \new_[9632]_ ;
  assign \new_[304]_  = \new_[9623]_  & \new_[9614]_ ;
  assign \new_[305]_  = \new_[9605]_  & \new_[9596]_ ;
  assign \new_[306]_  = \new_[9587]_  & \new_[9578]_ ;
  assign \new_[307]_  = \new_[9569]_  & \new_[9560]_ ;
  assign \new_[308]_  = \new_[9551]_  & \new_[9542]_ ;
  assign \new_[309]_  = \new_[9533]_  & \new_[9524]_ ;
  assign \new_[310]_  = \new_[9515]_  & \new_[9506]_ ;
  assign \new_[311]_  = \new_[9497]_  & \new_[9488]_ ;
  assign \new_[312]_  = \new_[9479]_  & \new_[9470]_ ;
  assign \new_[313]_  = \new_[9461]_  & \new_[9452]_ ;
  assign \new_[314]_  = \new_[9443]_  & \new_[9434]_ ;
  assign \new_[315]_  = \new_[9425]_  & \new_[9416]_ ;
  assign \new_[316]_  = \new_[9407]_  & \new_[9398]_ ;
  assign \new_[317]_  = \new_[9389]_  & \new_[9380]_ ;
  assign \new_[318]_  = \new_[9371]_  & \new_[9362]_ ;
  assign \new_[319]_  = \new_[9353]_  & \new_[9344]_ ;
  assign \new_[320]_  = \new_[9335]_  & \new_[9326]_ ;
  assign \new_[321]_  = \new_[9317]_  & \new_[9308]_ ;
  assign \new_[322]_  = \new_[9299]_  & \new_[9290]_ ;
  assign \new_[323]_  = \new_[9281]_  & \new_[9272]_ ;
  assign \new_[324]_  = \new_[9263]_  & \new_[9254]_ ;
  assign \new_[325]_  = \new_[9245]_  & \new_[9236]_ ;
  assign \new_[326]_  = \new_[9227]_  & \new_[9218]_ ;
  assign \new_[327]_  = \new_[9209]_  & \new_[9200]_ ;
  assign \new_[328]_  = \new_[9191]_  & \new_[9182]_ ;
  assign \new_[329]_  = \new_[9173]_  & \new_[9164]_ ;
  assign \new_[330]_  = \new_[9155]_  & \new_[9146]_ ;
  assign \new_[331]_  = \new_[9137]_  & \new_[9128]_ ;
  assign \new_[332]_  = \new_[9119]_  & \new_[9110]_ ;
  assign \new_[333]_  = \new_[9101]_  & \new_[9092]_ ;
  assign \new_[334]_  = \new_[9083]_  & \new_[9074]_ ;
  assign \new_[335]_  = \new_[9065]_  & \new_[9056]_ ;
  assign \new_[336]_  = \new_[9047]_  & \new_[9038]_ ;
  assign \new_[337]_  = \new_[9029]_  & \new_[9020]_ ;
  assign \new_[338]_  = \new_[9011]_  & \new_[9002]_ ;
  assign \new_[339]_  = \new_[8993]_  & \new_[8984]_ ;
  assign \new_[340]_  = \new_[8975]_  & \new_[8966]_ ;
  assign \new_[341]_  = \new_[8957]_  & \new_[8948]_ ;
  assign \new_[342]_  = \new_[8939]_  & \new_[8930]_ ;
  assign \new_[343]_  = \new_[8921]_  & \new_[8912]_ ;
  assign \new_[344]_  = \new_[8903]_  & \new_[8894]_ ;
  assign \new_[345]_  = \new_[8885]_  & \new_[8876]_ ;
  assign \new_[346]_  = \new_[8867]_  & \new_[8858]_ ;
  assign \new_[347]_  = \new_[8849]_  & \new_[8840]_ ;
  assign \new_[348]_  = \new_[8831]_  & \new_[8822]_ ;
  assign \new_[349]_  = \new_[8813]_  & \new_[8804]_ ;
  assign \new_[350]_  = \new_[8795]_  & \new_[8786]_ ;
  assign \new_[351]_  = \new_[8777]_  & \new_[8768]_ ;
  assign \new_[352]_  = \new_[8759]_  & \new_[8750]_ ;
  assign \new_[353]_  = \new_[8741]_  & \new_[8732]_ ;
  assign \new_[354]_  = \new_[8723]_  & \new_[8714]_ ;
  assign \new_[355]_  = \new_[8705]_  & \new_[8696]_ ;
  assign \new_[356]_  = \new_[8687]_  & \new_[8678]_ ;
  assign \new_[357]_  = \new_[8669]_  & \new_[8660]_ ;
  assign \new_[358]_  = \new_[8651]_  & \new_[8642]_ ;
  assign \new_[359]_  = \new_[8633]_  & \new_[8624]_ ;
  assign \new_[360]_  = \new_[8615]_  & \new_[8606]_ ;
  assign \new_[361]_  = \new_[8597]_  & \new_[8588]_ ;
  assign \new_[362]_  = \new_[8579]_  & \new_[8570]_ ;
  assign \new_[363]_  = \new_[8561]_  & \new_[8552]_ ;
  assign \new_[364]_  = \new_[8543]_  & \new_[8534]_ ;
  assign \new_[365]_  = \new_[8525]_  & \new_[8516]_ ;
  assign \new_[366]_  = \new_[8507]_  & \new_[8498]_ ;
  assign \new_[367]_  = \new_[8489]_  & \new_[8480]_ ;
  assign \new_[368]_  = \new_[8471]_  & \new_[8462]_ ;
  assign \new_[369]_  = \new_[8453]_  & \new_[8444]_ ;
  assign \new_[370]_  = \new_[8435]_  & \new_[8426]_ ;
  assign \new_[371]_  = \new_[8417]_  & \new_[8408]_ ;
  assign \new_[372]_  = \new_[8399]_  & \new_[8390]_ ;
  assign \new_[373]_  = \new_[8381]_  & \new_[8372]_ ;
  assign \new_[374]_  = \new_[8363]_  & \new_[8354]_ ;
  assign \new_[375]_  = \new_[8345]_  & \new_[8336]_ ;
  assign \new_[376]_  = \new_[8327]_  & \new_[8318]_ ;
  assign \new_[377]_  = \new_[8309]_  & \new_[8300]_ ;
  assign \new_[378]_  = \new_[8291]_  & \new_[8282]_ ;
  assign \new_[379]_  = \new_[8273]_  & \new_[8264]_ ;
  assign \new_[380]_  = \new_[8255]_  & \new_[8246]_ ;
  assign \new_[381]_  = \new_[8237]_  & \new_[8228]_ ;
  assign \new_[382]_  = \new_[8219]_  & \new_[8210]_ ;
  assign \new_[383]_  = \new_[8201]_  & \new_[8192]_ ;
  assign \new_[384]_  = \new_[8183]_  & \new_[8174]_ ;
  assign \new_[385]_  = \new_[8165]_  & \new_[8156]_ ;
  assign \new_[386]_  = \new_[8147]_  & \new_[8138]_ ;
  assign \new_[387]_  = \new_[8129]_  & \new_[8120]_ ;
  assign \new_[388]_  = \new_[8111]_  & \new_[8102]_ ;
  assign \new_[389]_  = \new_[8093]_  & \new_[8084]_ ;
  assign \new_[390]_  = \new_[8075]_  & \new_[8066]_ ;
  assign \new_[391]_  = \new_[8057]_  & \new_[8048]_ ;
  assign \new_[392]_  = \new_[8039]_  & \new_[8030]_ ;
  assign \new_[393]_  = \new_[8021]_  & \new_[8012]_ ;
  assign \new_[394]_  = \new_[8003]_  & \new_[7994]_ ;
  assign \new_[395]_  = \new_[7985]_  & \new_[7976]_ ;
  assign \new_[396]_  = \new_[7967]_  & \new_[7958]_ ;
  assign \new_[397]_  = \new_[7949]_  & \new_[7940]_ ;
  assign \new_[398]_  = \new_[7931]_  & \new_[7922]_ ;
  assign \new_[399]_  = \new_[7913]_  & \new_[7904]_ ;
  assign \new_[400]_  = \new_[7895]_  & \new_[7886]_ ;
  assign \new_[401]_  = \new_[7877]_  & \new_[7868]_ ;
  assign \new_[402]_  = \new_[7859]_  & \new_[7850]_ ;
  assign \new_[403]_  = \new_[7841]_  & \new_[7832]_ ;
  assign \new_[404]_  = \new_[7823]_  & \new_[7814]_ ;
  assign \new_[405]_  = \new_[7805]_  & \new_[7796]_ ;
  assign \new_[406]_  = \new_[7787]_  & \new_[7778]_ ;
  assign \new_[407]_  = \new_[7769]_  & \new_[7760]_ ;
  assign \new_[408]_  = \new_[7751]_  & \new_[7742]_ ;
  assign \new_[409]_  = \new_[7733]_  & \new_[7724]_ ;
  assign \new_[410]_  = \new_[7715]_  & \new_[7706]_ ;
  assign \new_[411]_  = \new_[7697]_  & \new_[7688]_ ;
  assign \new_[412]_  = \new_[7679]_  & \new_[7670]_ ;
  assign \new_[413]_  = \new_[7661]_  & \new_[7652]_ ;
  assign \new_[414]_  = \new_[7643]_  & \new_[7634]_ ;
  assign \new_[415]_  = \new_[7625]_  & \new_[7616]_ ;
  assign \new_[416]_  = \new_[7607]_  & \new_[7598]_ ;
  assign \new_[417]_  = \new_[7589]_  & \new_[7580]_ ;
  assign \new_[418]_  = \new_[7571]_  & \new_[7562]_ ;
  assign \new_[419]_  = \new_[7553]_  & \new_[7544]_ ;
  assign \new_[420]_  = \new_[7535]_  & \new_[7526]_ ;
  assign \new_[421]_  = \new_[7517]_  & \new_[7508]_ ;
  assign \new_[422]_  = \new_[7499]_  & \new_[7490]_ ;
  assign \new_[423]_  = \new_[7481]_  & \new_[7472]_ ;
  assign \new_[424]_  = \new_[7463]_  & \new_[7454]_ ;
  assign \new_[425]_  = \new_[7445]_  & \new_[7436]_ ;
  assign \new_[426]_  = \new_[7427]_  & \new_[7418]_ ;
  assign \new_[427]_  = \new_[7409]_  & \new_[7400]_ ;
  assign \new_[428]_  = \new_[7391]_  & \new_[7382]_ ;
  assign \new_[429]_  = \new_[7373]_  & \new_[7364]_ ;
  assign \new_[430]_  = \new_[7355]_  & \new_[7346]_ ;
  assign \new_[431]_  = \new_[7337]_  & \new_[7328]_ ;
  assign \new_[432]_  = \new_[7319]_  & \new_[7310]_ ;
  assign \new_[433]_  = \new_[7301]_  & \new_[7292]_ ;
  assign \new_[434]_  = \new_[7283]_  & \new_[7274]_ ;
  assign \new_[435]_  = \new_[7265]_  & \new_[7256]_ ;
  assign \new_[436]_  = \new_[7247]_  & \new_[7238]_ ;
  assign \new_[437]_  = \new_[7229]_  & \new_[7220]_ ;
  assign \new_[438]_  = \new_[7211]_  & \new_[7202]_ ;
  assign \new_[439]_  = \new_[7193]_  & \new_[7184]_ ;
  assign \new_[440]_  = \new_[7175]_  & \new_[7166]_ ;
  assign \new_[441]_  = \new_[7157]_  & \new_[7148]_ ;
  assign \new_[442]_  = \new_[7139]_  & \new_[7130]_ ;
  assign \new_[443]_  = \new_[7121]_  & \new_[7112]_ ;
  assign \new_[444]_  = \new_[7103]_  & \new_[7094]_ ;
  assign \new_[445]_  = \new_[7085]_  & \new_[7076]_ ;
  assign \new_[446]_  = \new_[7067]_  & \new_[7058]_ ;
  assign \new_[447]_  = \new_[7049]_  & \new_[7040]_ ;
  assign \new_[448]_  = \new_[7031]_  & \new_[7022]_ ;
  assign \new_[449]_  = \new_[7013]_  & \new_[7004]_ ;
  assign \new_[450]_  = \new_[6995]_  & \new_[6986]_ ;
  assign \new_[451]_  = \new_[6977]_  & \new_[6968]_ ;
  assign \new_[452]_  = \new_[6959]_  & \new_[6950]_ ;
  assign \new_[453]_  = \new_[6941]_  & \new_[6932]_ ;
  assign \new_[454]_  = \new_[6923]_  & \new_[6914]_ ;
  assign \new_[455]_  = \new_[6905]_  & \new_[6896]_ ;
  assign \new_[456]_  = \new_[6887]_  & \new_[6878]_ ;
  assign \new_[457]_  = \new_[6869]_  & \new_[6860]_ ;
  assign \new_[458]_  = \new_[6851]_  & \new_[6842]_ ;
  assign \new_[459]_  = \new_[6833]_  & \new_[6824]_ ;
  assign \new_[460]_  = \new_[6815]_  & \new_[6806]_ ;
  assign \new_[461]_  = \new_[6797]_  & \new_[6788]_ ;
  assign \new_[462]_  = \new_[6779]_  & \new_[6770]_ ;
  assign \new_[463]_  = \new_[6761]_  & \new_[6752]_ ;
  assign \new_[464]_  = \new_[6743]_  & \new_[6734]_ ;
  assign \new_[465]_  = \new_[6725]_  & \new_[6716]_ ;
  assign \new_[466]_  = \new_[6707]_  & \new_[6698]_ ;
  assign \new_[467]_  = \new_[6689]_  & \new_[6680]_ ;
  assign \new_[468]_  = \new_[6671]_  & \new_[6662]_ ;
  assign \new_[469]_  = \new_[6653]_  & \new_[6644]_ ;
  assign \new_[470]_  = \new_[6635]_  & \new_[6626]_ ;
  assign \new_[471]_  = \new_[6617]_  & \new_[6608]_ ;
  assign \new_[472]_  = \new_[6599]_  & \new_[6590]_ ;
  assign \new_[473]_  = \new_[6581]_  & \new_[6572]_ ;
  assign \new_[474]_  = \new_[6565]_  & \new_[6556]_ ;
  assign \new_[475]_  = \new_[6549]_  & \new_[6540]_ ;
  assign \new_[476]_  = \new_[6533]_  & \new_[6524]_ ;
  assign \new_[477]_  = \new_[6517]_  & \new_[6508]_ ;
  assign \new_[478]_  = \new_[6501]_  & \new_[6492]_ ;
  assign \new_[479]_  = \new_[6485]_  & \new_[6476]_ ;
  assign \new_[480]_  = \new_[6469]_  & \new_[6460]_ ;
  assign \new_[481]_  = \new_[6453]_  & \new_[6444]_ ;
  assign \new_[482]_  = \new_[6437]_  & \new_[6428]_ ;
  assign \new_[483]_  = \new_[6421]_  & \new_[6412]_ ;
  assign \new_[484]_  = \new_[6405]_  & \new_[6396]_ ;
  assign \new_[485]_  = \new_[6389]_  & \new_[6380]_ ;
  assign \new_[486]_  = \new_[6373]_  & \new_[6364]_ ;
  assign \new_[487]_  = \new_[6357]_  & \new_[6348]_ ;
  assign \new_[488]_  = \new_[6341]_  & \new_[6332]_ ;
  assign \new_[489]_  = \new_[6325]_  & \new_[6316]_ ;
  assign \new_[490]_  = \new_[6309]_  & \new_[6300]_ ;
  assign \new_[491]_  = \new_[6293]_  & \new_[6284]_ ;
  assign \new_[492]_  = \new_[6277]_  & \new_[6268]_ ;
  assign \new_[493]_  = \new_[6261]_  & \new_[6252]_ ;
  assign \new_[494]_  = \new_[6245]_  & \new_[6236]_ ;
  assign \new_[495]_  = \new_[6229]_  & \new_[6220]_ ;
  assign \new_[496]_  = \new_[6213]_  & \new_[6204]_ ;
  assign \new_[497]_  = \new_[6197]_  & \new_[6188]_ ;
  assign \new_[498]_  = \new_[6181]_  & \new_[6172]_ ;
  assign \new_[499]_  = \new_[6165]_  & \new_[6156]_ ;
  assign \new_[500]_  = \new_[6149]_  & \new_[6140]_ ;
  assign \new_[501]_  = \new_[6133]_  & \new_[6124]_ ;
  assign \new_[502]_  = \new_[6117]_  & \new_[6108]_ ;
  assign \new_[503]_  = \new_[6101]_  & \new_[6092]_ ;
  assign \new_[504]_  = \new_[6085]_  & \new_[6076]_ ;
  assign \new_[505]_  = \new_[6069]_  & \new_[6060]_ ;
  assign \new_[506]_  = \new_[6053]_  & \new_[6044]_ ;
  assign \new_[507]_  = \new_[6037]_  & \new_[6028]_ ;
  assign \new_[508]_  = \new_[6021]_  & \new_[6012]_ ;
  assign \new_[509]_  = \new_[6005]_  & \new_[5996]_ ;
  assign \new_[510]_  = \new_[5989]_  & \new_[5980]_ ;
  assign \new_[511]_  = \new_[5973]_  & \new_[5964]_ ;
  assign \new_[512]_  = \new_[5957]_  & \new_[5948]_ ;
  assign \new_[513]_  = \new_[5941]_  & \new_[5932]_ ;
  assign \new_[514]_  = \new_[5925]_  & \new_[5916]_ ;
  assign \new_[515]_  = \new_[5909]_  & \new_[5900]_ ;
  assign \new_[516]_  = \new_[5893]_  & \new_[5884]_ ;
  assign \new_[517]_  = \new_[5877]_  & \new_[5868]_ ;
  assign \new_[518]_  = \new_[5861]_  & \new_[5852]_ ;
  assign \new_[519]_  = \new_[5845]_  & \new_[5836]_ ;
  assign \new_[520]_  = \new_[5829]_  & \new_[5820]_ ;
  assign \new_[521]_  = \new_[5813]_  & \new_[5804]_ ;
  assign \new_[522]_  = \new_[5797]_  & \new_[5788]_ ;
  assign \new_[523]_  = \new_[5781]_  & \new_[5772]_ ;
  assign \new_[524]_  = \new_[5765]_  & \new_[5756]_ ;
  assign \new_[525]_  = \new_[5749]_  & \new_[5740]_ ;
  assign \new_[526]_  = \new_[5733]_  & \new_[5724]_ ;
  assign \new_[527]_  = \new_[5717]_  & \new_[5708]_ ;
  assign \new_[528]_  = \new_[5701]_  & \new_[5692]_ ;
  assign \new_[529]_  = \new_[5685]_  & \new_[5676]_ ;
  assign \new_[530]_  = \new_[5669]_  & \new_[5660]_ ;
  assign \new_[531]_  = \new_[5653]_  & \new_[5644]_ ;
  assign \new_[532]_  = \new_[5637]_  & \new_[5628]_ ;
  assign \new_[533]_  = \new_[5621]_  & \new_[5612]_ ;
  assign \new_[534]_  = \new_[5605]_  & \new_[5596]_ ;
  assign \new_[535]_  = \new_[5589]_  & \new_[5580]_ ;
  assign \new_[536]_  = \new_[5573]_  & \new_[5564]_ ;
  assign \new_[537]_  = \new_[5557]_  & \new_[5548]_ ;
  assign \new_[538]_  = \new_[5541]_  & \new_[5532]_ ;
  assign \new_[539]_  = \new_[5525]_  & \new_[5516]_ ;
  assign \new_[540]_  = \new_[5509]_  & \new_[5500]_ ;
  assign \new_[541]_  = \new_[5493]_  & \new_[5484]_ ;
  assign \new_[542]_  = \new_[5477]_  & \new_[5468]_ ;
  assign \new_[543]_  = \new_[5461]_  & \new_[5452]_ ;
  assign \new_[544]_  = \new_[5445]_  & \new_[5436]_ ;
  assign \new_[545]_  = \new_[5429]_  & \new_[5420]_ ;
  assign \new_[546]_  = \new_[5413]_  & \new_[5404]_ ;
  assign \new_[547]_  = \new_[5397]_  & \new_[5388]_ ;
  assign \new_[548]_  = \new_[5381]_  & \new_[5372]_ ;
  assign \new_[549]_  = \new_[5365]_  & \new_[5356]_ ;
  assign \new_[550]_  = \new_[5349]_  & \new_[5340]_ ;
  assign \new_[551]_  = \new_[5333]_  & \new_[5324]_ ;
  assign \new_[552]_  = \new_[5317]_  & \new_[5308]_ ;
  assign \new_[553]_  = \new_[5301]_  & \new_[5292]_ ;
  assign \new_[554]_  = \new_[5285]_  & \new_[5276]_ ;
  assign \new_[555]_  = \new_[5269]_  & \new_[5260]_ ;
  assign \new_[556]_  = \new_[5253]_  & \new_[5244]_ ;
  assign \new_[557]_  = \new_[5237]_  & \new_[5228]_ ;
  assign \new_[558]_  = \new_[5221]_  & \new_[5212]_ ;
  assign \new_[559]_  = \new_[5205]_  & \new_[5196]_ ;
  assign \new_[560]_  = \new_[5189]_  & \new_[5180]_ ;
  assign \new_[561]_  = \new_[5173]_  & \new_[5164]_ ;
  assign \new_[562]_  = \new_[5157]_  & \new_[5148]_ ;
  assign \new_[563]_  = \new_[5141]_  & \new_[5132]_ ;
  assign \new_[564]_  = \new_[5125]_  & \new_[5116]_ ;
  assign \new_[565]_  = \new_[5109]_  & \new_[5100]_ ;
  assign \new_[566]_  = \new_[5093]_  & \new_[5084]_ ;
  assign \new_[567]_  = \new_[5077]_  & \new_[5068]_ ;
  assign \new_[568]_  = \new_[5061]_  & \new_[5052]_ ;
  assign \new_[569]_  = \new_[5045]_  & \new_[5036]_ ;
  assign \new_[570]_  = \new_[5029]_  & \new_[5020]_ ;
  assign \new_[571]_  = \new_[5013]_  & \new_[5004]_ ;
  assign \new_[572]_  = \new_[4997]_  & \new_[4988]_ ;
  assign \new_[573]_  = \new_[4981]_  & \new_[4972]_ ;
  assign \new_[574]_  = \new_[4965]_  & \new_[4956]_ ;
  assign \new_[575]_  = \new_[4949]_  & \new_[4940]_ ;
  assign \new_[576]_  = \new_[4933]_  & \new_[4924]_ ;
  assign \new_[577]_  = \new_[4917]_  & \new_[4908]_ ;
  assign \new_[578]_  = \new_[4901]_  & \new_[4892]_ ;
  assign \new_[579]_  = \new_[4885]_  & \new_[4876]_ ;
  assign \new_[580]_  = \new_[4869]_  & \new_[4860]_ ;
  assign \new_[581]_  = \new_[4853]_  & \new_[4844]_ ;
  assign \new_[582]_  = \new_[4837]_  & \new_[4828]_ ;
  assign \new_[583]_  = \new_[4821]_  & \new_[4812]_ ;
  assign \new_[584]_  = \new_[4805]_  & \new_[4796]_ ;
  assign \new_[585]_  = \new_[4789]_  & \new_[4780]_ ;
  assign \new_[586]_  = \new_[4773]_  & \new_[4764]_ ;
  assign \new_[587]_  = \new_[4757]_  & \new_[4748]_ ;
  assign \new_[588]_  = \new_[4741]_  & \new_[4732]_ ;
  assign \new_[589]_  = \new_[4725]_  & \new_[4716]_ ;
  assign \new_[590]_  = \new_[4709]_  & \new_[4700]_ ;
  assign \new_[591]_  = \new_[4693]_  & \new_[4684]_ ;
  assign \new_[592]_  = \new_[4677]_  & \new_[4668]_ ;
  assign \new_[593]_  = \new_[4661]_  & \new_[4652]_ ;
  assign \new_[594]_  = \new_[4645]_  & \new_[4636]_ ;
  assign \new_[595]_  = \new_[4629]_  & \new_[4620]_ ;
  assign \new_[596]_  = \new_[4613]_  & \new_[4604]_ ;
  assign \new_[597]_  = \new_[4597]_  & \new_[4588]_ ;
  assign \new_[598]_  = \new_[4581]_  & \new_[4572]_ ;
  assign \new_[599]_  = \new_[4565]_  & \new_[4556]_ ;
  assign \new_[600]_  = \new_[4549]_  & \new_[4540]_ ;
  assign \new_[601]_  = \new_[4533]_  & \new_[4524]_ ;
  assign \new_[602]_  = \new_[4517]_  & \new_[4508]_ ;
  assign \new_[603]_  = \new_[4501]_  & \new_[4492]_ ;
  assign \new_[604]_  = \new_[4485]_  & \new_[4476]_ ;
  assign \new_[605]_  = \new_[4469]_  & \new_[4460]_ ;
  assign \new_[606]_  = \new_[4453]_  & \new_[4444]_ ;
  assign \new_[607]_  = \new_[4437]_  & \new_[4428]_ ;
  assign \new_[608]_  = \new_[4421]_  & \new_[4412]_ ;
  assign \new_[609]_  = \new_[4405]_  & \new_[4396]_ ;
  assign \new_[610]_  = \new_[4389]_  & \new_[4380]_ ;
  assign \new_[611]_  = \new_[4373]_  & \new_[4364]_ ;
  assign \new_[612]_  = \new_[4357]_  & \new_[4348]_ ;
  assign \new_[613]_  = \new_[4341]_  & \new_[4332]_ ;
  assign \new_[614]_  = \new_[4325]_  & \new_[4316]_ ;
  assign \new_[615]_  = \new_[4309]_  & \new_[4300]_ ;
  assign \new_[616]_  = \new_[4293]_  & \new_[4284]_ ;
  assign \new_[617]_  = \new_[4277]_  & \new_[4268]_ ;
  assign \new_[618]_  = \new_[4261]_  & \new_[4252]_ ;
  assign \new_[619]_  = \new_[4245]_  & \new_[4236]_ ;
  assign \new_[620]_  = \new_[4229]_  & \new_[4220]_ ;
  assign \new_[621]_  = \new_[4213]_  & \new_[4204]_ ;
  assign \new_[622]_  = \new_[4197]_  & \new_[4188]_ ;
  assign \new_[623]_  = \new_[4181]_  & \new_[4172]_ ;
  assign \new_[624]_  = \new_[4165]_  & \new_[4156]_ ;
  assign \new_[625]_  = \new_[4149]_  & \new_[4140]_ ;
  assign \new_[626]_  = \new_[4133]_  & \new_[4124]_ ;
  assign \new_[627]_  = \new_[4117]_  & \new_[4108]_ ;
  assign \new_[628]_  = \new_[4101]_  & \new_[4092]_ ;
  assign \new_[629]_  = \new_[4085]_  & \new_[4076]_ ;
  assign \new_[630]_  = \new_[4069]_  & \new_[4060]_ ;
  assign \new_[631]_  = \new_[4053]_  & \new_[4044]_ ;
  assign \new_[632]_  = \new_[4037]_  & \new_[4028]_ ;
  assign \new_[633]_  = \new_[4021]_  & \new_[4012]_ ;
  assign \new_[634]_  = \new_[4005]_  & \new_[3996]_ ;
  assign \new_[635]_  = \new_[3989]_  & \new_[3980]_ ;
  assign \new_[636]_  = \new_[3973]_  & \new_[3964]_ ;
  assign \new_[637]_  = \new_[3957]_  & \new_[3950]_ ;
  assign \new_[638]_  = \new_[3943]_  & \new_[3936]_ ;
  assign \new_[639]_  = \new_[3929]_  & \new_[3922]_ ;
  assign \new_[640]_  = \new_[3915]_  & \new_[3908]_ ;
  assign \new_[641]_  = \new_[3901]_  & \new_[3894]_ ;
  assign \new_[642]_  = \new_[3887]_  & \new_[3880]_ ;
  assign \new_[643]_  = \new_[3873]_  & \new_[3866]_ ;
  assign \new_[644]_  = \new_[3859]_  & \new_[3852]_ ;
  assign \new_[645]_  = \new_[3845]_  & \new_[3838]_ ;
  assign \new_[646]_  = \new_[3831]_  & \new_[3824]_ ;
  assign \new_[647]_  = \new_[3817]_  & \new_[3810]_ ;
  assign \new_[648]_  = \new_[3803]_  & \new_[3796]_ ;
  assign \new_[649]_  = \new_[3789]_  & \new_[3782]_ ;
  assign \new_[650]_  = \new_[3775]_  & \new_[3768]_ ;
  assign \new_[651]_  = \new_[3761]_  & \new_[3754]_ ;
  assign \new_[652]_  = \new_[3747]_  & \new_[3740]_ ;
  assign \new_[653]_  = \new_[3733]_  & \new_[3726]_ ;
  assign \new_[654]_  = \new_[3719]_  & \new_[3712]_ ;
  assign \new_[655]_  = \new_[3705]_  & \new_[3698]_ ;
  assign \new_[656]_  = \new_[3691]_  & \new_[3684]_ ;
  assign \new_[657]_  = \new_[3677]_  & \new_[3670]_ ;
  assign \new_[658]_  = \new_[3663]_  & \new_[3656]_ ;
  assign \new_[659]_  = \new_[3649]_  & \new_[3642]_ ;
  assign \new_[660]_  = \new_[3635]_  & \new_[3628]_ ;
  assign \new_[661]_  = \new_[3621]_  & \new_[3614]_ ;
  assign \new_[662]_  = \new_[3607]_  & \new_[3600]_ ;
  assign \new_[663]_  = \new_[3593]_  & \new_[3586]_ ;
  assign \new_[664]_  = \new_[3579]_  & \new_[3572]_ ;
  assign \new_[665]_  = \new_[3565]_  & \new_[3558]_ ;
  assign \new_[666]_  = \new_[3551]_  & \new_[3544]_ ;
  assign \new_[667]_  = \new_[3537]_  & \new_[3530]_ ;
  assign \new_[668]_  = \new_[3523]_  & \new_[3516]_ ;
  assign \new_[669]_  = \new_[3509]_  & \new_[3502]_ ;
  assign \new_[670]_  = \new_[3495]_  & \new_[3488]_ ;
  assign \new_[671]_  = \new_[3481]_  & \new_[3474]_ ;
  assign \new_[672]_  = \new_[3467]_  & \new_[3460]_ ;
  assign \new_[673]_  = \new_[3453]_  & \new_[3446]_ ;
  assign \new_[674]_  = \new_[3439]_  & \new_[3432]_ ;
  assign \new_[675]_  = \new_[3425]_  & \new_[3418]_ ;
  assign \new_[676]_  = \new_[3411]_  & \new_[3404]_ ;
  assign \new_[677]_  = \new_[3397]_  & \new_[3390]_ ;
  assign \new_[678]_  = \new_[3383]_  & \new_[3376]_ ;
  assign \new_[679]_  = \new_[3369]_  & \new_[3362]_ ;
  assign \new_[680]_  = \new_[3355]_  & \new_[3348]_ ;
  assign \new_[681]_  = \new_[3341]_  & \new_[3334]_ ;
  assign \new_[682]_  = \new_[3327]_  & \new_[3320]_ ;
  assign \new_[683]_  = \new_[3313]_  & \new_[3306]_ ;
  assign \new_[684]_  = \new_[3299]_  & \new_[3292]_ ;
  assign \new_[685]_  = \new_[3285]_  & \new_[3278]_ ;
  assign \new_[686]_  = \new_[3271]_  & \new_[3264]_ ;
  assign \new_[687]_  = \new_[3257]_  & \new_[3250]_ ;
  assign \new_[688]_  = \new_[3243]_  & \new_[3236]_ ;
  assign \new_[689]_  = \new_[3229]_  & \new_[3222]_ ;
  assign \new_[690]_  = \new_[3215]_  & \new_[3208]_ ;
  assign \new_[691]_  = \new_[3201]_  & \new_[3194]_ ;
  assign \new_[692]_  = \new_[3187]_  & \new_[3180]_ ;
  assign \new_[693]_  = \new_[3173]_  & \new_[3166]_ ;
  assign \new_[694]_  = \new_[3159]_  & \new_[3152]_ ;
  assign \new_[695]_  = \new_[3145]_  & \new_[3138]_ ;
  assign \new_[696]_  = \new_[3131]_  & \new_[3124]_ ;
  assign \new_[697]_  = \new_[3117]_  & \new_[3110]_ ;
  assign \new_[698]_  = \new_[3103]_  & \new_[3096]_ ;
  assign \new_[699]_  = \new_[3089]_  & \new_[3082]_ ;
  assign \new_[700]_  = \new_[3075]_  & \new_[3068]_ ;
  assign \new_[701]_  = \new_[3061]_  & \new_[3054]_ ;
  assign \new_[702]_  = \new_[3047]_  & \new_[3040]_ ;
  assign \new_[703]_  = \new_[3033]_  & \new_[3026]_ ;
  assign \new_[704]_  = \new_[3019]_  & \new_[3012]_ ;
  assign \new_[705]_  = \new_[3005]_  & \new_[2998]_ ;
  assign \new_[706]_  = \new_[2991]_  & \new_[2984]_ ;
  assign \new_[707]_  = \new_[2977]_  & \new_[2970]_ ;
  assign \new_[708]_  = \new_[2963]_  & \new_[2956]_ ;
  assign \new_[709]_  = \new_[2949]_  & \new_[2942]_ ;
  assign \new_[710]_  = \new_[2935]_  & \new_[2928]_ ;
  assign \new_[711]_  = \new_[2921]_  & \new_[2914]_ ;
  assign \new_[712]_  = \new_[2907]_  & \new_[2900]_ ;
  assign \new_[713]_  = \new_[2893]_  & \new_[2886]_ ;
  assign \new_[714]_  = \new_[2879]_  & \new_[2872]_ ;
  assign \new_[715]_  = \new_[2865]_  & \new_[2858]_ ;
  assign \new_[716]_  = \new_[2851]_  & \new_[2844]_ ;
  assign \new_[717]_  = \new_[2837]_  & \new_[2830]_ ;
  assign \new_[718]_  = \new_[2823]_  & \new_[2816]_ ;
  assign \new_[719]_  = \new_[2809]_  & \new_[2802]_ ;
  assign \new_[720]_  = \new_[2795]_  & \new_[2788]_ ;
  assign \new_[721]_  = \new_[2781]_  & \new_[2774]_ ;
  assign \new_[722]_  = \new_[2769]_  & \new_[2762]_ ;
  assign \new_[723]_  = \new_[2757]_  & \new_[2750]_ ;
  assign \new_[724]_  = \new_[2745]_  & \new_[2738]_ ;
  assign \new_[725]_  = \new_[2733]_  & \new_[2726]_ ;
  assign \new_[726]_  = \new_[2721]_  & \new_[2714]_ ;
  assign \new_[727]_  = \new_[2709]_  & \new_[2702]_ ;
  assign \new_[728]_  = \new_[2697]_  & \new_[2690]_ ;
  assign \new_[729]_  = \new_[2685]_  & \new_[2678]_ ;
  assign \new_[730]_  = \new_[2673]_  & \new_[2666]_ ;
  assign \new_[731]_  = \new_[2661]_  & \new_[2654]_ ;
  assign \new_[732]_  = \new_[2649]_  & \new_[2642]_ ;
  assign \new_[733]_  = \new_[2637]_  & \new_[2630]_ ;
  assign \new_[734]_  = \new_[2625]_  & \new_[2618]_ ;
  assign \new_[735]_  = \new_[2613]_  & \new_[2606]_ ;
  assign \new_[736]_  = \new_[2601]_  & \new_[2594]_ ;
  assign \new_[737]_  = \new_[2589]_  & \new_[2582]_ ;
  assign \new_[738]_  = \new_[2577]_  & \new_[2570]_ ;
  assign \new_[739]_  = \new_[2565]_  & \new_[2558]_ ;
  assign \new_[740]_  = \new_[2553]_  & \new_[2546]_ ;
  assign \new_[741]_  = \new_[2541]_  & \new_[2534]_ ;
  assign \new_[742]_  = \new_[2529]_  & \new_[2522]_ ;
  assign \new_[743]_  = \new_[2517]_  & \new_[2510]_ ;
  assign \new_[744]_  = \new_[2505]_  & \new_[2498]_ ;
  assign \new_[745]_  = \new_[2493]_  & \new_[2486]_ ;
  assign \new_[746]_  = \new_[2481]_  & \new_[2474]_ ;
  assign \new_[747]_  = \new_[2469]_  & \new_[2462]_ ;
  assign \new_[748]_  = \new_[2457]_  & \new_[2450]_ ;
  assign \new_[749]_  = \new_[2445]_  & \new_[2440]_ ;
  assign \new_[750]_  = \new_[2435]_  & \new_[2430]_ ;
  assign \new_[751]_  = \new_[2425]_  & \new_[2420]_ ;
  assign \new_[752]_  = \new_[2415]_  & \new_[2410]_ ;
  assign \new_[753]_  = \new_[2405]_  & \new_[2400]_ ;
  assign \new_[754]_  = \new_[2395]_  & \new_[2390]_ ;
  assign \new_[755]_  = \new_[2385]_  & \new_[2380]_ ;
  assign \new_[756]_  = \new_[2375]_  & \new_[2370]_ ;
  assign \new_[757]_  = \new_[2365]_  & \new_[2360]_ ;
  assign \new_[758]_  = \new_[2355]_  & \new_[2350]_ ;
  assign \new_[759]_  = \new_[2345]_  & \new_[2340]_ ;
  assign \new_[760]_  = \new_[2337]_  & \new_[2332]_ ;
  assign \new_[761]_  = \new_[2329]_  & \new_[2324]_ ;
  assign \new_[762]_  = \new_[2321]_  & \new_[2316]_ ;
  assign \new_[763]_  = \new_[2313]_  & \new_[2308]_ ;
  assign \new_[764]_  = \new_[2305]_  & \new_[2302]_ ;
  assign \new_[765]_  = \new_[2299]_  & \new_[2296]_ ;
  assign \new_[768]_  = \new_[764]_  | \new_[765]_ ;
  assign \new_[772]_  = \new_[761]_  | \new_[762]_ ;
  assign \new_[773]_  = \new_[763]_  | \new_[772]_ ;
  assign \new_[774]_  = \new_[773]_  | \new_[768]_ ;
  assign \new_[778]_  = \new_[758]_  | \new_[759]_ ;
  assign \new_[779]_  = \new_[760]_  | \new_[778]_ ;
  assign \new_[783]_  = \new_[755]_  | \new_[756]_ ;
  assign \new_[784]_  = \new_[757]_  | \new_[783]_ ;
  assign \new_[785]_  = \new_[784]_  | \new_[779]_ ;
  assign \new_[786]_  = \new_[785]_  | \new_[774]_ ;
  assign \new_[790]_  = \new_[752]_  | \new_[753]_ ;
  assign \new_[791]_  = \new_[754]_  | \new_[790]_ ;
  assign \new_[795]_  = \new_[749]_  | \new_[750]_ ;
  assign \new_[796]_  = \new_[751]_  | \new_[795]_ ;
  assign \new_[797]_  = \new_[796]_  | \new_[791]_ ;
  assign \new_[801]_  = \new_[746]_  | \new_[747]_ ;
  assign \new_[802]_  = \new_[748]_  | \new_[801]_ ;
  assign \new_[806]_  = \new_[743]_  | \new_[744]_ ;
  assign \new_[807]_  = \new_[745]_  | \new_[806]_ ;
  assign \new_[808]_  = \new_[807]_  | \new_[802]_ ;
  assign \new_[809]_  = \new_[808]_  | \new_[797]_ ;
  assign \new_[810]_  = \new_[809]_  | \new_[786]_ ;
  assign \new_[814]_  = \new_[740]_  | \new_[741]_ ;
  assign \new_[815]_  = \new_[742]_  | \new_[814]_ ;
  assign \new_[819]_  = \new_[737]_  | \new_[738]_ ;
  assign \new_[820]_  = \new_[739]_  | \new_[819]_ ;
  assign \new_[821]_  = \new_[820]_  | \new_[815]_ ;
  assign \new_[825]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[826]_  = \new_[736]_  | \new_[825]_ ;
  assign \new_[830]_  = \new_[731]_  | \new_[732]_ ;
  assign \new_[831]_  = \new_[733]_  | \new_[830]_ ;
  assign \new_[832]_  = \new_[831]_  | \new_[826]_ ;
  assign \new_[833]_  = \new_[832]_  | \new_[821]_ ;
  assign \new_[837]_  = \new_[728]_  | \new_[729]_ ;
  assign \new_[838]_  = \new_[730]_  | \new_[837]_ ;
  assign \new_[842]_  = \new_[725]_  | \new_[726]_ ;
  assign \new_[843]_  = \new_[727]_  | \new_[842]_ ;
  assign \new_[844]_  = \new_[843]_  | \new_[838]_ ;
  assign \new_[848]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[849]_  = \new_[724]_  | \new_[848]_ ;
  assign \new_[853]_  = \new_[719]_  | \new_[720]_ ;
  assign \new_[854]_  = \new_[721]_  | \new_[853]_ ;
  assign \new_[855]_  = \new_[854]_  | \new_[849]_ ;
  assign \new_[856]_  = \new_[855]_  | \new_[844]_ ;
  assign \new_[857]_  = \new_[856]_  | \new_[833]_ ;
  assign \new_[858]_  = \new_[857]_  | \new_[810]_ ;
  assign \new_[862]_  = \new_[716]_  | \new_[717]_ ;
  assign \new_[863]_  = \new_[718]_  | \new_[862]_ ;
  assign \new_[867]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[868]_  = \new_[715]_  | \new_[867]_ ;
  assign \new_[869]_  = \new_[868]_  | \new_[863]_ ;
  assign \new_[873]_  = \new_[710]_  | \new_[711]_ ;
  assign \new_[874]_  = \new_[712]_  | \new_[873]_ ;
  assign \new_[878]_  = \new_[707]_  | \new_[708]_ ;
  assign \new_[879]_  = \new_[709]_  | \new_[878]_ ;
  assign \new_[880]_  = \new_[879]_  | \new_[874]_ ;
  assign \new_[881]_  = \new_[880]_  | \new_[869]_ ;
  assign \new_[885]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[886]_  = \new_[706]_  | \new_[885]_ ;
  assign \new_[890]_  = \new_[701]_  | \new_[702]_ ;
  assign \new_[891]_  = \new_[703]_  | \new_[890]_ ;
  assign \new_[892]_  = \new_[891]_  | \new_[886]_ ;
  assign \new_[896]_  = \new_[698]_  | \new_[699]_ ;
  assign \new_[897]_  = \new_[700]_  | \new_[896]_ ;
  assign \new_[901]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[902]_  = \new_[697]_  | \new_[901]_ ;
  assign \new_[903]_  = \new_[902]_  | \new_[897]_ ;
  assign \new_[904]_  = \new_[903]_  | \new_[892]_ ;
  assign \new_[905]_  = \new_[904]_  | \new_[881]_ ;
  assign \new_[909]_  = \new_[692]_  | \new_[693]_ ;
  assign \new_[910]_  = \new_[694]_  | \new_[909]_ ;
  assign \new_[914]_  = \new_[689]_  | \new_[690]_ ;
  assign \new_[915]_  = \new_[691]_  | \new_[914]_ ;
  assign \new_[916]_  = \new_[915]_  | \new_[910]_ ;
  assign \new_[920]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[921]_  = \new_[688]_  | \new_[920]_ ;
  assign \new_[925]_  = \new_[683]_  | \new_[684]_ ;
  assign \new_[926]_  = \new_[685]_  | \new_[925]_ ;
  assign \new_[927]_  = \new_[926]_  | \new_[921]_ ;
  assign \new_[928]_  = \new_[927]_  | \new_[916]_ ;
  assign \new_[932]_  = \new_[680]_  | \new_[681]_ ;
  assign \new_[933]_  = \new_[682]_  | \new_[932]_ ;
  assign \new_[937]_  = \new_[677]_  | \new_[678]_ ;
  assign \new_[938]_  = \new_[679]_  | \new_[937]_ ;
  assign \new_[939]_  = \new_[938]_  | \new_[933]_ ;
  assign \new_[943]_  = \new_[674]_  | \new_[675]_ ;
  assign \new_[944]_  = \new_[676]_  | \new_[943]_ ;
  assign \new_[948]_  = \new_[671]_  | \new_[672]_ ;
  assign \new_[949]_  = \new_[673]_  | \new_[948]_ ;
  assign \new_[950]_  = \new_[949]_  | \new_[944]_ ;
  assign \new_[951]_  = \new_[950]_  | \new_[939]_ ;
  assign \new_[952]_  = \new_[951]_  | \new_[928]_ ;
  assign \new_[953]_  = \new_[952]_  | \new_[905]_ ;
  assign \new_[954]_  = \new_[953]_  | \new_[858]_ ;
  assign \new_[958]_  = \new_[668]_  | \new_[669]_ ;
  assign \new_[959]_  = \new_[670]_  | \new_[958]_ ;
  assign \new_[963]_  = \new_[665]_  | \new_[666]_ ;
  assign \new_[964]_  = \new_[667]_  | \new_[963]_ ;
  assign \new_[965]_  = \new_[964]_  | \new_[959]_ ;
  assign \new_[969]_  = \new_[662]_  | \new_[663]_ ;
  assign \new_[970]_  = \new_[664]_  | \new_[969]_ ;
  assign \new_[974]_  = \new_[659]_  | \new_[660]_ ;
  assign \new_[975]_  = \new_[661]_  | \new_[974]_ ;
  assign \new_[976]_  = \new_[975]_  | \new_[970]_ ;
  assign \new_[977]_  = \new_[976]_  | \new_[965]_ ;
  assign \new_[981]_  = \new_[656]_  | \new_[657]_ ;
  assign \new_[982]_  = \new_[658]_  | \new_[981]_ ;
  assign \new_[986]_  = \new_[653]_  | \new_[654]_ ;
  assign \new_[987]_  = \new_[655]_  | \new_[986]_ ;
  assign \new_[988]_  = \new_[987]_  | \new_[982]_ ;
  assign \new_[992]_  = \new_[650]_  | \new_[651]_ ;
  assign \new_[993]_  = \new_[652]_  | \new_[992]_ ;
  assign \new_[997]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[998]_  = \new_[649]_  | \new_[997]_ ;
  assign \new_[999]_  = \new_[998]_  | \new_[993]_ ;
  assign \new_[1000]_  = \new_[999]_  | \new_[988]_ ;
  assign \new_[1001]_  = \new_[1000]_  | \new_[977]_ ;
  assign \new_[1005]_  = \new_[644]_  | \new_[645]_ ;
  assign \new_[1006]_  = \new_[646]_  | \new_[1005]_ ;
  assign \new_[1010]_  = \new_[641]_  | \new_[642]_ ;
  assign \new_[1011]_  = \new_[643]_  | \new_[1010]_ ;
  assign \new_[1012]_  = \new_[1011]_  | \new_[1006]_ ;
  assign \new_[1016]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[1017]_  = \new_[640]_  | \new_[1016]_ ;
  assign \new_[1021]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[1022]_  = \new_[637]_  | \new_[1021]_ ;
  assign \new_[1023]_  = \new_[1022]_  | \new_[1017]_ ;
  assign \new_[1024]_  = \new_[1023]_  | \new_[1012]_ ;
  assign \new_[1028]_  = \new_[632]_  | \new_[633]_ ;
  assign \new_[1029]_  = \new_[634]_  | \new_[1028]_ ;
  assign \new_[1033]_  = \new_[629]_  | \new_[630]_ ;
  assign \new_[1034]_  = \new_[631]_  | \new_[1033]_ ;
  assign \new_[1035]_  = \new_[1034]_  | \new_[1029]_ ;
  assign \new_[1039]_  = \new_[626]_  | \new_[627]_ ;
  assign \new_[1040]_  = \new_[628]_  | \new_[1039]_ ;
  assign \new_[1044]_  = \new_[623]_  | \new_[624]_ ;
  assign \new_[1045]_  = \new_[625]_  | \new_[1044]_ ;
  assign \new_[1046]_  = \new_[1045]_  | \new_[1040]_ ;
  assign \new_[1047]_  = \new_[1046]_  | \new_[1035]_ ;
  assign \new_[1048]_  = \new_[1047]_  | \new_[1024]_ ;
  assign \new_[1049]_  = \new_[1048]_  | \new_[1001]_ ;
  assign \new_[1053]_  = \new_[620]_  | \new_[621]_ ;
  assign \new_[1054]_  = \new_[622]_  | \new_[1053]_ ;
  assign \new_[1058]_  = \new_[617]_  | \new_[618]_ ;
  assign \new_[1059]_  = \new_[619]_  | \new_[1058]_ ;
  assign \new_[1060]_  = \new_[1059]_  | \new_[1054]_ ;
  assign \new_[1064]_  = \new_[614]_  | \new_[615]_ ;
  assign \new_[1065]_  = \new_[616]_  | \new_[1064]_ ;
  assign \new_[1069]_  = \new_[611]_  | \new_[612]_ ;
  assign \new_[1070]_  = \new_[613]_  | \new_[1069]_ ;
  assign \new_[1071]_  = \new_[1070]_  | \new_[1065]_ ;
  assign \new_[1072]_  = \new_[1071]_  | \new_[1060]_ ;
  assign \new_[1076]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[1077]_  = \new_[610]_  | \new_[1076]_ ;
  assign \new_[1081]_  = \new_[605]_  | \new_[606]_ ;
  assign \new_[1082]_  = \new_[607]_  | \new_[1081]_ ;
  assign \new_[1083]_  = \new_[1082]_  | \new_[1077]_ ;
  assign \new_[1087]_  = \new_[602]_  | \new_[603]_ ;
  assign \new_[1088]_  = \new_[604]_  | \new_[1087]_ ;
  assign \new_[1092]_  = \new_[599]_  | \new_[600]_ ;
  assign \new_[1093]_  = \new_[601]_  | \new_[1092]_ ;
  assign \new_[1094]_  = \new_[1093]_  | \new_[1088]_ ;
  assign \new_[1095]_  = \new_[1094]_  | \new_[1083]_ ;
  assign \new_[1096]_  = \new_[1095]_  | \new_[1072]_ ;
  assign \new_[1100]_  = \new_[596]_  | \new_[597]_ ;
  assign \new_[1101]_  = \new_[598]_  | \new_[1100]_ ;
  assign \new_[1105]_  = \new_[593]_  | \new_[594]_ ;
  assign \new_[1106]_  = \new_[595]_  | \new_[1105]_ ;
  assign \new_[1107]_  = \new_[1106]_  | \new_[1101]_ ;
  assign \new_[1111]_  = \new_[590]_  | \new_[591]_ ;
  assign \new_[1112]_  = \new_[592]_  | \new_[1111]_ ;
  assign \new_[1116]_  = \new_[587]_  | \new_[588]_ ;
  assign \new_[1117]_  = \new_[589]_  | \new_[1116]_ ;
  assign \new_[1118]_  = \new_[1117]_  | \new_[1112]_ ;
  assign \new_[1119]_  = \new_[1118]_  | \new_[1107]_ ;
  assign \new_[1123]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[1124]_  = \new_[586]_  | \new_[1123]_ ;
  assign \new_[1128]_  = \new_[581]_  | \new_[582]_ ;
  assign \new_[1129]_  = \new_[583]_  | \new_[1128]_ ;
  assign \new_[1130]_  = \new_[1129]_  | \new_[1124]_ ;
  assign \new_[1134]_  = \new_[578]_  | \new_[579]_ ;
  assign \new_[1135]_  = \new_[580]_  | \new_[1134]_ ;
  assign \new_[1139]_  = \new_[575]_  | \new_[576]_ ;
  assign \new_[1140]_  = \new_[577]_  | \new_[1139]_ ;
  assign \new_[1141]_  = \new_[1140]_  | \new_[1135]_ ;
  assign \new_[1142]_  = \new_[1141]_  | \new_[1130]_ ;
  assign \new_[1143]_  = \new_[1142]_  | \new_[1119]_ ;
  assign \new_[1144]_  = \new_[1143]_  | \new_[1096]_ ;
  assign \new_[1145]_  = \new_[1144]_  | \new_[1049]_ ;
  assign \new_[1146]_  = \new_[1145]_  | \new_[954]_ ;
  assign \new_[1149]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[1153]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[1154]_  = \new_[572]_  | \new_[1153]_ ;
  assign \new_[1155]_  = \new_[1154]_  | \new_[1149]_ ;
  assign \new_[1159]_  = \new_[567]_  | \new_[568]_ ;
  assign \new_[1160]_  = \new_[569]_  | \new_[1159]_ ;
  assign \new_[1164]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[1165]_  = \new_[566]_  | \new_[1164]_ ;
  assign \new_[1166]_  = \new_[1165]_  | \new_[1160]_ ;
  assign \new_[1167]_  = \new_[1166]_  | \new_[1155]_ ;
  assign \new_[1171]_  = \new_[561]_  | \new_[562]_ ;
  assign \new_[1172]_  = \new_[563]_  | \new_[1171]_ ;
  assign \new_[1176]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[1177]_  = \new_[560]_  | \new_[1176]_ ;
  assign \new_[1178]_  = \new_[1177]_  | \new_[1172]_ ;
  assign \new_[1182]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[1183]_  = \new_[557]_  | \new_[1182]_ ;
  assign \new_[1187]_  = \new_[552]_  | \new_[553]_ ;
  assign \new_[1188]_  = \new_[554]_  | \new_[1187]_ ;
  assign \new_[1189]_  = \new_[1188]_  | \new_[1183]_ ;
  assign \new_[1190]_  = \new_[1189]_  | \new_[1178]_ ;
  assign \new_[1191]_  = \new_[1190]_  | \new_[1167]_ ;
  assign \new_[1195]_  = \new_[549]_  | \new_[550]_ ;
  assign \new_[1196]_  = \new_[551]_  | \new_[1195]_ ;
  assign \new_[1200]_  = \new_[546]_  | \new_[547]_ ;
  assign \new_[1201]_  = \new_[548]_  | \new_[1200]_ ;
  assign \new_[1202]_  = \new_[1201]_  | \new_[1196]_ ;
  assign \new_[1206]_  = \new_[543]_  | \new_[544]_ ;
  assign \new_[1207]_  = \new_[545]_  | \new_[1206]_ ;
  assign \new_[1211]_  = \new_[540]_  | \new_[541]_ ;
  assign \new_[1212]_  = \new_[542]_  | \new_[1211]_ ;
  assign \new_[1213]_  = \new_[1212]_  | \new_[1207]_ ;
  assign \new_[1214]_  = \new_[1213]_  | \new_[1202]_ ;
  assign \new_[1218]_  = \new_[537]_  | \new_[538]_ ;
  assign \new_[1219]_  = \new_[539]_  | \new_[1218]_ ;
  assign \new_[1223]_  = \new_[534]_  | \new_[535]_ ;
  assign \new_[1224]_  = \new_[536]_  | \new_[1223]_ ;
  assign \new_[1225]_  = \new_[1224]_  | \new_[1219]_ ;
  assign \new_[1229]_  = \new_[531]_  | \new_[532]_ ;
  assign \new_[1230]_  = \new_[533]_  | \new_[1229]_ ;
  assign \new_[1234]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[1235]_  = \new_[530]_  | \new_[1234]_ ;
  assign \new_[1236]_  = \new_[1235]_  | \new_[1230]_ ;
  assign \new_[1237]_  = \new_[1236]_  | \new_[1225]_ ;
  assign \new_[1238]_  = \new_[1237]_  | \new_[1214]_ ;
  assign \new_[1239]_  = \new_[1238]_  | \new_[1191]_ ;
  assign \new_[1243]_  = \new_[525]_  | \new_[526]_ ;
  assign \new_[1244]_  = \new_[527]_  | \new_[1243]_ ;
  assign \new_[1248]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[1249]_  = \new_[524]_  | \new_[1248]_ ;
  assign \new_[1250]_  = \new_[1249]_  | \new_[1244]_ ;
  assign \new_[1254]_  = \new_[519]_  | \new_[520]_ ;
  assign \new_[1255]_  = \new_[521]_  | \new_[1254]_ ;
  assign \new_[1259]_  = \new_[516]_  | \new_[517]_ ;
  assign \new_[1260]_  = \new_[518]_  | \new_[1259]_ ;
  assign \new_[1261]_  = \new_[1260]_  | \new_[1255]_ ;
  assign \new_[1262]_  = \new_[1261]_  | \new_[1250]_ ;
  assign \new_[1266]_  = \new_[513]_  | \new_[514]_ ;
  assign \new_[1267]_  = \new_[515]_  | \new_[1266]_ ;
  assign \new_[1271]_  = \new_[510]_  | \new_[511]_ ;
  assign \new_[1272]_  = \new_[512]_  | \new_[1271]_ ;
  assign \new_[1273]_  = \new_[1272]_  | \new_[1267]_ ;
  assign \new_[1277]_  = \new_[507]_  | \new_[508]_ ;
  assign \new_[1278]_  = \new_[509]_  | \new_[1277]_ ;
  assign \new_[1282]_  = \new_[504]_  | \new_[505]_ ;
  assign \new_[1283]_  = \new_[506]_  | \new_[1282]_ ;
  assign \new_[1284]_  = \new_[1283]_  | \new_[1278]_ ;
  assign \new_[1285]_  = \new_[1284]_  | \new_[1273]_ ;
  assign \new_[1286]_  = \new_[1285]_  | \new_[1262]_ ;
  assign \new_[1290]_  = \new_[501]_  | \new_[502]_ ;
  assign \new_[1291]_  = \new_[503]_  | \new_[1290]_ ;
  assign \new_[1295]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[1296]_  = \new_[500]_  | \new_[1295]_ ;
  assign \new_[1297]_  = \new_[1296]_  | \new_[1291]_ ;
  assign \new_[1301]_  = \new_[495]_  | \new_[496]_ ;
  assign \new_[1302]_  = \new_[497]_  | \new_[1301]_ ;
  assign \new_[1306]_  = \new_[492]_  | \new_[493]_ ;
  assign \new_[1307]_  = \new_[494]_  | \new_[1306]_ ;
  assign \new_[1308]_  = \new_[1307]_  | \new_[1302]_ ;
  assign \new_[1309]_  = \new_[1308]_  | \new_[1297]_ ;
  assign \new_[1313]_  = \new_[489]_  | \new_[490]_ ;
  assign \new_[1314]_  = \new_[491]_  | \new_[1313]_ ;
  assign \new_[1318]_  = \new_[486]_  | \new_[487]_ ;
  assign \new_[1319]_  = \new_[488]_  | \new_[1318]_ ;
  assign \new_[1320]_  = \new_[1319]_  | \new_[1314]_ ;
  assign \new_[1324]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[1325]_  = \new_[485]_  | \new_[1324]_ ;
  assign \new_[1329]_  = \new_[480]_  | \new_[481]_ ;
  assign \new_[1330]_  = \new_[482]_  | \new_[1329]_ ;
  assign \new_[1331]_  = \new_[1330]_  | \new_[1325]_ ;
  assign \new_[1332]_  = \new_[1331]_  | \new_[1320]_ ;
  assign \new_[1333]_  = \new_[1332]_  | \new_[1309]_ ;
  assign \new_[1334]_  = \new_[1333]_  | \new_[1286]_ ;
  assign \new_[1335]_  = \new_[1334]_  | \new_[1239]_ ;
  assign \new_[1339]_  = \new_[477]_  | \new_[478]_ ;
  assign \new_[1340]_  = \new_[479]_  | \new_[1339]_ ;
  assign \new_[1344]_  = \new_[474]_  | \new_[475]_ ;
  assign \new_[1345]_  = \new_[476]_  | \new_[1344]_ ;
  assign \new_[1346]_  = \new_[1345]_  | \new_[1340]_ ;
  assign \new_[1350]_  = \new_[471]_  | \new_[472]_ ;
  assign \new_[1351]_  = \new_[473]_  | \new_[1350]_ ;
  assign \new_[1355]_  = \new_[468]_  | \new_[469]_ ;
  assign \new_[1356]_  = \new_[470]_  | \new_[1355]_ ;
  assign \new_[1357]_  = \new_[1356]_  | \new_[1351]_ ;
  assign \new_[1358]_  = \new_[1357]_  | \new_[1346]_ ;
  assign \new_[1362]_  = \new_[465]_  | \new_[466]_ ;
  assign \new_[1363]_  = \new_[467]_  | \new_[1362]_ ;
  assign \new_[1367]_  = \new_[462]_  | \new_[463]_ ;
  assign \new_[1368]_  = \new_[464]_  | \new_[1367]_ ;
  assign \new_[1369]_  = \new_[1368]_  | \new_[1363]_ ;
  assign \new_[1373]_  = \new_[459]_  | \new_[460]_ ;
  assign \new_[1374]_  = \new_[461]_  | \new_[1373]_ ;
  assign \new_[1378]_  = \new_[456]_  | \new_[457]_ ;
  assign \new_[1379]_  = \new_[458]_  | \new_[1378]_ ;
  assign \new_[1380]_  = \new_[1379]_  | \new_[1374]_ ;
  assign \new_[1381]_  = \new_[1380]_  | \new_[1369]_ ;
  assign \new_[1382]_  = \new_[1381]_  | \new_[1358]_ ;
  assign \new_[1386]_  = \new_[453]_  | \new_[454]_ ;
  assign \new_[1387]_  = \new_[455]_  | \new_[1386]_ ;
  assign \new_[1391]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[1392]_  = \new_[452]_  | \new_[1391]_ ;
  assign \new_[1393]_  = \new_[1392]_  | \new_[1387]_ ;
  assign \new_[1397]_  = \new_[447]_  | \new_[448]_ ;
  assign \new_[1398]_  = \new_[449]_  | \new_[1397]_ ;
  assign \new_[1402]_  = \new_[444]_  | \new_[445]_ ;
  assign \new_[1403]_  = \new_[446]_  | \new_[1402]_ ;
  assign \new_[1404]_  = \new_[1403]_  | \new_[1398]_ ;
  assign \new_[1405]_  = \new_[1404]_  | \new_[1393]_ ;
  assign \new_[1409]_  = \new_[441]_  | \new_[442]_ ;
  assign \new_[1410]_  = \new_[443]_  | \new_[1409]_ ;
  assign \new_[1414]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[1415]_  = \new_[440]_  | \new_[1414]_ ;
  assign \new_[1416]_  = \new_[1415]_  | \new_[1410]_ ;
  assign \new_[1420]_  = \new_[435]_  | \new_[436]_ ;
  assign \new_[1421]_  = \new_[437]_  | \new_[1420]_ ;
  assign \new_[1425]_  = \new_[432]_  | \new_[433]_ ;
  assign \new_[1426]_  = \new_[434]_  | \new_[1425]_ ;
  assign \new_[1427]_  = \new_[1426]_  | \new_[1421]_ ;
  assign \new_[1428]_  = \new_[1427]_  | \new_[1416]_ ;
  assign \new_[1429]_  = \new_[1428]_  | \new_[1405]_ ;
  assign \new_[1430]_  = \new_[1429]_  | \new_[1382]_ ;
  assign \new_[1434]_  = \new_[429]_  | \new_[430]_ ;
  assign \new_[1435]_  = \new_[431]_  | \new_[1434]_ ;
  assign \new_[1439]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[1440]_  = \new_[428]_  | \new_[1439]_ ;
  assign \new_[1441]_  = \new_[1440]_  | \new_[1435]_ ;
  assign \new_[1445]_  = \new_[423]_  | \new_[424]_ ;
  assign \new_[1446]_  = \new_[425]_  | \new_[1445]_ ;
  assign \new_[1450]_  = \new_[420]_  | \new_[421]_ ;
  assign \new_[1451]_  = \new_[422]_  | \new_[1450]_ ;
  assign \new_[1452]_  = \new_[1451]_  | \new_[1446]_ ;
  assign \new_[1453]_  = \new_[1452]_  | \new_[1441]_ ;
  assign \new_[1457]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[1458]_  = \new_[419]_  | \new_[1457]_ ;
  assign \new_[1462]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[1463]_  = \new_[416]_  | \new_[1462]_ ;
  assign \new_[1464]_  = \new_[1463]_  | \new_[1458]_ ;
  assign \new_[1468]_  = \new_[411]_  | \new_[412]_ ;
  assign \new_[1469]_  = \new_[413]_  | \new_[1468]_ ;
  assign \new_[1473]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[1474]_  = \new_[410]_  | \new_[1473]_ ;
  assign \new_[1475]_  = \new_[1474]_  | \new_[1469]_ ;
  assign \new_[1476]_  = \new_[1475]_  | \new_[1464]_ ;
  assign \new_[1477]_  = \new_[1476]_  | \new_[1453]_ ;
  assign \new_[1481]_  = \new_[405]_  | \new_[406]_ ;
  assign \new_[1482]_  = \new_[407]_  | \new_[1481]_ ;
  assign \new_[1486]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[1487]_  = \new_[404]_  | \new_[1486]_ ;
  assign \new_[1488]_  = \new_[1487]_  | \new_[1482]_ ;
  assign \new_[1492]_  = \new_[399]_  | \new_[400]_ ;
  assign \new_[1493]_  = \new_[401]_  | \new_[1492]_ ;
  assign \new_[1497]_  = \new_[396]_  | \new_[397]_ ;
  assign \new_[1498]_  = \new_[398]_  | \new_[1497]_ ;
  assign \new_[1499]_  = \new_[1498]_  | \new_[1493]_ ;
  assign \new_[1500]_  = \new_[1499]_  | \new_[1488]_ ;
  assign \new_[1504]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[1505]_  = \new_[395]_  | \new_[1504]_ ;
  assign \new_[1509]_  = \new_[390]_  | \new_[391]_ ;
  assign \new_[1510]_  = \new_[392]_  | \new_[1509]_ ;
  assign \new_[1511]_  = \new_[1510]_  | \new_[1505]_ ;
  assign \new_[1515]_  = \new_[387]_  | \new_[388]_ ;
  assign \new_[1516]_  = \new_[389]_  | \new_[1515]_ ;
  assign \new_[1520]_  = \new_[384]_  | \new_[385]_ ;
  assign \new_[1521]_  = \new_[386]_  | \new_[1520]_ ;
  assign \new_[1522]_  = \new_[1521]_  | \new_[1516]_ ;
  assign \new_[1523]_  = \new_[1522]_  | \new_[1511]_ ;
  assign \new_[1524]_  = \new_[1523]_  | \new_[1500]_ ;
  assign \new_[1525]_  = \new_[1524]_  | \new_[1477]_ ;
  assign \new_[1526]_  = \new_[1525]_  | \new_[1430]_ ;
  assign \new_[1527]_  = \new_[1526]_  | \new_[1335]_ ;
  assign \new_[1528]_  = \new_[1527]_  | \new_[1146]_ ;
  assign \new_[1531]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[1535]_  = \new_[379]_  | \new_[380]_ ;
  assign \new_[1536]_  = \new_[381]_  | \new_[1535]_ ;
  assign \new_[1537]_  = \new_[1536]_  | \new_[1531]_ ;
  assign \new_[1541]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[1542]_  = \new_[378]_  | \new_[1541]_ ;
  assign \new_[1546]_  = \new_[373]_  | \new_[374]_ ;
  assign \new_[1547]_  = \new_[375]_  | \new_[1546]_ ;
  assign \new_[1548]_  = \new_[1547]_  | \new_[1542]_ ;
  assign \new_[1549]_  = \new_[1548]_  | \new_[1537]_ ;
  assign \new_[1553]_  = \new_[370]_  | \new_[371]_ ;
  assign \new_[1554]_  = \new_[372]_  | \new_[1553]_ ;
  assign \new_[1558]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[1559]_  = \new_[369]_  | \new_[1558]_ ;
  assign \new_[1560]_  = \new_[1559]_  | \new_[1554]_ ;
  assign \new_[1564]_  = \new_[364]_  | \new_[365]_ ;
  assign \new_[1565]_  = \new_[366]_  | \new_[1564]_ ;
  assign \new_[1569]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[1570]_  = \new_[363]_  | \new_[1569]_ ;
  assign \new_[1571]_  = \new_[1570]_  | \new_[1565]_ ;
  assign \new_[1572]_  = \new_[1571]_  | \new_[1560]_ ;
  assign \new_[1573]_  = \new_[1572]_  | \new_[1549]_ ;
  assign \new_[1577]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[1578]_  = \new_[360]_  | \new_[1577]_ ;
  assign \new_[1582]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[1583]_  = \new_[357]_  | \new_[1582]_ ;
  assign \new_[1584]_  = \new_[1583]_  | \new_[1578]_ ;
  assign \new_[1588]_  = \new_[352]_  | \new_[353]_ ;
  assign \new_[1589]_  = \new_[354]_  | \new_[1588]_ ;
  assign \new_[1593]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[1594]_  = \new_[351]_  | \new_[1593]_ ;
  assign \new_[1595]_  = \new_[1594]_  | \new_[1589]_ ;
  assign \new_[1596]_  = \new_[1595]_  | \new_[1584]_ ;
  assign \new_[1600]_  = \new_[346]_  | \new_[347]_ ;
  assign \new_[1601]_  = \new_[348]_  | \new_[1600]_ ;
  assign \new_[1605]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[1606]_  = \new_[345]_  | \new_[1605]_ ;
  assign \new_[1607]_  = \new_[1606]_  | \new_[1601]_ ;
  assign \new_[1611]_  = \new_[340]_  | \new_[341]_ ;
  assign \new_[1612]_  = \new_[342]_  | \new_[1611]_ ;
  assign \new_[1616]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[1617]_  = \new_[339]_  | \new_[1616]_ ;
  assign \new_[1618]_  = \new_[1617]_  | \new_[1612]_ ;
  assign \new_[1619]_  = \new_[1618]_  | \new_[1607]_ ;
  assign \new_[1620]_  = \new_[1619]_  | \new_[1596]_ ;
  assign \new_[1621]_  = \new_[1620]_  | \new_[1573]_ ;
  assign \new_[1625]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[1626]_  = \new_[336]_  | \new_[1625]_ ;
  assign \new_[1630]_  = \new_[331]_  | \new_[332]_ ;
  assign \new_[1631]_  = \new_[333]_  | \new_[1630]_ ;
  assign \new_[1632]_  = \new_[1631]_  | \new_[1626]_ ;
  assign \new_[1636]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[1637]_  = \new_[330]_  | \new_[1636]_ ;
  assign \new_[1641]_  = \new_[325]_  | \new_[326]_ ;
  assign \new_[1642]_  = \new_[327]_  | \new_[1641]_ ;
  assign \new_[1643]_  = \new_[1642]_  | \new_[1637]_ ;
  assign \new_[1644]_  = \new_[1643]_  | \new_[1632]_ ;
  assign \new_[1648]_  = \new_[322]_  | \new_[323]_ ;
  assign \new_[1649]_  = \new_[324]_  | \new_[1648]_ ;
  assign \new_[1653]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[1654]_  = \new_[321]_  | \new_[1653]_ ;
  assign \new_[1655]_  = \new_[1654]_  | \new_[1649]_ ;
  assign \new_[1659]_  = \new_[316]_  | \new_[317]_ ;
  assign \new_[1660]_  = \new_[318]_  | \new_[1659]_ ;
  assign \new_[1664]_  = \new_[313]_  | \new_[314]_ ;
  assign \new_[1665]_  = \new_[315]_  | \new_[1664]_ ;
  assign \new_[1666]_  = \new_[1665]_  | \new_[1660]_ ;
  assign \new_[1667]_  = \new_[1666]_  | \new_[1655]_ ;
  assign \new_[1668]_  = \new_[1667]_  | \new_[1644]_ ;
  assign \new_[1672]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[1673]_  = \new_[312]_  | \new_[1672]_ ;
  assign \new_[1677]_  = \new_[307]_  | \new_[308]_ ;
  assign \new_[1678]_  = \new_[309]_  | \new_[1677]_ ;
  assign \new_[1679]_  = \new_[1678]_  | \new_[1673]_ ;
  assign \new_[1683]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[1684]_  = \new_[306]_  | \new_[1683]_ ;
  assign \new_[1688]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[1689]_  = \new_[303]_  | \new_[1688]_ ;
  assign \new_[1690]_  = \new_[1689]_  | \new_[1684]_ ;
  assign \new_[1691]_  = \new_[1690]_  | \new_[1679]_ ;
  assign \new_[1695]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[1696]_  = \new_[300]_  | \new_[1695]_ ;
  assign \new_[1700]_  = \new_[295]_  | \new_[296]_ ;
  assign \new_[1701]_  = \new_[297]_  | \new_[1700]_ ;
  assign \new_[1702]_  = \new_[1701]_  | \new_[1696]_ ;
  assign \new_[1706]_  = \new_[292]_  | \new_[293]_ ;
  assign \new_[1707]_  = \new_[294]_  | \new_[1706]_ ;
  assign \new_[1711]_  = \new_[289]_  | \new_[290]_ ;
  assign \new_[1712]_  = \new_[291]_  | \new_[1711]_ ;
  assign \new_[1713]_  = \new_[1712]_  | \new_[1707]_ ;
  assign \new_[1714]_  = \new_[1713]_  | \new_[1702]_ ;
  assign \new_[1715]_  = \new_[1714]_  | \new_[1691]_ ;
  assign \new_[1716]_  = \new_[1715]_  | \new_[1668]_ ;
  assign \new_[1717]_  = \new_[1716]_  | \new_[1621]_ ;
  assign \new_[1721]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[1722]_  = \new_[288]_  | \new_[1721]_ ;
  assign \new_[1726]_  = \new_[283]_  | \new_[284]_ ;
  assign \new_[1727]_  = \new_[285]_  | \new_[1726]_ ;
  assign \new_[1728]_  = \new_[1727]_  | \new_[1722]_ ;
  assign \new_[1732]_  = \new_[280]_  | \new_[281]_ ;
  assign \new_[1733]_  = \new_[282]_  | \new_[1732]_ ;
  assign \new_[1737]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[1738]_  = \new_[279]_  | \new_[1737]_ ;
  assign \new_[1739]_  = \new_[1738]_  | \new_[1733]_ ;
  assign \new_[1740]_  = \new_[1739]_  | \new_[1728]_ ;
  assign \new_[1744]_  = \new_[274]_  | \new_[275]_ ;
  assign \new_[1745]_  = \new_[276]_  | \new_[1744]_ ;
  assign \new_[1749]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[1750]_  = \new_[273]_  | \new_[1749]_ ;
  assign \new_[1751]_  = \new_[1750]_  | \new_[1745]_ ;
  assign \new_[1755]_  = \new_[268]_  | \new_[269]_ ;
  assign \new_[1756]_  = \new_[270]_  | \new_[1755]_ ;
  assign \new_[1760]_  = \new_[265]_  | \new_[266]_ ;
  assign \new_[1761]_  = \new_[267]_  | \new_[1760]_ ;
  assign \new_[1762]_  = \new_[1761]_  | \new_[1756]_ ;
  assign \new_[1763]_  = \new_[1762]_  | \new_[1751]_ ;
  assign \new_[1764]_  = \new_[1763]_  | \new_[1740]_ ;
  assign \new_[1768]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[1769]_  = \new_[264]_  | \new_[1768]_ ;
  assign \new_[1773]_  = \new_[259]_  | \new_[260]_ ;
  assign \new_[1774]_  = \new_[261]_  | \new_[1773]_ ;
  assign \new_[1775]_  = \new_[1774]_  | \new_[1769]_ ;
  assign \new_[1779]_  = \new_[256]_  | \new_[257]_ ;
  assign \new_[1780]_  = \new_[258]_  | \new_[1779]_ ;
  assign \new_[1784]_  = \new_[253]_  | \new_[254]_ ;
  assign \new_[1785]_  = \new_[255]_  | \new_[1784]_ ;
  assign \new_[1786]_  = \new_[1785]_  | \new_[1780]_ ;
  assign \new_[1787]_  = \new_[1786]_  | \new_[1775]_ ;
  assign \new_[1791]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[1792]_  = \new_[252]_  | \new_[1791]_ ;
  assign \new_[1796]_  = \new_[247]_  | \new_[248]_ ;
  assign \new_[1797]_  = \new_[249]_  | \new_[1796]_ ;
  assign \new_[1798]_  = \new_[1797]_  | \new_[1792]_ ;
  assign \new_[1802]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[1803]_  = \new_[246]_  | \new_[1802]_ ;
  assign \new_[1807]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[1808]_  = \new_[243]_  | \new_[1807]_ ;
  assign \new_[1809]_  = \new_[1808]_  | \new_[1803]_ ;
  assign \new_[1810]_  = \new_[1809]_  | \new_[1798]_ ;
  assign \new_[1811]_  = \new_[1810]_  | \new_[1787]_ ;
  assign \new_[1812]_  = \new_[1811]_  | \new_[1764]_ ;
  assign \new_[1816]_  = \new_[238]_  | \new_[239]_ ;
  assign \new_[1817]_  = \new_[240]_  | \new_[1816]_ ;
  assign \new_[1821]_  = \new_[235]_  | \new_[236]_ ;
  assign \new_[1822]_  = \new_[237]_  | \new_[1821]_ ;
  assign \new_[1823]_  = \new_[1822]_  | \new_[1817]_ ;
  assign \new_[1827]_  = \new_[232]_  | \new_[233]_ ;
  assign \new_[1828]_  = \new_[234]_  | \new_[1827]_ ;
  assign \new_[1832]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[1833]_  = \new_[231]_  | \new_[1832]_ ;
  assign \new_[1834]_  = \new_[1833]_  | \new_[1828]_ ;
  assign \new_[1835]_  = \new_[1834]_  | \new_[1823]_ ;
  assign \new_[1839]_  = \new_[226]_  | \new_[227]_ ;
  assign \new_[1840]_  = \new_[228]_  | \new_[1839]_ ;
  assign \new_[1844]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[1845]_  = \new_[225]_  | \new_[1844]_ ;
  assign \new_[1846]_  = \new_[1845]_  | \new_[1840]_ ;
  assign \new_[1850]_  = \new_[220]_  | \new_[221]_ ;
  assign \new_[1851]_  = \new_[222]_  | \new_[1850]_ ;
  assign \new_[1855]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[1856]_  = \new_[219]_  | \new_[1855]_ ;
  assign \new_[1857]_  = \new_[1856]_  | \new_[1851]_ ;
  assign \new_[1858]_  = \new_[1857]_  | \new_[1846]_ ;
  assign \new_[1859]_  = \new_[1858]_  | \new_[1835]_ ;
  assign \new_[1863]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[1864]_  = \new_[216]_  | \new_[1863]_ ;
  assign \new_[1868]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[1869]_  = \new_[213]_  | \new_[1868]_ ;
  assign \new_[1870]_  = \new_[1869]_  | \new_[1864]_ ;
  assign \new_[1874]_  = \new_[208]_  | \new_[209]_ ;
  assign \new_[1875]_  = \new_[210]_  | \new_[1874]_ ;
  assign \new_[1879]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[1880]_  = \new_[207]_  | \new_[1879]_ ;
  assign \new_[1881]_  = \new_[1880]_  | \new_[1875]_ ;
  assign \new_[1882]_  = \new_[1881]_  | \new_[1870]_ ;
  assign \new_[1886]_  = \new_[202]_  | \new_[203]_ ;
  assign \new_[1887]_  = \new_[204]_  | \new_[1886]_ ;
  assign \new_[1891]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[1892]_  = \new_[201]_  | \new_[1891]_ ;
  assign \new_[1893]_  = \new_[1892]_  | \new_[1887]_ ;
  assign \new_[1897]_  = \new_[196]_  | \new_[197]_ ;
  assign \new_[1898]_  = \new_[198]_  | \new_[1897]_ ;
  assign \new_[1902]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[1903]_  = \new_[195]_  | \new_[1902]_ ;
  assign \new_[1904]_  = \new_[1903]_  | \new_[1898]_ ;
  assign \new_[1905]_  = \new_[1904]_  | \new_[1893]_ ;
  assign \new_[1906]_  = \new_[1905]_  | \new_[1882]_ ;
  assign \new_[1907]_  = \new_[1906]_  | \new_[1859]_ ;
  assign \new_[1908]_  = \new_[1907]_  | \new_[1812]_ ;
  assign \new_[1909]_  = \new_[1908]_  | \new_[1717]_ ;
  assign \new_[1913]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[1914]_  = \new_[192]_  | \new_[1913]_ ;
  assign \new_[1918]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[1919]_  = \new_[189]_  | \new_[1918]_ ;
  assign \new_[1920]_  = \new_[1919]_  | \new_[1914]_ ;
  assign \new_[1924]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[1925]_  = \new_[186]_  | \new_[1924]_ ;
  assign \new_[1929]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[1930]_  = \new_[183]_  | \new_[1929]_ ;
  assign \new_[1931]_  = \new_[1930]_  | \new_[1925]_ ;
  assign \new_[1932]_  = \new_[1931]_  | \new_[1920]_ ;
  assign \new_[1936]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[1937]_  = \new_[180]_  | \new_[1936]_ ;
  assign \new_[1941]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[1942]_  = \new_[177]_  | \new_[1941]_ ;
  assign \new_[1943]_  = \new_[1942]_  | \new_[1937]_ ;
  assign \new_[1947]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[1948]_  = \new_[174]_  | \new_[1947]_ ;
  assign \new_[1952]_  = \new_[169]_  | \new_[170]_ ;
  assign \new_[1953]_  = \new_[171]_  | \new_[1952]_ ;
  assign \new_[1954]_  = \new_[1953]_  | \new_[1948]_ ;
  assign \new_[1955]_  = \new_[1954]_  | \new_[1943]_ ;
  assign \new_[1956]_  = \new_[1955]_  | \new_[1932]_ ;
  assign \new_[1960]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[1961]_  = \new_[168]_  | \new_[1960]_ ;
  assign \new_[1965]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[1966]_  = \new_[165]_  | \new_[1965]_ ;
  assign \new_[1967]_  = \new_[1966]_  | \new_[1961]_ ;
  assign \new_[1971]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[1972]_  = \new_[162]_  | \new_[1971]_ ;
  assign \new_[1976]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[1977]_  = \new_[159]_  | \new_[1976]_ ;
  assign \new_[1978]_  = \new_[1977]_  | \new_[1972]_ ;
  assign \new_[1979]_  = \new_[1978]_  | \new_[1967]_ ;
  assign \new_[1983]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[1984]_  = \new_[156]_  | \new_[1983]_ ;
  assign \new_[1988]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[1989]_  = \new_[153]_  | \new_[1988]_ ;
  assign \new_[1990]_  = \new_[1989]_  | \new_[1984]_ ;
  assign \new_[1994]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[1995]_  = \new_[150]_  | \new_[1994]_ ;
  assign \new_[1999]_  = \new_[145]_  | \new_[146]_ ;
  assign \new_[2000]_  = \new_[147]_  | \new_[1999]_ ;
  assign \new_[2001]_  = \new_[2000]_  | \new_[1995]_ ;
  assign \new_[2002]_  = \new_[2001]_  | \new_[1990]_ ;
  assign \new_[2003]_  = \new_[2002]_  | \new_[1979]_ ;
  assign \new_[2004]_  = \new_[2003]_  | \new_[1956]_ ;
  assign \new_[2008]_  = \new_[142]_  | \new_[143]_ ;
  assign \new_[2009]_  = \new_[144]_  | \new_[2008]_ ;
  assign \new_[2013]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[2014]_  = \new_[141]_  | \new_[2013]_ ;
  assign \new_[2015]_  = \new_[2014]_  | \new_[2009]_ ;
  assign \new_[2019]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[2020]_  = \new_[138]_  | \new_[2019]_ ;
  assign \new_[2024]_  = \new_[133]_  | \new_[134]_ ;
  assign \new_[2025]_  = \new_[135]_  | \new_[2024]_ ;
  assign \new_[2026]_  = \new_[2025]_  | \new_[2020]_ ;
  assign \new_[2027]_  = \new_[2026]_  | \new_[2015]_ ;
  assign \new_[2031]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[2032]_  = \new_[132]_  | \new_[2031]_ ;
  assign \new_[2036]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[2037]_  = \new_[129]_  | \new_[2036]_ ;
  assign \new_[2038]_  = \new_[2037]_  | \new_[2032]_ ;
  assign \new_[2042]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[2043]_  = \new_[126]_  | \new_[2042]_ ;
  assign \new_[2047]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[2048]_  = \new_[123]_  | \new_[2047]_ ;
  assign \new_[2049]_  = \new_[2048]_  | \new_[2043]_ ;
  assign \new_[2050]_  = \new_[2049]_  | \new_[2038]_ ;
  assign \new_[2051]_  = \new_[2050]_  | \new_[2027]_ ;
  assign \new_[2055]_  = \new_[118]_  | \new_[119]_ ;
  assign \new_[2056]_  = \new_[120]_  | \new_[2055]_ ;
  assign \new_[2060]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[2061]_  = \new_[117]_  | \new_[2060]_ ;
  assign \new_[2062]_  = \new_[2061]_  | \new_[2056]_ ;
  assign \new_[2066]_  = \new_[112]_  | \new_[113]_ ;
  assign \new_[2067]_  = \new_[114]_  | \new_[2066]_ ;
  assign \new_[2071]_  = \new_[109]_  | \new_[110]_ ;
  assign \new_[2072]_  = \new_[111]_  | \new_[2071]_ ;
  assign \new_[2073]_  = \new_[2072]_  | \new_[2067]_ ;
  assign \new_[2074]_  = \new_[2073]_  | \new_[2062]_ ;
  assign \new_[2078]_  = \new_[106]_  | \new_[107]_ ;
  assign \new_[2079]_  = \new_[108]_  | \new_[2078]_ ;
  assign \new_[2083]_  = \new_[103]_  | \new_[104]_ ;
  assign \new_[2084]_  = \new_[105]_  | \new_[2083]_ ;
  assign \new_[2085]_  = \new_[2084]_  | \new_[2079]_ ;
  assign \new_[2089]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[2090]_  = \new_[102]_  | \new_[2089]_ ;
  assign \new_[2094]_  = \new_[97]_  | \new_[98]_ ;
  assign \new_[2095]_  = \new_[99]_  | \new_[2094]_ ;
  assign \new_[2096]_  = \new_[2095]_  | \new_[2090]_ ;
  assign \new_[2097]_  = \new_[2096]_  | \new_[2085]_ ;
  assign \new_[2098]_  = \new_[2097]_  | \new_[2074]_ ;
  assign \new_[2099]_  = \new_[2098]_  | \new_[2051]_ ;
  assign \new_[2100]_  = \new_[2099]_  | \new_[2004]_ ;
  assign \new_[2104]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[2105]_  = \new_[96]_  | \new_[2104]_ ;
  assign \new_[2109]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[2110]_  = \new_[93]_  | \new_[2109]_ ;
  assign \new_[2111]_  = \new_[2110]_  | \new_[2105]_ ;
  assign \new_[2115]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[2116]_  = \new_[90]_  | \new_[2115]_ ;
  assign \new_[2120]_  = \new_[85]_  | \new_[86]_ ;
  assign \new_[2121]_  = \new_[87]_  | \new_[2120]_ ;
  assign \new_[2122]_  = \new_[2121]_  | \new_[2116]_ ;
  assign \new_[2123]_  = \new_[2122]_  | \new_[2111]_ ;
  assign \new_[2127]_  = \new_[82]_  | \new_[83]_ ;
  assign \new_[2128]_  = \new_[84]_  | \new_[2127]_ ;
  assign \new_[2132]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[2133]_  = \new_[81]_  | \new_[2132]_ ;
  assign \new_[2134]_  = \new_[2133]_  | \new_[2128]_ ;
  assign \new_[2138]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[2139]_  = \new_[78]_  | \new_[2138]_ ;
  assign \new_[2143]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[2144]_  = \new_[75]_  | \new_[2143]_ ;
  assign \new_[2145]_  = \new_[2144]_  | \new_[2139]_ ;
  assign \new_[2146]_  = \new_[2145]_  | \new_[2134]_ ;
  assign \new_[2147]_  = \new_[2146]_  | \new_[2123]_ ;
  assign \new_[2151]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[2152]_  = \new_[72]_  | \new_[2151]_ ;
  assign \new_[2156]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[2157]_  = \new_[69]_  | \new_[2156]_ ;
  assign \new_[2158]_  = \new_[2157]_  | \new_[2152]_ ;
  assign \new_[2162]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[2163]_  = \new_[66]_  | \new_[2162]_ ;
  assign \new_[2167]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[2168]_  = \new_[63]_  | \new_[2167]_ ;
  assign \new_[2169]_  = \new_[2168]_  | \new_[2163]_ ;
  assign \new_[2170]_  = \new_[2169]_  | \new_[2158]_ ;
  assign \new_[2174]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[2175]_  = \new_[60]_  | \new_[2174]_ ;
  assign \new_[2179]_  = \new_[55]_  | \new_[56]_ ;
  assign \new_[2180]_  = \new_[57]_  | \new_[2179]_ ;
  assign \new_[2181]_  = \new_[2180]_  | \new_[2175]_ ;
  assign \new_[2185]_  = \new_[52]_  | \new_[53]_ ;
  assign \new_[2186]_  = \new_[54]_  | \new_[2185]_ ;
  assign \new_[2190]_  = \new_[49]_  | \new_[50]_ ;
  assign \new_[2191]_  = \new_[51]_  | \new_[2190]_ ;
  assign \new_[2192]_  = \new_[2191]_  | \new_[2186]_ ;
  assign \new_[2193]_  = \new_[2192]_  | \new_[2181]_ ;
  assign \new_[2194]_  = \new_[2193]_  | \new_[2170]_ ;
  assign \new_[2195]_  = \new_[2194]_  | \new_[2147]_ ;
  assign \new_[2199]_  = \new_[46]_  | \new_[47]_ ;
  assign \new_[2200]_  = \new_[48]_  | \new_[2199]_ ;
  assign \new_[2204]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[2205]_  = \new_[45]_  | \new_[2204]_ ;
  assign \new_[2206]_  = \new_[2205]_  | \new_[2200]_ ;
  assign \new_[2210]_  = \new_[40]_  | \new_[41]_ ;
  assign \new_[2211]_  = \new_[42]_  | \new_[2210]_ ;
  assign \new_[2215]_  = \new_[37]_  | \new_[38]_ ;
  assign \new_[2216]_  = \new_[39]_  | \new_[2215]_ ;
  assign \new_[2217]_  = \new_[2216]_  | \new_[2211]_ ;
  assign \new_[2218]_  = \new_[2217]_  | \new_[2206]_ ;
  assign \new_[2222]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[2223]_  = \new_[36]_  | \new_[2222]_ ;
  assign \new_[2227]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[2228]_  = \new_[33]_  | \new_[2227]_ ;
  assign \new_[2229]_  = \new_[2228]_  | \new_[2223]_ ;
  assign \new_[2233]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[2234]_  = \new_[30]_  | \new_[2233]_ ;
  assign \new_[2238]_  = \new_[25]_  | \new_[26]_ ;
  assign \new_[2239]_  = \new_[27]_  | \new_[2238]_ ;
  assign \new_[2240]_  = \new_[2239]_  | \new_[2234]_ ;
  assign \new_[2241]_  = \new_[2240]_  | \new_[2229]_ ;
  assign \new_[2242]_  = \new_[2241]_  | \new_[2218]_ ;
  assign \new_[2246]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[2247]_  = \new_[24]_  | \new_[2246]_ ;
  assign \new_[2251]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[2252]_  = \new_[21]_  | \new_[2251]_ ;
  assign \new_[2253]_  = \new_[2252]_  | \new_[2247]_ ;
  assign \new_[2257]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[2258]_  = \new_[18]_  | \new_[2257]_ ;
  assign \new_[2262]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[2263]_  = \new_[15]_  | \new_[2262]_ ;
  assign \new_[2264]_  = \new_[2263]_  | \new_[2258]_ ;
  assign \new_[2265]_  = \new_[2264]_  | \new_[2253]_ ;
  assign \new_[2269]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[2270]_  = \new_[12]_  | \new_[2269]_ ;
  assign \new_[2274]_  = \new_[7]_  | \new_[8]_ ;
  assign \new_[2275]_  = \new_[9]_  | \new_[2274]_ ;
  assign \new_[2276]_  = \new_[2275]_  | \new_[2270]_ ;
  assign \new_[2280]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[2281]_  = \new_[6]_  | \new_[2280]_ ;
  assign \new_[2285]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[2286]_  = \new_[3]_  | \new_[2285]_ ;
  assign \new_[2287]_  = \new_[2286]_  | \new_[2281]_ ;
  assign \new_[2288]_  = \new_[2287]_  | \new_[2276]_ ;
  assign \new_[2289]_  = \new_[2288]_  | \new_[2265]_ ;
  assign \new_[2290]_  = \new_[2289]_  | \new_[2242]_ ;
  assign \new_[2291]_  = \new_[2290]_  | \new_[2195]_ ;
  assign \new_[2292]_  = \new_[2291]_  | \new_[2100]_ ;
  assign \new_[2293]_  = \new_[2292]_  | \new_[1909]_ ;
  assign \new_[2296]_  = ~A167 & ~A169;
  assign \new_[2299]_  = A202 & ~A166;
  assign \new_[2302]_  = ~A169 & ~A170;
  assign \new_[2305]_  = A202 & ~A168;
  assign \new_[2308]_  = ~A167 & ~A169;
  assign \new_[2312]_  = A201 & A199;
  assign \new_[2313]_  = ~A166 & \new_[2312]_ ;
  assign \new_[2316]_  = ~A167 & ~A169;
  assign \new_[2320]_  = A201 & A200;
  assign \new_[2321]_  = ~A166 & \new_[2320]_ ;
  assign \new_[2324]_  = ~A168 & ~A169;
  assign \new_[2328]_  = A202 & A166;
  assign \new_[2329]_  = A167 & \new_[2328]_ ;
  assign \new_[2332]_  = ~A169 & ~A170;
  assign \new_[2336]_  = A201 & A199;
  assign \new_[2337]_  = ~A168 & \new_[2336]_ ;
  assign \new_[2340]_  = ~A169 & ~A170;
  assign \new_[2344]_  = A201 & A200;
  assign \new_[2345]_  = ~A168 & \new_[2344]_ ;
  assign \new_[2349]_  = ~A202 & ~A201;
  assign \new_[2350]_  = A169 & \new_[2349]_ ;
  assign \new_[2354]_  = A301 & A235;
  assign \new_[2355]_  = ~A203 & \new_[2354]_ ;
  assign \new_[2359]_  = ~A202 & ~A201;
  assign \new_[2360]_  = A169 & \new_[2359]_ ;
  assign \new_[2364]_  = A268 & A235;
  assign \new_[2365]_  = ~A203 & \new_[2364]_ ;
  assign \new_[2369]_  = ~A200 & ~A199;
  assign \new_[2370]_  = A169 & \new_[2369]_ ;
  assign \new_[2374]_  = A301 & A235;
  assign \new_[2375]_  = ~A202 & \new_[2374]_ ;
  assign \new_[2379]_  = ~A200 & ~A199;
  assign \new_[2380]_  = A169 & \new_[2379]_ ;
  assign \new_[2384]_  = A268 & A235;
  assign \new_[2385]_  = ~A202 & \new_[2384]_ ;
  assign \new_[2389]_  = ~A166 & ~A167;
  assign \new_[2390]_  = ~A169 & \new_[2389]_ ;
  assign \new_[2394]_  = A203 & A200;
  assign \new_[2395]_  = ~A199 & \new_[2394]_ ;
  assign \new_[2399]_  = ~A166 & ~A167;
  assign \new_[2400]_  = ~A169 & \new_[2399]_ ;
  assign \new_[2404]_  = A203 & ~A200;
  assign \new_[2405]_  = A199 & \new_[2404]_ ;
  assign \new_[2409]_  = A167 & ~A168;
  assign \new_[2410]_  = ~A169 & \new_[2409]_ ;
  assign \new_[2414]_  = A201 & A199;
  assign \new_[2415]_  = A166 & \new_[2414]_ ;
  assign \new_[2419]_  = A167 & ~A168;
  assign \new_[2420]_  = ~A169 & \new_[2419]_ ;
  assign \new_[2424]_  = A201 & A200;
  assign \new_[2425]_  = A166 & \new_[2424]_ ;
  assign \new_[2429]_  = ~A168 & ~A169;
  assign \new_[2430]_  = ~A170 & \new_[2429]_ ;
  assign \new_[2434]_  = A203 & A200;
  assign \new_[2435]_  = ~A199 & \new_[2434]_ ;
  assign \new_[2439]_  = ~A168 & ~A169;
  assign \new_[2440]_  = ~A170 & \new_[2439]_ ;
  assign \new_[2444]_  = A203 & ~A200;
  assign \new_[2445]_  = A199 & \new_[2444]_ ;
  assign \new_[2449]_  = ~A201 & A166;
  assign \new_[2450]_  = A168 & \new_[2449]_ ;
  assign \new_[2453]_  = ~A203 & ~A202;
  assign \new_[2456]_  = A301 & A235;
  assign \new_[2457]_  = \new_[2456]_  & \new_[2453]_ ;
  assign \new_[2461]_  = ~A201 & A166;
  assign \new_[2462]_  = A168 & \new_[2461]_ ;
  assign \new_[2465]_  = ~A203 & ~A202;
  assign \new_[2468]_  = A268 & A235;
  assign \new_[2469]_  = \new_[2468]_  & \new_[2465]_ ;
  assign \new_[2473]_  = ~A199 & A166;
  assign \new_[2474]_  = A168 & \new_[2473]_ ;
  assign \new_[2477]_  = ~A202 & ~A200;
  assign \new_[2480]_  = A301 & A235;
  assign \new_[2481]_  = \new_[2480]_  & \new_[2477]_ ;
  assign \new_[2485]_  = ~A199 & A166;
  assign \new_[2486]_  = A168 & \new_[2485]_ ;
  assign \new_[2489]_  = ~A202 & ~A200;
  assign \new_[2492]_  = A268 & A235;
  assign \new_[2493]_  = \new_[2492]_  & \new_[2489]_ ;
  assign \new_[2497]_  = ~A201 & A167;
  assign \new_[2498]_  = A168 & \new_[2497]_ ;
  assign \new_[2501]_  = ~A203 & ~A202;
  assign \new_[2504]_  = A301 & A235;
  assign \new_[2505]_  = \new_[2504]_  & \new_[2501]_ ;
  assign \new_[2509]_  = ~A201 & A167;
  assign \new_[2510]_  = A168 & \new_[2509]_ ;
  assign \new_[2513]_  = ~A203 & ~A202;
  assign \new_[2516]_  = A268 & A235;
  assign \new_[2517]_  = \new_[2516]_  & \new_[2513]_ ;
  assign \new_[2521]_  = ~A199 & A167;
  assign \new_[2522]_  = A168 & \new_[2521]_ ;
  assign \new_[2525]_  = ~A202 & ~A200;
  assign \new_[2528]_  = A301 & A235;
  assign \new_[2529]_  = \new_[2528]_  & \new_[2525]_ ;
  assign \new_[2533]_  = ~A199 & A167;
  assign \new_[2534]_  = A168 & \new_[2533]_ ;
  assign \new_[2537]_  = ~A202 & ~A200;
  assign \new_[2540]_  = A268 & A235;
  assign \new_[2541]_  = \new_[2540]_  & \new_[2537]_ ;
  assign \new_[2545]_  = ~A202 & ~A201;
  assign \new_[2546]_  = A169 & \new_[2545]_ ;
  assign \new_[2549]_  = A235 & ~A203;
  assign \new_[2552]_  = A300 & A299;
  assign \new_[2553]_  = \new_[2552]_  & \new_[2549]_ ;
  assign \new_[2557]_  = ~A202 & ~A201;
  assign \new_[2558]_  = A169 & \new_[2557]_ ;
  assign \new_[2561]_  = A235 & ~A203;
  assign \new_[2564]_  = A300 & A298;
  assign \new_[2565]_  = \new_[2564]_  & \new_[2561]_ ;
  assign \new_[2569]_  = ~A202 & ~A201;
  assign \new_[2570]_  = A169 & \new_[2569]_ ;
  assign \new_[2573]_  = A235 & ~A203;
  assign \new_[2576]_  = A267 & A265;
  assign \new_[2577]_  = \new_[2576]_  & \new_[2573]_ ;
  assign \new_[2581]_  = ~A202 & ~A201;
  assign \new_[2582]_  = A169 & \new_[2581]_ ;
  assign \new_[2585]_  = A235 & ~A203;
  assign \new_[2588]_  = A267 & A266;
  assign \new_[2589]_  = \new_[2588]_  & \new_[2585]_ ;
  assign \new_[2593]_  = ~A202 & ~A201;
  assign \new_[2594]_  = A169 & \new_[2593]_ ;
  assign \new_[2597]_  = A232 & ~A203;
  assign \new_[2600]_  = A301 & A234;
  assign \new_[2601]_  = \new_[2600]_  & \new_[2597]_ ;
  assign \new_[2605]_  = ~A202 & ~A201;
  assign \new_[2606]_  = A169 & \new_[2605]_ ;
  assign \new_[2609]_  = A232 & ~A203;
  assign \new_[2612]_  = A268 & A234;
  assign \new_[2613]_  = \new_[2612]_  & \new_[2609]_ ;
  assign \new_[2617]_  = ~A202 & ~A201;
  assign \new_[2618]_  = A169 & \new_[2617]_ ;
  assign \new_[2621]_  = A233 & ~A203;
  assign \new_[2624]_  = A301 & A234;
  assign \new_[2625]_  = \new_[2624]_  & \new_[2621]_ ;
  assign \new_[2629]_  = ~A202 & ~A201;
  assign \new_[2630]_  = A169 & \new_[2629]_ ;
  assign \new_[2633]_  = A233 & ~A203;
  assign \new_[2636]_  = A268 & A234;
  assign \new_[2637]_  = \new_[2636]_  & \new_[2633]_ ;
  assign \new_[2641]_  = A200 & A199;
  assign \new_[2642]_  = A169 & \new_[2641]_ ;
  assign \new_[2645]_  = ~A202 & ~A201;
  assign \new_[2648]_  = A301 & A235;
  assign \new_[2649]_  = \new_[2648]_  & \new_[2645]_ ;
  assign \new_[2653]_  = A200 & A199;
  assign \new_[2654]_  = A169 & \new_[2653]_ ;
  assign \new_[2657]_  = ~A202 & ~A201;
  assign \new_[2660]_  = A268 & A235;
  assign \new_[2661]_  = \new_[2660]_  & \new_[2657]_ ;
  assign \new_[2665]_  = ~A200 & ~A199;
  assign \new_[2666]_  = A169 & \new_[2665]_ ;
  assign \new_[2669]_  = A235 & ~A202;
  assign \new_[2672]_  = A300 & A299;
  assign \new_[2673]_  = \new_[2672]_  & \new_[2669]_ ;
  assign \new_[2677]_  = ~A200 & ~A199;
  assign \new_[2678]_  = A169 & \new_[2677]_ ;
  assign \new_[2681]_  = A235 & ~A202;
  assign \new_[2684]_  = A300 & A298;
  assign \new_[2685]_  = \new_[2684]_  & \new_[2681]_ ;
  assign \new_[2689]_  = ~A200 & ~A199;
  assign \new_[2690]_  = A169 & \new_[2689]_ ;
  assign \new_[2693]_  = A235 & ~A202;
  assign \new_[2696]_  = A267 & A265;
  assign \new_[2697]_  = \new_[2696]_  & \new_[2693]_ ;
  assign \new_[2701]_  = ~A200 & ~A199;
  assign \new_[2702]_  = A169 & \new_[2701]_ ;
  assign \new_[2705]_  = A235 & ~A202;
  assign \new_[2708]_  = A267 & A266;
  assign \new_[2709]_  = \new_[2708]_  & \new_[2705]_ ;
  assign \new_[2713]_  = ~A200 & ~A199;
  assign \new_[2714]_  = A169 & \new_[2713]_ ;
  assign \new_[2717]_  = A232 & ~A202;
  assign \new_[2720]_  = A301 & A234;
  assign \new_[2721]_  = \new_[2720]_  & \new_[2717]_ ;
  assign \new_[2725]_  = ~A200 & ~A199;
  assign \new_[2726]_  = A169 & \new_[2725]_ ;
  assign \new_[2729]_  = A232 & ~A202;
  assign \new_[2732]_  = A268 & A234;
  assign \new_[2733]_  = \new_[2732]_  & \new_[2729]_ ;
  assign \new_[2737]_  = ~A200 & ~A199;
  assign \new_[2738]_  = A169 & \new_[2737]_ ;
  assign \new_[2741]_  = A233 & ~A202;
  assign \new_[2744]_  = A301 & A234;
  assign \new_[2745]_  = \new_[2744]_  & \new_[2741]_ ;
  assign \new_[2749]_  = ~A200 & ~A199;
  assign \new_[2750]_  = A169 & \new_[2749]_ ;
  assign \new_[2753]_  = A233 & ~A202;
  assign \new_[2756]_  = A268 & A234;
  assign \new_[2757]_  = \new_[2756]_  & \new_[2753]_ ;
  assign \new_[2761]_  = A167 & ~A168;
  assign \new_[2762]_  = ~A169 & \new_[2761]_ ;
  assign \new_[2765]_  = ~A199 & A166;
  assign \new_[2768]_  = A203 & A200;
  assign \new_[2769]_  = \new_[2768]_  & \new_[2765]_ ;
  assign \new_[2773]_  = A167 & ~A168;
  assign \new_[2774]_  = ~A169 & \new_[2773]_ ;
  assign \new_[2777]_  = A199 & A166;
  assign \new_[2780]_  = A203 & ~A200;
  assign \new_[2781]_  = \new_[2780]_  & \new_[2777]_ ;
  assign \new_[2784]_  = A166 & A168;
  assign \new_[2787]_  = ~A202 & ~A201;
  assign \new_[2788]_  = \new_[2787]_  & \new_[2784]_ ;
  assign \new_[2791]_  = A235 & ~A203;
  assign \new_[2794]_  = A300 & A299;
  assign \new_[2795]_  = \new_[2794]_  & \new_[2791]_ ;
  assign \new_[2798]_  = A166 & A168;
  assign \new_[2801]_  = ~A202 & ~A201;
  assign \new_[2802]_  = \new_[2801]_  & \new_[2798]_ ;
  assign \new_[2805]_  = A235 & ~A203;
  assign \new_[2808]_  = A300 & A298;
  assign \new_[2809]_  = \new_[2808]_  & \new_[2805]_ ;
  assign \new_[2812]_  = A166 & A168;
  assign \new_[2815]_  = ~A202 & ~A201;
  assign \new_[2816]_  = \new_[2815]_  & \new_[2812]_ ;
  assign \new_[2819]_  = A235 & ~A203;
  assign \new_[2822]_  = A267 & A265;
  assign \new_[2823]_  = \new_[2822]_  & \new_[2819]_ ;
  assign \new_[2826]_  = A166 & A168;
  assign \new_[2829]_  = ~A202 & ~A201;
  assign \new_[2830]_  = \new_[2829]_  & \new_[2826]_ ;
  assign \new_[2833]_  = A235 & ~A203;
  assign \new_[2836]_  = A267 & A266;
  assign \new_[2837]_  = \new_[2836]_  & \new_[2833]_ ;
  assign \new_[2840]_  = A166 & A168;
  assign \new_[2843]_  = ~A202 & ~A201;
  assign \new_[2844]_  = \new_[2843]_  & \new_[2840]_ ;
  assign \new_[2847]_  = A232 & ~A203;
  assign \new_[2850]_  = A301 & A234;
  assign \new_[2851]_  = \new_[2850]_  & \new_[2847]_ ;
  assign \new_[2854]_  = A166 & A168;
  assign \new_[2857]_  = ~A202 & ~A201;
  assign \new_[2858]_  = \new_[2857]_  & \new_[2854]_ ;
  assign \new_[2861]_  = A232 & ~A203;
  assign \new_[2864]_  = A268 & A234;
  assign \new_[2865]_  = \new_[2864]_  & \new_[2861]_ ;
  assign \new_[2868]_  = A166 & A168;
  assign \new_[2871]_  = ~A202 & ~A201;
  assign \new_[2872]_  = \new_[2871]_  & \new_[2868]_ ;
  assign \new_[2875]_  = A233 & ~A203;
  assign \new_[2878]_  = A301 & A234;
  assign \new_[2879]_  = \new_[2878]_  & \new_[2875]_ ;
  assign \new_[2882]_  = A166 & A168;
  assign \new_[2885]_  = ~A202 & ~A201;
  assign \new_[2886]_  = \new_[2885]_  & \new_[2882]_ ;
  assign \new_[2889]_  = A233 & ~A203;
  assign \new_[2892]_  = A268 & A234;
  assign \new_[2893]_  = \new_[2892]_  & \new_[2889]_ ;
  assign \new_[2896]_  = A166 & A168;
  assign \new_[2899]_  = A200 & A199;
  assign \new_[2900]_  = \new_[2899]_  & \new_[2896]_ ;
  assign \new_[2903]_  = ~A202 & ~A201;
  assign \new_[2906]_  = A301 & A235;
  assign \new_[2907]_  = \new_[2906]_  & \new_[2903]_ ;
  assign \new_[2910]_  = A166 & A168;
  assign \new_[2913]_  = A200 & A199;
  assign \new_[2914]_  = \new_[2913]_  & \new_[2910]_ ;
  assign \new_[2917]_  = ~A202 & ~A201;
  assign \new_[2920]_  = A268 & A235;
  assign \new_[2921]_  = \new_[2920]_  & \new_[2917]_ ;
  assign \new_[2924]_  = A166 & A168;
  assign \new_[2927]_  = ~A200 & ~A199;
  assign \new_[2928]_  = \new_[2927]_  & \new_[2924]_ ;
  assign \new_[2931]_  = A235 & ~A202;
  assign \new_[2934]_  = A300 & A299;
  assign \new_[2935]_  = \new_[2934]_  & \new_[2931]_ ;
  assign \new_[2938]_  = A166 & A168;
  assign \new_[2941]_  = ~A200 & ~A199;
  assign \new_[2942]_  = \new_[2941]_  & \new_[2938]_ ;
  assign \new_[2945]_  = A235 & ~A202;
  assign \new_[2948]_  = A300 & A298;
  assign \new_[2949]_  = \new_[2948]_  & \new_[2945]_ ;
  assign \new_[2952]_  = A166 & A168;
  assign \new_[2955]_  = ~A200 & ~A199;
  assign \new_[2956]_  = \new_[2955]_  & \new_[2952]_ ;
  assign \new_[2959]_  = A235 & ~A202;
  assign \new_[2962]_  = A267 & A265;
  assign \new_[2963]_  = \new_[2962]_  & \new_[2959]_ ;
  assign \new_[2966]_  = A166 & A168;
  assign \new_[2969]_  = ~A200 & ~A199;
  assign \new_[2970]_  = \new_[2969]_  & \new_[2966]_ ;
  assign \new_[2973]_  = A235 & ~A202;
  assign \new_[2976]_  = A267 & A266;
  assign \new_[2977]_  = \new_[2976]_  & \new_[2973]_ ;
  assign \new_[2980]_  = A166 & A168;
  assign \new_[2983]_  = ~A200 & ~A199;
  assign \new_[2984]_  = \new_[2983]_  & \new_[2980]_ ;
  assign \new_[2987]_  = A232 & ~A202;
  assign \new_[2990]_  = A301 & A234;
  assign \new_[2991]_  = \new_[2990]_  & \new_[2987]_ ;
  assign \new_[2994]_  = A166 & A168;
  assign \new_[2997]_  = ~A200 & ~A199;
  assign \new_[2998]_  = \new_[2997]_  & \new_[2994]_ ;
  assign \new_[3001]_  = A232 & ~A202;
  assign \new_[3004]_  = A268 & A234;
  assign \new_[3005]_  = \new_[3004]_  & \new_[3001]_ ;
  assign \new_[3008]_  = A166 & A168;
  assign \new_[3011]_  = ~A200 & ~A199;
  assign \new_[3012]_  = \new_[3011]_  & \new_[3008]_ ;
  assign \new_[3015]_  = A233 & ~A202;
  assign \new_[3018]_  = A301 & A234;
  assign \new_[3019]_  = \new_[3018]_  & \new_[3015]_ ;
  assign \new_[3022]_  = A166 & A168;
  assign \new_[3025]_  = ~A200 & ~A199;
  assign \new_[3026]_  = \new_[3025]_  & \new_[3022]_ ;
  assign \new_[3029]_  = A233 & ~A202;
  assign \new_[3032]_  = A268 & A234;
  assign \new_[3033]_  = \new_[3032]_  & \new_[3029]_ ;
  assign \new_[3036]_  = A167 & A168;
  assign \new_[3039]_  = ~A202 & ~A201;
  assign \new_[3040]_  = \new_[3039]_  & \new_[3036]_ ;
  assign \new_[3043]_  = A235 & ~A203;
  assign \new_[3046]_  = A300 & A299;
  assign \new_[3047]_  = \new_[3046]_  & \new_[3043]_ ;
  assign \new_[3050]_  = A167 & A168;
  assign \new_[3053]_  = ~A202 & ~A201;
  assign \new_[3054]_  = \new_[3053]_  & \new_[3050]_ ;
  assign \new_[3057]_  = A235 & ~A203;
  assign \new_[3060]_  = A300 & A298;
  assign \new_[3061]_  = \new_[3060]_  & \new_[3057]_ ;
  assign \new_[3064]_  = A167 & A168;
  assign \new_[3067]_  = ~A202 & ~A201;
  assign \new_[3068]_  = \new_[3067]_  & \new_[3064]_ ;
  assign \new_[3071]_  = A235 & ~A203;
  assign \new_[3074]_  = A267 & A265;
  assign \new_[3075]_  = \new_[3074]_  & \new_[3071]_ ;
  assign \new_[3078]_  = A167 & A168;
  assign \new_[3081]_  = ~A202 & ~A201;
  assign \new_[3082]_  = \new_[3081]_  & \new_[3078]_ ;
  assign \new_[3085]_  = A235 & ~A203;
  assign \new_[3088]_  = A267 & A266;
  assign \new_[3089]_  = \new_[3088]_  & \new_[3085]_ ;
  assign \new_[3092]_  = A167 & A168;
  assign \new_[3095]_  = ~A202 & ~A201;
  assign \new_[3096]_  = \new_[3095]_  & \new_[3092]_ ;
  assign \new_[3099]_  = A232 & ~A203;
  assign \new_[3102]_  = A301 & A234;
  assign \new_[3103]_  = \new_[3102]_  & \new_[3099]_ ;
  assign \new_[3106]_  = A167 & A168;
  assign \new_[3109]_  = ~A202 & ~A201;
  assign \new_[3110]_  = \new_[3109]_  & \new_[3106]_ ;
  assign \new_[3113]_  = A232 & ~A203;
  assign \new_[3116]_  = A268 & A234;
  assign \new_[3117]_  = \new_[3116]_  & \new_[3113]_ ;
  assign \new_[3120]_  = A167 & A168;
  assign \new_[3123]_  = ~A202 & ~A201;
  assign \new_[3124]_  = \new_[3123]_  & \new_[3120]_ ;
  assign \new_[3127]_  = A233 & ~A203;
  assign \new_[3130]_  = A301 & A234;
  assign \new_[3131]_  = \new_[3130]_  & \new_[3127]_ ;
  assign \new_[3134]_  = A167 & A168;
  assign \new_[3137]_  = ~A202 & ~A201;
  assign \new_[3138]_  = \new_[3137]_  & \new_[3134]_ ;
  assign \new_[3141]_  = A233 & ~A203;
  assign \new_[3144]_  = A268 & A234;
  assign \new_[3145]_  = \new_[3144]_  & \new_[3141]_ ;
  assign \new_[3148]_  = A167 & A168;
  assign \new_[3151]_  = A200 & A199;
  assign \new_[3152]_  = \new_[3151]_  & \new_[3148]_ ;
  assign \new_[3155]_  = ~A202 & ~A201;
  assign \new_[3158]_  = A301 & A235;
  assign \new_[3159]_  = \new_[3158]_  & \new_[3155]_ ;
  assign \new_[3162]_  = A167 & A168;
  assign \new_[3165]_  = A200 & A199;
  assign \new_[3166]_  = \new_[3165]_  & \new_[3162]_ ;
  assign \new_[3169]_  = ~A202 & ~A201;
  assign \new_[3172]_  = A268 & A235;
  assign \new_[3173]_  = \new_[3172]_  & \new_[3169]_ ;
  assign \new_[3176]_  = A167 & A168;
  assign \new_[3179]_  = ~A200 & ~A199;
  assign \new_[3180]_  = \new_[3179]_  & \new_[3176]_ ;
  assign \new_[3183]_  = A235 & ~A202;
  assign \new_[3186]_  = A300 & A299;
  assign \new_[3187]_  = \new_[3186]_  & \new_[3183]_ ;
  assign \new_[3190]_  = A167 & A168;
  assign \new_[3193]_  = ~A200 & ~A199;
  assign \new_[3194]_  = \new_[3193]_  & \new_[3190]_ ;
  assign \new_[3197]_  = A235 & ~A202;
  assign \new_[3200]_  = A300 & A298;
  assign \new_[3201]_  = \new_[3200]_  & \new_[3197]_ ;
  assign \new_[3204]_  = A167 & A168;
  assign \new_[3207]_  = ~A200 & ~A199;
  assign \new_[3208]_  = \new_[3207]_  & \new_[3204]_ ;
  assign \new_[3211]_  = A235 & ~A202;
  assign \new_[3214]_  = A267 & A265;
  assign \new_[3215]_  = \new_[3214]_  & \new_[3211]_ ;
  assign \new_[3218]_  = A167 & A168;
  assign \new_[3221]_  = ~A200 & ~A199;
  assign \new_[3222]_  = \new_[3221]_  & \new_[3218]_ ;
  assign \new_[3225]_  = A235 & ~A202;
  assign \new_[3228]_  = A267 & A266;
  assign \new_[3229]_  = \new_[3228]_  & \new_[3225]_ ;
  assign \new_[3232]_  = A167 & A168;
  assign \new_[3235]_  = ~A200 & ~A199;
  assign \new_[3236]_  = \new_[3235]_  & \new_[3232]_ ;
  assign \new_[3239]_  = A232 & ~A202;
  assign \new_[3242]_  = A301 & A234;
  assign \new_[3243]_  = \new_[3242]_  & \new_[3239]_ ;
  assign \new_[3246]_  = A167 & A168;
  assign \new_[3249]_  = ~A200 & ~A199;
  assign \new_[3250]_  = \new_[3249]_  & \new_[3246]_ ;
  assign \new_[3253]_  = A232 & ~A202;
  assign \new_[3256]_  = A268 & A234;
  assign \new_[3257]_  = \new_[3256]_  & \new_[3253]_ ;
  assign \new_[3260]_  = A167 & A168;
  assign \new_[3263]_  = ~A200 & ~A199;
  assign \new_[3264]_  = \new_[3263]_  & \new_[3260]_ ;
  assign \new_[3267]_  = A233 & ~A202;
  assign \new_[3270]_  = A301 & A234;
  assign \new_[3271]_  = \new_[3270]_  & \new_[3267]_ ;
  assign \new_[3274]_  = A167 & A168;
  assign \new_[3277]_  = ~A200 & ~A199;
  assign \new_[3278]_  = \new_[3277]_  & \new_[3274]_ ;
  assign \new_[3281]_  = A233 & ~A202;
  assign \new_[3284]_  = A268 & A234;
  assign \new_[3285]_  = \new_[3284]_  & \new_[3281]_ ;
  assign \new_[3288]_  = A167 & A170;
  assign \new_[3291]_  = ~A201 & ~A166;
  assign \new_[3292]_  = \new_[3291]_  & \new_[3288]_ ;
  assign \new_[3295]_  = ~A203 & ~A202;
  assign \new_[3298]_  = A301 & A235;
  assign \new_[3299]_  = \new_[3298]_  & \new_[3295]_ ;
  assign \new_[3302]_  = A167 & A170;
  assign \new_[3305]_  = ~A201 & ~A166;
  assign \new_[3306]_  = \new_[3305]_  & \new_[3302]_ ;
  assign \new_[3309]_  = ~A203 & ~A202;
  assign \new_[3312]_  = A268 & A235;
  assign \new_[3313]_  = \new_[3312]_  & \new_[3309]_ ;
  assign \new_[3316]_  = A167 & A170;
  assign \new_[3319]_  = ~A199 & ~A166;
  assign \new_[3320]_  = \new_[3319]_  & \new_[3316]_ ;
  assign \new_[3323]_  = ~A202 & ~A200;
  assign \new_[3326]_  = A301 & A235;
  assign \new_[3327]_  = \new_[3326]_  & \new_[3323]_ ;
  assign \new_[3330]_  = A167 & A170;
  assign \new_[3333]_  = ~A199 & ~A166;
  assign \new_[3334]_  = \new_[3333]_  & \new_[3330]_ ;
  assign \new_[3337]_  = ~A202 & ~A200;
  assign \new_[3340]_  = A268 & A235;
  assign \new_[3341]_  = \new_[3340]_  & \new_[3337]_ ;
  assign \new_[3344]_  = ~A167 & A170;
  assign \new_[3347]_  = ~A201 & A166;
  assign \new_[3348]_  = \new_[3347]_  & \new_[3344]_ ;
  assign \new_[3351]_  = ~A203 & ~A202;
  assign \new_[3354]_  = A301 & A235;
  assign \new_[3355]_  = \new_[3354]_  & \new_[3351]_ ;
  assign \new_[3358]_  = ~A167 & A170;
  assign \new_[3361]_  = ~A201 & A166;
  assign \new_[3362]_  = \new_[3361]_  & \new_[3358]_ ;
  assign \new_[3365]_  = ~A203 & ~A202;
  assign \new_[3368]_  = A268 & A235;
  assign \new_[3369]_  = \new_[3368]_  & \new_[3365]_ ;
  assign \new_[3372]_  = ~A167 & A170;
  assign \new_[3375]_  = ~A199 & A166;
  assign \new_[3376]_  = \new_[3375]_  & \new_[3372]_ ;
  assign \new_[3379]_  = ~A202 & ~A200;
  assign \new_[3382]_  = A301 & A235;
  assign \new_[3383]_  = \new_[3382]_  & \new_[3379]_ ;
  assign \new_[3386]_  = ~A167 & A170;
  assign \new_[3389]_  = ~A199 & A166;
  assign \new_[3390]_  = \new_[3389]_  & \new_[3386]_ ;
  assign \new_[3393]_  = ~A202 & ~A200;
  assign \new_[3396]_  = A268 & A235;
  assign \new_[3397]_  = \new_[3396]_  & \new_[3393]_ ;
  assign \new_[3400]_  = ~A201 & A169;
  assign \new_[3403]_  = ~A203 & ~A202;
  assign \new_[3404]_  = \new_[3403]_  & \new_[3400]_ ;
  assign \new_[3407]_  = A298 & A235;
  assign \new_[3410]_  = A302 & ~A299;
  assign \new_[3411]_  = \new_[3410]_  & \new_[3407]_ ;
  assign \new_[3414]_  = ~A201 & A169;
  assign \new_[3417]_  = ~A203 & ~A202;
  assign \new_[3418]_  = \new_[3417]_  & \new_[3414]_ ;
  assign \new_[3421]_  = ~A298 & A235;
  assign \new_[3424]_  = A302 & A299;
  assign \new_[3425]_  = \new_[3424]_  & \new_[3421]_ ;
  assign \new_[3428]_  = ~A201 & A169;
  assign \new_[3431]_  = ~A203 & ~A202;
  assign \new_[3432]_  = \new_[3431]_  & \new_[3428]_ ;
  assign \new_[3435]_  = ~A265 & A235;
  assign \new_[3438]_  = A269 & A266;
  assign \new_[3439]_  = \new_[3438]_  & \new_[3435]_ ;
  assign \new_[3442]_  = ~A201 & A169;
  assign \new_[3445]_  = ~A203 & ~A202;
  assign \new_[3446]_  = \new_[3445]_  & \new_[3442]_ ;
  assign \new_[3449]_  = A265 & A235;
  assign \new_[3452]_  = A269 & ~A266;
  assign \new_[3453]_  = \new_[3452]_  & \new_[3449]_ ;
  assign \new_[3456]_  = ~A201 & A169;
  assign \new_[3459]_  = ~A203 & ~A202;
  assign \new_[3460]_  = \new_[3459]_  & \new_[3456]_ ;
  assign \new_[3463]_  = A234 & A232;
  assign \new_[3466]_  = A300 & A299;
  assign \new_[3467]_  = \new_[3466]_  & \new_[3463]_ ;
  assign \new_[3470]_  = ~A201 & A169;
  assign \new_[3473]_  = ~A203 & ~A202;
  assign \new_[3474]_  = \new_[3473]_  & \new_[3470]_ ;
  assign \new_[3477]_  = A234 & A232;
  assign \new_[3480]_  = A300 & A298;
  assign \new_[3481]_  = \new_[3480]_  & \new_[3477]_ ;
  assign \new_[3484]_  = ~A201 & A169;
  assign \new_[3487]_  = ~A203 & ~A202;
  assign \new_[3488]_  = \new_[3487]_  & \new_[3484]_ ;
  assign \new_[3491]_  = A234 & A232;
  assign \new_[3494]_  = A267 & A265;
  assign \new_[3495]_  = \new_[3494]_  & \new_[3491]_ ;
  assign \new_[3498]_  = ~A201 & A169;
  assign \new_[3501]_  = ~A203 & ~A202;
  assign \new_[3502]_  = \new_[3501]_  & \new_[3498]_ ;
  assign \new_[3505]_  = A234 & A232;
  assign \new_[3508]_  = A267 & A266;
  assign \new_[3509]_  = \new_[3508]_  & \new_[3505]_ ;
  assign \new_[3512]_  = ~A201 & A169;
  assign \new_[3515]_  = ~A203 & ~A202;
  assign \new_[3516]_  = \new_[3515]_  & \new_[3512]_ ;
  assign \new_[3519]_  = A234 & A233;
  assign \new_[3522]_  = A300 & A299;
  assign \new_[3523]_  = \new_[3522]_  & \new_[3519]_ ;
  assign \new_[3526]_  = ~A201 & A169;
  assign \new_[3529]_  = ~A203 & ~A202;
  assign \new_[3530]_  = \new_[3529]_  & \new_[3526]_ ;
  assign \new_[3533]_  = A234 & A233;
  assign \new_[3536]_  = A300 & A298;
  assign \new_[3537]_  = \new_[3536]_  & \new_[3533]_ ;
  assign \new_[3540]_  = ~A201 & A169;
  assign \new_[3543]_  = ~A203 & ~A202;
  assign \new_[3544]_  = \new_[3543]_  & \new_[3540]_ ;
  assign \new_[3547]_  = A234 & A233;
  assign \new_[3550]_  = A267 & A265;
  assign \new_[3551]_  = \new_[3550]_  & \new_[3547]_ ;
  assign \new_[3554]_  = ~A201 & A169;
  assign \new_[3557]_  = ~A203 & ~A202;
  assign \new_[3558]_  = \new_[3557]_  & \new_[3554]_ ;
  assign \new_[3561]_  = A234 & A233;
  assign \new_[3564]_  = A267 & A266;
  assign \new_[3565]_  = \new_[3564]_  & \new_[3561]_ ;
  assign \new_[3568]_  = ~A201 & A169;
  assign \new_[3571]_  = ~A203 & ~A202;
  assign \new_[3572]_  = \new_[3571]_  & \new_[3568]_ ;
  assign \new_[3575]_  = A233 & ~A232;
  assign \new_[3578]_  = A301 & A236;
  assign \new_[3579]_  = \new_[3578]_  & \new_[3575]_ ;
  assign \new_[3582]_  = ~A201 & A169;
  assign \new_[3585]_  = ~A203 & ~A202;
  assign \new_[3586]_  = \new_[3585]_  & \new_[3582]_ ;
  assign \new_[3589]_  = A233 & ~A232;
  assign \new_[3592]_  = A268 & A236;
  assign \new_[3593]_  = \new_[3592]_  & \new_[3589]_ ;
  assign \new_[3596]_  = ~A201 & A169;
  assign \new_[3599]_  = ~A203 & ~A202;
  assign \new_[3600]_  = \new_[3599]_  & \new_[3596]_ ;
  assign \new_[3603]_  = ~A233 & A232;
  assign \new_[3606]_  = A301 & A236;
  assign \new_[3607]_  = \new_[3606]_  & \new_[3603]_ ;
  assign \new_[3610]_  = ~A201 & A169;
  assign \new_[3613]_  = ~A203 & ~A202;
  assign \new_[3614]_  = \new_[3613]_  & \new_[3610]_ ;
  assign \new_[3617]_  = ~A233 & A232;
  assign \new_[3620]_  = A268 & A236;
  assign \new_[3621]_  = \new_[3620]_  & \new_[3617]_ ;
  assign \new_[3624]_  = A199 & A169;
  assign \new_[3627]_  = ~A201 & A200;
  assign \new_[3628]_  = \new_[3627]_  & \new_[3624]_ ;
  assign \new_[3631]_  = A235 & ~A202;
  assign \new_[3634]_  = A300 & A299;
  assign \new_[3635]_  = \new_[3634]_  & \new_[3631]_ ;
  assign \new_[3638]_  = A199 & A169;
  assign \new_[3641]_  = ~A201 & A200;
  assign \new_[3642]_  = \new_[3641]_  & \new_[3638]_ ;
  assign \new_[3645]_  = A235 & ~A202;
  assign \new_[3648]_  = A300 & A298;
  assign \new_[3649]_  = \new_[3648]_  & \new_[3645]_ ;
  assign \new_[3652]_  = A199 & A169;
  assign \new_[3655]_  = ~A201 & A200;
  assign \new_[3656]_  = \new_[3655]_  & \new_[3652]_ ;
  assign \new_[3659]_  = A235 & ~A202;
  assign \new_[3662]_  = A267 & A265;
  assign \new_[3663]_  = \new_[3662]_  & \new_[3659]_ ;
  assign \new_[3666]_  = A199 & A169;
  assign \new_[3669]_  = ~A201 & A200;
  assign \new_[3670]_  = \new_[3669]_  & \new_[3666]_ ;
  assign \new_[3673]_  = A235 & ~A202;
  assign \new_[3676]_  = A267 & A266;
  assign \new_[3677]_  = \new_[3676]_  & \new_[3673]_ ;
  assign \new_[3680]_  = A199 & A169;
  assign \new_[3683]_  = ~A201 & A200;
  assign \new_[3684]_  = \new_[3683]_  & \new_[3680]_ ;
  assign \new_[3687]_  = A232 & ~A202;
  assign \new_[3690]_  = A301 & A234;
  assign \new_[3691]_  = \new_[3690]_  & \new_[3687]_ ;
  assign \new_[3694]_  = A199 & A169;
  assign \new_[3697]_  = ~A201 & A200;
  assign \new_[3698]_  = \new_[3697]_  & \new_[3694]_ ;
  assign \new_[3701]_  = A232 & ~A202;
  assign \new_[3704]_  = A268 & A234;
  assign \new_[3705]_  = \new_[3704]_  & \new_[3701]_ ;
  assign \new_[3708]_  = A199 & A169;
  assign \new_[3711]_  = ~A201 & A200;
  assign \new_[3712]_  = \new_[3711]_  & \new_[3708]_ ;
  assign \new_[3715]_  = A233 & ~A202;
  assign \new_[3718]_  = A301 & A234;
  assign \new_[3719]_  = \new_[3718]_  & \new_[3715]_ ;
  assign \new_[3722]_  = A199 & A169;
  assign \new_[3725]_  = ~A201 & A200;
  assign \new_[3726]_  = \new_[3725]_  & \new_[3722]_ ;
  assign \new_[3729]_  = A233 & ~A202;
  assign \new_[3732]_  = A268 & A234;
  assign \new_[3733]_  = \new_[3732]_  & \new_[3729]_ ;
  assign \new_[3736]_  = ~A199 & A169;
  assign \new_[3739]_  = ~A202 & ~A200;
  assign \new_[3740]_  = \new_[3739]_  & \new_[3736]_ ;
  assign \new_[3743]_  = A298 & A235;
  assign \new_[3746]_  = A302 & ~A299;
  assign \new_[3747]_  = \new_[3746]_  & \new_[3743]_ ;
  assign \new_[3750]_  = ~A199 & A169;
  assign \new_[3753]_  = ~A202 & ~A200;
  assign \new_[3754]_  = \new_[3753]_  & \new_[3750]_ ;
  assign \new_[3757]_  = ~A298 & A235;
  assign \new_[3760]_  = A302 & A299;
  assign \new_[3761]_  = \new_[3760]_  & \new_[3757]_ ;
  assign \new_[3764]_  = ~A199 & A169;
  assign \new_[3767]_  = ~A202 & ~A200;
  assign \new_[3768]_  = \new_[3767]_  & \new_[3764]_ ;
  assign \new_[3771]_  = ~A265 & A235;
  assign \new_[3774]_  = A269 & A266;
  assign \new_[3775]_  = \new_[3774]_  & \new_[3771]_ ;
  assign \new_[3778]_  = ~A199 & A169;
  assign \new_[3781]_  = ~A202 & ~A200;
  assign \new_[3782]_  = \new_[3781]_  & \new_[3778]_ ;
  assign \new_[3785]_  = A265 & A235;
  assign \new_[3788]_  = A269 & ~A266;
  assign \new_[3789]_  = \new_[3788]_  & \new_[3785]_ ;
  assign \new_[3792]_  = ~A199 & A169;
  assign \new_[3795]_  = ~A202 & ~A200;
  assign \new_[3796]_  = \new_[3795]_  & \new_[3792]_ ;
  assign \new_[3799]_  = A234 & A232;
  assign \new_[3802]_  = A300 & A299;
  assign \new_[3803]_  = \new_[3802]_  & \new_[3799]_ ;
  assign \new_[3806]_  = ~A199 & A169;
  assign \new_[3809]_  = ~A202 & ~A200;
  assign \new_[3810]_  = \new_[3809]_  & \new_[3806]_ ;
  assign \new_[3813]_  = A234 & A232;
  assign \new_[3816]_  = A300 & A298;
  assign \new_[3817]_  = \new_[3816]_  & \new_[3813]_ ;
  assign \new_[3820]_  = ~A199 & A169;
  assign \new_[3823]_  = ~A202 & ~A200;
  assign \new_[3824]_  = \new_[3823]_  & \new_[3820]_ ;
  assign \new_[3827]_  = A234 & A232;
  assign \new_[3830]_  = A267 & A265;
  assign \new_[3831]_  = \new_[3830]_  & \new_[3827]_ ;
  assign \new_[3834]_  = ~A199 & A169;
  assign \new_[3837]_  = ~A202 & ~A200;
  assign \new_[3838]_  = \new_[3837]_  & \new_[3834]_ ;
  assign \new_[3841]_  = A234 & A232;
  assign \new_[3844]_  = A267 & A266;
  assign \new_[3845]_  = \new_[3844]_  & \new_[3841]_ ;
  assign \new_[3848]_  = ~A199 & A169;
  assign \new_[3851]_  = ~A202 & ~A200;
  assign \new_[3852]_  = \new_[3851]_  & \new_[3848]_ ;
  assign \new_[3855]_  = A234 & A233;
  assign \new_[3858]_  = A300 & A299;
  assign \new_[3859]_  = \new_[3858]_  & \new_[3855]_ ;
  assign \new_[3862]_  = ~A199 & A169;
  assign \new_[3865]_  = ~A202 & ~A200;
  assign \new_[3866]_  = \new_[3865]_  & \new_[3862]_ ;
  assign \new_[3869]_  = A234 & A233;
  assign \new_[3872]_  = A300 & A298;
  assign \new_[3873]_  = \new_[3872]_  & \new_[3869]_ ;
  assign \new_[3876]_  = ~A199 & A169;
  assign \new_[3879]_  = ~A202 & ~A200;
  assign \new_[3880]_  = \new_[3879]_  & \new_[3876]_ ;
  assign \new_[3883]_  = A234 & A233;
  assign \new_[3886]_  = A267 & A265;
  assign \new_[3887]_  = \new_[3886]_  & \new_[3883]_ ;
  assign \new_[3890]_  = ~A199 & A169;
  assign \new_[3893]_  = ~A202 & ~A200;
  assign \new_[3894]_  = \new_[3893]_  & \new_[3890]_ ;
  assign \new_[3897]_  = A234 & A233;
  assign \new_[3900]_  = A267 & A266;
  assign \new_[3901]_  = \new_[3900]_  & \new_[3897]_ ;
  assign \new_[3904]_  = ~A199 & A169;
  assign \new_[3907]_  = ~A202 & ~A200;
  assign \new_[3908]_  = \new_[3907]_  & \new_[3904]_ ;
  assign \new_[3911]_  = A233 & ~A232;
  assign \new_[3914]_  = A301 & A236;
  assign \new_[3915]_  = \new_[3914]_  & \new_[3911]_ ;
  assign \new_[3918]_  = ~A199 & A169;
  assign \new_[3921]_  = ~A202 & ~A200;
  assign \new_[3922]_  = \new_[3921]_  & \new_[3918]_ ;
  assign \new_[3925]_  = A233 & ~A232;
  assign \new_[3928]_  = A268 & A236;
  assign \new_[3929]_  = \new_[3928]_  & \new_[3925]_ ;
  assign \new_[3932]_  = ~A199 & A169;
  assign \new_[3935]_  = ~A202 & ~A200;
  assign \new_[3936]_  = \new_[3935]_  & \new_[3932]_ ;
  assign \new_[3939]_  = ~A233 & A232;
  assign \new_[3942]_  = A301 & A236;
  assign \new_[3943]_  = \new_[3942]_  & \new_[3939]_ ;
  assign \new_[3946]_  = ~A199 & A169;
  assign \new_[3949]_  = ~A202 & ~A200;
  assign \new_[3950]_  = \new_[3949]_  & \new_[3946]_ ;
  assign \new_[3953]_  = ~A233 & A232;
  assign \new_[3956]_  = A268 & A236;
  assign \new_[3957]_  = \new_[3956]_  & \new_[3953]_ ;
  assign \new_[3960]_  = A166 & A168;
  assign \new_[3963]_  = ~A202 & ~A201;
  assign \new_[3964]_  = \new_[3963]_  & \new_[3960]_ ;
  assign \new_[3967]_  = A235 & ~A203;
  assign \new_[3971]_  = A302 & ~A299;
  assign \new_[3972]_  = A298 & \new_[3971]_ ;
  assign \new_[3973]_  = \new_[3972]_  & \new_[3967]_ ;
  assign \new_[3976]_  = A166 & A168;
  assign \new_[3979]_  = ~A202 & ~A201;
  assign \new_[3980]_  = \new_[3979]_  & \new_[3976]_ ;
  assign \new_[3983]_  = A235 & ~A203;
  assign \new_[3987]_  = A302 & A299;
  assign \new_[3988]_  = ~A298 & \new_[3987]_ ;
  assign \new_[3989]_  = \new_[3988]_  & \new_[3983]_ ;
  assign \new_[3992]_  = A166 & A168;
  assign \new_[3995]_  = ~A202 & ~A201;
  assign \new_[3996]_  = \new_[3995]_  & \new_[3992]_ ;
  assign \new_[3999]_  = A235 & ~A203;
  assign \new_[4003]_  = A269 & A266;
  assign \new_[4004]_  = ~A265 & \new_[4003]_ ;
  assign \new_[4005]_  = \new_[4004]_  & \new_[3999]_ ;
  assign \new_[4008]_  = A166 & A168;
  assign \new_[4011]_  = ~A202 & ~A201;
  assign \new_[4012]_  = \new_[4011]_  & \new_[4008]_ ;
  assign \new_[4015]_  = A235 & ~A203;
  assign \new_[4019]_  = A269 & ~A266;
  assign \new_[4020]_  = A265 & \new_[4019]_ ;
  assign \new_[4021]_  = \new_[4020]_  & \new_[4015]_ ;
  assign \new_[4024]_  = A166 & A168;
  assign \new_[4027]_  = ~A202 & ~A201;
  assign \new_[4028]_  = \new_[4027]_  & \new_[4024]_ ;
  assign \new_[4031]_  = A232 & ~A203;
  assign \new_[4035]_  = A300 & A299;
  assign \new_[4036]_  = A234 & \new_[4035]_ ;
  assign \new_[4037]_  = \new_[4036]_  & \new_[4031]_ ;
  assign \new_[4040]_  = A166 & A168;
  assign \new_[4043]_  = ~A202 & ~A201;
  assign \new_[4044]_  = \new_[4043]_  & \new_[4040]_ ;
  assign \new_[4047]_  = A232 & ~A203;
  assign \new_[4051]_  = A300 & A298;
  assign \new_[4052]_  = A234 & \new_[4051]_ ;
  assign \new_[4053]_  = \new_[4052]_  & \new_[4047]_ ;
  assign \new_[4056]_  = A166 & A168;
  assign \new_[4059]_  = ~A202 & ~A201;
  assign \new_[4060]_  = \new_[4059]_  & \new_[4056]_ ;
  assign \new_[4063]_  = A232 & ~A203;
  assign \new_[4067]_  = A267 & A265;
  assign \new_[4068]_  = A234 & \new_[4067]_ ;
  assign \new_[4069]_  = \new_[4068]_  & \new_[4063]_ ;
  assign \new_[4072]_  = A166 & A168;
  assign \new_[4075]_  = ~A202 & ~A201;
  assign \new_[4076]_  = \new_[4075]_  & \new_[4072]_ ;
  assign \new_[4079]_  = A232 & ~A203;
  assign \new_[4083]_  = A267 & A266;
  assign \new_[4084]_  = A234 & \new_[4083]_ ;
  assign \new_[4085]_  = \new_[4084]_  & \new_[4079]_ ;
  assign \new_[4088]_  = A166 & A168;
  assign \new_[4091]_  = ~A202 & ~A201;
  assign \new_[4092]_  = \new_[4091]_  & \new_[4088]_ ;
  assign \new_[4095]_  = A233 & ~A203;
  assign \new_[4099]_  = A300 & A299;
  assign \new_[4100]_  = A234 & \new_[4099]_ ;
  assign \new_[4101]_  = \new_[4100]_  & \new_[4095]_ ;
  assign \new_[4104]_  = A166 & A168;
  assign \new_[4107]_  = ~A202 & ~A201;
  assign \new_[4108]_  = \new_[4107]_  & \new_[4104]_ ;
  assign \new_[4111]_  = A233 & ~A203;
  assign \new_[4115]_  = A300 & A298;
  assign \new_[4116]_  = A234 & \new_[4115]_ ;
  assign \new_[4117]_  = \new_[4116]_  & \new_[4111]_ ;
  assign \new_[4120]_  = A166 & A168;
  assign \new_[4123]_  = ~A202 & ~A201;
  assign \new_[4124]_  = \new_[4123]_  & \new_[4120]_ ;
  assign \new_[4127]_  = A233 & ~A203;
  assign \new_[4131]_  = A267 & A265;
  assign \new_[4132]_  = A234 & \new_[4131]_ ;
  assign \new_[4133]_  = \new_[4132]_  & \new_[4127]_ ;
  assign \new_[4136]_  = A166 & A168;
  assign \new_[4139]_  = ~A202 & ~A201;
  assign \new_[4140]_  = \new_[4139]_  & \new_[4136]_ ;
  assign \new_[4143]_  = A233 & ~A203;
  assign \new_[4147]_  = A267 & A266;
  assign \new_[4148]_  = A234 & \new_[4147]_ ;
  assign \new_[4149]_  = \new_[4148]_  & \new_[4143]_ ;
  assign \new_[4152]_  = A166 & A168;
  assign \new_[4155]_  = ~A202 & ~A201;
  assign \new_[4156]_  = \new_[4155]_  & \new_[4152]_ ;
  assign \new_[4159]_  = ~A232 & ~A203;
  assign \new_[4163]_  = A301 & A236;
  assign \new_[4164]_  = A233 & \new_[4163]_ ;
  assign \new_[4165]_  = \new_[4164]_  & \new_[4159]_ ;
  assign \new_[4168]_  = A166 & A168;
  assign \new_[4171]_  = ~A202 & ~A201;
  assign \new_[4172]_  = \new_[4171]_  & \new_[4168]_ ;
  assign \new_[4175]_  = ~A232 & ~A203;
  assign \new_[4179]_  = A268 & A236;
  assign \new_[4180]_  = A233 & \new_[4179]_ ;
  assign \new_[4181]_  = \new_[4180]_  & \new_[4175]_ ;
  assign \new_[4184]_  = A166 & A168;
  assign \new_[4187]_  = ~A202 & ~A201;
  assign \new_[4188]_  = \new_[4187]_  & \new_[4184]_ ;
  assign \new_[4191]_  = A232 & ~A203;
  assign \new_[4195]_  = A301 & A236;
  assign \new_[4196]_  = ~A233 & \new_[4195]_ ;
  assign \new_[4197]_  = \new_[4196]_  & \new_[4191]_ ;
  assign \new_[4200]_  = A166 & A168;
  assign \new_[4203]_  = ~A202 & ~A201;
  assign \new_[4204]_  = \new_[4203]_  & \new_[4200]_ ;
  assign \new_[4207]_  = A232 & ~A203;
  assign \new_[4211]_  = A268 & A236;
  assign \new_[4212]_  = ~A233 & \new_[4211]_ ;
  assign \new_[4213]_  = \new_[4212]_  & \new_[4207]_ ;
  assign \new_[4216]_  = A166 & A168;
  assign \new_[4219]_  = A200 & A199;
  assign \new_[4220]_  = \new_[4219]_  & \new_[4216]_ ;
  assign \new_[4223]_  = ~A202 & ~A201;
  assign \new_[4227]_  = A300 & A299;
  assign \new_[4228]_  = A235 & \new_[4227]_ ;
  assign \new_[4229]_  = \new_[4228]_  & \new_[4223]_ ;
  assign \new_[4232]_  = A166 & A168;
  assign \new_[4235]_  = A200 & A199;
  assign \new_[4236]_  = \new_[4235]_  & \new_[4232]_ ;
  assign \new_[4239]_  = ~A202 & ~A201;
  assign \new_[4243]_  = A300 & A298;
  assign \new_[4244]_  = A235 & \new_[4243]_ ;
  assign \new_[4245]_  = \new_[4244]_  & \new_[4239]_ ;
  assign \new_[4248]_  = A166 & A168;
  assign \new_[4251]_  = A200 & A199;
  assign \new_[4252]_  = \new_[4251]_  & \new_[4248]_ ;
  assign \new_[4255]_  = ~A202 & ~A201;
  assign \new_[4259]_  = A267 & A265;
  assign \new_[4260]_  = A235 & \new_[4259]_ ;
  assign \new_[4261]_  = \new_[4260]_  & \new_[4255]_ ;
  assign \new_[4264]_  = A166 & A168;
  assign \new_[4267]_  = A200 & A199;
  assign \new_[4268]_  = \new_[4267]_  & \new_[4264]_ ;
  assign \new_[4271]_  = ~A202 & ~A201;
  assign \new_[4275]_  = A267 & A266;
  assign \new_[4276]_  = A235 & \new_[4275]_ ;
  assign \new_[4277]_  = \new_[4276]_  & \new_[4271]_ ;
  assign \new_[4280]_  = A166 & A168;
  assign \new_[4283]_  = A200 & A199;
  assign \new_[4284]_  = \new_[4283]_  & \new_[4280]_ ;
  assign \new_[4287]_  = ~A202 & ~A201;
  assign \new_[4291]_  = A301 & A234;
  assign \new_[4292]_  = A232 & \new_[4291]_ ;
  assign \new_[4293]_  = \new_[4292]_  & \new_[4287]_ ;
  assign \new_[4296]_  = A166 & A168;
  assign \new_[4299]_  = A200 & A199;
  assign \new_[4300]_  = \new_[4299]_  & \new_[4296]_ ;
  assign \new_[4303]_  = ~A202 & ~A201;
  assign \new_[4307]_  = A268 & A234;
  assign \new_[4308]_  = A232 & \new_[4307]_ ;
  assign \new_[4309]_  = \new_[4308]_  & \new_[4303]_ ;
  assign \new_[4312]_  = A166 & A168;
  assign \new_[4315]_  = A200 & A199;
  assign \new_[4316]_  = \new_[4315]_  & \new_[4312]_ ;
  assign \new_[4319]_  = ~A202 & ~A201;
  assign \new_[4323]_  = A301 & A234;
  assign \new_[4324]_  = A233 & \new_[4323]_ ;
  assign \new_[4325]_  = \new_[4324]_  & \new_[4319]_ ;
  assign \new_[4328]_  = A166 & A168;
  assign \new_[4331]_  = A200 & A199;
  assign \new_[4332]_  = \new_[4331]_  & \new_[4328]_ ;
  assign \new_[4335]_  = ~A202 & ~A201;
  assign \new_[4339]_  = A268 & A234;
  assign \new_[4340]_  = A233 & \new_[4339]_ ;
  assign \new_[4341]_  = \new_[4340]_  & \new_[4335]_ ;
  assign \new_[4344]_  = A166 & A168;
  assign \new_[4347]_  = ~A200 & ~A199;
  assign \new_[4348]_  = \new_[4347]_  & \new_[4344]_ ;
  assign \new_[4351]_  = A235 & ~A202;
  assign \new_[4355]_  = A302 & ~A299;
  assign \new_[4356]_  = A298 & \new_[4355]_ ;
  assign \new_[4357]_  = \new_[4356]_  & \new_[4351]_ ;
  assign \new_[4360]_  = A166 & A168;
  assign \new_[4363]_  = ~A200 & ~A199;
  assign \new_[4364]_  = \new_[4363]_  & \new_[4360]_ ;
  assign \new_[4367]_  = A235 & ~A202;
  assign \new_[4371]_  = A302 & A299;
  assign \new_[4372]_  = ~A298 & \new_[4371]_ ;
  assign \new_[4373]_  = \new_[4372]_  & \new_[4367]_ ;
  assign \new_[4376]_  = A166 & A168;
  assign \new_[4379]_  = ~A200 & ~A199;
  assign \new_[4380]_  = \new_[4379]_  & \new_[4376]_ ;
  assign \new_[4383]_  = A235 & ~A202;
  assign \new_[4387]_  = A269 & A266;
  assign \new_[4388]_  = ~A265 & \new_[4387]_ ;
  assign \new_[4389]_  = \new_[4388]_  & \new_[4383]_ ;
  assign \new_[4392]_  = A166 & A168;
  assign \new_[4395]_  = ~A200 & ~A199;
  assign \new_[4396]_  = \new_[4395]_  & \new_[4392]_ ;
  assign \new_[4399]_  = A235 & ~A202;
  assign \new_[4403]_  = A269 & ~A266;
  assign \new_[4404]_  = A265 & \new_[4403]_ ;
  assign \new_[4405]_  = \new_[4404]_  & \new_[4399]_ ;
  assign \new_[4408]_  = A166 & A168;
  assign \new_[4411]_  = ~A200 & ~A199;
  assign \new_[4412]_  = \new_[4411]_  & \new_[4408]_ ;
  assign \new_[4415]_  = A232 & ~A202;
  assign \new_[4419]_  = A300 & A299;
  assign \new_[4420]_  = A234 & \new_[4419]_ ;
  assign \new_[4421]_  = \new_[4420]_  & \new_[4415]_ ;
  assign \new_[4424]_  = A166 & A168;
  assign \new_[4427]_  = ~A200 & ~A199;
  assign \new_[4428]_  = \new_[4427]_  & \new_[4424]_ ;
  assign \new_[4431]_  = A232 & ~A202;
  assign \new_[4435]_  = A300 & A298;
  assign \new_[4436]_  = A234 & \new_[4435]_ ;
  assign \new_[4437]_  = \new_[4436]_  & \new_[4431]_ ;
  assign \new_[4440]_  = A166 & A168;
  assign \new_[4443]_  = ~A200 & ~A199;
  assign \new_[4444]_  = \new_[4443]_  & \new_[4440]_ ;
  assign \new_[4447]_  = A232 & ~A202;
  assign \new_[4451]_  = A267 & A265;
  assign \new_[4452]_  = A234 & \new_[4451]_ ;
  assign \new_[4453]_  = \new_[4452]_  & \new_[4447]_ ;
  assign \new_[4456]_  = A166 & A168;
  assign \new_[4459]_  = ~A200 & ~A199;
  assign \new_[4460]_  = \new_[4459]_  & \new_[4456]_ ;
  assign \new_[4463]_  = A232 & ~A202;
  assign \new_[4467]_  = A267 & A266;
  assign \new_[4468]_  = A234 & \new_[4467]_ ;
  assign \new_[4469]_  = \new_[4468]_  & \new_[4463]_ ;
  assign \new_[4472]_  = A166 & A168;
  assign \new_[4475]_  = ~A200 & ~A199;
  assign \new_[4476]_  = \new_[4475]_  & \new_[4472]_ ;
  assign \new_[4479]_  = A233 & ~A202;
  assign \new_[4483]_  = A300 & A299;
  assign \new_[4484]_  = A234 & \new_[4483]_ ;
  assign \new_[4485]_  = \new_[4484]_  & \new_[4479]_ ;
  assign \new_[4488]_  = A166 & A168;
  assign \new_[4491]_  = ~A200 & ~A199;
  assign \new_[4492]_  = \new_[4491]_  & \new_[4488]_ ;
  assign \new_[4495]_  = A233 & ~A202;
  assign \new_[4499]_  = A300 & A298;
  assign \new_[4500]_  = A234 & \new_[4499]_ ;
  assign \new_[4501]_  = \new_[4500]_  & \new_[4495]_ ;
  assign \new_[4504]_  = A166 & A168;
  assign \new_[4507]_  = ~A200 & ~A199;
  assign \new_[4508]_  = \new_[4507]_  & \new_[4504]_ ;
  assign \new_[4511]_  = A233 & ~A202;
  assign \new_[4515]_  = A267 & A265;
  assign \new_[4516]_  = A234 & \new_[4515]_ ;
  assign \new_[4517]_  = \new_[4516]_  & \new_[4511]_ ;
  assign \new_[4520]_  = A166 & A168;
  assign \new_[4523]_  = ~A200 & ~A199;
  assign \new_[4524]_  = \new_[4523]_  & \new_[4520]_ ;
  assign \new_[4527]_  = A233 & ~A202;
  assign \new_[4531]_  = A267 & A266;
  assign \new_[4532]_  = A234 & \new_[4531]_ ;
  assign \new_[4533]_  = \new_[4532]_  & \new_[4527]_ ;
  assign \new_[4536]_  = A166 & A168;
  assign \new_[4539]_  = ~A200 & ~A199;
  assign \new_[4540]_  = \new_[4539]_  & \new_[4536]_ ;
  assign \new_[4543]_  = ~A232 & ~A202;
  assign \new_[4547]_  = A301 & A236;
  assign \new_[4548]_  = A233 & \new_[4547]_ ;
  assign \new_[4549]_  = \new_[4548]_  & \new_[4543]_ ;
  assign \new_[4552]_  = A166 & A168;
  assign \new_[4555]_  = ~A200 & ~A199;
  assign \new_[4556]_  = \new_[4555]_  & \new_[4552]_ ;
  assign \new_[4559]_  = ~A232 & ~A202;
  assign \new_[4563]_  = A268 & A236;
  assign \new_[4564]_  = A233 & \new_[4563]_ ;
  assign \new_[4565]_  = \new_[4564]_  & \new_[4559]_ ;
  assign \new_[4568]_  = A166 & A168;
  assign \new_[4571]_  = ~A200 & ~A199;
  assign \new_[4572]_  = \new_[4571]_  & \new_[4568]_ ;
  assign \new_[4575]_  = A232 & ~A202;
  assign \new_[4579]_  = A301 & A236;
  assign \new_[4580]_  = ~A233 & \new_[4579]_ ;
  assign \new_[4581]_  = \new_[4580]_  & \new_[4575]_ ;
  assign \new_[4584]_  = A166 & A168;
  assign \new_[4587]_  = ~A200 & ~A199;
  assign \new_[4588]_  = \new_[4587]_  & \new_[4584]_ ;
  assign \new_[4591]_  = A232 & ~A202;
  assign \new_[4595]_  = A268 & A236;
  assign \new_[4596]_  = ~A233 & \new_[4595]_ ;
  assign \new_[4597]_  = \new_[4596]_  & \new_[4591]_ ;
  assign \new_[4600]_  = A167 & A168;
  assign \new_[4603]_  = ~A202 & ~A201;
  assign \new_[4604]_  = \new_[4603]_  & \new_[4600]_ ;
  assign \new_[4607]_  = A235 & ~A203;
  assign \new_[4611]_  = A302 & ~A299;
  assign \new_[4612]_  = A298 & \new_[4611]_ ;
  assign \new_[4613]_  = \new_[4612]_  & \new_[4607]_ ;
  assign \new_[4616]_  = A167 & A168;
  assign \new_[4619]_  = ~A202 & ~A201;
  assign \new_[4620]_  = \new_[4619]_  & \new_[4616]_ ;
  assign \new_[4623]_  = A235 & ~A203;
  assign \new_[4627]_  = A302 & A299;
  assign \new_[4628]_  = ~A298 & \new_[4627]_ ;
  assign \new_[4629]_  = \new_[4628]_  & \new_[4623]_ ;
  assign \new_[4632]_  = A167 & A168;
  assign \new_[4635]_  = ~A202 & ~A201;
  assign \new_[4636]_  = \new_[4635]_  & \new_[4632]_ ;
  assign \new_[4639]_  = A235 & ~A203;
  assign \new_[4643]_  = A269 & A266;
  assign \new_[4644]_  = ~A265 & \new_[4643]_ ;
  assign \new_[4645]_  = \new_[4644]_  & \new_[4639]_ ;
  assign \new_[4648]_  = A167 & A168;
  assign \new_[4651]_  = ~A202 & ~A201;
  assign \new_[4652]_  = \new_[4651]_  & \new_[4648]_ ;
  assign \new_[4655]_  = A235 & ~A203;
  assign \new_[4659]_  = A269 & ~A266;
  assign \new_[4660]_  = A265 & \new_[4659]_ ;
  assign \new_[4661]_  = \new_[4660]_  & \new_[4655]_ ;
  assign \new_[4664]_  = A167 & A168;
  assign \new_[4667]_  = ~A202 & ~A201;
  assign \new_[4668]_  = \new_[4667]_  & \new_[4664]_ ;
  assign \new_[4671]_  = A232 & ~A203;
  assign \new_[4675]_  = A300 & A299;
  assign \new_[4676]_  = A234 & \new_[4675]_ ;
  assign \new_[4677]_  = \new_[4676]_  & \new_[4671]_ ;
  assign \new_[4680]_  = A167 & A168;
  assign \new_[4683]_  = ~A202 & ~A201;
  assign \new_[4684]_  = \new_[4683]_  & \new_[4680]_ ;
  assign \new_[4687]_  = A232 & ~A203;
  assign \new_[4691]_  = A300 & A298;
  assign \new_[4692]_  = A234 & \new_[4691]_ ;
  assign \new_[4693]_  = \new_[4692]_  & \new_[4687]_ ;
  assign \new_[4696]_  = A167 & A168;
  assign \new_[4699]_  = ~A202 & ~A201;
  assign \new_[4700]_  = \new_[4699]_  & \new_[4696]_ ;
  assign \new_[4703]_  = A232 & ~A203;
  assign \new_[4707]_  = A267 & A265;
  assign \new_[4708]_  = A234 & \new_[4707]_ ;
  assign \new_[4709]_  = \new_[4708]_  & \new_[4703]_ ;
  assign \new_[4712]_  = A167 & A168;
  assign \new_[4715]_  = ~A202 & ~A201;
  assign \new_[4716]_  = \new_[4715]_  & \new_[4712]_ ;
  assign \new_[4719]_  = A232 & ~A203;
  assign \new_[4723]_  = A267 & A266;
  assign \new_[4724]_  = A234 & \new_[4723]_ ;
  assign \new_[4725]_  = \new_[4724]_  & \new_[4719]_ ;
  assign \new_[4728]_  = A167 & A168;
  assign \new_[4731]_  = ~A202 & ~A201;
  assign \new_[4732]_  = \new_[4731]_  & \new_[4728]_ ;
  assign \new_[4735]_  = A233 & ~A203;
  assign \new_[4739]_  = A300 & A299;
  assign \new_[4740]_  = A234 & \new_[4739]_ ;
  assign \new_[4741]_  = \new_[4740]_  & \new_[4735]_ ;
  assign \new_[4744]_  = A167 & A168;
  assign \new_[4747]_  = ~A202 & ~A201;
  assign \new_[4748]_  = \new_[4747]_  & \new_[4744]_ ;
  assign \new_[4751]_  = A233 & ~A203;
  assign \new_[4755]_  = A300 & A298;
  assign \new_[4756]_  = A234 & \new_[4755]_ ;
  assign \new_[4757]_  = \new_[4756]_  & \new_[4751]_ ;
  assign \new_[4760]_  = A167 & A168;
  assign \new_[4763]_  = ~A202 & ~A201;
  assign \new_[4764]_  = \new_[4763]_  & \new_[4760]_ ;
  assign \new_[4767]_  = A233 & ~A203;
  assign \new_[4771]_  = A267 & A265;
  assign \new_[4772]_  = A234 & \new_[4771]_ ;
  assign \new_[4773]_  = \new_[4772]_  & \new_[4767]_ ;
  assign \new_[4776]_  = A167 & A168;
  assign \new_[4779]_  = ~A202 & ~A201;
  assign \new_[4780]_  = \new_[4779]_  & \new_[4776]_ ;
  assign \new_[4783]_  = A233 & ~A203;
  assign \new_[4787]_  = A267 & A266;
  assign \new_[4788]_  = A234 & \new_[4787]_ ;
  assign \new_[4789]_  = \new_[4788]_  & \new_[4783]_ ;
  assign \new_[4792]_  = A167 & A168;
  assign \new_[4795]_  = ~A202 & ~A201;
  assign \new_[4796]_  = \new_[4795]_  & \new_[4792]_ ;
  assign \new_[4799]_  = ~A232 & ~A203;
  assign \new_[4803]_  = A301 & A236;
  assign \new_[4804]_  = A233 & \new_[4803]_ ;
  assign \new_[4805]_  = \new_[4804]_  & \new_[4799]_ ;
  assign \new_[4808]_  = A167 & A168;
  assign \new_[4811]_  = ~A202 & ~A201;
  assign \new_[4812]_  = \new_[4811]_  & \new_[4808]_ ;
  assign \new_[4815]_  = ~A232 & ~A203;
  assign \new_[4819]_  = A268 & A236;
  assign \new_[4820]_  = A233 & \new_[4819]_ ;
  assign \new_[4821]_  = \new_[4820]_  & \new_[4815]_ ;
  assign \new_[4824]_  = A167 & A168;
  assign \new_[4827]_  = ~A202 & ~A201;
  assign \new_[4828]_  = \new_[4827]_  & \new_[4824]_ ;
  assign \new_[4831]_  = A232 & ~A203;
  assign \new_[4835]_  = A301 & A236;
  assign \new_[4836]_  = ~A233 & \new_[4835]_ ;
  assign \new_[4837]_  = \new_[4836]_  & \new_[4831]_ ;
  assign \new_[4840]_  = A167 & A168;
  assign \new_[4843]_  = ~A202 & ~A201;
  assign \new_[4844]_  = \new_[4843]_  & \new_[4840]_ ;
  assign \new_[4847]_  = A232 & ~A203;
  assign \new_[4851]_  = A268 & A236;
  assign \new_[4852]_  = ~A233 & \new_[4851]_ ;
  assign \new_[4853]_  = \new_[4852]_  & \new_[4847]_ ;
  assign \new_[4856]_  = A167 & A168;
  assign \new_[4859]_  = A200 & A199;
  assign \new_[4860]_  = \new_[4859]_  & \new_[4856]_ ;
  assign \new_[4863]_  = ~A202 & ~A201;
  assign \new_[4867]_  = A300 & A299;
  assign \new_[4868]_  = A235 & \new_[4867]_ ;
  assign \new_[4869]_  = \new_[4868]_  & \new_[4863]_ ;
  assign \new_[4872]_  = A167 & A168;
  assign \new_[4875]_  = A200 & A199;
  assign \new_[4876]_  = \new_[4875]_  & \new_[4872]_ ;
  assign \new_[4879]_  = ~A202 & ~A201;
  assign \new_[4883]_  = A300 & A298;
  assign \new_[4884]_  = A235 & \new_[4883]_ ;
  assign \new_[4885]_  = \new_[4884]_  & \new_[4879]_ ;
  assign \new_[4888]_  = A167 & A168;
  assign \new_[4891]_  = A200 & A199;
  assign \new_[4892]_  = \new_[4891]_  & \new_[4888]_ ;
  assign \new_[4895]_  = ~A202 & ~A201;
  assign \new_[4899]_  = A267 & A265;
  assign \new_[4900]_  = A235 & \new_[4899]_ ;
  assign \new_[4901]_  = \new_[4900]_  & \new_[4895]_ ;
  assign \new_[4904]_  = A167 & A168;
  assign \new_[4907]_  = A200 & A199;
  assign \new_[4908]_  = \new_[4907]_  & \new_[4904]_ ;
  assign \new_[4911]_  = ~A202 & ~A201;
  assign \new_[4915]_  = A267 & A266;
  assign \new_[4916]_  = A235 & \new_[4915]_ ;
  assign \new_[4917]_  = \new_[4916]_  & \new_[4911]_ ;
  assign \new_[4920]_  = A167 & A168;
  assign \new_[4923]_  = A200 & A199;
  assign \new_[4924]_  = \new_[4923]_  & \new_[4920]_ ;
  assign \new_[4927]_  = ~A202 & ~A201;
  assign \new_[4931]_  = A301 & A234;
  assign \new_[4932]_  = A232 & \new_[4931]_ ;
  assign \new_[4933]_  = \new_[4932]_  & \new_[4927]_ ;
  assign \new_[4936]_  = A167 & A168;
  assign \new_[4939]_  = A200 & A199;
  assign \new_[4940]_  = \new_[4939]_  & \new_[4936]_ ;
  assign \new_[4943]_  = ~A202 & ~A201;
  assign \new_[4947]_  = A268 & A234;
  assign \new_[4948]_  = A232 & \new_[4947]_ ;
  assign \new_[4949]_  = \new_[4948]_  & \new_[4943]_ ;
  assign \new_[4952]_  = A167 & A168;
  assign \new_[4955]_  = A200 & A199;
  assign \new_[4956]_  = \new_[4955]_  & \new_[4952]_ ;
  assign \new_[4959]_  = ~A202 & ~A201;
  assign \new_[4963]_  = A301 & A234;
  assign \new_[4964]_  = A233 & \new_[4963]_ ;
  assign \new_[4965]_  = \new_[4964]_  & \new_[4959]_ ;
  assign \new_[4968]_  = A167 & A168;
  assign \new_[4971]_  = A200 & A199;
  assign \new_[4972]_  = \new_[4971]_  & \new_[4968]_ ;
  assign \new_[4975]_  = ~A202 & ~A201;
  assign \new_[4979]_  = A268 & A234;
  assign \new_[4980]_  = A233 & \new_[4979]_ ;
  assign \new_[4981]_  = \new_[4980]_  & \new_[4975]_ ;
  assign \new_[4984]_  = A167 & A168;
  assign \new_[4987]_  = ~A200 & ~A199;
  assign \new_[4988]_  = \new_[4987]_  & \new_[4984]_ ;
  assign \new_[4991]_  = A235 & ~A202;
  assign \new_[4995]_  = A302 & ~A299;
  assign \new_[4996]_  = A298 & \new_[4995]_ ;
  assign \new_[4997]_  = \new_[4996]_  & \new_[4991]_ ;
  assign \new_[5000]_  = A167 & A168;
  assign \new_[5003]_  = ~A200 & ~A199;
  assign \new_[5004]_  = \new_[5003]_  & \new_[5000]_ ;
  assign \new_[5007]_  = A235 & ~A202;
  assign \new_[5011]_  = A302 & A299;
  assign \new_[5012]_  = ~A298 & \new_[5011]_ ;
  assign \new_[5013]_  = \new_[5012]_  & \new_[5007]_ ;
  assign \new_[5016]_  = A167 & A168;
  assign \new_[5019]_  = ~A200 & ~A199;
  assign \new_[5020]_  = \new_[5019]_  & \new_[5016]_ ;
  assign \new_[5023]_  = A235 & ~A202;
  assign \new_[5027]_  = A269 & A266;
  assign \new_[5028]_  = ~A265 & \new_[5027]_ ;
  assign \new_[5029]_  = \new_[5028]_  & \new_[5023]_ ;
  assign \new_[5032]_  = A167 & A168;
  assign \new_[5035]_  = ~A200 & ~A199;
  assign \new_[5036]_  = \new_[5035]_  & \new_[5032]_ ;
  assign \new_[5039]_  = A235 & ~A202;
  assign \new_[5043]_  = A269 & ~A266;
  assign \new_[5044]_  = A265 & \new_[5043]_ ;
  assign \new_[5045]_  = \new_[5044]_  & \new_[5039]_ ;
  assign \new_[5048]_  = A167 & A168;
  assign \new_[5051]_  = ~A200 & ~A199;
  assign \new_[5052]_  = \new_[5051]_  & \new_[5048]_ ;
  assign \new_[5055]_  = A232 & ~A202;
  assign \new_[5059]_  = A300 & A299;
  assign \new_[5060]_  = A234 & \new_[5059]_ ;
  assign \new_[5061]_  = \new_[5060]_  & \new_[5055]_ ;
  assign \new_[5064]_  = A167 & A168;
  assign \new_[5067]_  = ~A200 & ~A199;
  assign \new_[5068]_  = \new_[5067]_  & \new_[5064]_ ;
  assign \new_[5071]_  = A232 & ~A202;
  assign \new_[5075]_  = A300 & A298;
  assign \new_[5076]_  = A234 & \new_[5075]_ ;
  assign \new_[5077]_  = \new_[5076]_  & \new_[5071]_ ;
  assign \new_[5080]_  = A167 & A168;
  assign \new_[5083]_  = ~A200 & ~A199;
  assign \new_[5084]_  = \new_[5083]_  & \new_[5080]_ ;
  assign \new_[5087]_  = A232 & ~A202;
  assign \new_[5091]_  = A267 & A265;
  assign \new_[5092]_  = A234 & \new_[5091]_ ;
  assign \new_[5093]_  = \new_[5092]_  & \new_[5087]_ ;
  assign \new_[5096]_  = A167 & A168;
  assign \new_[5099]_  = ~A200 & ~A199;
  assign \new_[5100]_  = \new_[5099]_  & \new_[5096]_ ;
  assign \new_[5103]_  = A232 & ~A202;
  assign \new_[5107]_  = A267 & A266;
  assign \new_[5108]_  = A234 & \new_[5107]_ ;
  assign \new_[5109]_  = \new_[5108]_  & \new_[5103]_ ;
  assign \new_[5112]_  = A167 & A168;
  assign \new_[5115]_  = ~A200 & ~A199;
  assign \new_[5116]_  = \new_[5115]_  & \new_[5112]_ ;
  assign \new_[5119]_  = A233 & ~A202;
  assign \new_[5123]_  = A300 & A299;
  assign \new_[5124]_  = A234 & \new_[5123]_ ;
  assign \new_[5125]_  = \new_[5124]_  & \new_[5119]_ ;
  assign \new_[5128]_  = A167 & A168;
  assign \new_[5131]_  = ~A200 & ~A199;
  assign \new_[5132]_  = \new_[5131]_  & \new_[5128]_ ;
  assign \new_[5135]_  = A233 & ~A202;
  assign \new_[5139]_  = A300 & A298;
  assign \new_[5140]_  = A234 & \new_[5139]_ ;
  assign \new_[5141]_  = \new_[5140]_  & \new_[5135]_ ;
  assign \new_[5144]_  = A167 & A168;
  assign \new_[5147]_  = ~A200 & ~A199;
  assign \new_[5148]_  = \new_[5147]_  & \new_[5144]_ ;
  assign \new_[5151]_  = A233 & ~A202;
  assign \new_[5155]_  = A267 & A265;
  assign \new_[5156]_  = A234 & \new_[5155]_ ;
  assign \new_[5157]_  = \new_[5156]_  & \new_[5151]_ ;
  assign \new_[5160]_  = A167 & A168;
  assign \new_[5163]_  = ~A200 & ~A199;
  assign \new_[5164]_  = \new_[5163]_  & \new_[5160]_ ;
  assign \new_[5167]_  = A233 & ~A202;
  assign \new_[5171]_  = A267 & A266;
  assign \new_[5172]_  = A234 & \new_[5171]_ ;
  assign \new_[5173]_  = \new_[5172]_  & \new_[5167]_ ;
  assign \new_[5176]_  = A167 & A168;
  assign \new_[5179]_  = ~A200 & ~A199;
  assign \new_[5180]_  = \new_[5179]_  & \new_[5176]_ ;
  assign \new_[5183]_  = ~A232 & ~A202;
  assign \new_[5187]_  = A301 & A236;
  assign \new_[5188]_  = A233 & \new_[5187]_ ;
  assign \new_[5189]_  = \new_[5188]_  & \new_[5183]_ ;
  assign \new_[5192]_  = A167 & A168;
  assign \new_[5195]_  = ~A200 & ~A199;
  assign \new_[5196]_  = \new_[5195]_  & \new_[5192]_ ;
  assign \new_[5199]_  = ~A232 & ~A202;
  assign \new_[5203]_  = A268 & A236;
  assign \new_[5204]_  = A233 & \new_[5203]_ ;
  assign \new_[5205]_  = \new_[5204]_  & \new_[5199]_ ;
  assign \new_[5208]_  = A167 & A168;
  assign \new_[5211]_  = ~A200 & ~A199;
  assign \new_[5212]_  = \new_[5211]_  & \new_[5208]_ ;
  assign \new_[5215]_  = A232 & ~A202;
  assign \new_[5219]_  = A301 & A236;
  assign \new_[5220]_  = ~A233 & \new_[5219]_ ;
  assign \new_[5221]_  = \new_[5220]_  & \new_[5215]_ ;
  assign \new_[5224]_  = A167 & A168;
  assign \new_[5227]_  = ~A200 & ~A199;
  assign \new_[5228]_  = \new_[5227]_  & \new_[5224]_ ;
  assign \new_[5231]_  = A232 & ~A202;
  assign \new_[5235]_  = A268 & A236;
  assign \new_[5236]_  = ~A233 & \new_[5235]_ ;
  assign \new_[5237]_  = \new_[5236]_  & \new_[5231]_ ;
  assign \new_[5240]_  = A167 & A170;
  assign \new_[5243]_  = ~A201 & ~A166;
  assign \new_[5244]_  = \new_[5243]_  & \new_[5240]_ ;
  assign \new_[5247]_  = ~A203 & ~A202;
  assign \new_[5251]_  = A300 & A299;
  assign \new_[5252]_  = A235 & \new_[5251]_ ;
  assign \new_[5253]_  = \new_[5252]_  & \new_[5247]_ ;
  assign \new_[5256]_  = A167 & A170;
  assign \new_[5259]_  = ~A201 & ~A166;
  assign \new_[5260]_  = \new_[5259]_  & \new_[5256]_ ;
  assign \new_[5263]_  = ~A203 & ~A202;
  assign \new_[5267]_  = A300 & A298;
  assign \new_[5268]_  = A235 & \new_[5267]_ ;
  assign \new_[5269]_  = \new_[5268]_  & \new_[5263]_ ;
  assign \new_[5272]_  = A167 & A170;
  assign \new_[5275]_  = ~A201 & ~A166;
  assign \new_[5276]_  = \new_[5275]_  & \new_[5272]_ ;
  assign \new_[5279]_  = ~A203 & ~A202;
  assign \new_[5283]_  = A267 & A265;
  assign \new_[5284]_  = A235 & \new_[5283]_ ;
  assign \new_[5285]_  = \new_[5284]_  & \new_[5279]_ ;
  assign \new_[5288]_  = A167 & A170;
  assign \new_[5291]_  = ~A201 & ~A166;
  assign \new_[5292]_  = \new_[5291]_  & \new_[5288]_ ;
  assign \new_[5295]_  = ~A203 & ~A202;
  assign \new_[5299]_  = A267 & A266;
  assign \new_[5300]_  = A235 & \new_[5299]_ ;
  assign \new_[5301]_  = \new_[5300]_  & \new_[5295]_ ;
  assign \new_[5304]_  = A167 & A170;
  assign \new_[5307]_  = ~A201 & ~A166;
  assign \new_[5308]_  = \new_[5307]_  & \new_[5304]_ ;
  assign \new_[5311]_  = ~A203 & ~A202;
  assign \new_[5315]_  = A301 & A234;
  assign \new_[5316]_  = A232 & \new_[5315]_ ;
  assign \new_[5317]_  = \new_[5316]_  & \new_[5311]_ ;
  assign \new_[5320]_  = A167 & A170;
  assign \new_[5323]_  = ~A201 & ~A166;
  assign \new_[5324]_  = \new_[5323]_  & \new_[5320]_ ;
  assign \new_[5327]_  = ~A203 & ~A202;
  assign \new_[5331]_  = A268 & A234;
  assign \new_[5332]_  = A232 & \new_[5331]_ ;
  assign \new_[5333]_  = \new_[5332]_  & \new_[5327]_ ;
  assign \new_[5336]_  = A167 & A170;
  assign \new_[5339]_  = ~A201 & ~A166;
  assign \new_[5340]_  = \new_[5339]_  & \new_[5336]_ ;
  assign \new_[5343]_  = ~A203 & ~A202;
  assign \new_[5347]_  = A301 & A234;
  assign \new_[5348]_  = A233 & \new_[5347]_ ;
  assign \new_[5349]_  = \new_[5348]_  & \new_[5343]_ ;
  assign \new_[5352]_  = A167 & A170;
  assign \new_[5355]_  = ~A201 & ~A166;
  assign \new_[5356]_  = \new_[5355]_  & \new_[5352]_ ;
  assign \new_[5359]_  = ~A203 & ~A202;
  assign \new_[5363]_  = A268 & A234;
  assign \new_[5364]_  = A233 & \new_[5363]_ ;
  assign \new_[5365]_  = \new_[5364]_  & \new_[5359]_ ;
  assign \new_[5368]_  = A167 & A170;
  assign \new_[5371]_  = A199 & ~A166;
  assign \new_[5372]_  = \new_[5371]_  & \new_[5368]_ ;
  assign \new_[5375]_  = ~A201 & A200;
  assign \new_[5379]_  = A301 & A235;
  assign \new_[5380]_  = ~A202 & \new_[5379]_ ;
  assign \new_[5381]_  = \new_[5380]_  & \new_[5375]_ ;
  assign \new_[5384]_  = A167 & A170;
  assign \new_[5387]_  = A199 & ~A166;
  assign \new_[5388]_  = \new_[5387]_  & \new_[5384]_ ;
  assign \new_[5391]_  = ~A201 & A200;
  assign \new_[5395]_  = A268 & A235;
  assign \new_[5396]_  = ~A202 & \new_[5395]_ ;
  assign \new_[5397]_  = \new_[5396]_  & \new_[5391]_ ;
  assign \new_[5400]_  = A167 & A170;
  assign \new_[5403]_  = ~A199 & ~A166;
  assign \new_[5404]_  = \new_[5403]_  & \new_[5400]_ ;
  assign \new_[5407]_  = ~A202 & ~A200;
  assign \new_[5411]_  = A300 & A299;
  assign \new_[5412]_  = A235 & \new_[5411]_ ;
  assign \new_[5413]_  = \new_[5412]_  & \new_[5407]_ ;
  assign \new_[5416]_  = A167 & A170;
  assign \new_[5419]_  = ~A199 & ~A166;
  assign \new_[5420]_  = \new_[5419]_  & \new_[5416]_ ;
  assign \new_[5423]_  = ~A202 & ~A200;
  assign \new_[5427]_  = A300 & A298;
  assign \new_[5428]_  = A235 & \new_[5427]_ ;
  assign \new_[5429]_  = \new_[5428]_  & \new_[5423]_ ;
  assign \new_[5432]_  = A167 & A170;
  assign \new_[5435]_  = ~A199 & ~A166;
  assign \new_[5436]_  = \new_[5435]_  & \new_[5432]_ ;
  assign \new_[5439]_  = ~A202 & ~A200;
  assign \new_[5443]_  = A267 & A265;
  assign \new_[5444]_  = A235 & \new_[5443]_ ;
  assign \new_[5445]_  = \new_[5444]_  & \new_[5439]_ ;
  assign \new_[5448]_  = A167 & A170;
  assign \new_[5451]_  = ~A199 & ~A166;
  assign \new_[5452]_  = \new_[5451]_  & \new_[5448]_ ;
  assign \new_[5455]_  = ~A202 & ~A200;
  assign \new_[5459]_  = A267 & A266;
  assign \new_[5460]_  = A235 & \new_[5459]_ ;
  assign \new_[5461]_  = \new_[5460]_  & \new_[5455]_ ;
  assign \new_[5464]_  = A167 & A170;
  assign \new_[5467]_  = ~A199 & ~A166;
  assign \new_[5468]_  = \new_[5467]_  & \new_[5464]_ ;
  assign \new_[5471]_  = ~A202 & ~A200;
  assign \new_[5475]_  = A301 & A234;
  assign \new_[5476]_  = A232 & \new_[5475]_ ;
  assign \new_[5477]_  = \new_[5476]_  & \new_[5471]_ ;
  assign \new_[5480]_  = A167 & A170;
  assign \new_[5483]_  = ~A199 & ~A166;
  assign \new_[5484]_  = \new_[5483]_  & \new_[5480]_ ;
  assign \new_[5487]_  = ~A202 & ~A200;
  assign \new_[5491]_  = A268 & A234;
  assign \new_[5492]_  = A232 & \new_[5491]_ ;
  assign \new_[5493]_  = \new_[5492]_  & \new_[5487]_ ;
  assign \new_[5496]_  = A167 & A170;
  assign \new_[5499]_  = ~A199 & ~A166;
  assign \new_[5500]_  = \new_[5499]_  & \new_[5496]_ ;
  assign \new_[5503]_  = ~A202 & ~A200;
  assign \new_[5507]_  = A301 & A234;
  assign \new_[5508]_  = A233 & \new_[5507]_ ;
  assign \new_[5509]_  = \new_[5508]_  & \new_[5503]_ ;
  assign \new_[5512]_  = A167 & A170;
  assign \new_[5515]_  = ~A199 & ~A166;
  assign \new_[5516]_  = \new_[5515]_  & \new_[5512]_ ;
  assign \new_[5519]_  = ~A202 & ~A200;
  assign \new_[5523]_  = A268 & A234;
  assign \new_[5524]_  = A233 & \new_[5523]_ ;
  assign \new_[5525]_  = \new_[5524]_  & \new_[5519]_ ;
  assign \new_[5528]_  = ~A167 & A170;
  assign \new_[5531]_  = ~A201 & A166;
  assign \new_[5532]_  = \new_[5531]_  & \new_[5528]_ ;
  assign \new_[5535]_  = ~A203 & ~A202;
  assign \new_[5539]_  = A300 & A299;
  assign \new_[5540]_  = A235 & \new_[5539]_ ;
  assign \new_[5541]_  = \new_[5540]_  & \new_[5535]_ ;
  assign \new_[5544]_  = ~A167 & A170;
  assign \new_[5547]_  = ~A201 & A166;
  assign \new_[5548]_  = \new_[5547]_  & \new_[5544]_ ;
  assign \new_[5551]_  = ~A203 & ~A202;
  assign \new_[5555]_  = A300 & A298;
  assign \new_[5556]_  = A235 & \new_[5555]_ ;
  assign \new_[5557]_  = \new_[5556]_  & \new_[5551]_ ;
  assign \new_[5560]_  = ~A167 & A170;
  assign \new_[5563]_  = ~A201 & A166;
  assign \new_[5564]_  = \new_[5563]_  & \new_[5560]_ ;
  assign \new_[5567]_  = ~A203 & ~A202;
  assign \new_[5571]_  = A267 & A265;
  assign \new_[5572]_  = A235 & \new_[5571]_ ;
  assign \new_[5573]_  = \new_[5572]_  & \new_[5567]_ ;
  assign \new_[5576]_  = ~A167 & A170;
  assign \new_[5579]_  = ~A201 & A166;
  assign \new_[5580]_  = \new_[5579]_  & \new_[5576]_ ;
  assign \new_[5583]_  = ~A203 & ~A202;
  assign \new_[5587]_  = A267 & A266;
  assign \new_[5588]_  = A235 & \new_[5587]_ ;
  assign \new_[5589]_  = \new_[5588]_  & \new_[5583]_ ;
  assign \new_[5592]_  = ~A167 & A170;
  assign \new_[5595]_  = ~A201 & A166;
  assign \new_[5596]_  = \new_[5595]_  & \new_[5592]_ ;
  assign \new_[5599]_  = ~A203 & ~A202;
  assign \new_[5603]_  = A301 & A234;
  assign \new_[5604]_  = A232 & \new_[5603]_ ;
  assign \new_[5605]_  = \new_[5604]_  & \new_[5599]_ ;
  assign \new_[5608]_  = ~A167 & A170;
  assign \new_[5611]_  = ~A201 & A166;
  assign \new_[5612]_  = \new_[5611]_  & \new_[5608]_ ;
  assign \new_[5615]_  = ~A203 & ~A202;
  assign \new_[5619]_  = A268 & A234;
  assign \new_[5620]_  = A232 & \new_[5619]_ ;
  assign \new_[5621]_  = \new_[5620]_  & \new_[5615]_ ;
  assign \new_[5624]_  = ~A167 & A170;
  assign \new_[5627]_  = ~A201 & A166;
  assign \new_[5628]_  = \new_[5627]_  & \new_[5624]_ ;
  assign \new_[5631]_  = ~A203 & ~A202;
  assign \new_[5635]_  = A301 & A234;
  assign \new_[5636]_  = A233 & \new_[5635]_ ;
  assign \new_[5637]_  = \new_[5636]_  & \new_[5631]_ ;
  assign \new_[5640]_  = ~A167 & A170;
  assign \new_[5643]_  = ~A201 & A166;
  assign \new_[5644]_  = \new_[5643]_  & \new_[5640]_ ;
  assign \new_[5647]_  = ~A203 & ~A202;
  assign \new_[5651]_  = A268 & A234;
  assign \new_[5652]_  = A233 & \new_[5651]_ ;
  assign \new_[5653]_  = \new_[5652]_  & \new_[5647]_ ;
  assign \new_[5656]_  = ~A167 & A170;
  assign \new_[5659]_  = A199 & A166;
  assign \new_[5660]_  = \new_[5659]_  & \new_[5656]_ ;
  assign \new_[5663]_  = ~A201 & A200;
  assign \new_[5667]_  = A301 & A235;
  assign \new_[5668]_  = ~A202 & \new_[5667]_ ;
  assign \new_[5669]_  = \new_[5668]_  & \new_[5663]_ ;
  assign \new_[5672]_  = ~A167 & A170;
  assign \new_[5675]_  = A199 & A166;
  assign \new_[5676]_  = \new_[5675]_  & \new_[5672]_ ;
  assign \new_[5679]_  = ~A201 & A200;
  assign \new_[5683]_  = A268 & A235;
  assign \new_[5684]_  = ~A202 & \new_[5683]_ ;
  assign \new_[5685]_  = \new_[5684]_  & \new_[5679]_ ;
  assign \new_[5688]_  = ~A167 & A170;
  assign \new_[5691]_  = ~A199 & A166;
  assign \new_[5692]_  = \new_[5691]_  & \new_[5688]_ ;
  assign \new_[5695]_  = ~A202 & ~A200;
  assign \new_[5699]_  = A300 & A299;
  assign \new_[5700]_  = A235 & \new_[5699]_ ;
  assign \new_[5701]_  = \new_[5700]_  & \new_[5695]_ ;
  assign \new_[5704]_  = ~A167 & A170;
  assign \new_[5707]_  = ~A199 & A166;
  assign \new_[5708]_  = \new_[5707]_  & \new_[5704]_ ;
  assign \new_[5711]_  = ~A202 & ~A200;
  assign \new_[5715]_  = A300 & A298;
  assign \new_[5716]_  = A235 & \new_[5715]_ ;
  assign \new_[5717]_  = \new_[5716]_  & \new_[5711]_ ;
  assign \new_[5720]_  = ~A167 & A170;
  assign \new_[5723]_  = ~A199 & A166;
  assign \new_[5724]_  = \new_[5723]_  & \new_[5720]_ ;
  assign \new_[5727]_  = ~A202 & ~A200;
  assign \new_[5731]_  = A267 & A265;
  assign \new_[5732]_  = A235 & \new_[5731]_ ;
  assign \new_[5733]_  = \new_[5732]_  & \new_[5727]_ ;
  assign \new_[5736]_  = ~A167 & A170;
  assign \new_[5739]_  = ~A199 & A166;
  assign \new_[5740]_  = \new_[5739]_  & \new_[5736]_ ;
  assign \new_[5743]_  = ~A202 & ~A200;
  assign \new_[5747]_  = A267 & A266;
  assign \new_[5748]_  = A235 & \new_[5747]_ ;
  assign \new_[5749]_  = \new_[5748]_  & \new_[5743]_ ;
  assign \new_[5752]_  = ~A167 & A170;
  assign \new_[5755]_  = ~A199 & A166;
  assign \new_[5756]_  = \new_[5755]_  & \new_[5752]_ ;
  assign \new_[5759]_  = ~A202 & ~A200;
  assign \new_[5763]_  = A301 & A234;
  assign \new_[5764]_  = A232 & \new_[5763]_ ;
  assign \new_[5765]_  = \new_[5764]_  & \new_[5759]_ ;
  assign \new_[5768]_  = ~A167 & A170;
  assign \new_[5771]_  = ~A199 & A166;
  assign \new_[5772]_  = \new_[5771]_  & \new_[5768]_ ;
  assign \new_[5775]_  = ~A202 & ~A200;
  assign \new_[5779]_  = A268 & A234;
  assign \new_[5780]_  = A232 & \new_[5779]_ ;
  assign \new_[5781]_  = \new_[5780]_  & \new_[5775]_ ;
  assign \new_[5784]_  = ~A167 & A170;
  assign \new_[5787]_  = ~A199 & A166;
  assign \new_[5788]_  = \new_[5787]_  & \new_[5784]_ ;
  assign \new_[5791]_  = ~A202 & ~A200;
  assign \new_[5795]_  = A301 & A234;
  assign \new_[5796]_  = A233 & \new_[5795]_ ;
  assign \new_[5797]_  = \new_[5796]_  & \new_[5791]_ ;
  assign \new_[5800]_  = ~A167 & A170;
  assign \new_[5803]_  = ~A199 & A166;
  assign \new_[5804]_  = \new_[5803]_  & \new_[5800]_ ;
  assign \new_[5807]_  = ~A202 & ~A200;
  assign \new_[5811]_  = A268 & A234;
  assign \new_[5812]_  = A233 & \new_[5811]_ ;
  assign \new_[5813]_  = \new_[5812]_  & \new_[5807]_ ;
  assign \new_[5816]_  = ~A201 & A169;
  assign \new_[5819]_  = ~A203 & ~A202;
  assign \new_[5820]_  = \new_[5819]_  & \new_[5816]_ ;
  assign \new_[5823]_  = A234 & A232;
  assign \new_[5827]_  = A302 & ~A299;
  assign \new_[5828]_  = A298 & \new_[5827]_ ;
  assign \new_[5829]_  = \new_[5828]_  & \new_[5823]_ ;
  assign \new_[5832]_  = ~A201 & A169;
  assign \new_[5835]_  = ~A203 & ~A202;
  assign \new_[5836]_  = \new_[5835]_  & \new_[5832]_ ;
  assign \new_[5839]_  = A234 & A232;
  assign \new_[5843]_  = A302 & A299;
  assign \new_[5844]_  = ~A298 & \new_[5843]_ ;
  assign \new_[5845]_  = \new_[5844]_  & \new_[5839]_ ;
  assign \new_[5848]_  = ~A201 & A169;
  assign \new_[5851]_  = ~A203 & ~A202;
  assign \new_[5852]_  = \new_[5851]_  & \new_[5848]_ ;
  assign \new_[5855]_  = A234 & A232;
  assign \new_[5859]_  = A269 & A266;
  assign \new_[5860]_  = ~A265 & \new_[5859]_ ;
  assign \new_[5861]_  = \new_[5860]_  & \new_[5855]_ ;
  assign \new_[5864]_  = ~A201 & A169;
  assign \new_[5867]_  = ~A203 & ~A202;
  assign \new_[5868]_  = \new_[5867]_  & \new_[5864]_ ;
  assign \new_[5871]_  = A234 & A232;
  assign \new_[5875]_  = A269 & ~A266;
  assign \new_[5876]_  = A265 & \new_[5875]_ ;
  assign \new_[5877]_  = \new_[5876]_  & \new_[5871]_ ;
  assign \new_[5880]_  = ~A201 & A169;
  assign \new_[5883]_  = ~A203 & ~A202;
  assign \new_[5884]_  = \new_[5883]_  & \new_[5880]_ ;
  assign \new_[5887]_  = A234 & A233;
  assign \new_[5891]_  = A302 & ~A299;
  assign \new_[5892]_  = A298 & \new_[5891]_ ;
  assign \new_[5893]_  = \new_[5892]_  & \new_[5887]_ ;
  assign \new_[5896]_  = ~A201 & A169;
  assign \new_[5899]_  = ~A203 & ~A202;
  assign \new_[5900]_  = \new_[5899]_  & \new_[5896]_ ;
  assign \new_[5903]_  = A234 & A233;
  assign \new_[5907]_  = A302 & A299;
  assign \new_[5908]_  = ~A298 & \new_[5907]_ ;
  assign \new_[5909]_  = \new_[5908]_  & \new_[5903]_ ;
  assign \new_[5912]_  = ~A201 & A169;
  assign \new_[5915]_  = ~A203 & ~A202;
  assign \new_[5916]_  = \new_[5915]_  & \new_[5912]_ ;
  assign \new_[5919]_  = A234 & A233;
  assign \new_[5923]_  = A269 & A266;
  assign \new_[5924]_  = ~A265 & \new_[5923]_ ;
  assign \new_[5925]_  = \new_[5924]_  & \new_[5919]_ ;
  assign \new_[5928]_  = ~A201 & A169;
  assign \new_[5931]_  = ~A203 & ~A202;
  assign \new_[5932]_  = \new_[5931]_  & \new_[5928]_ ;
  assign \new_[5935]_  = A234 & A233;
  assign \new_[5939]_  = A269 & ~A266;
  assign \new_[5940]_  = A265 & \new_[5939]_ ;
  assign \new_[5941]_  = \new_[5940]_  & \new_[5935]_ ;
  assign \new_[5944]_  = ~A201 & A169;
  assign \new_[5947]_  = ~A203 & ~A202;
  assign \new_[5948]_  = \new_[5947]_  & \new_[5944]_ ;
  assign \new_[5951]_  = A233 & ~A232;
  assign \new_[5955]_  = A300 & A299;
  assign \new_[5956]_  = A236 & \new_[5955]_ ;
  assign \new_[5957]_  = \new_[5956]_  & \new_[5951]_ ;
  assign \new_[5960]_  = ~A201 & A169;
  assign \new_[5963]_  = ~A203 & ~A202;
  assign \new_[5964]_  = \new_[5963]_  & \new_[5960]_ ;
  assign \new_[5967]_  = A233 & ~A232;
  assign \new_[5971]_  = A300 & A298;
  assign \new_[5972]_  = A236 & \new_[5971]_ ;
  assign \new_[5973]_  = \new_[5972]_  & \new_[5967]_ ;
  assign \new_[5976]_  = ~A201 & A169;
  assign \new_[5979]_  = ~A203 & ~A202;
  assign \new_[5980]_  = \new_[5979]_  & \new_[5976]_ ;
  assign \new_[5983]_  = A233 & ~A232;
  assign \new_[5987]_  = A267 & A265;
  assign \new_[5988]_  = A236 & \new_[5987]_ ;
  assign \new_[5989]_  = \new_[5988]_  & \new_[5983]_ ;
  assign \new_[5992]_  = ~A201 & A169;
  assign \new_[5995]_  = ~A203 & ~A202;
  assign \new_[5996]_  = \new_[5995]_  & \new_[5992]_ ;
  assign \new_[5999]_  = A233 & ~A232;
  assign \new_[6003]_  = A267 & A266;
  assign \new_[6004]_  = A236 & \new_[6003]_ ;
  assign \new_[6005]_  = \new_[6004]_  & \new_[5999]_ ;
  assign \new_[6008]_  = ~A201 & A169;
  assign \new_[6011]_  = ~A203 & ~A202;
  assign \new_[6012]_  = \new_[6011]_  & \new_[6008]_ ;
  assign \new_[6015]_  = ~A233 & A232;
  assign \new_[6019]_  = A300 & A299;
  assign \new_[6020]_  = A236 & \new_[6019]_ ;
  assign \new_[6021]_  = \new_[6020]_  & \new_[6015]_ ;
  assign \new_[6024]_  = ~A201 & A169;
  assign \new_[6027]_  = ~A203 & ~A202;
  assign \new_[6028]_  = \new_[6027]_  & \new_[6024]_ ;
  assign \new_[6031]_  = ~A233 & A232;
  assign \new_[6035]_  = A300 & A298;
  assign \new_[6036]_  = A236 & \new_[6035]_ ;
  assign \new_[6037]_  = \new_[6036]_  & \new_[6031]_ ;
  assign \new_[6040]_  = ~A201 & A169;
  assign \new_[6043]_  = ~A203 & ~A202;
  assign \new_[6044]_  = \new_[6043]_  & \new_[6040]_ ;
  assign \new_[6047]_  = ~A233 & A232;
  assign \new_[6051]_  = A267 & A265;
  assign \new_[6052]_  = A236 & \new_[6051]_ ;
  assign \new_[6053]_  = \new_[6052]_  & \new_[6047]_ ;
  assign \new_[6056]_  = ~A201 & A169;
  assign \new_[6059]_  = ~A203 & ~A202;
  assign \new_[6060]_  = \new_[6059]_  & \new_[6056]_ ;
  assign \new_[6063]_  = ~A233 & A232;
  assign \new_[6067]_  = A267 & A266;
  assign \new_[6068]_  = A236 & \new_[6067]_ ;
  assign \new_[6069]_  = \new_[6068]_  & \new_[6063]_ ;
  assign \new_[6072]_  = A199 & A169;
  assign \new_[6075]_  = ~A201 & A200;
  assign \new_[6076]_  = \new_[6075]_  & \new_[6072]_ ;
  assign \new_[6079]_  = A235 & ~A202;
  assign \new_[6083]_  = A302 & ~A299;
  assign \new_[6084]_  = A298 & \new_[6083]_ ;
  assign \new_[6085]_  = \new_[6084]_  & \new_[6079]_ ;
  assign \new_[6088]_  = A199 & A169;
  assign \new_[6091]_  = ~A201 & A200;
  assign \new_[6092]_  = \new_[6091]_  & \new_[6088]_ ;
  assign \new_[6095]_  = A235 & ~A202;
  assign \new_[6099]_  = A302 & A299;
  assign \new_[6100]_  = ~A298 & \new_[6099]_ ;
  assign \new_[6101]_  = \new_[6100]_  & \new_[6095]_ ;
  assign \new_[6104]_  = A199 & A169;
  assign \new_[6107]_  = ~A201 & A200;
  assign \new_[6108]_  = \new_[6107]_  & \new_[6104]_ ;
  assign \new_[6111]_  = A235 & ~A202;
  assign \new_[6115]_  = A269 & A266;
  assign \new_[6116]_  = ~A265 & \new_[6115]_ ;
  assign \new_[6117]_  = \new_[6116]_  & \new_[6111]_ ;
  assign \new_[6120]_  = A199 & A169;
  assign \new_[6123]_  = ~A201 & A200;
  assign \new_[6124]_  = \new_[6123]_  & \new_[6120]_ ;
  assign \new_[6127]_  = A235 & ~A202;
  assign \new_[6131]_  = A269 & ~A266;
  assign \new_[6132]_  = A265 & \new_[6131]_ ;
  assign \new_[6133]_  = \new_[6132]_  & \new_[6127]_ ;
  assign \new_[6136]_  = A199 & A169;
  assign \new_[6139]_  = ~A201 & A200;
  assign \new_[6140]_  = \new_[6139]_  & \new_[6136]_ ;
  assign \new_[6143]_  = A232 & ~A202;
  assign \new_[6147]_  = A300 & A299;
  assign \new_[6148]_  = A234 & \new_[6147]_ ;
  assign \new_[6149]_  = \new_[6148]_  & \new_[6143]_ ;
  assign \new_[6152]_  = A199 & A169;
  assign \new_[6155]_  = ~A201 & A200;
  assign \new_[6156]_  = \new_[6155]_  & \new_[6152]_ ;
  assign \new_[6159]_  = A232 & ~A202;
  assign \new_[6163]_  = A300 & A298;
  assign \new_[6164]_  = A234 & \new_[6163]_ ;
  assign \new_[6165]_  = \new_[6164]_  & \new_[6159]_ ;
  assign \new_[6168]_  = A199 & A169;
  assign \new_[6171]_  = ~A201 & A200;
  assign \new_[6172]_  = \new_[6171]_  & \new_[6168]_ ;
  assign \new_[6175]_  = A232 & ~A202;
  assign \new_[6179]_  = A267 & A265;
  assign \new_[6180]_  = A234 & \new_[6179]_ ;
  assign \new_[6181]_  = \new_[6180]_  & \new_[6175]_ ;
  assign \new_[6184]_  = A199 & A169;
  assign \new_[6187]_  = ~A201 & A200;
  assign \new_[6188]_  = \new_[6187]_  & \new_[6184]_ ;
  assign \new_[6191]_  = A232 & ~A202;
  assign \new_[6195]_  = A267 & A266;
  assign \new_[6196]_  = A234 & \new_[6195]_ ;
  assign \new_[6197]_  = \new_[6196]_  & \new_[6191]_ ;
  assign \new_[6200]_  = A199 & A169;
  assign \new_[6203]_  = ~A201 & A200;
  assign \new_[6204]_  = \new_[6203]_  & \new_[6200]_ ;
  assign \new_[6207]_  = A233 & ~A202;
  assign \new_[6211]_  = A300 & A299;
  assign \new_[6212]_  = A234 & \new_[6211]_ ;
  assign \new_[6213]_  = \new_[6212]_  & \new_[6207]_ ;
  assign \new_[6216]_  = A199 & A169;
  assign \new_[6219]_  = ~A201 & A200;
  assign \new_[6220]_  = \new_[6219]_  & \new_[6216]_ ;
  assign \new_[6223]_  = A233 & ~A202;
  assign \new_[6227]_  = A300 & A298;
  assign \new_[6228]_  = A234 & \new_[6227]_ ;
  assign \new_[6229]_  = \new_[6228]_  & \new_[6223]_ ;
  assign \new_[6232]_  = A199 & A169;
  assign \new_[6235]_  = ~A201 & A200;
  assign \new_[6236]_  = \new_[6235]_  & \new_[6232]_ ;
  assign \new_[6239]_  = A233 & ~A202;
  assign \new_[6243]_  = A267 & A265;
  assign \new_[6244]_  = A234 & \new_[6243]_ ;
  assign \new_[6245]_  = \new_[6244]_  & \new_[6239]_ ;
  assign \new_[6248]_  = A199 & A169;
  assign \new_[6251]_  = ~A201 & A200;
  assign \new_[6252]_  = \new_[6251]_  & \new_[6248]_ ;
  assign \new_[6255]_  = A233 & ~A202;
  assign \new_[6259]_  = A267 & A266;
  assign \new_[6260]_  = A234 & \new_[6259]_ ;
  assign \new_[6261]_  = \new_[6260]_  & \new_[6255]_ ;
  assign \new_[6264]_  = A199 & A169;
  assign \new_[6267]_  = ~A201 & A200;
  assign \new_[6268]_  = \new_[6267]_  & \new_[6264]_ ;
  assign \new_[6271]_  = ~A232 & ~A202;
  assign \new_[6275]_  = A301 & A236;
  assign \new_[6276]_  = A233 & \new_[6275]_ ;
  assign \new_[6277]_  = \new_[6276]_  & \new_[6271]_ ;
  assign \new_[6280]_  = A199 & A169;
  assign \new_[6283]_  = ~A201 & A200;
  assign \new_[6284]_  = \new_[6283]_  & \new_[6280]_ ;
  assign \new_[6287]_  = ~A232 & ~A202;
  assign \new_[6291]_  = A268 & A236;
  assign \new_[6292]_  = A233 & \new_[6291]_ ;
  assign \new_[6293]_  = \new_[6292]_  & \new_[6287]_ ;
  assign \new_[6296]_  = A199 & A169;
  assign \new_[6299]_  = ~A201 & A200;
  assign \new_[6300]_  = \new_[6299]_  & \new_[6296]_ ;
  assign \new_[6303]_  = A232 & ~A202;
  assign \new_[6307]_  = A301 & A236;
  assign \new_[6308]_  = ~A233 & \new_[6307]_ ;
  assign \new_[6309]_  = \new_[6308]_  & \new_[6303]_ ;
  assign \new_[6312]_  = A199 & A169;
  assign \new_[6315]_  = ~A201 & A200;
  assign \new_[6316]_  = \new_[6315]_  & \new_[6312]_ ;
  assign \new_[6319]_  = A232 & ~A202;
  assign \new_[6323]_  = A268 & A236;
  assign \new_[6324]_  = ~A233 & \new_[6323]_ ;
  assign \new_[6325]_  = \new_[6324]_  & \new_[6319]_ ;
  assign \new_[6328]_  = ~A199 & A169;
  assign \new_[6331]_  = ~A202 & ~A200;
  assign \new_[6332]_  = \new_[6331]_  & \new_[6328]_ ;
  assign \new_[6335]_  = A234 & A232;
  assign \new_[6339]_  = A302 & ~A299;
  assign \new_[6340]_  = A298 & \new_[6339]_ ;
  assign \new_[6341]_  = \new_[6340]_  & \new_[6335]_ ;
  assign \new_[6344]_  = ~A199 & A169;
  assign \new_[6347]_  = ~A202 & ~A200;
  assign \new_[6348]_  = \new_[6347]_  & \new_[6344]_ ;
  assign \new_[6351]_  = A234 & A232;
  assign \new_[6355]_  = A302 & A299;
  assign \new_[6356]_  = ~A298 & \new_[6355]_ ;
  assign \new_[6357]_  = \new_[6356]_  & \new_[6351]_ ;
  assign \new_[6360]_  = ~A199 & A169;
  assign \new_[6363]_  = ~A202 & ~A200;
  assign \new_[6364]_  = \new_[6363]_  & \new_[6360]_ ;
  assign \new_[6367]_  = A234 & A232;
  assign \new_[6371]_  = A269 & A266;
  assign \new_[6372]_  = ~A265 & \new_[6371]_ ;
  assign \new_[6373]_  = \new_[6372]_  & \new_[6367]_ ;
  assign \new_[6376]_  = ~A199 & A169;
  assign \new_[6379]_  = ~A202 & ~A200;
  assign \new_[6380]_  = \new_[6379]_  & \new_[6376]_ ;
  assign \new_[6383]_  = A234 & A232;
  assign \new_[6387]_  = A269 & ~A266;
  assign \new_[6388]_  = A265 & \new_[6387]_ ;
  assign \new_[6389]_  = \new_[6388]_  & \new_[6383]_ ;
  assign \new_[6392]_  = ~A199 & A169;
  assign \new_[6395]_  = ~A202 & ~A200;
  assign \new_[6396]_  = \new_[6395]_  & \new_[6392]_ ;
  assign \new_[6399]_  = A234 & A233;
  assign \new_[6403]_  = A302 & ~A299;
  assign \new_[6404]_  = A298 & \new_[6403]_ ;
  assign \new_[6405]_  = \new_[6404]_  & \new_[6399]_ ;
  assign \new_[6408]_  = ~A199 & A169;
  assign \new_[6411]_  = ~A202 & ~A200;
  assign \new_[6412]_  = \new_[6411]_  & \new_[6408]_ ;
  assign \new_[6415]_  = A234 & A233;
  assign \new_[6419]_  = A302 & A299;
  assign \new_[6420]_  = ~A298 & \new_[6419]_ ;
  assign \new_[6421]_  = \new_[6420]_  & \new_[6415]_ ;
  assign \new_[6424]_  = ~A199 & A169;
  assign \new_[6427]_  = ~A202 & ~A200;
  assign \new_[6428]_  = \new_[6427]_  & \new_[6424]_ ;
  assign \new_[6431]_  = A234 & A233;
  assign \new_[6435]_  = A269 & A266;
  assign \new_[6436]_  = ~A265 & \new_[6435]_ ;
  assign \new_[6437]_  = \new_[6436]_  & \new_[6431]_ ;
  assign \new_[6440]_  = ~A199 & A169;
  assign \new_[6443]_  = ~A202 & ~A200;
  assign \new_[6444]_  = \new_[6443]_  & \new_[6440]_ ;
  assign \new_[6447]_  = A234 & A233;
  assign \new_[6451]_  = A269 & ~A266;
  assign \new_[6452]_  = A265 & \new_[6451]_ ;
  assign \new_[6453]_  = \new_[6452]_  & \new_[6447]_ ;
  assign \new_[6456]_  = ~A199 & A169;
  assign \new_[6459]_  = ~A202 & ~A200;
  assign \new_[6460]_  = \new_[6459]_  & \new_[6456]_ ;
  assign \new_[6463]_  = A233 & ~A232;
  assign \new_[6467]_  = A300 & A299;
  assign \new_[6468]_  = A236 & \new_[6467]_ ;
  assign \new_[6469]_  = \new_[6468]_  & \new_[6463]_ ;
  assign \new_[6472]_  = ~A199 & A169;
  assign \new_[6475]_  = ~A202 & ~A200;
  assign \new_[6476]_  = \new_[6475]_  & \new_[6472]_ ;
  assign \new_[6479]_  = A233 & ~A232;
  assign \new_[6483]_  = A300 & A298;
  assign \new_[6484]_  = A236 & \new_[6483]_ ;
  assign \new_[6485]_  = \new_[6484]_  & \new_[6479]_ ;
  assign \new_[6488]_  = ~A199 & A169;
  assign \new_[6491]_  = ~A202 & ~A200;
  assign \new_[6492]_  = \new_[6491]_  & \new_[6488]_ ;
  assign \new_[6495]_  = A233 & ~A232;
  assign \new_[6499]_  = A267 & A265;
  assign \new_[6500]_  = A236 & \new_[6499]_ ;
  assign \new_[6501]_  = \new_[6500]_  & \new_[6495]_ ;
  assign \new_[6504]_  = ~A199 & A169;
  assign \new_[6507]_  = ~A202 & ~A200;
  assign \new_[6508]_  = \new_[6507]_  & \new_[6504]_ ;
  assign \new_[6511]_  = A233 & ~A232;
  assign \new_[6515]_  = A267 & A266;
  assign \new_[6516]_  = A236 & \new_[6515]_ ;
  assign \new_[6517]_  = \new_[6516]_  & \new_[6511]_ ;
  assign \new_[6520]_  = ~A199 & A169;
  assign \new_[6523]_  = ~A202 & ~A200;
  assign \new_[6524]_  = \new_[6523]_  & \new_[6520]_ ;
  assign \new_[6527]_  = ~A233 & A232;
  assign \new_[6531]_  = A300 & A299;
  assign \new_[6532]_  = A236 & \new_[6531]_ ;
  assign \new_[6533]_  = \new_[6532]_  & \new_[6527]_ ;
  assign \new_[6536]_  = ~A199 & A169;
  assign \new_[6539]_  = ~A202 & ~A200;
  assign \new_[6540]_  = \new_[6539]_  & \new_[6536]_ ;
  assign \new_[6543]_  = ~A233 & A232;
  assign \new_[6547]_  = A300 & A298;
  assign \new_[6548]_  = A236 & \new_[6547]_ ;
  assign \new_[6549]_  = \new_[6548]_  & \new_[6543]_ ;
  assign \new_[6552]_  = ~A199 & A169;
  assign \new_[6555]_  = ~A202 & ~A200;
  assign \new_[6556]_  = \new_[6555]_  & \new_[6552]_ ;
  assign \new_[6559]_  = ~A233 & A232;
  assign \new_[6563]_  = A267 & A265;
  assign \new_[6564]_  = A236 & \new_[6563]_ ;
  assign \new_[6565]_  = \new_[6564]_  & \new_[6559]_ ;
  assign \new_[6568]_  = ~A199 & A169;
  assign \new_[6571]_  = ~A202 & ~A200;
  assign \new_[6572]_  = \new_[6571]_  & \new_[6568]_ ;
  assign \new_[6575]_  = ~A233 & A232;
  assign \new_[6579]_  = A267 & A266;
  assign \new_[6580]_  = A236 & \new_[6579]_ ;
  assign \new_[6581]_  = \new_[6580]_  & \new_[6575]_ ;
  assign \new_[6584]_  = A166 & A168;
  assign \new_[6588]_  = ~A203 & ~A202;
  assign \new_[6589]_  = ~A201 & \new_[6588]_ ;
  assign \new_[6590]_  = \new_[6589]_  & \new_[6584]_ ;
  assign \new_[6593]_  = A234 & A232;
  assign \new_[6597]_  = A302 & ~A299;
  assign \new_[6598]_  = A298 & \new_[6597]_ ;
  assign \new_[6599]_  = \new_[6598]_  & \new_[6593]_ ;
  assign \new_[6602]_  = A166 & A168;
  assign \new_[6606]_  = ~A203 & ~A202;
  assign \new_[6607]_  = ~A201 & \new_[6606]_ ;
  assign \new_[6608]_  = \new_[6607]_  & \new_[6602]_ ;
  assign \new_[6611]_  = A234 & A232;
  assign \new_[6615]_  = A302 & A299;
  assign \new_[6616]_  = ~A298 & \new_[6615]_ ;
  assign \new_[6617]_  = \new_[6616]_  & \new_[6611]_ ;
  assign \new_[6620]_  = A166 & A168;
  assign \new_[6624]_  = ~A203 & ~A202;
  assign \new_[6625]_  = ~A201 & \new_[6624]_ ;
  assign \new_[6626]_  = \new_[6625]_  & \new_[6620]_ ;
  assign \new_[6629]_  = A234 & A232;
  assign \new_[6633]_  = A269 & A266;
  assign \new_[6634]_  = ~A265 & \new_[6633]_ ;
  assign \new_[6635]_  = \new_[6634]_  & \new_[6629]_ ;
  assign \new_[6638]_  = A166 & A168;
  assign \new_[6642]_  = ~A203 & ~A202;
  assign \new_[6643]_  = ~A201 & \new_[6642]_ ;
  assign \new_[6644]_  = \new_[6643]_  & \new_[6638]_ ;
  assign \new_[6647]_  = A234 & A232;
  assign \new_[6651]_  = A269 & ~A266;
  assign \new_[6652]_  = A265 & \new_[6651]_ ;
  assign \new_[6653]_  = \new_[6652]_  & \new_[6647]_ ;
  assign \new_[6656]_  = A166 & A168;
  assign \new_[6660]_  = ~A203 & ~A202;
  assign \new_[6661]_  = ~A201 & \new_[6660]_ ;
  assign \new_[6662]_  = \new_[6661]_  & \new_[6656]_ ;
  assign \new_[6665]_  = A234 & A233;
  assign \new_[6669]_  = A302 & ~A299;
  assign \new_[6670]_  = A298 & \new_[6669]_ ;
  assign \new_[6671]_  = \new_[6670]_  & \new_[6665]_ ;
  assign \new_[6674]_  = A166 & A168;
  assign \new_[6678]_  = ~A203 & ~A202;
  assign \new_[6679]_  = ~A201 & \new_[6678]_ ;
  assign \new_[6680]_  = \new_[6679]_  & \new_[6674]_ ;
  assign \new_[6683]_  = A234 & A233;
  assign \new_[6687]_  = A302 & A299;
  assign \new_[6688]_  = ~A298 & \new_[6687]_ ;
  assign \new_[6689]_  = \new_[6688]_  & \new_[6683]_ ;
  assign \new_[6692]_  = A166 & A168;
  assign \new_[6696]_  = ~A203 & ~A202;
  assign \new_[6697]_  = ~A201 & \new_[6696]_ ;
  assign \new_[6698]_  = \new_[6697]_  & \new_[6692]_ ;
  assign \new_[6701]_  = A234 & A233;
  assign \new_[6705]_  = A269 & A266;
  assign \new_[6706]_  = ~A265 & \new_[6705]_ ;
  assign \new_[6707]_  = \new_[6706]_  & \new_[6701]_ ;
  assign \new_[6710]_  = A166 & A168;
  assign \new_[6714]_  = ~A203 & ~A202;
  assign \new_[6715]_  = ~A201 & \new_[6714]_ ;
  assign \new_[6716]_  = \new_[6715]_  & \new_[6710]_ ;
  assign \new_[6719]_  = A234 & A233;
  assign \new_[6723]_  = A269 & ~A266;
  assign \new_[6724]_  = A265 & \new_[6723]_ ;
  assign \new_[6725]_  = \new_[6724]_  & \new_[6719]_ ;
  assign \new_[6728]_  = A166 & A168;
  assign \new_[6732]_  = ~A203 & ~A202;
  assign \new_[6733]_  = ~A201 & \new_[6732]_ ;
  assign \new_[6734]_  = \new_[6733]_  & \new_[6728]_ ;
  assign \new_[6737]_  = A233 & ~A232;
  assign \new_[6741]_  = A300 & A299;
  assign \new_[6742]_  = A236 & \new_[6741]_ ;
  assign \new_[6743]_  = \new_[6742]_  & \new_[6737]_ ;
  assign \new_[6746]_  = A166 & A168;
  assign \new_[6750]_  = ~A203 & ~A202;
  assign \new_[6751]_  = ~A201 & \new_[6750]_ ;
  assign \new_[6752]_  = \new_[6751]_  & \new_[6746]_ ;
  assign \new_[6755]_  = A233 & ~A232;
  assign \new_[6759]_  = A300 & A298;
  assign \new_[6760]_  = A236 & \new_[6759]_ ;
  assign \new_[6761]_  = \new_[6760]_  & \new_[6755]_ ;
  assign \new_[6764]_  = A166 & A168;
  assign \new_[6768]_  = ~A203 & ~A202;
  assign \new_[6769]_  = ~A201 & \new_[6768]_ ;
  assign \new_[6770]_  = \new_[6769]_  & \new_[6764]_ ;
  assign \new_[6773]_  = A233 & ~A232;
  assign \new_[6777]_  = A267 & A265;
  assign \new_[6778]_  = A236 & \new_[6777]_ ;
  assign \new_[6779]_  = \new_[6778]_  & \new_[6773]_ ;
  assign \new_[6782]_  = A166 & A168;
  assign \new_[6786]_  = ~A203 & ~A202;
  assign \new_[6787]_  = ~A201 & \new_[6786]_ ;
  assign \new_[6788]_  = \new_[6787]_  & \new_[6782]_ ;
  assign \new_[6791]_  = A233 & ~A232;
  assign \new_[6795]_  = A267 & A266;
  assign \new_[6796]_  = A236 & \new_[6795]_ ;
  assign \new_[6797]_  = \new_[6796]_  & \new_[6791]_ ;
  assign \new_[6800]_  = A166 & A168;
  assign \new_[6804]_  = ~A203 & ~A202;
  assign \new_[6805]_  = ~A201 & \new_[6804]_ ;
  assign \new_[6806]_  = \new_[6805]_  & \new_[6800]_ ;
  assign \new_[6809]_  = ~A233 & A232;
  assign \new_[6813]_  = A300 & A299;
  assign \new_[6814]_  = A236 & \new_[6813]_ ;
  assign \new_[6815]_  = \new_[6814]_  & \new_[6809]_ ;
  assign \new_[6818]_  = A166 & A168;
  assign \new_[6822]_  = ~A203 & ~A202;
  assign \new_[6823]_  = ~A201 & \new_[6822]_ ;
  assign \new_[6824]_  = \new_[6823]_  & \new_[6818]_ ;
  assign \new_[6827]_  = ~A233 & A232;
  assign \new_[6831]_  = A300 & A298;
  assign \new_[6832]_  = A236 & \new_[6831]_ ;
  assign \new_[6833]_  = \new_[6832]_  & \new_[6827]_ ;
  assign \new_[6836]_  = A166 & A168;
  assign \new_[6840]_  = ~A203 & ~A202;
  assign \new_[6841]_  = ~A201 & \new_[6840]_ ;
  assign \new_[6842]_  = \new_[6841]_  & \new_[6836]_ ;
  assign \new_[6845]_  = ~A233 & A232;
  assign \new_[6849]_  = A267 & A265;
  assign \new_[6850]_  = A236 & \new_[6849]_ ;
  assign \new_[6851]_  = \new_[6850]_  & \new_[6845]_ ;
  assign \new_[6854]_  = A166 & A168;
  assign \new_[6858]_  = ~A203 & ~A202;
  assign \new_[6859]_  = ~A201 & \new_[6858]_ ;
  assign \new_[6860]_  = \new_[6859]_  & \new_[6854]_ ;
  assign \new_[6863]_  = ~A233 & A232;
  assign \new_[6867]_  = A267 & A266;
  assign \new_[6868]_  = A236 & \new_[6867]_ ;
  assign \new_[6869]_  = \new_[6868]_  & \new_[6863]_ ;
  assign \new_[6872]_  = A166 & A168;
  assign \new_[6876]_  = ~A201 & A200;
  assign \new_[6877]_  = A199 & \new_[6876]_ ;
  assign \new_[6878]_  = \new_[6877]_  & \new_[6872]_ ;
  assign \new_[6881]_  = A235 & ~A202;
  assign \new_[6885]_  = A302 & ~A299;
  assign \new_[6886]_  = A298 & \new_[6885]_ ;
  assign \new_[6887]_  = \new_[6886]_  & \new_[6881]_ ;
  assign \new_[6890]_  = A166 & A168;
  assign \new_[6894]_  = ~A201 & A200;
  assign \new_[6895]_  = A199 & \new_[6894]_ ;
  assign \new_[6896]_  = \new_[6895]_  & \new_[6890]_ ;
  assign \new_[6899]_  = A235 & ~A202;
  assign \new_[6903]_  = A302 & A299;
  assign \new_[6904]_  = ~A298 & \new_[6903]_ ;
  assign \new_[6905]_  = \new_[6904]_  & \new_[6899]_ ;
  assign \new_[6908]_  = A166 & A168;
  assign \new_[6912]_  = ~A201 & A200;
  assign \new_[6913]_  = A199 & \new_[6912]_ ;
  assign \new_[6914]_  = \new_[6913]_  & \new_[6908]_ ;
  assign \new_[6917]_  = A235 & ~A202;
  assign \new_[6921]_  = A269 & A266;
  assign \new_[6922]_  = ~A265 & \new_[6921]_ ;
  assign \new_[6923]_  = \new_[6922]_  & \new_[6917]_ ;
  assign \new_[6926]_  = A166 & A168;
  assign \new_[6930]_  = ~A201 & A200;
  assign \new_[6931]_  = A199 & \new_[6930]_ ;
  assign \new_[6932]_  = \new_[6931]_  & \new_[6926]_ ;
  assign \new_[6935]_  = A235 & ~A202;
  assign \new_[6939]_  = A269 & ~A266;
  assign \new_[6940]_  = A265 & \new_[6939]_ ;
  assign \new_[6941]_  = \new_[6940]_  & \new_[6935]_ ;
  assign \new_[6944]_  = A166 & A168;
  assign \new_[6948]_  = ~A201 & A200;
  assign \new_[6949]_  = A199 & \new_[6948]_ ;
  assign \new_[6950]_  = \new_[6949]_  & \new_[6944]_ ;
  assign \new_[6953]_  = A232 & ~A202;
  assign \new_[6957]_  = A300 & A299;
  assign \new_[6958]_  = A234 & \new_[6957]_ ;
  assign \new_[6959]_  = \new_[6958]_  & \new_[6953]_ ;
  assign \new_[6962]_  = A166 & A168;
  assign \new_[6966]_  = ~A201 & A200;
  assign \new_[6967]_  = A199 & \new_[6966]_ ;
  assign \new_[6968]_  = \new_[6967]_  & \new_[6962]_ ;
  assign \new_[6971]_  = A232 & ~A202;
  assign \new_[6975]_  = A300 & A298;
  assign \new_[6976]_  = A234 & \new_[6975]_ ;
  assign \new_[6977]_  = \new_[6976]_  & \new_[6971]_ ;
  assign \new_[6980]_  = A166 & A168;
  assign \new_[6984]_  = ~A201 & A200;
  assign \new_[6985]_  = A199 & \new_[6984]_ ;
  assign \new_[6986]_  = \new_[6985]_  & \new_[6980]_ ;
  assign \new_[6989]_  = A232 & ~A202;
  assign \new_[6993]_  = A267 & A265;
  assign \new_[6994]_  = A234 & \new_[6993]_ ;
  assign \new_[6995]_  = \new_[6994]_  & \new_[6989]_ ;
  assign \new_[6998]_  = A166 & A168;
  assign \new_[7002]_  = ~A201 & A200;
  assign \new_[7003]_  = A199 & \new_[7002]_ ;
  assign \new_[7004]_  = \new_[7003]_  & \new_[6998]_ ;
  assign \new_[7007]_  = A232 & ~A202;
  assign \new_[7011]_  = A267 & A266;
  assign \new_[7012]_  = A234 & \new_[7011]_ ;
  assign \new_[7013]_  = \new_[7012]_  & \new_[7007]_ ;
  assign \new_[7016]_  = A166 & A168;
  assign \new_[7020]_  = ~A201 & A200;
  assign \new_[7021]_  = A199 & \new_[7020]_ ;
  assign \new_[7022]_  = \new_[7021]_  & \new_[7016]_ ;
  assign \new_[7025]_  = A233 & ~A202;
  assign \new_[7029]_  = A300 & A299;
  assign \new_[7030]_  = A234 & \new_[7029]_ ;
  assign \new_[7031]_  = \new_[7030]_  & \new_[7025]_ ;
  assign \new_[7034]_  = A166 & A168;
  assign \new_[7038]_  = ~A201 & A200;
  assign \new_[7039]_  = A199 & \new_[7038]_ ;
  assign \new_[7040]_  = \new_[7039]_  & \new_[7034]_ ;
  assign \new_[7043]_  = A233 & ~A202;
  assign \new_[7047]_  = A300 & A298;
  assign \new_[7048]_  = A234 & \new_[7047]_ ;
  assign \new_[7049]_  = \new_[7048]_  & \new_[7043]_ ;
  assign \new_[7052]_  = A166 & A168;
  assign \new_[7056]_  = ~A201 & A200;
  assign \new_[7057]_  = A199 & \new_[7056]_ ;
  assign \new_[7058]_  = \new_[7057]_  & \new_[7052]_ ;
  assign \new_[7061]_  = A233 & ~A202;
  assign \new_[7065]_  = A267 & A265;
  assign \new_[7066]_  = A234 & \new_[7065]_ ;
  assign \new_[7067]_  = \new_[7066]_  & \new_[7061]_ ;
  assign \new_[7070]_  = A166 & A168;
  assign \new_[7074]_  = ~A201 & A200;
  assign \new_[7075]_  = A199 & \new_[7074]_ ;
  assign \new_[7076]_  = \new_[7075]_  & \new_[7070]_ ;
  assign \new_[7079]_  = A233 & ~A202;
  assign \new_[7083]_  = A267 & A266;
  assign \new_[7084]_  = A234 & \new_[7083]_ ;
  assign \new_[7085]_  = \new_[7084]_  & \new_[7079]_ ;
  assign \new_[7088]_  = A166 & A168;
  assign \new_[7092]_  = ~A201 & A200;
  assign \new_[7093]_  = A199 & \new_[7092]_ ;
  assign \new_[7094]_  = \new_[7093]_  & \new_[7088]_ ;
  assign \new_[7097]_  = ~A232 & ~A202;
  assign \new_[7101]_  = A301 & A236;
  assign \new_[7102]_  = A233 & \new_[7101]_ ;
  assign \new_[7103]_  = \new_[7102]_  & \new_[7097]_ ;
  assign \new_[7106]_  = A166 & A168;
  assign \new_[7110]_  = ~A201 & A200;
  assign \new_[7111]_  = A199 & \new_[7110]_ ;
  assign \new_[7112]_  = \new_[7111]_  & \new_[7106]_ ;
  assign \new_[7115]_  = ~A232 & ~A202;
  assign \new_[7119]_  = A268 & A236;
  assign \new_[7120]_  = A233 & \new_[7119]_ ;
  assign \new_[7121]_  = \new_[7120]_  & \new_[7115]_ ;
  assign \new_[7124]_  = A166 & A168;
  assign \new_[7128]_  = ~A201 & A200;
  assign \new_[7129]_  = A199 & \new_[7128]_ ;
  assign \new_[7130]_  = \new_[7129]_  & \new_[7124]_ ;
  assign \new_[7133]_  = A232 & ~A202;
  assign \new_[7137]_  = A301 & A236;
  assign \new_[7138]_  = ~A233 & \new_[7137]_ ;
  assign \new_[7139]_  = \new_[7138]_  & \new_[7133]_ ;
  assign \new_[7142]_  = A166 & A168;
  assign \new_[7146]_  = ~A201 & A200;
  assign \new_[7147]_  = A199 & \new_[7146]_ ;
  assign \new_[7148]_  = \new_[7147]_  & \new_[7142]_ ;
  assign \new_[7151]_  = A232 & ~A202;
  assign \new_[7155]_  = A268 & A236;
  assign \new_[7156]_  = ~A233 & \new_[7155]_ ;
  assign \new_[7157]_  = \new_[7156]_  & \new_[7151]_ ;
  assign \new_[7160]_  = A166 & A168;
  assign \new_[7164]_  = ~A202 & ~A200;
  assign \new_[7165]_  = ~A199 & \new_[7164]_ ;
  assign \new_[7166]_  = \new_[7165]_  & \new_[7160]_ ;
  assign \new_[7169]_  = A234 & A232;
  assign \new_[7173]_  = A302 & ~A299;
  assign \new_[7174]_  = A298 & \new_[7173]_ ;
  assign \new_[7175]_  = \new_[7174]_  & \new_[7169]_ ;
  assign \new_[7178]_  = A166 & A168;
  assign \new_[7182]_  = ~A202 & ~A200;
  assign \new_[7183]_  = ~A199 & \new_[7182]_ ;
  assign \new_[7184]_  = \new_[7183]_  & \new_[7178]_ ;
  assign \new_[7187]_  = A234 & A232;
  assign \new_[7191]_  = A302 & A299;
  assign \new_[7192]_  = ~A298 & \new_[7191]_ ;
  assign \new_[7193]_  = \new_[7192]_  & \new_[7187]_ ;
  assign \new_[7196]_  = A166 & A168;
  assign \new_[7200]_  = ~A202 & ~A200;
  assign \new_[7201]_  = ~A199 & \new_[7200]_ ;
  assign \new_[7202]_  = \new_[7201]_  & \new_[7196]_ ;
  assign \new_[7205]_  = A234 & A232;
  assign \new_[7209]_  = A269 & A266;
  assign \new_[7210]_  = ~A265 & \new_[7209]_ ;
  assign \new_[7211]_  = \new_[7210]_  & \new_[7205]_ ;
  assign \new_[7214]_  = A166 & A168;
  assign \new_[7218]_  = ~A202 & ~A200;
  assign \new_[7219]_  = ~A199 & \new_[7218]_ ;
  assign \new_[7220]_  = \new_[7219]_  & \new_[7214]_ ;
  assign \new_[7223]_  = A234 & A232;
  assign \new_[7227]_  = A269 & ~A266;
  assign \new_[7228]_  = A265 & \new_[7227]_ ;
  assign \new_[7229]_  = \new_[7228]_  & \new_[7223]_ ;
  assign \new_[7232]_  = A166 & A168;
  assign \new_[7236]_  = ~A202 & ~A200;
  assign \new_[7237]_  = ~A199 & \new_[7236]_ ;
  assign \new_[7238]_  = \new_[7237]_  & \new_[7232]_ ;
  assign \new_[7241]_  = A234 & A233;
  assign \new_[7245]_  = A302 & ~A299;
  assign \new_[7246]_  = A298 & \new_[7245]_ ;
  assign \new_[7247]_  = \new_[7246]_  & \new_[7241]_ ;
  assign \new_[7250]_  = A166 & A168;
  assign \new_[7254]_  = ~A202 & ~A200;
  assign \new_[7255]_  = ~A199 & \new_[7254]_ ;
  assign \new_[7256]_  = \new_[7255]_  & \new_[7250]_ ;
  assign \new_[7259]_  = A234 & A233;
  assign \new_[7263]_  = A302 & A299;
  assign \new_[7264]_  = ~A298 & \new_[7263]_ ;
  assign \new_[7265]_  = \new_[7264]_  & \new_[7259]_ ;
  assign \new_[7268]_  = A166 & A168;
  assign \new_[7272]_  = ~A202 & ~A200;
  assign \new_[7273]_  = ~A199 & \new_[7272]_ ;
  assign \new_[7274]_  = \new_[7273]_  & \new_[7268]_ ;
  assign \new_[7277]_  = A234 & A233;
  assign \new_[7281]_  = A269 & A266;
  assign \new_[7282]_  = ~A265 & \new_[7281]_ ;
  assign \new_[7283]_  = \new_[7282]_  & \new_[7277]_ ;
  assign \new_[7286]_  = A166 & A168;
  assign \new_[7290]_  = ~A202 & ~A200;
  assign \new_[7291]_  = ~A199 & \new_[7290]_ ;
  assign \new_[7292]_  = \new_[7291]_  & \new_[7286]_ ;
  assign \new_[7295]_  = A234 & A233;
  assign \new_[7299]_  = A269 & ~A266;
  assign \new_[7300]_  = A265 & \new_[7299]_ ;
  assign \new_[7301]_  = \new_[7300]_  & \new_[7295]_ ;
  assign \new_[7304]_  = A166 & A168;
  assign \new_[7308]_  = ~A202 & ~A200;
  assign \new_[7309]_  = ~A199 & \new_[7308]_ ;
  assign \new_[7310]_  = \new_[7309]_  & \new_[7304]_ ;
  assign \new_[7313]_  = A233 & ~A232;
  assign \new_[7317]_  = A300 & A299;
  assign \new_[7318]_  = A236 & \new_[7317]_ ;
  assign \new_[7319]_  = \new_[7318]_  & \new_[7313]_ ;
  assign \new_[7322]_  = A166 & A168;
  assign \new_[7326]_  = ~A202 & ~A200;
  assign \new_[7327]_  = ~A199 & \new_[7326]_ ;
  assign \new_[7328]_  = \new_[7327]_  & \new_[7322]_ ;
  assign \new_[7331]_  = A233 & ~A232;
  assign \new_[7335]_  = A300 & A298;
  assign \new_[7336]_  = A236 & \new_[7335]_ ;
  assign \new_[7337]_  = \new_[7336]_  & \new_[7331]_ ;
  assign \new_[7340]_  = A166 & A168;
  assign \new_[7344]_  = ~A202 & ~A200;
  assign \new_[7345]_  = ~A199 & \new_[7344]_ ;
  assign \new_[7346]_  = \new_[7345]_  & \new_[7340]_ ;
  assign \new_[7349]_  = A233 & ~A232;
  assign \new_[7353]_  = A267 & A265;
  assign \new_[7354]_  = A236 & \new_[7353]_ ;
  assign \new_[7355]_  = \new_[7354]_  & \new_[7349]_ ;
  assign \new_[7358]_  = A166 & A168;
  assign \new_[7362]_  = ~A202 & ~A200;
  assign \new_[7363]_  = ~A199 & \new_[7362]_ ;
  assign \new_[7364]_  = \new_[7363]_  & \new_[7358]_ ;
  assign \new_[7367]_  = A233 & ~A232;
  assign \new_[7371]_  = A267 & A266;
  assign \new_[7372]_  = A236 & \new_[7371]_ ;
  assign \new_[7373]_  = \new_[7372]_  & \new_[7367]_ ;
  assign \new_[7376]_  = A166 & A168;
  assign \new_[7380]_  = ~A202 & ~A200;
  assign \new_[7381]_  = ~A199 & \new_[7380]_ ;
  assign \new_[7382]_  = \new_[7381]_  & \new_[7376]_ ;
  assign \new_[7385]_  = ~A233 & A232;
  assign \new_[7389]_  = A300 & A299;
  assign \new_[7390]_  = A236 & \new_[7389]_ ;
  assign \new_[7391]_  = \new_[7390]_  & \new_[7385]_ ;
  assign \new_[7394]_  = A166 & A168;
  assign \new_[7398]_  = ~A202 & ~A200;
  assign \new_[7399]_  = ~A199 & \new_[7398]_ ;
  assign \new_[7400]_  = \new_[7399]_  & \new_[7394]_ ;
  assign \new_[7403]_  = ~A233 & A232;
  assign \new_[7407]_  = A300 & A298;
  assign \new_[7408]_  = A236 & \new_[7407]_ ;
  assign \new_[7409]_  = \new_[7408]_  & \new_[7403]_ ;
  assign \new_[7412]_  = A166 & A168;
  assign \new_[7416]_  = ~A202 & ~A200;
  assign \new_[7417]_  = ~A199 & \new_[7416]_ ;
  assign \new_[7418]_  = \new_[7417]_  & \new_[7412]_ ;
  assign \new_[7421]_  = ~A233 & A232;
  assign \new_[7425]_  = A267 & A265;
  assign \new_[7426]_  = A236 & \new_[7425]_ ;
  assign \new_[7427]_  = \new_[7426]_  & \new_[7421]_ ;
  assign \new_[7430]_  = A166 & A168;
  assign \new_[7434]_  = ~A202 & ~A200;
  assign \new_[7435]_  = ~A199 & \new_[7434]_ ;
  assign \new_[7436]_  = \new_[7435]_  & \new_[7430]_ ;
  assign \new_[7439]_  = ~A233 & A232;
  assign \new_[7443]_  = A267 & A266;
  assign \new_[7444]_  = A236 & \new_[7443]_ ;
  assign \new_[7445]_  = \new_[7444]_  & \new_[7439]_ ;
  assign \new_[7448]_  = A167 & A168;
  assign \new_[7452]_  = ~A203 & ~A202;
  assign \new_[7453]_  = ~A201 & \new_[7452]_ ;
  assign \new_[7454]_  = \new_[7453]_  & \new_[7448]_ ;
  assign \new_[7457]_  = A234 & A232;
  assign \new_[7461]_  = A302 & ~A299;
  assign \new_[7462]_  = A298 & \new_[7461]_ ;
  assign \new_[7463]_  = \new_[7462]_  & \new_[7457]_ ;
  assign \new_[7466]_  = A167 & A168;
  assign \new_[7470]_  = ~A203 & ~A202;
  assign \new_[7471]_  = ~A201 & \new_[7470]_ ;
  assign \new_[7472]_  = \new_[7471]_  & \new_[7466]_ ;
  assign \new_[7475]_  = A234 & A232;
  assign \new_[7479]_  = A302 & A299;
  assign \new_[7480]_  = ~A298 & \new_[7479]_ ;
  assign \new_[7481]_  = \new_[7480]_  & \new_[7475]_ ;
  assign \new_[7484]_  = A167 & A168;
  assign \new_[7488]_  = ~A203 & ~A202;
  assign \new_[7489]_  = ~A201 & \new_[7488]_ ;
  assign \new_[7490]_  = \new_[7489]_  & \new_[7484]_ ;
  assign \new_[7493]_  = A234 & A232;
  assign \new_[7497]_  = A269 & A266;
  assign \new_[7498]_  = ~A265 & \new_[7497]_ ;
  assign \new_[7499]_  = \new_[7498]_  & \new_[7493]_ ;
  assign \new_[7502]_  = A167 & A168;
  assign \new_[7506]_  = ~A203 & ~A202;
  assign \new_[7507]_  = ~A201 & \new_[7506]_ ;
  assign \new_[7508]_  = \new_[7507]_  & \new_[7502]_ ;
  assign \new_[7511]_  = A234 & A232;
  assign \new_[7515]_  = A269 & ~A266;
  assign \new_[7516]_  = A265 & \new_[7515]_ ;
  assign \new_[7517]_  = \new_[7516]_  & \new_[7511]_ ;
  assign \new_[7520]_  = A167 & A168;
  assign \new_[7524]_  = ~A203 & ~A202;
  assign \new_[7525]_  = ~A201 & \new_[7524]_ ;
  assign \new_[7526]_  = \new_[7525]_  & \new_[7520]_ ;
  assign \new_[7529]_  = A234 & A233;
  assign \new_[7533]_  = A302 & ~A299;
  assign \new_[7534]_  = A298 & \new_[7533]_ ;
  assign \new_[7535]_  = \new_[7534]_  & \new_[7529]_ ;
  assign \new_[7538]_  = A167 & A168;
  assign \new_[7542]_  = ~A203 & ~A202;
  assign \new_[7543]_  = ~A201 & \new_[7542]_ ;
  assign \new_[7544]_  = \new_[7543]_  & \new_[7538]_ ;
  assign \new_[7547]_  = A234 & A233;
  assign \new_[7551]_  = A302 & A299;
  assign \new_[7552]_  = ~A298 & \new_[7551]_ ;
  assign \new_[7553]_  = \new_[7552]_  & \new_[7547]_ ;
  assign \new_[7556]_  = A167 & A168;
  assign \new_[7560]_  = ~A203 & ~A202;
  assign \new_[7561]_  = ~A201 & \new_[7560]_ ;
  assign \new_[7562]_  = \new_[7561]_  & \new_[7556]_ ;
  assign \new_[7565]_  = A234 & A233;
  assign \new_[7569]_  = A269 & A266;
  assign \new_[7570]_  = ~A265 & \new_[7569]_ ;
  assign \new_[7571]_  = \new_[7570]_  & \new_[7565]_ ;
  assign \new_[7574]_  = A167 & A168;
  assign \new_[7578]_  = ~A203 & ~A202;
  assign \new_[7579]_  = ~A201 & \new_[7578]_ ;
  assign \new_[7580]_  = \new_[7579]_  & \new_[7574]_ ;
  assign \new_[7583]_  = A234 & A233;
  assign \new_[7587]_  = A269 & ~A266;
  assign \new_[7588]_  = A265 & \new_[7587]_ ;
  assign \new_[7589]_  = \new_[7588]_  & \new_[7583]_ ;
  assign \new_[7592]_  = A167 & A168;
  assign \new_[7596]_  = ~A203 & ~A202;
  assign \new_[7597]_  = ~A201 & \new_[7596]_ ;
  assign \new_[7598]_  = \new_[7597]_  & \new_[7592]_ ;
  assign \new_[7601]_  = A233 & ~A232;
  assign \new_[7605]_  = A300 & A299;
  assign \new_[7606]_  = A236 & \new_[7605]_ ;
  assign \new_[7607]_  = \new_[7606]_  & \new_[7601]_ ;
  assign \new_[7610]_  = A167 & A168;
  assign \new_[7614]_  = ~A203 & ~A202;
  assign \new_[7615]_  = ~A201 & \new_[7614]_ ;
  assign \new_[7616]_  = \new_[7615]_  & \new_[7610]_ ;
  assign \new_[7619]_  = A233 & ~A232;
  assign \new_[7623]_  = A300 & A298;
  assign \new_[7624]_  = A236 & \new_[7623]_ ;
  assign \new_[7625]_  = \new_[7624]_  & \new_[7619]_ ;
  assign \new_[7628]_  = A167 & A168;
  assign \new_[7632]_  = ~A203 & ~A202;
  assign \new_[7633]_  = ~A201 & \new_[7632]_ ;
  assign \new_[7634]_  = \new_[7633]_  & \new_[7628]_ ;
  assign \new_[7637]_  = A233 & ~A232;
  assign \new_[7641]_  = A267 & A265;
  assign \new_[7642]_  = A236 & \new_[7641]_ ;
  assign \new_[7643]_  = \new_[7642]_  & \new_[7637]_ ;
  assign \new_[7646]_  = A167 & A168;
  assign \new_[7650]_  = ~A203 & ~A202;
  assign \new_[7651]_  = ~A201 & \new_[7650]_ ;
  assign \new_[7652]_  = \new_[7651]_  & \new_[7646]_ ;
  assign \new_[7655]_  = A233 & ~A232;
  assign \new_[7659]_  = A267 & A266;
  assign \new_[7660]_  = A236 & \new_[7659]_ ;
  assign \new_[7661]_  = \new_[7660]_  & \new_[7655]_ ;
  assign \new_[7664]_  = A167 & A168;
  assign \new_[7668]_  = ~A203 & ~A202;
  assign \new_[7669]_  = ~A201 & \new_[7668]_ ;
  assign \new_[7670]_  = \new_[7669]_  & \new_[7664]_ ;
  assign \new_[7673]_  = ~A233 & A232;
  assign \new_[7677]_  = A300 & A299;
  assign \new_[7678]_  = A236 & \new_[7677]_ ;
  assign \new_[7679]_  = \new_[7678]_  & \new_[7673]_ ;
  assign \new_[7682]_  = A167 & A168;
  assign \new_[7686]_  = ~A203 & ~A202;
  assign \new_[7687]_  = ~A201 & \new_[7686]_ ;
  assign \new_[7688]_  = \new_[7687]_  & \new_[7682]_ ;
  assign \new_[7691]_  = ~A233 & A232;
  assign \new_[7695]_  = A300 & A298;
  assign \new_[7696]_  = A236 & \new_[7695]_ ;
  assign \new_[7697]_  = \new_[7696]_  & \new_[7691]_ ;
  assign \new_[7700]_  = A167 & A168;
  assign \new_[7704]_  = ~A203 & ~A202;
  assign \new_[7705]_  = ~A201 & \new_[7704]_ ;
  assign \new_[7706]_  = \new_[7705]_  & \new_[7700]_ ;
  assign \new_[7709]_  = ~A233 & A232;
  assign \new_[7713]_  = A267 & A265;
  assign \new_[7714]_  = A236 & \new_[7713]_ ;
  assign \new_[7715]_  = \new_[7714]_  & \new_[7709]_ ;
  assign \new_[7718]_  = A167 & A168;
  assign \new_[7722]_  = ~A203 & ~A202;
  assign \new_[7723]_  = ~A201 & \new_[7722]_ ;
  assign \new_[7724]_  = \new_[7723]_  & \new_[7718]_ ;
  assign \new_[7727]_  = ~A233 & A232;
  assign \new_[7731]_  = A267 & A266;
  assign \new_[7732]_  = A236 & \new_[7731]_ ;
  assign \new_[7733]_  = \new_[7732]_  & \new_[7727]_ ;
  assign \new_[7736]_  = A167 & A168;
  assign \new_[7740]_  = ~A201 & A200;
  assign \new_[7741]_  = A199 & \new_[7740]_ ;
  assign \new_[7742]_  = \new_[7741]_  & \new_[7736]_ ;
  assign \new_[7745]_  = A235 & ~A202;
  assign \new_[7749]_  = A302 & ~A299;
  assign \new_[7750]_  = A298 & \new_[7749]_ ;
  assign \new_[7751]_  = \new_[7750]_  & \new_[7745]_ ;
  assign \new_[7754]_  = A167 & A168;
  assign \new_[7758]_  = ~A201 & A200;
  assign \new_[7759]_  = A199 & \new_[7758]_ ;
  assign \new_[7760]_  = \new_[7759]_  & \new_[7754]_ ;
  assign \new_[7763]_  = A235 & ~A202;
  assign \new_[7767]_  = A302 & A299;
  assign \new_[7768]_  = ~A298 & \new_[7767]_ ;
  assign \new_[7769]_  = \new_[7768]_  & \new_[7763]_ ;
  assign \new_[7772]_  = A167 & A168;
  assign \new_[7776]_  = ~A201 & A200;
  assign \new_[7777]_  = A199 & \new_[7776]_ ;
  assign \new_[7778]_  = \new_[7777]_  & \new_[7772]_ ;
  assign \new_[7781]_  = A235 & ~A202;
  assign \new_[7785]_  = A269 & A266;
  assign \new_[7786]_  = ~A265 & \new_[7785]_ ;
  assign \new_[7787]_  = \new_[7786]_  & \new_[7781]_ ;
  assign \new_[7790]_  = A167 & A168;
  assign \new_[7794]_  = ~A201 & A200;
  assign \new_[7795]_  = A199 & \new_[7794]_ ;
  assign \new_[7796]_  = \new_[7795]_  & \new_[7790]_ ;
  assign \new_[7799]_  = A235 & ~A202;
  assign \new_[7803]_  = A269 & ~A266;
  assign \new_[7804]_  = A265 & \new_[7803]_ ;
  assign \new_[7805]_  = \new_[7804]_  & \new_[7799]_ ;
  assign \new_[7808]_  = A167 & A168;
  assign \new_[7812]_  = ~A201 & A200;
  assign \new_[7813]_  = A199 & \new_[7812]_ ;
  assign \new_[7814]_  = \new_[7813]_  & \new_[7808]_ ;
  assign \new_[7817]_  = A232 & ~A202;
  assign \new_[7821]_  = A300 & A299;
  assign \new_[7822]_  = A234 & \new_[7821]_ ;
  assign \new_[7823]_  = \new_[7822]_  & \new_[7817]_ ;
  assign \new_[7826]_  = A167 & A168;
  assign \new_[7830]_  = ~A201 & A200;
  assign \new_[7831]_  = A199 & \new_[7830]_ ;
  assign \new_[7832]_  = \new_[7831]_  & \new_[7826]_ ;
  assign \new_[7835]_  = A232 & ~A202;
  assign \new_[7839]_  = A300 & A298;
  assign \new_[7840]_  = A234 & \new_[7839]_ ;
  assign \new_[7841]_  = \new_[7840]_  & \new_[7835]_ ;
  assign \new_[7844]_  = A167 & A168;
  assign \new_[7848]_  = ~A201 & A200;
  assign \new_[7849]_  = A199 & \new_[7848]_ ;
  assign \new_[7850]_  = \new_[7849]_  & \new_[7844]_ ;
  assign \new_[7853]_  = A232 & ~A202;
  assign \new_[7857]_  = A267 & A265;
  assign \new_[7858]_  = A234 & \new_[7857]_ ;
  assign \new_[7859]_  = \new_[7858]_  & \new_[7853]_ ;
  assign \new_[7862]_  = A167 & A168;
  assign \new_[7866]_  = ~A201 & A200;
  assign \new_[7867]_  = A199 & \new_[7866]_ ;
  assign \new_[7868]_  = \new_[7867]_  & \new_[7862]_ ;
  assign \new_[7871]_  = A232 & ~A202;
  assign \new_[7875]_  = A267 & A266;
  assign \new_[7876]_  = A234 & \new_[7875]_ ;
  assign \new_[7877]_  = \new_[7876]_  & \new_[7871]_ ;
  assign \new_[7880]_  = A167 & A168;
  assign \new_[7884]_  = ~A201 & A200;
  assign \new_[7885]_  = A199 & \new_[7884]_ ;
  assign \new_[7886]_  = \new_[7885]_  & \new_[7880]_ ;
  assign \new_[7889]_  = A233 & ~A202;
  assign \new_[7893]_  = A300 & A299;
  assign \new_[7894]_  = A234 & \new_[7893]_ ;
  assign \new_[7895]_  = \new_[7894]_  & \new_[7889]_ ;
  assign \new_[7898]_  = A167 & A168;
  assign \new_[7902]_  = ~A201 & A200;
  assign \new_[7903]_  = A199 & \new_[7902]_ ;
  assign \new_[7904]_  = \new_[7903]_  & \new_[7898]_ ;
  assign \new_[7907]_  = A233 & ~A202;
  assign \new_[7911]_  = A300 & A298;
  assign \new_[7912]_  = A234 & \new_[7911]_ ;
  assign \new_[7913]_  = \new_[7912]_  & \new_[7907]_ ;
  assign \new_[7916]_  = A167 & A168;
  assign \new_[7920]_  = ~A201 & A200;
  assign \new_[7921]_  = A199 & \new_[7920]_ ;
  assign \new_[7922]_  = \new_[7921]_  & \new_[7916]_ ;
  assign \new_[7925]_  = A233 & ~A202;
  assign \new_[7929]_  = A267 & A265;
  assign \new_[7930]_  = A234 & \new_[7929]_ ;
  assign \new_[7931]_  = \new_[7930]_  & \new_[7925]_ ;
  assign \new_[7934]_  = A167 & A168;
  assign \new_[7938]_  = ~A201 & A200;
  assign \new_[7939]_  = A199 & \new_[7938]_ ;
  assign \new_[7940]_  = \new_[7939]_  & \new_[7934]_ ;
  assign \new_[7943]_  = A233 & ~A202;
  assign \new_[7947]_  = A267 & A266;
  assign \new_[7948]_  = A234 & \new_[7947]_ ;
  assign \new_[7949]_  = \new_[7948]_  & \new_[7943]_ ;
  assign \new_[7952]_  = A167 & A168;
  assign \new_[7956]_  = ~A201 & A200;
  assign \new_[7957]_  = A199 & \new_[7956]_ ;
  assign \new_[7958]_  = \new_[7957]_  & \new_[7952]_ ;
  assign \new_[7961]_  = ~A232 & ~A202;
  assign \new_[7965]_  = A301 & A236;
  assign \new_[7966]_  = A233 & \new_[7965]_ ;
  assign \new_[7967]_  = \new_[7966]_  & \new_[7961]_ ;
  assign \new_[7970]_  = A167 & A168;
  assign \new_[7974]_  = ~A201 & A200;
  assign \new_[7975]_  = A199 & \new_[7974]_ ;
  assign \new_[7976]_  = \new_[7975]_  & \new_[7970]_ ;
  assign \new_[7979]_  = ~A232 & ~A202;
  assign \new_[7983]_  = A268 & A236;
  assign \new_[7984]_  = A233 & \new_[7983]_ ;
  assign \new_[7985]_  = \new_[7984]_  & \new_[7979]_ ;
  assign \new_[7988]_  = A167 & A168;
  assign \new_[7992]_  = ~A201 & A200;
  assign \new_[7993]_  = A199 & \new_[7992]_ ;
  assign \new_[7994]_  = \new_[7993]_  & \new_[7988]_ ;
  assign \new_[7997]_  = A232 & ~A202;
  assign \new_[8001]_  = A301 & A236;
  assign \new_[8002]_  = ~A233 & \new_[8001]_ ;
  assign \new_[8003]_  = \new_[8002]_  & \new_[7997]_ ;
  assign \new_[8006]_  = A167 & A168;
  assign \new_[8010]_  = ~A201 & A200;
  assign \new_[8011]_  = A199 & \new_[8010]_ ;
  assign \new_[8012]_  = \new_[8011]_  & \new_[8006]_ ;
  assign \new_[8015]_  = A232 & ~A202;
  assign \new_[8019]_  = A268 & A236;
  assign \new_[8020]_  = ~A233 & \new_[8019]_ ;
  assign \new_[8021]_  = \new_[8020]_  & \new_[8015]_ ;
  assign \new_[8024]_  = A167 & A168;
  assign \new_[8028]_  = ~A202 & ~A200;
  assign \new_[8029]_  = ~A199 & \new_[8028]_ ;
  assign \new_[8030]_  = \new_[8029]_  & \new_[8024]_ ;
  assign \new_[8033]_  = A234 & A232;
  assign \new_[8037]_  = A302 & ~A299;
  assign \new_[8038]_  = A298 & \new_[8037]_ ;
  assign \new_[8039]_  = \new_[8038]_  & \new_[8033]_ ;
  assign \new_[8042]_  = A167 & A168;
  assign \new_[8046]_  = ~A202 & ~A200;
  assign \new_[8047]_  = ~A199 & \new_[8046]_ ;
  assign \new_[8048]_  = \new_[8047]_  & \new_[8042]_ ;
  assign \new_[8051]_  = A234 & A232;
  assign \new_[8055]_  = A302 & A299;
  assign \new_[8056]_  = ~A298 & \new_[8055]_ ;
  assign \new_[8057]_  = \new_[8056]_  & \new_[8051]_ ;
  assign \new_[8060]_  = A167 & A168;
  assign \new_[8064]_  = ~A202 & ~A200;
  assign \new_[8065]_  = ~A199 & \new_[8064]_ ;
  assign \new_[8066]_  = \new_[8065]_  & \new_[8060]_ ;
  assign \new_[8069]_  = A234 & A232;
  assign \new_[8073]_  = A269 & A266;
  assign \new_[8074]_  = ~A265 & \new_[8073]_ ;
  assign \new_[8075]_  = \new_[8074]_  & \new_[8069]_ ;
  assign \new_[8078]_  = A167 & A168;
  assign \new_[8082]_  = ~A202 & ~A200;
  assign \new_[8083]_  = ~A199 & \new_[8082]_ ;
  assign \new_[8084]_  = \new_[8083]_  & \new_[8078]_ ;
  assign \new_[8087]_  = A234 & A232;
  assign \new_[8091]_  = A269 & ~A266;
  assign \new_[8092]_  = A265 & \new_[8091]_ ;
  assign \new_[8093]_  = \new_[8092]_  & \new_[8087]_ ;
  assign \new_[8096]_  = A167 & A168;
  assign \new_[8100]_  = ~A202 & ~A200;
  assign \new_[8101]_  = ~A199 & \new_[8100]_ ;
  assign \new_[8102]_  = \new_[8101]_  & \new_[8096]_ ;
  assign \new_[8105]_  = A234 & A233;
  assign \new_[8109]_  = A302 & ~A299;
  assign \new_[8110]_  = A298 & \new_[8109]_ ;
  assign \new_[8111]_  = \new_[8110]_  & \new_[8105]_ ;
  assign \new_[8114]_  = A167 & A168;
  assign \new_[8118]_  = ~A202 & ~A200;
  assign \new_[8119]_  = ~A199 & \new_[8118]_ ;
  assign \new_[8120]_  = \new_[8119]_  & \new_[8114]_ ;
  assign \new_[8123]_  = A234 & A233;
  assign \new_[8127]_  = A302 & A299;
  assign \new_[8128]_  = ~A298 & \new_[8127]_ ;
  assign \new_[8129]_  = \new_[8128]_  & \new_[8123]_ ;
  assign \new_[8132]_  = A167 & A168;
  assign \new_[8136]_  = ~A202 & ~A200;
  assign \new_[8137]_  = ~A199 & \new_[8136]_ ;
  assign \new_[8138]_  = \new_[8137]_  & \new_[8132]_ ;
  assign \new_[8141]_  = A234 & A233;
  assign \new_[8145]_  = A269 & A266;
  assign \new_[8146]_  = ~A265 & \new_[8145]_ ;
  assign \new_[8147]_  = \new_[8146]_  & \new_[8141]_ ;
  assign \new_[8150]_  = A167 & A168;
  assign \new_[8154]_  = ~A202 & ~A200;
  assign \new_[8155]_  = ~A199 & \new_[8154]_ ;
  assign \new_[8156]_  = \new_[8155]_  & \new_[8150]_ ;
  assign \new_[8159]_  = A234 & A233;
  assign \new_[8163]_  = A269 & ~A266;
  assign \new_[8164]_  = A265 & \new_[8163]_ ;
  assign \new_[8165]_  = \new_[8164]_  & \new_[8159]_ ;
  assign \new_[8168]_  = A167 & A168;
  assign \new_[8172]_  = ~A202 & ~A200;
  assign \new_[8173]_  = ~A199 & \new_[8172]_ ;
  assign \new_[8174]_  = \new_[8173]_  & \new_[8168]_ ;
  assign \new_[8177]_  = A233 & ~A232;
  assign \new_[8181]_  = A300 & A299;
  assign \new_[8182]_  = A236 & \new_[8181]_ ;
  assign \new_[8183]_  = \new_[8182]_  & \new_[8177]_ ;
  assign \new_[8186]_  = A167 & A168;
  assign \new_[8190]_  = ~A202 & ~A200;
  assign \new_[8191]_  = ~A199 & \new_[8190]_ ;
  assign \new_[8192]_  = \new_[8191]_  & \new_[8186]_ ;
  assign \new_[8195]_  = A233 & ~A232;
  assign \new_[8199]_  = A300 & A298;
  assign \new_[8200]_  = A236 & \new_[8199]_ ;
  assign \new_[8201]_  = \new_[8200]_  & \new_[8195]_ ;
  assign \new_[8204]_  = A167 & A168;
  assign \new_[8208]_  = ~A202 & ~A200;
  assign \new_[8209]_  = ~A199 & \new_[8208]_ ;
  assign \new_[8210]_  = \new_[8209]_  & \new_[8204]_ ;
  assign \new_[8213]_  = A233 & ~A232;
  assign \new_[8217]_  = A267 & A265;
  assign \new_[8218]_  = A236 & \new_[8217]_ ;
  assign \new_[8219]_  = \new_[8218]_  & \new_[8213]_ ;
  assign \new_[8222]_  = A167 & A168;
  assign \new_[8226]_  = ~A202 & ~A200;
  assign \new_[8227]_  = ~A199 & \new_[8226]_ ;
  assign \new_[8228]_  = \new_[8227]_  & \new_[8222]_ ;
  assign \new_[8231]_  = A233 & ~A232;
  assign \new_[8235]_  = A267 & A266;
  assign \new_[8236]_  = A236 & \new_[8235]_ ;
  assign \new_[8237]_  = \new_[8236]_  & \new_[8231]_ ;
  assign \new_[8240]_  = A167 & A168;
  assign \new_[8244]_  = ~A202 & ~A200;
  assign \new_[8245]_  = ~A199 & \new_[8244]_ ;
  assign \new_[8246]_  = \new_[8245]_  & \new_[8240]_ ;
  assign \new_[8249]_  = ~A233 & A232;
  assign \new_[8253]_  = A300 & A299;
  assign \new_[8254]_  = A236 & \new_[8253]_ ;
  assign \new_[8255]_  = \new_[8254]_  & \new_[8249]_ ;
  assign \new_[8258]_  = A167 & A168;
  assign \new_[8262]_  = ~A202 & ~A200;
  assign \new_[8263]_  = ~A199 & \new_[8262]_ ;
  assign \new_[8264]_  = \new_[8263]_  & \new_[8258]_ ;
  assign \new_[8267]_  = ~A233 & A232;
  assign \new_[8271]_  = A300 & A298;
  assign \new_[8272]_  = A236 & \new_[8271]_ ;
  assign \new_[8273]_  = \new_[8272]_  & \new_[8267]_ ;
  assign \new_[8276]_  = A167 & A168;
  assign \new_[8280]_  = ~A202 & ~A200;
  assign \new_[8281]_  = ~A199 & \new_[8280]_ ;
  assign \new_[8282]_  = \new_[8281]_  & \new_[8276]_ ;
  assign \new_[8285]_  = ~A233 & A232;
  assign \new_[8289]_  = A267 & A265;
  assign \new_[8290]_  = A236 & \new_[8289]_ ;
  assign \new_[8291]_  = \new_[8290]_  & \new_[8285]_ ;
  assign \new_[8294]_  = A167 & A168;
  assign \new_[8298]_  = ~A202 & ~A200;
  assign \new_[8299]_  = ~A199 & \new_[8298]_ ;
  assign \new_[8300]_  = \new_[8299]_  & \new_[8294]_ ;
  assign \new_[8303]_  = ~A233 & A232;
  assign \new_[8307]_  = A267 & A266;
  assign \new_[8308]_  = A236 & \new_[8307]_ ;
  assign \new_[8309]_  = \new_[8308]_  & \new_[8303]_ ;
  assign \new_[8312]_  = A167 & A170;
  assign \new_[8316]_  = ~A202 & ~A201;
  assign \new_[8317]_  = ~A166 & \new_[8316]_ ;
  assign \new_[8318]_  = \new_[8317]_  & \new_[8312]_ ;
  assign \new_[8321]_  = A235 & ~A203;
  assign \new_[8325]_  = A302 & ~A299;
  assign \new_[8326]_  = A298 & \new_[8325]_ ;
  assign \new_[8327]_  = \new_[8326]_  & \new_[8321]_ ;
  assign \new_[8330]_  = A167 & A170;
  assign \new_[8334]_  = ~A202 & ~A201;
  assign \new_[8335]_  = ~A166 & \new_[8334]_ ;
  assign \new_[8336]_  = \new_[8335]_  & \new_[8330]_ ;
  assign \new_[8339]_  = A235 & ~A203;
  assign \new_[8343]_  = A302 & A299;
  assign \new_[8344]_  = ~A298 & \new_[8343]_ ;
  assign \new_[8345]_  = \new_[8344]_  & \new_[8339]_ ;
  assign \new_[8348]_  = A167 & A170;
  assign \new_[8352]_  = ~A202 & ~A201;
  assign \new_[8353]_  = ~A166 & \new_[8352]_ ;
  assign \new_[8354]_  = \new_[8353]_  & \new_[8348]_ ;
  assign \new_[8357]_  = A235 & ~A203;
  assign \new_[8361]_  = A269 & A266;
  assign \new_[8362]_  = ~A265 & \new_[8361]_ ;
  assign \new_[8363]_  = \new_[8362]_  & \new_[8357]_ ;
  assign \new_[8366]_  = A167 & A170;
  assign \new_[8370]_  = ~A202 & ~A201;
  assign \new_[8371]_  = ~A166 & \new_[8370]_ ;
  assign \new_[8372]_  = \new_[8371]_  & \new_[8366]_ ;
  assign \new_[8375]_  = A235 & ~A203;
  assign \new_[8379]_  = A269 & ~A266;
  assign \new_[8380]_  = A265 & \new_[8379]_ ;
  assign \new_[8381]_  = \new_[8380]_  & \new_[8375]_ ;
  assign \new_[8384]_  = A167 & A170;
  assign \new_[8388]_  = ~A202 & ~A201;
  assign \new_[8389]_  = ~A166 & \new_[8388]_ ;
  assign \new_[8390]_  = \new_[8389]_  & \new_[8384]_ ;
  assign \new_[8393]_  = A232 & ~A203;
  assign \new_[8397]_  = A300 & A299;
  assign \new_[8398]_  = A234 & \new_[8397]_ ;
  assign \new_[8399]_  = \new_[8398]_  & \new_[8393]_ ;
  assign \new_[8402]_  = A167 & A170;
  assign \new_[8406]_  = ~A202 & ~A201;
  assign \new_[8407]_  = ~A166 & \new_[8406]_ ;
  assign \new_[8408]_  = \new_[8407]_  & \new_[8402]_ ;
  assign \new_[8411]_  = A232 & ~A203;
  assign \new_[8415]_  = A300 & A298;
  assign \new_[8416]_  = A234 & \new_[8415]_ ;
  assign \new_[8417]_  = \new_[8416]_  & \new_[8411]_ ;
  assign \new_[8420]_  = A167 & A170;
  assign \new_[8424]_  = ~A202 & ~A201;
  assign \new_[8425]_  = ~A166 & \new_[8424]_ ;
  assign \new_[8426]_  = \new_[8425]_  & \new_[8420]_ ;
  assign \new_[8429]_  = A232 & ~A203;
  assign \new_[8433]_  = A267 & A265;
  assign \new_[8434]_  = A234 & \new_[8433]_ ;
  assign \new_[8435]_  = \new_[8434]_  & \new_[8429]_ ;
  assign \new_[8438]_  = A167 & A170;
  assign \new_[8442]_  = ~A202 & ~A201;
  assign \new_[8443]_  = ~A166 & \new_[8442]_ ;
  assign \new_[8444]_  = \new_[8443]_  & \new_[8438]_ ;
  assign \new_[8447]_  = A232 & ~A203;
  assign \new_[8451]_  = A267 & A266;
  assign \new_[8452]_  = A234 & \new_[8451]_ ;
  assign \new_[8453]_  = \new_[8452]_  & \new_[8447]_ ;
  assign \new_[8456]_  = A167 & A170;
  assign \new_[8460]_  = ~A202 & ~A201;
  assign \new_[8461]_  = ~A166 & \new_[8460]_ ;
  assign \new_[8462]_  = \new_[8461]_  & \new_[8456]_ ;
  assign \new_[8465]_  = A233 & ~A203;
  assign \new_[8469]_  = A300 & A299;
  assign \new_[8470]_  = A234 & \new_[8469]_ ;
  assign \new_[8471]_  = \new_[8470]_  & \new_[8465]_ ;
  assign \new_[8474]_  = A167 & A170;
  assign \new_[8478]_  = ~A202 & ~A201;
  assign \new_[8479]_  = ~A166 & \new_[8478]_ ;
  assign \new_[8480]_  = \new_[8479]_  & \new_[8474]_ ;
  assign \new_[8483]_  = A233 & ~A203;
  assign \new_[8487]_  = A300 & A298;
  assign \new_[8488]_  = A234 & \new_[8487]_ ;
  assign \new_[8489]_  = \new_[8488]_  & \new_[8483]_ ;
  assign \new_[8492]_  = A167 & A170;
  assign \new_[8496]_  = ~A202 & ~A201;
  assign \new_[8497]_  = ~A166 & \new_[8496]_ ;
  assign \new_[8498]_  = \new_[8497]_  & \new_[8492]_ ;
  assign \new_[8501]_  = A233 & ~A203;
  assign \new_[8505]_  = A267 & A265;
  assign \new_[8506]_  = A234 & \new_[8505]_ ;
  assign \new_[8507]_  = \new_[8506]_  & \new_[8501]_ ;
  assign \new_[8510]_  = A167 & A170;
  assign \new_[8514]_  = ~A202 & ~A201;
  assign \new_[8515]_  = ~A166 & \new_[8514]_ ;
  assign \new_[8516]_  = \new_[8515]_  & \new_[8510]_ ;
  assign \new_[8519]_  = A233 & ~A203;
  assign \new_[8523]_  = A267 & A266;
  assign \new_[8524]_  = A234 & \new_[8523]_ ;
  assign \new_[8525]_  = \new_[8524]_  & \new_[8519]_ ;
  assign \new_[8528]_  = A167 & A170;
  assign \new_[8532]_  = ~A202 & ~A201;
  assign \new_[8533]_  = ~A166 & \new_[8532]_ ;
  assign \new_[8534]_  = \new_[8533]_  & \new_[8528]_ ;
  assign \new_[8537]_  = ~A232 & ~A203;
  assign \new_[8541]_  = A301 & A236;
  assign \new_[8542]_  = A233 & \new_[8541]_ ;
  assign \new_[8543]_  = \new_[8542]_  & \new_[8537]_ ;
  assign \new_[8546]_  = A167 & A170;
  assign \new_[8550]_  = ~A202 & ~A201;
  assign \new_[8551]_  = ~A166 & \new_[8550]_ ;
  assign \new_[8552]_  = \new_[8551]_  & \new_[8546]_ ;
  assign \new_[8555]_  = ~A232 & ~A203;
  assign \new_[8559]_  = A268 & A236;
  assign \new_[8560]_  = A233 & \new_[8559]_ ;
  assign \new_[8561]_  = \new_[8560]_  & \new_[8555]_ ;
  assign \new_[8564]_  = A167 & A170;
  assign \new_[8568]_  = ~A202 & ~A201;
  assign \new_[8569]_  = ~A166 & \new_[8568]_ ;
  assign \new_[8570]_  = \new_[8569]_  & \new_[8564]_ ;
  assign \new_[8573]_  = A232 & ~A203;
  assign \new_[8577]_  = A301 & A236;
  assign \new_[8578]_  = ~A233 & \new_[8577]_ ;
  assign \new_[8579]_  = \new_[8578]_  & \new_[8573]_ ;
  assign \new_[8582]_  = A167 & A170;
  assign \new_[8586]_  = ~A202 & ~A201;
  assign \new_[8587]_  = ~A166 & \new_[8586]_ ;
  assign \new_[8588]_  = \new_[8587]_  & \new_[8582]_ ;
  assign \new_[8591]_  = A232 & ~A203;
  assign \new_[8595]_  = A268 & A236;
  assign \new_[8596]_  = ~A233 & \new_[8595]_ ;
  assign \new_[8597]_  = \new_[8596]_  & \new_[8591]_ ;
  assign \new_[8600]_  = A167 & A170;
  assign \new_[8604]_  = A200 & A199;
  assign \new_[8605]_  = ~A166 & \new_[8604]_ ;
  assign \new_[8606]_  = \new_[8605]_  & \new_[8600]_ ;
  assign \new_[8609]_  = ~A202 & ~A201;
  assign \new_[8613]_  = A300 & A299;
  assign \new_[8614]_  = A235 & \new_[8613]_ ;
  assign \new_[8615]_  = \new_[8614]_  & \new_[8609]_ ;
  assign \new_[8618]_  = A167 & A170;
  assign \new_[8622]_  = A200 & A199;
  assign \new_[8623]_  = ~A166 & \new_[8622]_ ;
  assign \new_[8624]_  = \new_[8623]_  & \new_[8618]_ ;
  assign \new_[8627]_  = ~A202 & ~A201;
  assign \new_[8631]_  = A300 & A298;
  assign \new_[8632]_  = A235 & \new_[8631]_ ;
  assign \new_[8633]_  = \new_[8632]_  & \new_[8627]_ ;
  assign \new_[8636]_  = A167 & A170;
  assign \new_[8640]_  = A200 & A199;
  assign \new_[8641]_  = ~A166 & \new_[8640]_ ;
  assign \new_[8642]_  = \new_[8641]_  & \new_[8636]_ ;
  assign \new_[8645]_  = ~A202 & ~A201;
  assign \new_[8649]_  = A267 & A265;
  assign \new_[8650]_  = A235 & \new_[8649]_ ;
  assign \new_[8651]_  = \new_[8650]_  & \new_[8645]_ ;
  assign \new_[8654]_  = A167 & A170;
  assign \new_[8658]_  = A200 & A199;
  assign \new_[8659]_  = ~A166 & \new_[8658]_ ;
  assign \new_[8660]_  = \new_[8659]_  & \new_[8654]_ ;
  assign \new_[8663]_  = ~A202 & ~A201;
  assign \new_[8667]_  = A267 & A266;
  assign \new_[8668]_  = A235 & \new_[8667]_ ;
  assign \new_[8669]_  = \new_[8668]_  & \new_[8663]_ ;
  assign \new_[8672]_  = A167 & A170;
  assign \new_[8676]_  = A200 & A199;
  assign \new_[8677]_  = ~A166 & \new_[8676]_ ;
  assign \new_[8678]_  = \new_[8677]_  & \new_[8672]_ ;
  assign \new_[8681]_  = ~A202 & ~A201;
  assign \new_[8685]_  = A301 & A234;
  assign \new_[8686]_  = A232 & \new_[8685]_ ;
  assign \new_[8687]_  = \new_[8686]_  & \new_[8681]_ ;
  assign \new_[8690]_  = A167 & A170;
  assign \new_[8694]_  = A200 & A199;
  assign \new_[8695]_  = ~A166 & \new_[8694]_ ;
  assign \new_[8696]_  = \new_[8695]_  & \new_[8690]_ ;
  assign \new_[8699]_  = ~A202 & ~A201;
  assign \new_[8703]_  = A268 & A234;
  assign \new_[8704]_  = A232 & \new_[8703]_ ;
  assign \new_[8705]_  = \new_[8704]_  & \new_[8699]_ ;
  assign \new_[8708]_  = A167 & A170;
  assign \new_[8712]_  = A200 & A199;
  assign \new_[8713]_  = ~A166 & \new_[8712]_ ;
  assign \new_[8714]_  = \new_[8713]_  & \new_[8708]_ ;
  assign \new_[8717]_  = ~A202 & ~A201;
  assign \new_[8721]_  = A301 & A234;
  assign \new_[8722]_  = A233 & \new_[8721]_ ;
  assign \new_[8723]_  = \new_[8722]_  & \new_[8717]_ ;
  assign \new_[8726]_  = A167 & A170;
  assign \new_[8730]_  = A200 & A199;
  assign \new_[8731]_  = ~A166 & \new_[8730]_ ;
  assign \new_[8732]_  = \new_[8731]_  & \new_[8726]_ ;
  assign \new_[8735]_  = ~A202 & ~A201;
  assign \new_[8739]_  = A268 & A234;
  assign \new_[8740]_  = A233 & \new_[8739]_ ;
  assign \new_[8741]_  = \new_[8740]_  & \new_[8735]_ ;
  assign \new_[8744]_  = A167 & A170;
  assign \new_[8748]_  = ~A200 & ~A199;
  assign \new_[8749]_  = ~A166 & \new_[8748]_ ;
  assign \new_[8750]_  = \new_[8749]_  & \new_[8744]_ ;
  assign \new_[8753]_  = A235 & ~A202;
  assign \new_[8757]_  = A302 & ~A299;
  assign \new_[8758]_  = A298 & \new_[8757]_ ;
  assign \new_[8759]_  = \new_[8758]_  & \new_[8753]_ ;
  assign \new_[8762]_  = A167 & A170;
  assign \new_[8766]_  = ~A200 & ~A199;
  assign \new_[8767]_  = ~A166 & \new_[8766]_ ;
  assign \new_[8768]_  = \new_[8767]_  & \new_[8762]_ ;
  assign \new_[8771]_  = A235 & ~A202;
  assign \new_[8775]_  = A302 & A299;
  assign \new_[8776]_  = ~A298 & \new_[8775]_ ;
  assign \new_[8777]_  = \new_[8776]_  & \new_[8771]_ ;
  assign \new_[8780]_  = A167 & A170;
  assign \new_[8784]_  = ~A200 & ~A199;
  assign \new_[8785]_  = ~A166 & \new_[8784]_ ;
  assign \new_[8786]_  = \new_[8785]_  & \new_[8780]_ ;
  assign \new_[8789]_  = A235 & ~A202;
  assign \new_[8793]_  = A269 & A266;
  assign \new_[8794]_  = ~A265 & \new_[8793]_ ;
  assign \new_[8795]_  = \new_[8794]_  & \new_[8789]_ ;
  assign \new_[8798]_  = A167 & A170;
  assign \new_[8802]_  = ~A200 & ~A199;
  assign \new_[8803]_  = ~A166 & \new_[8802]_ ;
  assign \new_[8804]_  = \new_[8803]_  & \new_[8798]_ ;
  assign \new_[8807]_  = A235 & ~A202;
  assign \new_[8811]_  = A269 & ~A266;
  assign \new_[8812]_  = A265 & \new_[8811]_ ;
  assign \new_[8813]_  = \new_[8812]_  & \new_[8807]_ ;
  assign \new_[8816]_  = A167 & A170;
  assign \new_[8820]_  = ~A200 & ~A199;
  assign \new_[8821]_  = ~A166 & \new_[8820]_ ;
  assign \new_[8822]_  = \new_[8821]_  & \new_[8816]_ ;
  assign \new_[8825]_  = A232 & ~A202;
  assign \new_[8829]_  = A300 & A299;
  assign \new_[8830]_  = A234 & \new_[8829]_ ;
  assign \new_[8831]_  = \new_[8830]_  & \new_[8825]_ ;
  assign \new_[8834]_  = A167 & A170;
  assign \new_[8838]_  = ~A200 & ~A199;
  assign \new_[8839]_  = ~A166 & \new_[8838]_ ;
  assign \new_[8840]_  = \new_[8839]_  & \new_[8834]_ ;
  assign \new_[8843]_  = A232 & ~A202;
  assign \new_[8847]_  = A300 & A298;
  assign \new_[8848]_  = A234 & \new_[8847]_ ;
  assign \new_[8849]_  = \new_[8848]_  & \new_[8843]_ ;
  assign \new_[8852]_  = A167 & A170;
  assign \new_[8856]_  = ~A200 & ~A199;
  assign \new_[8857]_  = ~A166 & \new_[8856]_ ;
  assign \new_[8858]_  = \new_[8857]_  & \new_[8852]_ ;
  assign \new_[8861]_  = A232 & ~A202;
  assign \new_[8865]_  = A267 & A265;
  assign \new_[8866]_  = A234 & \new_[8865]_ ;
  assign \new_[8867]_  = \new_[8866]_  & \new_[8861]_ ;
  assign \new_[8870]_  = A167 & A170;
  assign \new_[8874]_  = ~A200 & ~A199;
  assign \new_[8875]_  = ~A166 & \new_[8874]_ ;
  assign \new_[8876]_  = \new_[8875]_  & \new_[8870]_ ;
  assign \new_[8879]_  = A232 & ~A202;
  assign \new_[8883]_  = A267 & A266;
  assign \new_[8884]_  = A234 & \new_[8883]_ ;
  assign \new_[8885]_  = \new_[8884]_  & \new_[8879]_ ;
  assign \new_[8888]_  = A167 & A170;
  assign \new_[8892]_  = ~A200 & ~A199;
  assign \new_[8893]_  = ~A166 & \new_[8892]_ ;
  assign \new_[8894]_  = \new_[8893]_  & \new_[8888]_ ;
  assign \new_[8897]_  = A233 & ~A202;
  assign \new_[8901]_  = A300 & A299;
  assign \new_[8902]_  = A234 & \new_[8901]_ ;
  assign \new_[8903]_  = \new_[8902]_  & \new_[8897]_ ;
  assign \new_[8906]_  = A167 & A170;
  assign \new_[8910]_  = ~A200 & ~A199;
  assign \new_[8911]_  = ~A166 & \new_[8910]_ ;
  assign \new_[8912]_  = \new_[8911]_  & \new_[8906]_ ;
  assign \new_[8915]_  = A233 & ~A202;
  assign \new_[8919]_  = A300 & A298;
  assign \new_[8920]_  = A234 & \new_[8919]_ ;
  assign \new_[8921]_  = \new_[8920]_  & \new_[8915]_ ;
  assign \new_[8924]_  = A167 & A170;
  assign \new_[8928]_  = ~A200 & ~A199;
  assign \new_[8929]_  = ~A166 & \new_[8928]_ ;
  assign \new_[8930]_  = \new_[8929]_  & \new_[8924]_ ;
  assign \new_[8933]_  = A233 & ~A202;
  assign \new_[8937]_  = A267 & A265;
  assign \new_[8938]_  = A234 & \new_[8937]_ ;
  assign \new_[8939]_  = \new_[8938]_  & \new_[8933]_ ;
  assign \new_[8942]_  = A167 & A170;
  assign \new_[8946]_  = ~A200 & ~A199;
  assign \new_[8947]_  = ~A166 & \new_[8946]_ ;
  assign \new_[8948]_  = \new_[8947]_  & \new_[8942]_ ;
  assign \new_[8951]_  = A233 & ~A202;
  assign \new_[8955]_  = A267 & A266;
  assign \new_[8956]_  = A234 & \new_[8955]_ ;
  assign \new_[8957]_  = \new_[8956]_  & \new_[8951]_ ;
  assign \new_[8960]_  = A167 & A170;
  assign \new_[8964]_  = ~A200 & ~A199;
  assign \new_[8965]_  = ~A166 & \new_[8964]_ ;
  assign \new_[8966]_  = \new_[8965]_  & \new_[8960]_ ;
  assign \new_[8969]_  = ~A232 & ~A202;
  assign \new_[8973]_  = A301 & A236;
  assign \new_[8974]_  = A233 & \new_[8973]_ ;
  assign \new_[8975]_  = \new_[8974]_  & \new_[8969]_ ;
  assign \new_[8978]_  = A167 & A170;
  assign \new_[8982]_  = ~A200 & ~A199;
  assign \new_[8983]_  = ~A166 & \new_[8982]_ ;
  assign \new_[8984]_  = \new_[8983]_  & \new_[8978]_ ;
  assign \new_[8987]_  = ~A232 & ~A202;
  assign \new_[8991]_  = A268 & A236;
  assign \new_[8992]_  = A233 & \new_[8991]_ ;
  assign \new_[8993]_  = \new_[8992]_  & \new_[8987]_ ;
  assign \new_[8996]_  = A167 & A170;
  assign \new_[9000]_  = ~A200 & ~A199;
  assign \new_[9001]_  = ~A166 & \new_[9000]_ ;
  assign \new_[9002]_  = \new_[9001]_  & \new_[8996]_ ;
  assign \new_[9005]_  = A232 & ~A202;
  assign \new_[9009]_  = A301 & A236;
  assign \new_[9010]_  = ~A233 & \new_[9009]_ ;
  assign \new_[9011]_  = \new_[9010]_  & \new_[9005]_ ;
  assign \new_[9014]_  = A167 & A170;
  assign \new_[9018]_  = ~A200 & ~A199;
  assign \new_[9019]_  = ~A166 & \new_[9018]_ ;
  assign \new_[9020]_  = \new_[9019]_  & \new_[9014]_ ;
  assign \new_[9023]_  = A232 & ~A202;
  assign \new_[9027]_  = A268 & A236;
  assign \new_[9028]_  = ~A233 & \new_[9027]_ ;
  assign \new_[9029]_  = \new_[9028]_  & \new_[9023]_ ;
  assign \new_[9032]_  = ~A167 & A170;
  assign \new_[9036]_  = ~A202 & ~A201;
  assign \new_[9037]_  = A166 & \new_[9036]_ ;
  assign \new_[9038]_  = \new_[9037]_  & \new_[9032]_ ;
  assign \new_[9041]_  = A235 & ~A203;
  assign \new_[9045]_  = A302 & ~A299;
  assign \new_[9046]_  = A298 & \new_[9045]_ ;
  assign \new_[9047]_  = \new_[9046]_  & \new_[9041]_ ;
  assign \new_[9050]_  = ~A167 & A170;
  assign \new_[9054]_  = ~A202 & ~A201;
  assign \new_[9055]_  = A166 & \new_[9054]_ ;
  assign \new_[9056]_  = \new_[9055]_  & \new_[9050]_ ;
  assign \new_[9059]_  = A235 & ~A203;
  assign \new_[9063]_  = A302 & A299;
  assign \new_[9064]_  = ~A298 & \new_[9063]_ ;
  assign \new_[9065]_  = \new_[9064]_  & \new_[9059]_ ;
  assign \new_[9068]_  = ~A167 & A170;
  assign \new_[9072]_  = ~A202 & ~A201;
  assign \new_[9073]_  = A166 & \new_[9072]_ ;
  assign \new_[9074]_  = \new_[9073]_  & \new_[9068]_ ;
  assign \new_[9077]_  = A235 & ~A203;
  assign \new_[9081]_  = A269 & A266;
  assign \new_[9082]_  = ~A265 & \new_[9081]_ ;
  assign \new_[9083]_  = \new_[9082]_  & \new_[9077]_ ;
  assign \new_[9086]_  = ~A167 & A170;
  assign \new_[9090]_  = ~A202 & ~A201;
  assign \new_[9091]_  = A166 & \new_[9090]_ ;
  assign \new_[9092]_  = \new_[9091]_  & \new_[9086]_ ;
  assign \new_[9095]_  = A235 & ~A203;
  assign \new_[9099]_  = A269 & ~A266;
  assign \new_[9100]_  = A265 & \new_[9099]_ ;
  assign \new_[9101]_  = \new_[9100]_  & \new_[9095]_ ;
  assign \new_[9104]_  = ~A167 & A170;
  assign \new_[9108]_  = ~A202 & ~A201;
  assign \new_[9109]_  = A166 & \new_[9108]_ ;
  assign \new_[9110]_  = \new_[9109]_  & \new_[9104]_ ;
  assign \new_[9113]_  = A232 & ~A203;
  assign \new_[9117]_  = A300 & A299;
  assign \new_[9118]_  = A234 & \new_[9117]_ ;
  assign \new_[9119]_  = \new_[9118]_  & \new_[9113]_ ;
  assign \new_[9122]_  = ~A167 & A170;
  assign \new_[9126]_  = ~A202 & ~A201;
  assign \new_[9127]_  = A166 & \new_[9126]_ ;
  assign \new_[9128]_  = \new_[9127]_  & \new_[9122]_ ;
  assign \new_[9131]_  = A232 & ~A203;
  assign \new_[9135]_  = A300 & A298;
  assign \new_[9136]_  = A234 & \new_[9135]_ ;
  assign \new_[9137]_  = \new_[9136]_  & \new_[9131]_ ;
  assign \new_[9140]_  = ~A167 & A170;
  assign \new_[9144]_  = ~A202 & ~A201;
  assign \new_[9145]_  = A166 & \new_[9144]_ ;
  assign \new_[9146]_  = \new_[9145]_  & \new_[9140]_ ;
  assign \new_[9149]_  = A232 & ~A203;
  assign \new_[9153]_  = A267 & A265;
  assign \new_[9154]_  = A234 & \new_[9153]_ ;
  assign \new_[9155]_  = \new_[9154]_  & \new_[9149]_ ;
  assign \new_[9158]_  = ~A167 & A170;
  assign \new_[9162]_  = ~A202 & ~A201;
  assign \new_[9163]_  = A166 & \new_[9162]_ ;
  assign \new_[9164]_  = \new_[9163]_  & \new_[9158]_ ;
  assign \new_[9167]_  = A232 & ~A203;
  assign \new_[9171]_  = A267 & A266;
  assign \new_[9172]_  = A234 & \new_[9171]_ ;
  assign \new_[9173]_  = \new_[9172]_  & \new_[9167]_ ;
  assign \new_[9176]_  = ~A167 & A170;
  assign \new_[9180]_  = ~A202 & ~A201;
  assign \new_[9181]_  = A166 & \new_[9180]_ ;
  assign \new_[9182]_  = \new_[9181]_  & \new_[9176]_ ;
  assign \new_[9185]_  = A233 & ~A203;
  assign \new_[9189]_  = A300 & A299;
  assign \new_[9190]_  = A234 & \new_[9189]_ ;
  assign \new_[9191]_  = \new_[9190]_  & \new_[9185]_ ;
  assign \new_[9194]_  = ~A167 & A170;
  assign \new_[9198]_  = ~A202 & ~A201;
  assign \new_[9199]_  = A166 & \new_[9198]_ ;
  assign \new_[9200]_  = \new_[9199]_  & \new_[9194]_ ;
  assign \new_[9203]_  = A233 & ~A203;
  assign \new_[9207]_  = A300 & A298;
  assign \new_[9208]_  = A234 & \new_[9207]_ ;
  assign \new_[9209]_  = \new_[9208]_  & \new_[9203]_ ;
  assign \new_[9212]_  = ~A167 & A170;
  assign \new_[9216]_  = ~A202 & ~A201;
  assign \new_[9217]_  = A166 & \new_[9216]_ ;
  assign \new_[9218]_  = \new_[9217]_  & \new_[9212]_ ;
  assign \new_[9221]_  = A233 & ~A203;
  assign \new_[9225]_  = A267 & A265;
  assign \new_[9226]_  = A234 & \new_[9225]_ ;
  assign \new_[9227]_  = \new_[9226]_  & \new_[9221]_ ;
  assign \new_[9230]_  = ~A167 & A170;
  assign \new_[9234]_  = ~A202 & ~A201;
  assign \new_[9235]_  = A166 & \new_[9234]_ ;
  assign \new_[9236]_  = \new_[9235]_  & \new_[9230]_ ;
  assign \new_[9239]_  = A233 & ~A203;
  assign \new_[9243]_  = A267 & A266;
  assign \new_[9244]_  = A234 & \new_[9243]_ ;
  assign \new_[9245]_  = \new_[9244]_  & \new_[9239]_ ;
  assign \new_[9248]_  = ~A167 & A170;
  assign \new_[9252]_  = ~A202 & ~A201;
  assign \new_[9253]_  = A166 & \new_[9252]_ ;
  assign \new_[9254]_  = \new_[9253]_  & \new_[9248]_ ;
  assign \new_[9257]_  = ~A232 & ~A203;
  assign \new_[9261]_  = A301 & A236;
  assign \new_[9262]_  = A233 & \new_[9261]_ ;
  assign \new_[9263]_  = \new_[9262]_  & \new_[9257]_ ;
  assign \new_[9266]_  = ~A167 & A170;
  assign \new_[9270]_  = ~A202 & ~A201;
  assign \new_[9271]_  = A166 & \new_[9270]_ ;
  assign \new_[9272]_  = \new_[9271]_  & \new_[9266]_ ;
  assign \new_[9275]_  = ~A232 & ~A203;
  assign \new_[9279]_  = A268 & A236;
  assign \new_[9280]_  = A233 & \new_[9279]_ ;
  assign \new_[9281]_  = \new_[9280]_  & \new_[9275]_ ;
  assign \new_[9284]_  = ~A167 & A170;
  assign \new_[9288]_  = ~A202 & ~A201;
  assign \new_[9289]_  = A166 & \new_[9288]_ ;
  assign \new_[9290]_  = \new_[9289]_  & \new_[9284]_ ;
  assign \new_[9293]_  = A232 & ~A203;
  assign \new_[9297]_  = A301 & A236;
  assign \new_[9298]_  = ~A233 & \new_[9297]_ ;
  assign \new_[9299]_  = \new_[9298]_  & \new_[9293]_ ;
  assign \new_[9302]_  = ~A167 & A170;
  assign \new_[9306]_  = ~A202 & ~A201;
  assign \new_[9307]_  = A166 & \new_[9306]_ ;
  assign \new_[9308]_  = \new_[9307]_  & \new_[9302]_ ;
  assign \new_[9311]_  = A232 & ~A203;
  assign \new_[9315]_  = A268 & A236;
  assign \new_[9316]_  = ~A233 & \new_[9315]_ ;
  assign \new_[9317]_  = \new_[9316]_  & \new_[9311]_ ;
  assign \new_[9320]_  = ~A167 & A170;
  assign \new_[9324]_  = A200 & A199;
  assign \new_[9325]_  = A166 & \new_[9324]_ ;
  assign \new_[9326]_  = \new_[9325]_  & \new_[9320]_ ;
  assign \new_[9329]_  = ~A202 & ~A201;
  assign \new_[9333]_  = A300 & A299;
  assign \new_[9334]_  = A235 & \new_[9333]_ ;
  assign \new_[9335]_  = \new_[9334]_  & \new_[9329]_ ;
  assign \new_[9338]_  = ~A167 & A170;
  assign \new_[9342]_  = A200 & A199;
  assign \new_[9343]_  = A166 & \new_[9342]_ ;
  assign \new_[9344]_  = \new_[9343]_  & \new_[9338]_ ;
  assign \new_[9347]_  = ~A202 & ~A201;
  assign \new_[9351]_  = A300 & A298;
  assign \new_[9352]_  = A235 & \new_[9351]_ ;
  assign \new_[9353]_  = \new_[9352]_  & \new_[9347]_ ;
  assign \new_[9356]_  = ~A167 & A170;
  assign \new_[9360]_  = A200 & A199;
  assign \new_[9361]_  = A166 & \new_[9360]_ ;
  assign \new_[9362]_  = \new_[9361]_  & \new_[9356]_ ;
  assign \new_[9365]_  = ~A202 & ~A201;
  assign \new_[9369]_  = A267 & A265;
  assign \new_[9370]_  = A235 & \new_[9369]_ ;
  assign \new_[9371]_  = \new_[9370]_  & \new_[9365]_ ;
  assign \new_[9374]_  = ~A167 & A170;
  assign \new_[9378]_  = A200 & A199;
  assign \new_[9379]_  = A166 & \new_[9378]_ ;
  assign \new_[9380]_  = \new_[9379]_  & \new_[9374]_ ;
  assign \new_[9383]_  = ~A202 & ~A201;
  assign \new_[9387]_  = A267 & A266;
  assign \new_[9388]_  = A235 & \new_[9387]_ ;
  assign \new_[9389]_  = \new_[9388]_  & \new_[9383]_ ;
  assign \new_[9392]_  = ~A167 & A170;
  assign \new_[9396]_  = A200 & A199;
  assign \new_[9397]_  = A166 & \new_[9396]_ ;
  assign \new_[9398]_  = \new_[9397]_  & \new_[9392]_ ;
  assign \new_[9401]_  = ~A202 & ~A201;
  assign \new_[9405]_  = A301 & A234;
  assign \new_[9406]_  = A232 & \new_[9405]_ ;
  assign \new_[9407]_  = \new_[9406]_  & \new_[9401]_ ;
  assign \new_[9410]_  = ~A167 & A170;
  assign \new_[9414]_  = A200 & A199;
  assign \new_[9415]_  = A166 & \new_[9414]_ ;
  assign \new_[9416]_  = \new_[9415]_  & \new_[9410]_ ;
  assign \new_[9419]_  = ~A202 & ~A201;
  assign \new_[9423]_  = A268 & A234;
  assign \new_[9424]_  = A232 & \new_[9423]_ ;
  assign \new_[9425]_  = \new_[9424]_  & \new_[9419]_ ;
  assign \new_[9428]_  = ~A167 & A170;
  assign \new_[9432]_  = A200 & A199;
  assign \new_[9433]_  = A166 & \new_[9432]_ ;
  assign \new_[9434]_  = \new_[9433]_  & \new_[9428]_ ;
  assign \new_[9437]_  = ~A202 & ~A201;
  assign \new_[9441]_  = A301 & A234;
  assign \new_[9442]_  = A233 & \new_[9441]_ ;
  assign \new_[9443]_  = \new_[9442]_  & \new_[9437]_ ;
  assign \new_[9446]_  = ~A167 & A170;
  assign \new_[9450]_  = A200 & A199;
  assign \new_[9451]_  = A166 & \new_[9450]_ ;
  assign \new_[9452]_  = \new_[9451]_  & \new_[9446]_ ;
  assign \new_[9455]_  = ~A202 & ~A201;
  assign \new_[9459]_  = A268 & A234;
  assign \new_[9460]_  = A233 & \new_[9459]_ ;
  assign \new_[9461]_  = \new_[9460]_  & \new_[9455]_ ;
  assign \new_[9464]_  = ~A167 & A170;
  assign \new_[9468]_  = ~A200 & ~A199;
  assign \new_[9469]_  = A166 & \new_[9468]_ ;
  assign \new_[9470]_  = \new_[9469]_  & \new_[9464]_ ;
  assign \new_[9473]_  = A235 & ~A202;
  assign \new_[9477]_  = A302 & ~A299;
  assign \new_[9478]_  = A298 & \new_[9477]_ ;
  assign \new_[9479]_  = \new_[9478]_  & \new_[9473]_ ;
  assign \new_[9482]_  = ~A167 & A170;
  assign \new_[9486]_  = ~A200 & ~A199;
  assign \new_[9487]_  = A166 & \new_[9486]_ ;
  assign \new_[9488]_  = \new_[9487]_  & \new_[9482]_ ;
  assign \new_[9491]_  = A235 & ~A202;
  assign \new_[9495]_  = A302 & A299;
  assign \new_[9496]_  = ~A298 & \new_[9495]_ ;
  assign \new_[9497]_  = \new_[9496]_  & \new_[9491]_ ;
  assign \new_[9500]_  = ~A167 & A170;
  assign \new_[9504]_  = ~A200 & ~A199;
  assign \new_[9505]_  = A166 & \new_[9504]_ ;
  assign \new_[9506]_  = \new_[9505]_  & \new_[9500]_ ;
  assign \new_[9509]_  = A235 & ~A202;
  assign \new_[9513]_  = A269 & A266;
  assign \new_[9514]_  = ~A265 & \new_[9513]_ ;
  assign \new_[9515]_  = \new_[9514]_  & \new_[9509]_ ;
  assign \new_[9518]_  = ~A167 & A170;
  assign \new_[9522]_  = ~A200 & ~A199;
  assign \new_[9523]_  = A166 & \new_[9522]_ ;
  assign \new_[9524]_  = \new_[9523]_  & \new_[9518]_ ;
  assign \new_[9527]_  = A235 & ~A202;
  assign \new_[9531]_  = A269 & ~A266;
  assign \new_[9532]_  = A265 & \new_[9531]_ ;
  assign \new_[9533]_  = \new_[9532]_  & \new_[9527]_ ;
  assign \new_[9536]_  = ~A167 & A170;
  assign \new_[9540]_  = ~A200 & ~A199;
  assign \new_[9541]_  = A166 & \new_[9540]_ ;
  assign \new_[9542]_  = \new_[9541]_  & \new_[9536]_ ;
  assign \new_[9545]_  = A232 & ~A202;
  assign \new_[9549]_  = A300 & A299;
  assign \new_[9550]_  = A234 & \new_[9549]_ ;
  assign \new_[9551]_  = \new_[9550]_  & \new_[9545]_ ;
  assign \new_[9554]_  = ~A167 & A170;
  assign \new_[9558]_  = ~A200 & ~A199;
  assign \new_[9559]_  = A166 & \new_[9558]_ ;
  assign \new_[9560]_  = \new_[9559]_  & \new_[9554]_ ;
  assign \new_[9563]_  = A232 & ~A202;
  assign \new_[9567]_  = A300 & A298;
  assign \new_[9568]_  = A234 & \new_[9567]_ ;
  assign \new_[9569]_  = \new_[9568]_  & \new_[9563]_ ;
  assign \new_[9572]_  = ~A167 & A170;
  assign \new_[9576]_  = ~A200 & ~A199;
  assign \new_[9577]_  = A166 & \new_[9576]_ ;
  assign \new_[9578]_  = \new_[9577]_  & \new_[9572]_ ;
  assign \new_[9581]_  = A232 & ~A202;
  assign \new_[9585]_  = A267 & A265;
  assign \new_[9586]_  = A234 & \new_[9585]_ ;
  assign \new_[9587]_  = \new_[9586]_  & \new_[9581]_ ;
  assign \new_[9590]_  = ~A167 & A170;
  assign \new_[9594]_  = ~A200 & ~A199;
  assign \new_[9595]_  = A166 & \new_[9594]_ ;
  assign \new_[9596]_  = \new_[9595]_  & \new_[9590]_ ;
  assign \new_[9599]_  = A232 & ~A202;
  assign \new_[9603]_  = A267 & A266;
  assign \new_[9604]_  = A234 & \new_[9603]_ ;
  assign \new_[9605]_  = \new_[9604]_  & \new_[9599]_ ;
  assign \new_[9608]_  = ~A167 & A170;
  assign \new_[9612]_  = ~A200 & ~A199;
  assign \new_[9613]_  = A166 & \new_[9612]_ ;
  assign \new_[9614]_  = \new_[9613]_  & \new_[9608]_ ;
  assign \new_[9617]_  = A233 & ~A202;
  assign \new_[9621]_  = A300 & A299;
  assign \new_[9622]_  = A234 & \new_[9621]_ ;
  assign \new_[9623]_  = \new_[9622]_  & \new_[9617]_ ;
  assign \new_[9626]_  = ~A167 & A170;
  assign \new_[9630]_  = ~A200 & ~A199;
  assign \new_[9631]_  = A166 & \new_[9630]_ ;
  assign \new_[9632]_  = \new_[9631]_  & \new_[9626]_ ;
  assign \new_[9635]_  = A233 & ~A202;
  assign \new_[9639]_  = A300 & A298;
  assign \new_[9640]_  = A234 & \new_[9639]_ ;
  assign \new_[9641]_  = \new_[9640]_  & \new_[9635]_ ;
  assign \new_[9644]_  = ~A167 & A170;
  assign \new_[9648]_  = ~A200 & ~A199;
  assign \new_[9649]_  = A166 & \new_[9648]_ ;
  assign \new_[9650]_  = \new_[9649]_  & \new_[9644]_ ;
  assign \new_[9653]_  = A233 & ~A202;
  assign \new_[9657]_  = A267 & A265;
  assign \new_[9658]_  = A234 & \new_[9657]_ ;
  assign \new_[9659]_  = \new_[9658]_  & \new_[9653]_ ;
  assign \new_[9662]_  = ~A167 & A170;
  assign \new_[9666]_  = ~A200 & ~A199;
  assign \new_[9667]_  = A166 & \new_[9666]_ ;
  assign \new_[9668]_  = \new_[9667]_  & \new_[9662]_ ;
  assign \new_[9671]_  = A233 & ~A202;
  assign \new_[9675]_  = A267 & A266;
  assign \new_[9676]_  = A234 & \new_[9675]_ ;
  assign \new_[9677]_  = \new_[9676]_  & \new_[9671]_ ;
  assign \new_[9680]_  = ~A167 & A170;
  assign \new_[9684]_  = ~A200 & ~A199;
  assign \new_[9685]_  = A166 & \new_[9684]_ ;
  assign \new_[9686]_  = \new_[9685]_  & \new_[9680]_ ;
  assign \new_[9689]_  = ~A232 & ~A202;
  assign \new_[9693]_  = A301 & A236;
  assign \new_[9694]_  = A233 & \new_[9693]_ ;
  assign \new_[9695]_  = \new_[9694]_  & \new_[9689]_ ;
  assign \new_[9698]_  = ~A167 & A170;
  assign \new_[9702]_  = ~A200 & ~A199;
  assign \new_[9703]_  = A166 & \new_[9702]_ ;
  assign \new_[9704]_  = \new_[9703]_  & \new_[9698]_ ;
  assign \new_[9707]_  = ~A232 & ~A202;
  assign \new_[9711]_  = A268 & A236;
  assign \new_[9712]_  = A233 & \new_[9711]_ ;
  assign \new_[9713]_  = \new_[9712]_  & \new_[9707]_ ;
  assign \new_[9716]_  = ~A167 & A170;
  assign \new_[9720]_  = ~A200 & ~A199;
  assign \new_[9721]_  = A166 & \new_[9720]_ ;
  assign \new_[9722]_  = \new_[9721]_  & \new_[9716]_ ;
  assign \new_[9725]_  = A232 & ~A202;
  assign \new_[9729]_  = A301 & A236;
  assign \new_[9730]_  = ~A233 & \new_[9729]_ ;
  assign \new_[9731]_  = \new_[9730]_  & \new_[9725]_ ;
  assign \new_[9734]_  = ~A167 & A170;
  assign \new_[9738]_  = ~A200 & ~A199;
  assign \new_[9739]_  = A166 & \new_[9738]_ ;
  assign \new_[9740]_  = \new_[9739]_  & \new_[9734]_ ;
  assign \new_[9743]_  = A232 & ~A202;
  assign \new_[9747]_  = A268 & A236;
  assign \new_[9748]_  = ~A233 & \new_[9747]_ ;
  assign \new_[9749]_  = \new_[9748]_  & \new_[9743]_ ;
  assign \new_[9752]_  = ~A201 & A169;
  assign \new_[9756]_  = ~A232 & ~A203;
  assign \new_[9757]_  = ~A202 & \new_[9756]_ ;
  assign \new_[9758]_  = \new_[9757]_  & \new_[9752]_ ;
  assign \new_[9761]_  = A236 & A233;
  assign \new_[9765]_  = A302 & ~A299;
  assign \new_[9766]_  = A298 & \new_[9765]_ ;
  assign \new_[9767]_  = \new_[9766]_  & \new_[9761]_ ;
  assign \new_[9770]_  = ~A201 & A169;
  assign \new_[9774]_  = ~A232 & ~A203;
  assign \new_[9775]_  = ~A202 & \new_[9774]_ ;
  assign \new_[9776]_  = \new_[9775]_  & \new_[9770]_ ;
  assign \new_[9779]_  = A236 & A233;
  assign \new_[9783]_  = A302 & A299;
  assign \new_[9784]_  = ~A298 & \new_[9783]_ ;
  assign \new_[9785]_  = \new_[9784]_  & \new_[9779]_ ;
  assign \new_[9788]_  = ~A201 & A169;
  assign \new_[9792]_  = ~A232 & ~A203;
  assign \new_[9793]_  = ~A202 & \new_[9792]_ ;
  assign \new_[9794]_  = \new_[9793]_  & \new_[9788]_ ;
  assign \new_[9797]_  = A236 & A233;
  assign \new_[9801]_  = A269 & A266;
  assign \new_[9802]_  = ~A265 & \new_[9801]_ ;
  assign \new_[9803]_  = \new_[9802]_  & \new_[9797]_ ;
  assign \new_[9806]_  = ~A201 & A169;
  assign \new_[9810]_  = ~A232 & ~A203;
  assign \new_[9811]_  = ~A202 & \new_[9810]_ ;
  assign \new_[9812]_  = \new_[9811]_  & \new_[9806]_ ;
  assign \new_[9815]_  = A236 & A233;
  assign \new_[9819]_  = A269 & ~A266;
  assign \new_[9820]_  = A265 & \new_[9819]_ ;
  assign \new_[9821]_  = \new_[9820]_  & \new_[9815]_ ;
  assign \new_[9824]_  = ~A201 & A169;
  assign \new_[9828]_  = A232 & ~A203;
  assign \new_[9829]_  = ~A202 & \new_[9828]_ ;
  assign \new_[9830]_  = \new_[9829]_  & \new_[9824]_ ;
  assign \new_[9833]_  = A236 & ~A233;
  assign \new_[9837]_  = A302 & ~A299;
  assign \new_[9838]_  = A298 & \new_[9837]_ ;
  assign \new_[9839]_  = \new_[9838]_  & \new_[9833]_ ;
  assign \new_[9842]_  = ~A201 & A169;
  assign \new_[9846]_  = A232 & ~A203;
  assign \new_[9847]_  = ~A202 & \new_[9846]_ ;
  assign \new_[9848]_  = \new_[9847]_  & \new_[9842]_ ;
  assign \new_[9851]_  = A236 & ~A233;
  assign \new_[9855]_  = A302 & A299;
  assign \new_[9856]_  = ~A298 & \new_[9855]_ ;
  assign \new_[9857]_  = \new_[9856]_  & \new_[9851]_ ;
  assign \new_[9860]_  = ~A201 & A169;
  assign \new_[9864]_  = A232 & ~A203;
  assign \new_[9865]_  = ~A202 & \new_[9864]_ ;
  assign \new_[9866]_  = \new_[9865]_  & \new_[9860]_ ;
  assign \new_[9869]_  = A236 & ~A233;
  assign \new_[9873]_  = A269 & A266;
  assign \new_[9874]_  = ~A265 & \new_[9873]_ ;
  assign \new_[9875]_  = \new_[9874]_  & \new_[9869]_ ;
  assign \new_[9878]_  = ~A201 & A169;
  assign \new_[9882]_  = A232 & ~A203;
  assign \new_[9883]_  = ~A202 & \new_[9882]_ ;
  assign \new_[9884]_  = \new_[9883]_  & \new_[9878]_ ;
  assign \new_[9887]_  = A236 & ~A233;
  assign \new_[9891]_  = A269 & ~A266;
  assign \new_[9892]_  = A265 & \new_[9891]_ ;
  assign \new_[9893]_  = \new_[9892]_  & \new_[9887]_ ;
  assign \new_[9896]_  = A199 & A169;
  assign \new_[9900]_  = ~A202 & ~A201;
  assign \new_[9901]_  = A200 & \new_[9900]_ ;
  assign \new_[9902]_  = \new_[9901]_  & \new_[9896]_ ;
  assign \new_[9905]_  = A234 & A232;
  assign \new_[9909]_  = A302 & ~A299;
  assign \new_[9910]_  = A298 & \new_[9909]_ ;
  assign \new_[9911]_  = \new_[9910]_  & \new_[9905]_ ;
  assign \new_[9914]_  = A199 & A169;
  assign \new_[9918]_  = ~A202 & ~A201;
  assign \new_[9919]_  = A200 & \new_[9918]_ ;
  assign \new_[9920]_  = \new_[9919]_  & \new_[9914]_ ;
  assign \new_[9923]_  = A234 & A232;
  assign \new_[9927]_  = A302 & A299;
  assign \new_[9928]_  = ~A298 & \new_[9927]_ ;
  assign \new_[9929]_  = \new_[9928]_  & \new_[9923]_ ;
  assign \new_[9932]_  = A199 & A169;
  assign \new_[9936]_  = ~A202 & ~A201;
  assign \new_[9937]_  = A200 & \new_[9936]_ ;
  assign \new_[9938]_  = \new_[9937]_  & \new_[9932]_ ;
  assign \new_[9941]_  = A234 & A232;
  assign \new_[9945]_  = A269 & A266;
  assign \new_[9946]_  = ~A265 & \new_[9945]_ ;
  assign \new_[9947]_  = \new_[9946]_  & \new_[9941]_ ;
  assign \new_[9950]_  = A199 & A169;
  assign \new_[9954]_  = ~A202 & ~A201;
  assign \new_[9955]_  = A200 & \new_[9954]_ ;
  assign \new_[9956]_  = \new_[9955]_  & \new_[9950]_ ;
  assign \new_[9959]_  = A234 & A232;
  assign \new_[9963]_  = A269 & ~A266;
  assign \new_[9964]_  = A265 & \new_[9963]_ ;
  assign \new_[9965]_  = \new_[9964]_  & \new_[9959]_ ;
  assign \new_[9968]_  = A199 & A169;
  assign \new_[9972]_  = ~A202 & ~A201;
  assign \new_[9973]_  = A200 & \new_[9972]_ ;
  assign \new_[9974]_  = \new_[9973]_  & \new_[9968]_ ;
  assign \new_[9977]_  = A234 & A233;
  assign \new_[9981]_  = A302 & ~A299;
  assign \new_[9982]_  = A298 & \new_[9981]_ ;
  assign \new_[9983]_  = \new_[9982]_  & \new_[9977]_ ;
  assign \new_[9986]_  = A199 & A169;
  assign \new_[9990]_  = ~A202 & ~A201;
  assign \new_[9991]_  = A200 & \new_[9990]_ ;
  assign \new_[9992]_  = \new_[9991]_  & \new_[9986]_ ;
  assign \new_[9995]_  = A234 & A233;
  assign \new_[9999]_  = A302 & A299;
  assign \new_[10000]_  = ~A298 & \new_[9999]_ ;
  assign \new_[10001]_  = \new_[10000]_  & \new_[9995]_ ;
  assign \new_[10004]_  = A199 & A169;
  assign \new_[10008]_  = ~A202 & ~A201;
  assign \new_[10009]_  = A200 & \new_[10008]_ ;
  assign \new_[10010]_  = \new_[10009]_  & \new_[10004]_ ;
  assign \new_[10013]_  = A234 & A233;
  assign \new_[10017]_  = A269 & A266;
  assign \new_[10018]_  = ~A265 & \new_[10017]_ ;
  assign \new_[10019]_  = \new_[10018]_  & \new_[10013]_ ;
  assign \new_[10022]_  = A199 & A169;
  assign \new_[10026]_  = ~A202 & ~A201;
  assign \new_[10027]_  = A200 & \new_[10026]_ ;
  assign \new_[10028]_  = \new_[10027]_  & \new_[10022]_ ;
  assign \new_[10031]_  = A234 & A233;
  assign \new_[10035]_  = A269 & ~A266;
  assign \new_[10036]_  = A265 & \new_[10035]_ ;
  assign \new_[10037]_  = \new_[10036]_  & \new_[10031]_ ;
  assign \new_[10040]_  = A199 & A169;
  assign \new_[10044]_  = ~A202 & ~A201;
  assign \new_[10045]_  = A200 & \new_[10044]_ ;
  assign \new_[10046]_  = \new_[10045]_  & \new_[10040]_ ;
  assign \new_[10049]_  = A233 & ~A232;
  assign \new_[10053]_  = A300 & A299;
  assign \new_[10054]_  = A236 & \new_[10053]_ ;
  assign \new_[10055]_  = \new_[10054]_  & \new_[10049]_ ;
  assign \new_[10058]_  = A199 & A169;
  assign \new_[10062]_  = ~A202 & ~A201;
  assign \new_[10063]_  = A200 & \new_[10062]_ ;
  assign \new_[10064]_  = \new_[10063]_  & \new_[10058]_ ;
  assign \new_[10067]_  = A233 & ~A232;
  assign \new_[10071]_  = A300 & A298;
  assign \new_[10072]_  = A236 & \new_[10071]_ ;
  assign \new_[10073]_  = \new_[10072]_  & \new_[10067]_ ;
  assign \new_[10076]_  = A199 & A169;
  assign \new_[10080]_  = ~A202 & ~A201;
  assign \new_[10081]_  = A200 & \new_[10080]_ ;
  assign \new_[10082]_  = \new_[10081]_  & \new_[10076]_ ;
  assign \new_[10085]_  = A233 & ~A232;
  assign \new_[10089]_  = A267 & A265;
  assign \new_[10090]_  = A236 & \new_[10089]_ ;
  assign \new_[10091]_  = \new_[10090]_  & \new_[10085]_ ;
  assign \new_[10094]_  = A199 & A169;
  assign \new_[10098]_  = ~A202 & ~A201;
  assign \new_[10099]_  = A200 & \new_[10098]_ ;
  assign \new_[10100]_  = \new_[10099]_  & \new_[10094]_ ;
  assign \new_[10103]_  = A233 & ~A232;
  assign \new_[10107]_  = A267 & A266;
  assign \new_[10108]_  = A236 & \new_[10107]_ ;
  assign \new_[10109]_  = \new_[10108]_  & \new_[10103]_ ;
  assign \new_[10112]_  = A199 & A169;
  assign \new_[10116]_  = ~A202 & ~A201;
  assign \new_[10117]_  = A200 & \new_[10116]_ ;
  assign \new_[10118]_  = \new_[10117]_  & \new_[10112]_ ;
  assign \new_[10121]_  = ~A233 & A232;
  assign \new_[10125]_  = A300 & A299;
  assign \new_[10126]_  = A236 & \new_[10125]_ ;
  assign \new_[10127]_  = \new_[10126]_  & \new_[10121]_ ;
  assign \new_[10130]_  = A199 & A169;
  assign \new_[10134]_  = ~A202 & ~A201;
  assign \new_[10135]_  = A200 & \new_[10134]_ ;
  assign \new_[10136]_  = \new_[10135]_  & \new_[10130]_ ;
  assign \new_[10139]_  = ~A233 & A232;
  assign \new_[10143]_  = A300 & A298;
  assign \new_[10144]_  = A236 & \new_[10143]_ ;
  assign \new_[10145]_  = \new_[10144]_  & \new_[10139]_ ;
  assign \new_[10148]_  = A199 & A169;
  assign \new_[10152]_  = ~A202 & ~A201;
  assign \new_[10153]_  = A200 & \new_[10152]_ ;
  assign \new_[10154]_  = \new_[10153]_  & \new_[10148]_ ;
  assign \new_[10157]_  = ~A233 & A232;
  assign \new_[10161]_  = A267 & A265;
  assign \new_[10162]_  = A236 & \new_[10161]_ ;
  assign \new_[10163]_  = \new_[10162]_  & \new_[10157]_ ;
  assign \new_[10166]_  = A199 & A169;
  assign \new_[10170]_  = ~A202 & ~A201;
  assign \new_[10171]_  = A200 & \new_[10170]_ ;
  assign \new_[10172]_  = \new_[10171]_  & \new_[10166]_ ;
  assign \new_[10175]_  = ~A233 & A232;
  assign \new_[10179]_  = A267 & A266;
  assign \new_[10180]_  = A236 & \new_[10179]_ ;
  assign \new_[10181]_  = \new_[10180]_  & \new_[10175]_ ;
  assign \new_[10184]_  = ~A199 & A169;
  assign \new_[10188]_  = ~A232 & ~A202;
  assign \new_[10189]_  = ~A200 & \new_[10188]_ ;
  assign \new_[10190]_  = \new_[10189]_  & \new_[10184]_ ;
  assign \new_[10193]_  = A236 & A233;
  assign \new_[10197]_  = A302 & ~A299;
  assign \new_[10198]_  = A298 & \new_[10197]_ ;
  assign \new_[10199]_  = \new_[10198]_  & \new_[10193]_ ;
  assign \new_[10202]_  = ~A199 & A169;
  assign \new_[10206]_  = ~A232 & ~A202;
  assign \new_[10207]_  = ~A200 & \new_[10206]_ ;
  assign \new_[10208]_  = \new_[10207]_  & \new_[10202]_ ;
  assign \new_[10211]_  = A236 & A233;
  assign \new_[10215]_  = A302 & A299;
  assign \new_[10216]_  = ~A298 & \new_[10215]_ ;
  assign \new_[10217]_  = \new_[10216]_  & \new_[10211]_ ;
  assign \new_[10220]_  = ~A199 & A169;
  assign \new_[10224]_  = ~A232 & ~A202;
  assign \new_[10225]_  = ~A200 & \new_[10224]_ ;
  assign \new_[10226]_  = \new_[10225]_  & \new_[10220]_ ;
  assign \new_[10229]_  = A236 & A233;
  assign \new_[10233]_  = A269 & A266;
  assign \new_[10234]_  = ~A265 & \new_[10233]_ ;
  assign \new_[10235]_  = \new_[10234]_  & \new_[10229]_ ;
  assign \new_[10238]_  = ~A199 & A169;
  assign \new_[10242]_  = ~A232 & ~A202;
  assign \new_[10243]_  = ~A200 & \new_[10242]_ ;
  assign \new_[10244]_  = \new_[10243]_  & \new_[10238]_ ;
  assign \new_[10247]_  = A236 & A233;
  assign \new_[10251]_  = A269 & ~A266;
  assign \new_[10252]_  = A265 & \new_[10251]_ ;
  assign \new_[10253]_  = \new_[10252]_  & \new_[10247]_ ;
  assign \new_[10256]_  = ~A199 & A169;
  assign \new_[10260]_  = A232 & ~A202;
  assign \new_[10261]_  = ~A200 & \new_[10260]_ ;
  assign \new_[10262]_  = \new_[10261]_  & \new_[10256]_ ;
  assign \new_[10265]_  = A236 & ~A233;
  assign \new_[10269]_  = A302 & ~A299;
  assign \new_[10270]_  = A298 & \new_[10269]_ ;
  assign \new_[10271]_  = \new_[10270]_  & \new_[10265]_ ;
  assign \new_[10274]_  = ~A199 & A169;
  assign \new_[10278]_  = A232 & ~A202;
  assign \new_[10279]_  = ~A200 & \new_[10278]_ ;
  assign \new_[10280]_  = \new_[10279]_  & \new_[10274]_ ;
  assign \new_[10283]_  = A236 & ~A233;
  assign \new_[10287]_  = A302 & A299;
  assign \new_[10288]_  = ~A298 & \new_[10287]_ ;
  assign \new_[10289]_  = \new_[10288]_  & \new_[10283]_ ;
  assign \new_[10292]_  = ~A199 & A169;
  assign \new_[10296]_  = A232 & ~A202;
  assign \new_[10297]_  = ~A200 & \new_[10296]_ ;
  assign \new_[10298]_  = \new_[10297]_  & \new_[10292]_ ;
  assign \new_[10301]_  = A236 & ~A233;
  assign \new_[10305]_  = A269 & A266;
  assign \new_[10306]_  = ~A265 & \new_[10305]_ ;
  assign \new_[10307]_  = \new_[10306]_  & \new_[10301]_ ;
  assign \new_[10310]_  = ~A199 & A169;
  assign \new_[10314]_  = A232 & ~A202;
  assign \new_[10315]_  = ~A200 & \new_[10314]_ ;
  assign \new_[10316]_  = \new_[10315]_  & \new_[10310]_ ;
  assign \new_[10319]_  = A236 & ~A233;
  assign \new_[10323]_  = A269 & ~A266;
  assign \new_[10324]_  = A265 & \new_[10323]_ ;
  assign \new_[10325]_  = \new_[10324]_  & \new_[10319]_ ;
  assign \new_[10328]_  = A166 & A168;
  assign \new_[10332]_  = ~A203 & ~A202;
  assign \new_[10333]_  = ~A201 & \new_[10332]_ ;
  assign \new_[10334]_  = \new_[10333]_  & \new_[10328]_ ;
  assign \new_[10338]_  = A236 & A233;
  assign \new_[10339]_  = ~A232 & \new_[10338]_ ;
  assign \new_[10343]_  = A302 & ~A299;
  assign \new_[10344]_  = A298 & \new_[10343]_ ;
  assign \new_[10345]_  = \new_[10344]_  & \new_[10339]_ ;
  assign \new_[10348]_  = A166 & A168;
  assign \new_[10352]_  = ~A203 & ~A202;
  assign \new_[10353]_  = ~A201 & \new_[10352]_ ;
  assign \new_[10354]_  = \new_[10353]_  & \new_[10348]_ ;
  assign \new_[10358]_  = A236 & A233;
  assign \new_[10359]_  = ~A232 & \new_[10358]_ ;
  assign \new_[10363]_  = A302 & A299;
  assign \new_[10364]_  = ~A298 & \new_[10363]_ ;
  assign \new_[10365]_  = \new_[10364]_  & \new_[10359]_ ;
  assign \new_[10368]_  = A166 & A168;
  assign \new_[10372]_  = ~A203 & ~A202;
  assign \new_[10373]_  = ~A201 & \new_[10372]_ ;
  assign \new_[10374]_  = \new_[10373]_  & \new_[10368]_ ;
  assign \new_[10378]_  = A236 & A233;
  assign \new_[10379]_  = ~A232 & \new_[10378]_ ;
  assign \new_[10383]_  = A269 & A266;
  assign \new_[10384]_  = ~A265 & \new_[10383]_ ;
  assign \new_[10385]_  = \new_[10384]_  & \new_[10379]_ ;
  assign \new_[10388]_  = A166 & A168;
  assign \new_[10392]_  = ~A203 & ~A202;
  assign \new_[10393]_  = ~A201 & \new_[10392]_ ;
  assign \new_[10394]_  = \new_[10393]_  & \new_[10388]_ ;
  assign \new_[10398]_  = A236 & A233;
  assign \new_[10399]_  = ~A232 & \new_[10398]_ ;
  assign \new_[10403]_  = A269 & ~A266;
  assign \new_[10404]_  = A265 & \new_[10403]_ ;
  assign \new_[10405]_  = \new_[10404]_  & \new_[10399]_ ;
  assign \new_[10408]_  = A166 & A168;
  assign \new_[10412]_  = ~A203 & ~A202;
  assign \new_[10413]_  = ~A201 & \new_[10412]_ ;
  assign \new_[10414]_  = \new_[10413]_  & \new_[10408]_ ;
  assign \new_[10418]_  = A236 & ~A233;
  assign \new_[10419]_  = A232 & \new_[10418]_ ;
  assign \new_[10423]_  = A302 & ~A299;
  assign \new_[10424]_  = A298 & \new_[10423]_ ;
  assign \new_[10425]_  = \new_[10424]_  & \new_[10419]_ ;
  assign \new_[10428]_  = A166 & A168;
  assign \new_[10432]_  = ~A203 & ~A202;
  assign \new_[10433]_  = ~A201 & \new_[10432]_ ;
  assign \new_[10434]_  = \new_[10433]_  & \new_[10428]_ ;
  assign \new_[10438]_  = A236 & ~A233;
  assign \new_[10439]_  = A232 & \new_[10438]_ ;
  assign \new_[10443]_  = A302 & A299;
  assign \new_[10444]_  = ~A298 & \new_[10443]_ ;
  assign \new_[10445]_  = \new_[10444]_  & \new_[10439]_ ;
  assign \new_[10448]_  = A166 & A168;
  assign \new_[10452]_  = ~A203 & ~A202;
  assign \new_[10453]_  = ~A201 & \new_[10452]_ ;
  assign \new_[10454]_  = \new_[10453]_  & \new_[10448]_ ;
  assign \new_[10458]_  = A236 & ~A233;
  assign \new_[10459]_  = A232 & \new_[10458]_ ;
  assign \new_[10463]_  = A269 & A266;
  assign \new_[10464]_  = ~A265 & \new_[10463]_ ;
  assign \new_[10465]_  = \new_[10464]_  & \new_[10459]_ ;
  assign \new_[10468]_  = A166 & A168;
  assign \new_[10472]_  = ~A203 & ~A202;
  assign \new_[10473]_  = ~A201 & \new_[10472]_ ;
  assign \new_[10474]_  = \new_[10473]_  & \new_[10468]_ ;
  assign \new_[10478]_  = A236 & ~A233;
  assign \new_[10479]_  = A232 & \new_[10478]_ ;
  assign \new_[10483]_  = A269 & ~A266;
  assign \new_[10484]_  = A265 & \new_[10483]_ ;
  assign \new_[10485]_  = \new_[10484]_  & \new_[10479]_ ;
  assign \new_[10488]_  = A166 & A168;
  assign \new_[10492]_  = ~A201 & A200;
  assign \new_[10493]_  = A199 & \new_[10492]_ ;
  assign \new_[10494]_  = \new_[10493]_  & \new_[10488]_ ;
  assign \new_[10498]_  = A234 & A232;
  assign \new_[10499]_  = ~A202 & \new_[10498]_ ;
  assign \new_[10503]_  = A302 & ~A299;
  assign \new_[10504]_  = A298 & \new_[10503]_ ;
  assign \new_[10505]_  = \new_[10504]_  & \new_[10499]_ ;
  assign \new_[10508]_  = A166 & A168;
  assign \new_[10512]_  = ~A201 & A200;
  assign \new_[10513]_  = A199 & \new_[10512]_ ;
  assign \new_[10514]_  = \new_[10513]_  & \new_[10508]_ ;
  assign \new_[10518]_  = A234 & A232;
  assign \new_[10519]_  = ~A202 & \new_[10518]_ ;
  assign \new_[10523]_  = A302 & A299;
  assign \new_[10524]_  = ~A298 & \new_[10523]_ ;
  assign \new_[10525]_  = \new_[10524]_  & \new_[10519]_ ;
  assign \new_[10528]_  = A166 & A168;
  assign \new_[10532]_  = ~A201 & A200;
  assign \new_[10533]_  = A199 & \new_[10532]_ ;
  assign \new_[10534]_  = \new_[10533]_  & \new_[10528]_ ;
  assign \new_[10538]_  = A234 & A232;
  assign \new_[10539]_  = ~A202 & \new_[10538]_ ;
  assign \new_[10543]_  = A269 & A266;
  assign \new_[10544]_  = ~A265 & \new_[10543]_ ;
  assign \new_[10545]_  = \new_[10544]_  & \new_[10539]_ ;
  assign \new_[10548]_  = A166 & A168;
  assign \new_[10552]_  = ~A201 & A200;
  assign \new_[10553]_  = A199 & \new_[10552]_ ;
  assign \new_[10554]_  = \new_[10553]_  & \new_[10548]_ ;
  assign \new_[10558]_  = A234 & A232;
  assign \new_[10559]_  = ~A202 & \new_[10558]_ ;
  assign \new_[10563]_  = A269 & ~A266;
  assign \new_[10564]_  = A265 & \new_[10563]_ ;
  assign \new_[10565]_  = \new_[10564]_  & \new_[10559]_ ;
  assign \new_[10568]_  = A166 & A168;
  assign \new_[10572]_  = ~A201 & A200;
  assign \new_[10573]_  = A199 & \new_[10572]_ ;
  assign \new_[10574]_  = \new_[10573]_  & \new_[10568]_ ;
  assign \new_[10578]_  = A234 & A233;
  assign \new_[10579]_  = ~A202 & \new_[10578]_ ;
  assign \new_[10583]_  = A302 & ~A299;
  assign \new_[10584]_  = A298 & \new_[10583]_ ;
  assign \new_[10585]_  = \new_[10584]_  & \new_[10579]_ ;
  assign \new_[10588]_  = A166 & A168;
  assign \new_[10592]_  = ~A201 & A200;
  assign \new_[10593]_  = A199 & \new_[10592]_ ;
  assign \new_[10594]_  = \new_[10593]_  & \new_[10588]_ ;
  assign \new_[10598]_  = A234 & A233;
  assign \new_[10599]_  = ~A202 & \new_[10598]_ ;
  assign \new_[10603]_  = A302 & A299;
  assign \new_[10604]_  = ~A298 & \new_[10603]_ ;
  assign \new_[10605]_  = \new_[10604]_  & \new_[10599]_ ;
  assign \new_[10608]_  = A166 & A168;
  assign \new_[10612]_  = ~A201 & A200;
  assign \new_[10613]_  = A199 & \new_[10612]_ ;
  assign \new_[10614]_  = \new_[10613]_  & \new_[10608]_ ;
  assign \new_[10618]_  = A234 & A233;
  assign \new_[10619]_  = ~A202 & \new_[10618]_ ;
  assign \new_[10623]_  = A269 & A266;
  assign \new_[10624]_  = ~A265 & \new_[10623]_ ;
  assign \new_[10625]_  = \new_[10624]_  & \new_[10619]_ ;
  assign \new_[10628]_  = A166 & A168;
  assign \new_[10632]_  = ~A201 & A200;
  assign \new_[10633]_  = A199 & \new_[10632]_ ;
  assign \new_[10634]_  = \new_[10633]_  & \new_[10628]_ ;
  assign \new_[10638]_  = A234 & A233;
  assign \new_[10639]_  = ~A202 & \new_[10638]_ ;
  assign \new_[10643]_  = A269 & ~A266;
  assign \new_[10644]_  = A265 & \new_[10643]_ ;
  assign \new_[10645]_  = \new_[10644]_  & \new_[10639]_ ;
  assign \new_[10648]_  = A166 & A168;
  assign \new_[10652]_  = ~A201 & A200;
  assign \new_[10653]_  = A199 & \new_[10652]_ ;
  assign \new_[10654]_  = \new_[10653]_  & \new_[10648]_ ;
  assign \new_[10658]_  = A233 & ~A232;
  assign \new_[10659]_  = ~A202 & \new_[10658]_ ;
  assign \new_[10663]_  = A300 & A299;
  assign \new_[10664]_  = A236 & \new_[10663]_ ;
  assign \new_[10665]_  = \new_[10664]_  & \new_[10659]_ ;
  assign \new_[10668]_  = A166 & A168;
  assign \new_[10672]_  = ~A201 & A200;
  assign \new_[10673]_  = A199 & \new_[10672]_ ;
  assign \new_[10674]_  = \new_[10673]_  & \new_[10668]_ ;
  assign \new_[10678]_  = A233 & ~A232;
  assign \new_[10679]_  = ~A202 & \new_[10678]_ ;
  assign \new_[10683]_  = A300 & A298;
  assign \new_[10684]_  = A236 & \new_[10683]_ ;
  assign \new_[10685]_  = \new_[10684]_  & \new_[10679]_ ;
  assign \new_[10688]_  = A166 & A168;
  assign \new_[10692]_  = ~A201 & A200;
  assign \new_[10693]_  = A199 & \new_[10692]_ ;
  assign \new_[10694]_  = \new_[10693]_  & \new_[10688]_ ;
  assign \new_[10698]_  = A233 & ~A232;
  assign \new_[10699]_  = ~A202 & \new_[10698]_ ;
  assign \new_[10703]_  = A267 & A265;
  assign \new_[10704]_  = A236 & \new_[10703]_ ;
  assign \new_[10705]_  = \new_[10704]_  & \new_[10699]_ ;
  assign \new_[10708]_  = A166 & A168;
  assign \new_[10712]_  = ~A201 & A200;
  assign \new_[10713]_  = A199 & \new_[10712]_ ;
  assign \new_[10714]_  = \new_[10713]_  & \new_[10708]_ ;
  assign \new_[10718]_  = A233 & ~A232;
  assign \new_[10719]_  = ~A202 & \new_[10718]_ ;
  assign \new_[10723]_  = A267 & A266;
  assign \new_[10724]_  = A236 & \new_[10723]_ ;
  assign \new_[10725]_  = \new_[10724]_  & \new_[10719]_ ;
  assign \new_[10728]_  = A166 & A168;
  assign \new_[10732]_  = ~A201 & A200;
  assign \new_[10733]_  = A199 & \new_[10732]_ ;
  assign \new_[10734]_  = \new_[10733]_  & \new_[10728]_ ;
  assign \new_[10738]_  = ~A233 & A232;
  assign \new_[10739]_  = ~A202 & \new_[10738]_ ;
  assign \new_[10743]_  = A300 & A299;
  assign \new_[10744]_  = A236 & \new_[10743]_ ;
  assign \new_[10745]_  = \new_[10744]_  & \new_[10739]_ ;
  assign \new_[10748]_  = A166 & A168;
  assign \new_[10752]_  = ~A201 & A200;
  assign \new_[10753]_  = A199 & \new_[10752]_ ;
  assign \new_[10754]_  = \new_[10753]_  & \new_[10748]_ ;
  assign \new_[10758]_  = ~A233 & A232;
  assign \new_[10759]_  = ~A202 & \new_[10758]_ ;
  assign \new_[10763]_  = A300 & A298;
  assign \new_[10764]_  = A236 & \new_[10763]_ ;
  assign \new_[10765]_  = \new_[10764]_  & \new_[10759]_ ;
  assign \new_[10768]_  = A166 & A168;
  assign \new_[10772]_  = ~A201 & A200;
  assign \new_[10773]_  = A199 & \new_[10772]_ ;
  assign \new_[10774]_  = \new_[10773]_  & \new_[10768]_ ;
  assign \new_[10778]_  = ~A233 & A232;
  assign \new_[10779]_  = ~A202 & \new_[10778]_ ;
  assign \new_[10783]_  = A267 & A265;
  assign \new_[10784]_  = A236 & \new_[10783]_ ;
  assign \new_[10785]_  = \new_[10784]_  & \new_[10779]_ ;
  assign \new_[10788]_  = A166 & A168;
  assign \new_[10792]_  = ~A201 & A200;
  assign \new_[10793]_  = A199 & \new_[10792]_ ;
  assign \new_[10794]_  = \new_[10793]_  & \new_[10788]_ ;
  assign \new_[10798]_  = ~A233 & A232;
  assign \new_[10799]_  = ~A202 & \new_[10798]_ ;
  assign \new_[10803]_  = A267 & A266;
  assign \new_[10804]_  = A236 & \new_[10803]_ ;
  assign \new_[10805]_  = \new_[10804]_  & \new_[10799]_ ;
  assign \new_[10808]_  = A166 & A168;
  assign \new_[10812]_  = ~A202 & ~A200;
  assign \new_[10813]_  = ~A199 & \new_[10812]_ ;
  assign \new_[10814]_  = \new_[10813]_  & \new_[10808]_ ;
  assign \new_[10818]_  = A236 & A233;
  assign \new_[10819]_  = ~A232 & \new_[10818]_ ;
  assign \new_[10823]_  = A302 & ~A299;
  assign \new_[10824]_  = A298 & \new_[10823]_ ;
  assign \new_[10825]_  = \new_[10824]_  & \new_[10819]_ ;
  assign \new_[10828]_  = A166 & A168;
  assign \new_[10832]_  = ~A202 & ~A200;
  assign \new_[10833]_  = ~A199 & \new_[10832]_ ;
  assign \new_[10834]_  = \new_[10833]_  & \new_[10828]_ ;
  assign \new_[10838]_  = A236 & A233;
  assign \new_[10839]_  = ~A232 & \new_[10838]_ ;
  assign \new_[10843]_  = A302 & A299;
  assign \new_[10844]_  = ~A298 & \new_[10843]_ ;
  assign \new_[10845]_  = \new_[10844]_  & \new_[10839]_ ;
  assign \new_[10848]_  = A166 & A168;
  assign \new_[10852]_  = ~A202 & ~A200;
  assign \new_[10853]_  = ~A199 & \new_[10852]_ ;
  assign \new_[10854]_  = \new_[10853]_  & \new_[10848]_ ;
  assign \new_[10858]_  = A236 & A233;
  assign \new_[10859]_  = ~A232 & \new_[10858]_ ;
  assign \new_[10863]_  = A269 & A266;
  assign \new_[10864]_  = ~A265 & \new_[10863]_ ;
  assign \new_[10865]_  = \new_[10864]_  & \new_[10859]_ ;
  assign \new_[10868]_  = A166 & A168;
  assign \new_[10872]_  = ~A202 & ~A200;
  assign \new_[10873]_  = ~A199 & \new_[10872]_ ;
  assign \new_[10874]_  = \new_[10873]_  & \new_[10868]_ ;
  assign \new_[10878]_  = A236 & A233;
  assign \new_[10879]_  = ~A232 & \new_[10878]_ ;
  assign \new_[10883]_  = A269 & ~A266;
  assign \new_[10884]_  = A265 & \new_[10883]_ ;
  assign \new_[10885]_  = \new_[10884]_  & \new_[10879]_ ;
  assign \new_[10888]_  = A166 & A168;
  assign \new_[10892]_  = ~A202 & ~A200;
  assign \new_[10893]_  = ~A199 & \new_[10892]_ ;
  assign \new_[10894]_  = \new_[10893]_  & \new_[10888]_ ;
  assign \new_[10898]_  = A236 & ~A233;
  assign \new_[10899]_  = A232 & \new_[10898]_ ;
  assign \new_[10903]_  = A302 & ~A299;
  assign \new_[10904]_  = A298 & \new_[10903]_ ;
  assign \new_[10905]_  = \new_[10904]_  & \new_[10899]_ ;
  assign \new_[10908]_  = A166 & A168;
  assign \new_[10912]_  = ~A202 & ~A200;
  assign \new_[10913]_  = ~A199 & \new_[10912]_ ;
  assign \new_[10914]_  = \new_[10913]_  & \new_[10908]_ ;
  assign \new_[10918]_  = A236 & ~A233;
  assign \new_[10919]_  = A232 & \new_[10918]_ ;
  assign \new_[10923]_  = A302 & A299;
  assign \new_[10924]_  = ~A298 & \new_[10923]_ ;
  assign \new_[10925]_  = \new_[10924]_  & \new_[10919]_ ;
  assign \new_[10928]_  = A166 & A168;
  assign \new_[10932]_  = ~A202 & ~A200;
  assign \new_[10933]_  = ~A199 & \new_[10932]_ ;
  assign \new_[10934]_  = \new_[10933]_  & \new_[10928]_ ;
  assign \new_[10938]_  = A236 & ~A233;
  assign \new_[10939]_  = A232 & \new_[10938]_ ;
  assign \new_[10943]_  = A269 & A266;
  assign \new_[10944]_  = ~A265 & \new_[10943]_ ;
  assign \new_[10945]_  = \new_[10944]_  & \new_[10939]_ ;
  assign \new_[10948]_  = A166 & A168;
  assign \new_[10952]_  = ~A202 & ~A200;
  assign \new_[10953]_  = ~A199 & \new_[10952]_ ;
  assign \new_[10954]_  = \new_[10953]_  & \new_[10948]_ ;
  assign \new_[10958]_  = A236 & ~A233;
  assign \new_[10959]_  = A232 & \new_[10958]_ ;
  assign \new_[10963]_  = A269 & ~A266;
  assign \new_[10964]_  = A265 & \new_[10963]_ ;
  assign \new_[10965]_  = \new_[10964]_  & \new_[10959]_ ;
  assign \new_[10968]_  = A167 & A168;
  assign \new_[10972]_  = ~A203 & ~A202;
  assign \new_[10973]_  = ~A201 & \new_[10972]_ ;
  assign \new_[10974]_  = \new_[10973]_  & \new_[10968]_ ;
  assign \new_[10978]_  = A236 & A233;
  assign \new_[10979]_  = ~A232 & \new_[10978]_ ;
  assign \new_[10983]_  = A302 & ~A299;
  assign \new_[10984]_  = A298 & \new_[10983]_ ;
  assign \new_[10985]_  = \new_[10984]_  & \new_[10979]_ ;
  assign \new_[10988]_  = A167 & A168;
  assign \new_[10992]_  = ~A203 & ~A202;
  assign \new_[10993]_  = ~A201 & \new_[10992]_ ;
  assign \new_[10994]_  = \new_[10993]_  & \new_[10988]_ ;
  assign \new_[10998]_  = A236 & A233;
  assign \new_[10999]_  = ~A232 & \new_[10998]_ ;
  assign \new_[11003]_  = A302 & A299;
  assign \new_[11004]_  = ~A298 & \new_[11003]_ ;
  assign \new_[11005]_  = \new_[11004]_  & \new_[10999]_ ;
  assign \new_[11008]_  = A167 & A168;
  assign \new_[11012]_  = ~A203 & ~A202;
  assign \new_[11013]_  = ~A201 & \new_[11012]_ ;
  assign \new_[11014]_  = \new_[11013]_  & \new_[11008]_ ;
  assign \new_[11018]_  = A236 & A233;
  assign \new_[11019]_  = ~A232 & \new_[11018]_ ;
  assign \new_[11023]_  = A269 & A266;
  assign \new_[11024]_  = ~A265 & \new_[11023]_ ;
  assign \new_[11025]_  = \new_[11024]_  & \new_[11019]_ ;
  assign \new_[11028]_  = A167 & A168;
  assign \new_[11032]_  = ~A203 & ~A202;
  assign \new_[11033]_  = ~A201 & \new_[11032]_ ;
  assign \new_[11034]_  = \new_[11033]_  & \new_[11028]_ ;
  assign \new_[11038]_  = A236 & A233;
  assign \new_[11039]_  = ~A232 & \new_[11038]_ ;
  assign \new_[11043]_  = A269 & ~A266;
  assign \new_[11044]_  = A265 & \new_[11043]_ ;
  assign \new_[11045]_  = \new_[11044]_  & \new_[11039]_ ;
  assign \new_[11048]_  = A167 & A168;
  assign \new_[11052]_  = ~A203 & ~A202;
  assign \new_[11053]_  = ~A201 & \new_[11052]_ ;
  assign \new_[11054]_  = \new_[11053]_  & \new_[11048]_ ;
  assign \new_[11058]_  = A236 & ~A233;
  assign \new_[11059]_  = A232 & \new_[11058]_ ;
  assign \new_[11063]_  = A302 & ~A299;
  assign \new_[11064]_  = A298 & \new_[11063]_ ;
  assign \new_[11065]_  = \new_[11064]_  & \new_[11059]_ ;
  assign \new_[11068]_  = A167 & A168;
  assign \new_[11072]_  = ~A203 & ~A202;
  assign \new_[11073]_  = ~A201 & \new_[11072]_ ;
  assign \new_[11074]_  = \new_[11073]_  & \new_[11068]_ ;
  assign \new_[11078]_  = A236 & ~A233;
  assign \new_[11079]_  = A232 & \new_[11078]_ ;
  assign \new_[11083]_  = A302 & A299;
  assign \new_[11084]_  = ~A298 & \new_[11083]_ ;
  assign \new_[11085]_  = \new_[11084]_  & \new_[11079]_ ;
  assign \new_[11088]_  = A167 & A168;
  assign \new_[11092]_  = ~A203 & ~A202;
  assign \new_[11093]_  = ~A201 & \new_[11092]_ ;
  assign \new_[11094]_  = \new_[11093]_  & \new_[11088]_ ;
  assign \new_[11098]_  = A236 & ~A233;
  assign \new_[11099]_  = A232 & \new_[11098]_ ;
  assign \new_[11103]_  = A269 & A266;
  assign \new_[11104]_  = ~A265 & \new_[11103]_ ;
  assign \new_[11105]_  = \new_[11104]_  & \new_[11099]_ ;
  assign \new_[11108]_  = A167 & A168;
  assign \new_[11112]_  = ~A203 & ~A202;
  assign \new_[11113]_  = ~A201 & \new_[11112]_ ;
  assign \new_[11114]_  = \new_[11113]_  & \new_[11108]_ ;
  assign \new_[11118]_  = A236 & ~A233;
  assign \new_[11119]_  = A232 & \new_[11118]_ ;
  assign \new_[11123]_  = A269 & ~A266;
  assign \new_[11124]_  = A265 & \new_[11123]_ ;
  assign \new_[11125]_  = \new_[11124]_  & \new_[11119]_ ;
  assign \new_[11128]_  = A167 & A168;
  assign \new_[11132]_  = ~A201 & A200;
  assign \new_[11133]_  = A199 & \new_[11132]_ ;
  assign \new_[11134]_  = \new_[11133]_  & \new_[11128]_ ;
  assign \new_[11138]_  = A234 & A232;
  assign \new_[11139]_  = ~A202 & \new_[11138]_ ;
  assign \new_[11143]_  = A302 & ~A299;
  assign \new_[11144]_  = A298 & \new_[11143]_ ;
  assign \new_[11145]_  = \new_[11144]_  & \new_[11139]_ ;
  assign \new_[11148]_  = A167 & A168;
  assign \new_[11152]_  = ~A201 & A200;
  assign \new_[11153]_  = A199 & \new_[11152]_ ;
  assign \new_[11154]_  = \new_[11153]_  & \new_[11148]_ ;
  assign \new_[11158]_  = A234 & A232;
  assign \new_[11159]_  = ~A202 & \new_[11158]_ ;
  assign \new_[11163]_  = A302 & A299;
  assign \new_[11164]_  = ~A298 & \new_[11163]_ ;
  assign \new_[11165]_  = \new_[11164]_  & \new_[11159]_ ;
  assign \new_[11168]_  = A167 & A168;
  assign \new_[11172]_  = ~A201 & A200;
  assign \new_[11173]_  = A199 & \new_[11172]_ ;
  assign \new_[11174]_  = \new_[11173]_  & \new_[11168]_ ;
  assign \new_[11178]_  = A234 & A232;
  assign \new_[11179]_  = ~A202 & \new_[11178]_ ;
  assign \new_[11183]_  = A269 & A266;
  assign \new_[11184]_  = ~A265 & \new_[11183]_ ;
  assign \new_[11185]_  = \new_[11184]_  & \new_[11179]_ ;
  assign \new_[11188]_  = A167 & A168;
  assign \new_[11192]_  = ~A201 & A200;
  assign \new_[11193]_  = A199 & \new_[11192]_ ;
  assign \new_[11194]_  = \new_[11193]_  & \new_[11188]_ ;
  assign \new_[11198]_  = A234 & A232;
  assign \new_[11199]_  = ~A202 & \new_[11198]_ ;
  assign \new_[11203]_  = A269 & ~A266;
  assign \new_[11204]_  = A265 & \new_[11203]_ ;
  assign \new_[11205]_  = \new_[11204]_  & \new_[11199]_ ;
  assign \new_[11208]_  = A167 & A168;
  assign \new_[11212]_  = ~A201 & A200;
  assign \new_[11213]_  = A199 & \new_[11212]_ ;
  assign \new_[11214]_  = \new_[11213]_  & \new_[11208]_ ;
  assign \new_[11218]_  = A234 & A233;
  assign \new_[11219]_  = ~A202 & \new_[11218]_ ;
  assign \new_[11223]_  = A302 & ~A299;
  assign \new_[11224]_  = A298 & \new_[11223]_ ;
  assign \new_[11225]_  = \new_[11224]_  & \new_[11219]_ ;
  assign \new_[11228]_  = A167 & A168;
  assign \new_[11232]_  = ~A201 & A200;
  assign \new_[11233]_  = A199 & \new_[11232]_ ;
  assign \new_[11234]_  = \new_[11233]_  & \new_[11228]_ ;
  assign \new_[11238]_  = A234 & A233;
  assign \new_[11239]_  = ~A202 & \new_[11238]_ ;
  assign \new_[11243]_  = A302 & A299;
  assign \new_[11244]_  = ~A298 & \new_[11243]_ ;
  assign \new_[11245]_  = \new_[11244]_  & \new_[11239]_ ;
  assign \new_[11248]_  = A167 & A168;
  assign \new_[11252]_  = ~A201 & A200;
  assign \new_[11253]_  = A199 & \new_[11252]_ ;
  assign \new_[11254]_  = \new_[11253]_  & \new_[11248]_ ;
  assign \new_[11258]_  = A234 & A233;
  assign \new_[11259]_  = ~A202 & \new_[11258]_ ;
  assign \new_[11263]_  = A269 & A266;
  assign \new_[11264]_  = ~A265 & \new_[11263]_ ;
  assign \new_[11265]_  = \new_[11264]_  & \new_[11259]_ ;
  assign \new_[11268]_  = A167 & A168;
  assign \new_[11272]_  = ~A201 & A200;
  assign \new_[11273]_  = A199 & \new_[11272]_ ;
  assign \new_[11274]_  = \new_[11273]_  & \new_[11268]_ ;
  assign \new_[11278]_  = A234 & A233;
  assign \new_[11279]_  = ~A202 & \new_[11278]_ ;
  assign \new_[11283]_  = A269 & ~A266;
  assign \new_[11284]_  = A265 & \new_[11283]_ ;
  assign \new_[11285]_  = \new_[11284]_  & \new_[11279]_ ;
  assign \new_[11288]_  = A167 & A168;
  assign \new_[11292]_  = ~A201 & A200;
  assign \new_[11293]_  = A199 & \new_[11292]_ ;
  assign \new_[11294]_  = \new_[11293]_  & \new_[11288]_ ;
  assign \new_[11298]_  = A233 & ~A232;
  assign \new_[11299]_  = ~A202 & \new_[11298]_ ;
  assign \new_[11303]_  = A300 & A299;
  assign \new_[11304]_  = A236 & \new_[11303]_ ;
  assign \new_[11305]_  = \new_[11304]_  & \new_[11299]_ ;
  assign \new_[11308]_  = A167 & A168;
  assign \new_[11312]_  = ~A201 & A200;
  assign \new_[11313]_  = A199 & \new_[11312]_ ;
  assign \new_[11314]_  = \new_[11313]_  & \new_[11308]_ ;
  assign \new_[11318]_  = A233 & ~A232;
  assign \new_[11319]_  = ~A202 & \new_[11318]_ ;
  assign \new_[11323]_  = A300 & A298;
  assign \new_[11324]_  = A236 & \new_[11323]_ ;
  assign \new_[11325]_  = \new_[11324]_  & \new_[11319]_ ;
  assign \new_[11328]_  = A167 & A168;
  assign \new_[11332]_  = ~A201 & A200;
  assign \new_[11333]_  = A199 & \new_[11332]_ ;
  assign \new_[11334]_  = \new_[11333]_  & \new_[11328]_ ;
  assign \new_[11338]_  = A233 & ~A232;
  assign \new_[11339]_  = ~A202 & \new_[11338]_ ;
  assign \new_[11343]_  = A267 & A265;
  assign \new_[11344]_  = A236 & \new_[11343]_ ;
  assign \new_[11345]_  = \new_[11344]_  & \new_[11339]_ ;
  assign \new_[11348]_  = A167 & A168;
  assign \new_[11352]_  = ~A201 & A200;
  assign \new_[11353]_  = A199 & \new_[11352]_ ;
  assign \new_[11354]_  = \new_[11353]_  & \new_[11348]_ ;
  assign \new_[11358]_  = A233 & ~A232;
  assign \new_[11359]_  = ~A202 & \new_[11358]_ ;
  assign \new_[11363]_  = A267 & A266;
  assign \new_[11364]_  = A236 & \new_[11363]_ ;
  assign \new_[11365]_  = \new_[11364]_  & \new_[11359]_ ;
  assign \new_[11368]_  = A167 & A168;
  assign \new_[11372]_  = ~A201 & A200;
  assign \new_[11373]_  = A199 & \new_[11372]_ ;
  assign \new_[11374]_  = \new_[11373]_  & \new_[11368]_ ;
  assign \new_[11378]_  = ~A233 & A232;
  assign \new_[11379]_  = ~A202 & \new_[11378]_ ;
  assign \new_[11383]_  = A300 & A299;
  assign \new_[11384]_  = A236 & \new_[11383]_ ;
  assign \new_[11385]_  = \new_[11384]_  & \new_[11379]_ ;
  assign \new_[11388]_  = A167 & A168;
  assign \new_[11392]_  = ~A201 & A200;
  assign \new_[11393]_  = A199 & \new_[11392]_ ;
  assign \new_[11394]_  = \new_[11393]_  & \new_[11388]_ ;
  assign \new_[11398]_  = ~A233 & A232;
  assign \new_[11399]_  = ~A202 & \new_[11398]_ ;
  assign \new_[11403]_  = A300 & A298;
  assign \new_[11404]_  = A236 & \new_[11403]_ ;
  assign \new_[11405]_  = \new_[11404]_  & \new_[11399]_ ;
  assign \new_[11408]_  = A167 & A168;
  assign \new_[11412]_  = ~A201 & A200;
  assign \new_[11413]_  = A199 & \new_[11412]_ ;
  assign \new_[11414]_  = \new_[11413]_  & \new_[11408]_ ;
  assign \new_[11418]_  = ~A233 & A232;
  assign \new_[11419]_  = ~A202 & \new_[11418]_ ;
  assign \new_[11423]_  = A267 & A265;
  assign \new_[11424]_  = A236 & \new_[11423]_ ;
  assign \new_[11425]_  = \new_[11424]_  & \new_[11419]_ ;
  assign \new_[11428]_  = A167 & A168;
  assign \new_[11432]_  = ~A201 & A200;
  assign \new_[11433]_  = A199 & \new_[11432]_ ;
  assign \new_[11434]_  = \new_[11433]_  & \new_[11428]_ ;
  assign \new_[11438]_  = ~A233 & A232;
  assign \new_[11439]_  = ~A202 & \new_[11438]_ ;
  assign \new_[11443]_  = A267 & A266;
  assign \new_[11444]_  = A236 & \new_[11443]_ ;
  assign \new_[11445]_  = \new_[11444]_  & \new_[11439]_ ;
  assign \new_[11448]_  = A167 & A168;
  assign \new_[11452]_  = ~A202 & ~A200;
  assign \new_[11453]_  = ~A199 & \new_[11452]_ ;
  assign \new_[11454]_  = \new_[11453]_  & \new_[11448]_ ;
  assign \new_[11458]_  = A236 & A233;
  assign \new_[11459]_  = ~A232 & \new_[11458]_ ;
  assign \new_[11463]_  = A302 & ~A299;
  assign \new_[11464]_  = A298 & \new_[11463]_ ;
  assign \new_[11465]_  = \new_[11464]_  & \new_[11459]_ ;
  assign \new_[11468]_  = A167 & A168;
  assign \new_[11472]_  = ~A202 & ~A200;
  assign \new_[11473]_  = ~A199 & \new_[11472]_ ;
  assign \new_[11474]_  = \new_[11473]_  & \new_[11468]_ ;
  assign \new_[11478]_  = A236 & A233;
  assign \new_[11479]_  = ~A232 & \new_[11478]_ ;
  assign \new_[11483]_  = A302 & A299;
  assign \new_[11484]_  = ~A298 & \new_[11483]_ ;
  assign \new_[11485]_  = \new_[11484]_  & \new_[11479]_ ;
  assign \new_[11488]_  = A167 & A168;
  assign \new_[11492]_  = ~A202 & ~A200;
  assign \new_[11493]_  = ~A199 & \new_[11492]_ ;
  assign \new_[11494]_  = \new_[11493]_  & \new_[11488]_ ;
  assign \new_[11498]_  = A236 & A233;
  assign \new_[11499]_  = ~A232 & \new_[11498]_ ;
  assign \new_[11503]_  = A269 & A266;
  assign \new_[11504]_  = ~A265 & \new_[11503]_ ;
  assign \new_[11505]_  = \new_[11504]_  & \new_[11499]_ ;
  assign \new_[11508]_  = A167 & A168;
  assign \new_[11512]_  = ~A202 & ~A200;
  assign \new_[11513]_  = ~A199 & \new_[11512]_ ;
  assign \new_[11514]_  = \new_[11513]_  & \new_[11508]_ ;
  assign \new_[11518]_  = A236 & A233;
  assign \new_[11519]_  = ~A232 & \new_[11518]_ ;
  assign \new_[11523]_  = A269 & ~A266;
  assign \new_[11524]_  = A265 & \new_[11523]_ ;
  assign \new_[11525]_  = \new_[11524]_  & \new_[11519]_ ;
  assign \new_[11528]_  = A167 & A168;
  assign \new_[11532]_  = ~A202 & ~A200;
  assign \new_[11533]_  = ~A199 & \new_[11532]_ ;
  assign \new_[11534]_  = \new_[11533]_  & \new_[11528]_ ;
  assign \new_[11538]_  = A236 & ~A233;
  assign \new_[11539]_  = A232 & \new_[11538]_ ;
  assign \new_[11543]_  = A302 & ~A299;
  assign \new_[11544]_  = A298 & \new_[11543]_ ;
  assign \new_[11545]_  = \new_[11544]_  & \new_[11539]_ ;
  assign \new_[11548]_  = A167 & A168;
  assign \new_[11552]_  = ~A202 & ~A200;
  assign \new_[11553]_  = ~A199 & \new_[11552]_ ;
  assign \new_[11554]_  = \new_[11553]_  & \new_[11548]_ ;
  assign \new_[11558]_  = A236 & ~A233;
  assign \new_[11559]_  = A232 & \new_[11558]_ ;
  assign \new_[11563]_  = A302 & A299;
  assign \new_[11564]_  = ~A298 & \new_[11563]_ ;
  assign \new_[11565]_  = \new_[11564]_  & \new_[11559]_ ;
  assign \new_[11568]_  = A167 & A168;
  assign \new_[11572]_  = ~A202 & ~A200;
  assign \new_[11573]_  = ~A199 & \new_[11572]_ ;
  assign \new_[11574]_  = \new_[11573]_  & \new_[11568]_ ;
  assign \new_[11578]_  = A236 & ~A233;
  assign \new_[11579]_  = A232 & \new_[11578]_ ;
  assign \new_[11583]_  = A269 & A266;
  assign \new_[11584]_  = ~A265 & \new_[11583]_ ;
  assign \new_[11585]_  = \new_[11584]_  & \new_[11579]_ ;
  assign \new_[11588]_  = A167 & A168;
  assign \new_[11592]_  = ~A202 & ~A200;
  assign \new_[11593]_  = ~A199 & \new_[11592]_ ;
  assign \new_[11594]_  = \new_[11593]_  & \new_[11588]_ ;
  assign \new_[11598]_  = A236 & ~A233;
  assign \new_[11599]_  = A232 & \new_[11598]_ ;
  assign \new_[11603]_  = A269 & ~A266;
  assign \new_[11604]_  = A265 & \new_[11603]_ ;
  assign \new_[11605]_  = \new_[11604]_  & \new_[11599]_ ;
  assign \new_[11608]_  = A167 & A170;
  assign \new_[11612]_  = ~A202 & ~A201;
  assign \new_[11613]_  = ~A166 & \new_[11612]_ ;
  assign \new_[11614]_  = \new_[11613]_  & \new_[11608]_ ;
  assign \new_[11618]_  = A234 & A232;
  assign \new_[11619]_  = ~A203 & \new_[11618]_ ;
  assign \new_[11623]_  = A302 & ~A299;
  assign \new_[11624]_  = A298 & \new_[11623]_ ;
  assign \new_[11625]_  = \new_[11624]_  & \new_[11619]_ ;
  assign \new_[11628]_  = A167 & A170;
  assign \new_[11632]_  = ~A202 & ~A201;
  assign \new_[11633]_  = ~A166 & \new_[11632]_ ;
  assign \new_[11634]_  = \new_[11633]_  & \new_[11628]_ ;
  assign \new_[11638]_  = A234 & A232;
  assign \new_[11639]_  = ~A203 & \new_[11638]_ ;
  assign \new_[11643]_  = A302 & A299;
  assign \new_[11644]_  = ~A298 & \new_[11643]_ ;
  assign \new_[11645]_  = \new_[11644]_  & \new_[11639]_ ;
  assign \new_[11648]_  = A167 & A170;
  assign \new_[11652]_  = ~A202 & ~A201;
  assign \new_[11653]_  = ~A166 & \new_[11652]_ ;
  assign \new_[11654]_  = \new_[11653]_  & \new_[11648]_ ;
  assign \new_[11658]_  = A234 & A232;
  assign \new_[11659]_  = ~A203 & \new_[11658]_ ;
  assign \new_[11663]_  = A269 & A266;
  assign \new_[11664]_  = ~A265 & \new_[11663]_ ;
  assign \new_[11665]_  = \new_[11664]_  & \new_[11659]_ ;
  assign \new_[11668]_  = A167 & A170;
  assign \new_[11672]_  = ~A202 & ~A201;
  assign \new_[11673]_  = ~A166 & \new_[11672]_ ;
  assign \new_[11674]_  = \new_[11673]_  & \new_[11668]_ ;
  assign \new_[11678]_  = A234 & A232;
  assign \new_[11679]_  = ~A203 & \new_[11678]_ ;
  assign \new_[11683]_  = A269 & ~A266;
  assign \new_[11684]_  = A265 & \new_[11683]_ ;
  assign \new_[11685]_  = \new_[11684]_  & \new_[11679]_ ;
  assign \new_[11688]_  = A167 & A170;
  assign \new_[11692]_  = ~A202 & ~A201;
  assign \new_[11693]_  = ~A166 & \new_[11692]_ ;
  assign \new_[11694]_  = \new_[11693]_  & \new_[11688]_ ;
  assign \new_[11698]_  = A234 & A233;
  assign \new_[11699]_  = ~A203 & \new_[11698]_ ;
  assign \new_[11703]_  = A302 & ~A299;
  assign \new_[11704]_  = A298 & \new_[11703]_ ;
  assign \new_[11705]_  = \new_[11704]_  & \new_[11699]_ ;
  assign \new_[11708]_  = A167 & A170;
  assign \new_[11712]_  = ~A202 & ~A201;
  assign \new_[11713]_  = ~A166 & \new_[11712]_ ;
  assign \new_[11714]_  = \new_[11713]_  & \new_[11708]_ ;
  assign \new_[11718]_  = A234 & A233;
  assign \new_[11719]_  = ~A203 & \new_[11718]_ ;
  assign \new_[11723]_  = A302 & A299;
  assign \new_[11724]_  = ~A298 & \new_[11723]_ ;
  assign \new_[11725]_  = \new_[11724]_  & \new_[11719]_ ;
  assign \new_[11728]_  = A167 & A170;
  assign \new_[11732]_  = ~A202 & ~A201;
  assign \new_[11733]_  = ~A166 & \new_[11732]_ ;
  assign \new_[11734]_  = \new_[11733]_  & \new_[11728]_ ;
  assign \new_[11738]_  = A234 & A233;
  assign \new_[11739]_  = ~A203 & \new_[11738]_ ;
  assign \new_[11743]_  = A269 & A266;
  assign \new_[11744]_  = ~A265 & \new_[11743]_ ;
  assign \new_[11745]_  = \new_[11744]_  & \new_[11739]_ ;
  assign \new_[11748]_  = A167 & A170;
  assign \new_[11752]_  = ~A202 & ~A201;
  assign \new_[11753]_  = ~A166 & \new_[11752]_ ;
  assign \new_[11754]_  = \new_[11753]_  & \new_[11748]_ ;
  assign \new_[11758]_  = A234 & A233;
  assign \new_[11759]_  = ~A203 & \new_[11758]_ ;
  assign \new_[11763]_  = A269 & ~A266;
  assign \new_[11764]_  = A265 & \new_[11763]_ ;
  assign \new_[11765]_  = \new_[11764]_  & \new_[11759]_ ;
  assign \new_[11768]_  = A167 & A170;
  assign \new_[11772]_  = ~A202 & ~A201;
  assign \new_[11773]_  = ~A166 & \new_[11772]_ ;
  assign \new_[11774]_  = \new_[11773]_  & \new_[11768]_ ;
  assign \new_[11778]_  = A233 & ~A232;
  assign \new_[11779]_  = ~A203 & \new_[11778]_ ;
  assign \new_[11783]_  = A300 & A299;
  assign \new_[11784]_  = A236 & \new_[11783]_ ;
  assign \new_[11785]_  = \new_[11784]_  & \new_[11779]_ ;
  assign \new_[11788]_  = A167 & A170;
  assign \new_[11792]_  = ~A202 & ~A201;
  assign \new_[11793]_  = ~A166 & \new_[11792]_ ;
  assign \new_[11794]_  = \new_[11793]_  & \new_[11788]_ ;
  assign \new_[11798]_  = A233 & ~A232;
  assign \new_[11799]_  = ~A203 & \new_[11798]_ ;
  assign \new_[11803]_  = A300 & A298;
  assign \new_[11804]_  = A236 & \new_[11803]_ ;
  assign \new_[11805]_  = \new_[11804]_  & \new_[11799]_ ;
  assign \new_[11808]_  = A167 & A170;
  assign \new_[11812]_  = ~A202 & ~A201;
  assign \new_[11813]_  = ~A166 & \new_[11812]_ ;
  assign \new_[11814]_  = \new_[11813]_  & \new_[11808]_ ;
  assign \new_[11818]_  = A233 & ~A232;
  assign \new_[11819]_  = ~A203 & \new_[11818]_ ;
  assign \new_[11823]_  = A267 & A265;
  assign \new_[11824]_  = A236 & \new_[11823]_ ;
  assign \new_[11825]_  = \new_[11824]_  & \new_[11819]_ ;
  assign \new_[11828]_  = A167 & A170;
  assign \new_[11832]_  = ~A202 & ~A201;
  assign \new_[11833]_  = ~A166 & \new_[11832]_ ;
  assign \new_[11834]_  = \new_[11833]_  & \new_[11828]_ ;
  assign \new_[11838]_  = A233 & ~A232;
  assign \new_[11839]_  = ~A203 & \new_[11838]_ ;
  assign \new_[11843]_  = A267 & A266;
  assign \new_[11844]_  = A236 & \new_[11843]_ ;
  assign \new_[11845]_  = \new_[11844]_  & \new_[11839]_ ;
  assign \new_[11848]_  = A167 & A170;
  assign \new_[11852]_  = ~A202 & ~A201;
  assign \new_[11853]_  = ~A166 & \new_[11852]_ ;
  assign \new_[11854]_  = \new_[11853]_  & \new_[11848]_ ;
  assign \new_[11858]_  = ~A233 & A232;
  assign \new_[11859]_  = ~A203 & \new_[11858]_ ;
  assign \new_[11863]_  = A300 & A299;
  assign \new_[11864]_  = A236 & \new_[11863]_ ;
  assign \new_[11865]_  = \new_[11864]_  & \new_[11859]_ ;
  assign \new_[11868]_  = A167 & A170;
  assign \new_[11872]_  = ~A202 & ~A201;
  assign \new_[11873]_  = ~A166 & \new_[11872]_ ;
  assign \new_[11874]_  = \new_[11873]_  & \new_[11868]_ ;
  assign \new_[11878]_  = ~A233 & A232;
  assign \new_[11879]_  = ~A203 & \new_[11878]_ ;
  assign \new_[11883]_  = A300 & A298;
  assign \new_[11884]_  = A236 & \new_[11883]_ ;
  assign \new_[11885]_  = \new_[11884]_  & \new_[11879]_ ;
  assign \new_[11888]_  = A167 & A170;
  assign \new_[11892]_  = ~A202 & ~A201;
  assign \new_[11893]_  = ~A166 & \new_[11892]_ ;
  assign \new_[11894]_  = \new_[11893]_  & \new_[11888]_ ;
  assign \new_[11898]_  = ~A233 & A232;
  assign \new_[11899]_  = ~A203 & \new_[11898]_ ;
  assign \new_[11903]_  = A267 & A265;
  assign \new_[11904]_  = A236 & \new_[11903]_ ;
  assign \new_[11905]_  = \new_[11904]_  & \new_[11899]_ ;
  assign \new_[11908]_  = A167 & A170;
  assign \new_[11912]_  = ~A202 & ~A201;
  assign \new_[11913]_  = ~A166 & \new_[11912]_ ;
  assign \new_[11914]_  = \new_[11913]_  & \new_[11908]_ ;
  assign \new_[11918]_  = ~A233 & A232;
  assign \new_[11919]_  = ~A203 & \new_[11918]_ ;
  assign \new_[11923]_  = A267 & A266;
  assign \new_[11924]_  = A236 & \new_[11923]_ ;
  assign \new_[11925]_  = \new_[11924]_  & \new_[11919]_ ;
  assign \new_[11928]_  = A167 & A170;
  assign \new_[11932]_  = A200 & A199;
  assign \new_[11933]_  = ~A166 & \new_[11932]_ ;
  assign \new_[11934]_  = \new_[11933]_  & \new_[11928]_ ;
  assign \new_[11938]_  = A235 & ~A202;
  assign \new_[11939]_  = ~A201 & \new_[11938]_ ;
  assign \new_[11943]_  = A302 & ~A299;
  assign \new_[11944]_  = A298 & \new_[11943]_ ;
  assign \new_[11945]_  = \new_[11944]_  & \new_[11939]_ ;
  assign \new_[11948]_  = A167 & A170;
  assign \new_[11952]_  = A200 & A199;
  assign \new_[11953]_  = ~A166 & \new_[11952]_ ;
  assign \new_[11954]_  = \new_[11953]_  & \new_[11948]_ ;
  assign \new_[11958]_  = A235 & ~A202;
  assign \new_[11959]_  = ~A201 & \new_[11958]_ ;
  assign \new_[11963]_  = A302 & A299;
  assign \new_[11964]_  = ~A298 & \new_[11963]_ ;
  assign \new_[11965]_  = \new_[11964]_  & \new_[11959]_ ;
  assign \new_[11968]_  = A167 & A170;
  assign \new_[11972]_  = A200 & A199;
  assign \new_[11973]_  = ~A166 & \new_[11972]_ ;
  assign \new_[11974]_  = \new_[11973]_  & \new_[11968]_ ;
  assign \new_[11978]_  = A235 & ~A202;
  assign \new_[11979]_  = ~A201 & \new_[11978]_ ;
  assign \new_[11983]_  = A269 & A266;
  assign \new_[11984]_  = ~A265 & \new_[11983]_ ;
  assign \new_[11985]_  = \new_[11984]_  & \new_[11979]_ ;
  assign \new_[11988]_  = A167 & A170;
  assign \new_[11992]_  = A200 & A199;
  assign \new_[11993]_  = ~A166 & \new_[11992]_ ;
  assign \new_[11994]_  = \new_[11993]_  & \new_[11988]_ ;
  assign \new_[11998]_  = A235 & ~A202;
  assign \new_[11999]_  = ~A201 & \new_[11998]_ ;
  assign \new_[12003]_  = A269 & ~A266;
  assign \new_[12004]_  = A265 & \new_[12003]_ ;
  assign \new_[12005]_  = \new_[12004]_  & \new_[11999]_ ;
  assign \new_[12008]_  = A167 & A170;
  assign \new_[12012]_  = A200 & A199;
  assign \new_[12013]_  = ~A166 & \new_[12012]_ ;
  assign \new_[12014]_  = \new_[12013]_  & \new_[12008]_ ;
  assign \new_[12018]_  = A232 & ~A202;
  assign \new_[12019]_  = ~A201 & \new_[12018]_ ;
  assign \new_[12023]_  = A300 & A299;
  assign \new_[12024]_  = A234 & \new_[12023]_ ;
  assign \new_[12025]_  = \new_[12024]_  & \new_[12019]_ ;
  assign \new_[12028]_  = A167 & A170;
  assign \new_[12032]_  = A200 & A199;
  assign \new_[12033]_  = ~A166 & \new_[12032]_ ;
  assign \new_[12034]_  = \new_[12033]_  & \new_[12028]_ ;
  assign \new_[12038]_  = A232 & ~A202;
  assign \new_[12039]_  = ~A201 & \new_[12038]_ ;
  assign \new_[12043]_  = A300 & A298;
  assign \new_[12044]_  = A234 & \new_[12043]_ ;
  assign \new_[12045]_  = \new_[12044]_  & \new_[12039]_ ;
  assign \new_[12048]_  = A167 & A170;
  assign \new_[12052]_  = A200 & A199;
  assign \new_[12053]_  = ~A166 & \new_[12052]_ ;
  assign \new_[12054]_  = \new_[12053]_  & \new_[12048]_ ;
  assign \new_[12058]_  = A232 & ~A202;
  assign \new_[12059]_  = ~A201 & \new_[12058]_ ;
  assign \new_[12063]_  = A267 & A265;
  assign \new_[12064]_  = A234 & \new_[12063]_ ;
  assign \new_[12065]_  = \new_[12064]_  & \new_[12059]_ ;
  assign \new_[12068]_  = A167 & A170;
  assign \new_[12072]_  = A200 & A199;
  assign \new_[12073]_  = ~A166 & \new_[12072]_ ;
  assign \new_[12074]_  = \new_[12073]_  & \new_[12068]_ ;
  assign \new_[12078]_  = A232 & ~A202;
  assign \new_[12079]_  = ~A201 & \new_[12078]_ ;
  assign \new_[12083]_  = A267 & A266;
  assign \new_[12084]_  = A234 & \new_[12083]_ ;
  assign \new_[12085]_  = \new_[12084]_  & \new_[12079]_ ;
  assign \new_[12088]_  = A167 & A170;
  assign \new_[12092]_  = A200 & A199;
  assign \new_[12093]_  = ~A166 & \new_[12092]_ ;
  assign \new_[12094]_  = \new_[12093]_  & \new_[12088]_ ;
  assign \new_[12098]_  = A233 & ~A202;
  assign \new_[12099]_  = ~A201 & \new_[12098]_ ;
  assign \new_[12103]_  = A300 & A299;
  assign \new_[12104]_  = A234 & \new_[12103]_ ;
  assign \new_[12105]_  = \new_[12104]_  & \new_[12099]_ ;
  assign \new_[12108]_  = A167 & A170;
  assign \new_[12112]_  = A200 & A199;
  assign \new_[12113]_  = ~A166 & \new_[12112]_ ;
  assign \new_[12114]_  = \new_[12113]_  & \new_[12108]_ ;
  assign \new_[12118]_  = A233 & ~A202;
  assign \new_[12119]_  = ~A201 & \new_[12118]_ ;
  assign \new_[12123]_  = A300 & A298;
  assign \new_[12124]_  = A234 & \new_[12123]_ ;
  assign \new_[12125]_  = \new_[12124]_  & \new_[12119]_ ;
  assign \new_[12128]_  = A167 & A170;
  assign \new_[12132]_  = A200 & A199;
  assign \new_[12133]_  = ~A166 & \new_[12132]_ ;
  assign \new_[12134]_  = \new_[12133]_  & \new_[12128]_ ;
  assign \new_[12138]_  = A233 & ~A202;
  assign \new_[12139]_  = ~A201 & \new_[12138]_ ;
  assign \new_[12143]_  = A267 & A265;
  assign \new_[12144]_  = A234 & \new_[12143]_ ;
  assign \new_[12145]_  = \new_[12144]_  & \new_[12139]_ ;
  assign \new_[12148]_  = A167 & A170;
  assign \new_[12152]_  = A200 & A199;
  assign \new_[12153]_  = ~A166 & \new_[12152]_ ;
  assign \new_[12154]_  = \new_[12153]_  & \new_[12148]_ ;
  assign \new_[12158]_  = A233 & ~A202;
  assign \new_[12159]_  = ~A201 & \new_[12158]_ ;
  assign \new_[12163]_  = A267 & A266;
  assign \new_[12164]_  = A234 & \new_[12163]_ ;
  assign \new_[12165]_  = \new_[12164]_  & \new_[12159]_ ;
  assign \new_[12168]_  = A167 & A170;
  assign \new_[12172]_  = A200 & A199;
  assign \new_[12173]_  = ~A166 & \new_[12172]_ ;
  assign \new_[12174]_  = \new_[12173]_  & \new_[12168]_ ;
  assign \new_[12178]_  = ~A232 & ~A202;
  assign \new_[12179]_  = ~A201 & \new_[12178]_ ;
  assign \new_[12183]_  = A301 & A236;
  assign \new_[12184]_  = A233 & \new_[12183]_ ;
  assign \new_[12185]_  = \new_[12184]_  & \new_[12179]_ ;
  assign \new_[12188]_  = A167 & A170;
  assign \new_[12192]_  = A200 & A199;
  assign \new_[12193]_  = ~A166 & \new_[12192]_ ;
  assign \new_[12194]_  = \new_[12193]_  & \new_[12188]_ ;
  assign \new_[12198]_  = ~A232 & ~A202;
  assign \new_[12199]_  = ~A201 & \new_[12198]_ ;
  assign \new_[12203]_  = A268 & A236;
  assign \new_[12204]_  = A233 & \new_[12203]_ ;
  assign \new_[12205]_  = \new_[12204]_  & \new_[12199]_ ;
  assign \new_[12208]_  = A167 & A170;
  assign \new_[12212]_  = A200 & A199;
  assign \new_[12213]_  = ~A166 & \new_[12212]_ ;
  assign \new_[12214]_  = \new_[12213]_  & \new_[12208]_ ;
  assign \new_[12218]_  = A232 & ~A202;
  assign \new_[12219]_  = ~A201 & \new_[12218]_ ;
  assign \new_[12223]_  = A301 & A236;
  assign \new_[12224]_  = ~A233 & \new_[12223]_ ;
  assign \new_[12225]_  = \new_[12224]_  & \new_[12219]_ ;
  assign \new_[12228]_  = A167 & A170;
  assign \new_[12232]_  = A200 & A199;
  assign \new_[12233]_  = ~A166 & \new_[12232]_ ;
  assign \new_[12234]_  = \new_[12233]_  & \new_[12228]_ ;
  assign \new_[12238]_  = A232 & ~A202;
  assign \new_[12239]_  = ~A201 & \new_[12238]_ ;
  assign \new_[12243]_  = A268 & A236;
  assign \new_[12244]_  = ~A233 & \new_[12243]_ ;
  assign \new_[12245]_  = \new_[12244]_  & \new_[12239]_ ;
  assign \new_[12248]_  = A167 & A170;
  assign \new_[12252]_  = ~A200 & ~A199;
  assign \new_[12253]_  = ~A166 & \new_[12252]_ ;
  assign \new_[12254]_  = \new_[12253]_  & \new_[12248]_ ;
  assign \new_[12258]_  = A234 & A232;
  assign \new_[12259]_  = ~A202 & \new_[12258]_ ;
  assign \new_[12263]_  = A302 & ~A299;
  assign \new_[12264]_  = A298 & \new_[12263]_ ;
  assign \new_[12265]_  = \new_[12264]_  & \new_[12259]_ ;
  assign \new_[12268]_  = A167 & A170;
  assign \new_[12272]_  = ~A200 & ~A199;
  assign \new_[12273]_  = ~A166 & \new_[12272]_ ;
  assign \new_[12274]_  = \new_[12273]_  & \new_[12268]_ ;
  assign \new_[12278]_  = A234 & A232;
  assign \new_[12279]_  = ~A202 & \new_[12278]_ ;
  assign \new_[12283]_  = A302 & A299;
  assign \new_[12284]_  = ~A298 & \new_[12283]_ ;
  assign \new_[12285]_  = \new_[12284]_  & \new_[12279]_ ;
  assign \new_[12288]_  = A167 & A170;
  assign \new_[12292]_  = ~A200 & ~A199;
  assign \new_[12293]_  = ~A166 & \new_[12292]_ ;
  assign \new_[12294]_  = \new_[12293]_  & \new_[12288]_ ;
  assign \new_[12298]_  = A234 & A232;
  assign \new_[12299]_  = ~A202 & \new_[12298]_ ;
  assign \new_[12303]_  = A269 & A266;
  assign \new_[12304]_  = ~A265 & \new_[12303]_ ;
  assign \new_[12305]_  = \new_[12304]_  & \new_[12299]_ ;
  assign \new_[12308]_  = A167 & A170;
  assign \new_[12312]_  = ~A200 & ~A199;
  assign \new_[12313]_  = ~A166 & \new_[12312]_ ;
  assign \new_[12314]_  = \new_[12313]_  & \new_[12308]_ ;
  assign \new_[12318]_  = A234 & A232;
  assign \new_[12319]_  = ~A202 & \new_[12318]_ ;
  assign \new_[12323]_  = A269 & ~A266;
  assign \new_[12324]_  = A265 & \new_[12323]_ ;
  assign \new_[12325]_  = \new_[12324]_  & \new_[12319]_ ;
  assign \new_[12328]_  = A167 & A170;
  assign \new_[12332]_  = ~A200 & ~A199;
  assign \new_[12333]_  = ~A166 & \new_[12332]_ ;
  assign \new_[12334]_  = \new_[12333]_  & \new_[12328]_ ;
  assign \new_[12338]_  = A234 & A233;
  assign \new_[12339]_  = ~A202 & \new_[12338]_ ;
  assign \new_[12343]_  = A302 & ~A299;
  assign \new_[12344]_  = A298 & \new_[12343]_ ;
  assign \new_[12345]_  = \new_[12344]_  & \new_[12339]_ ;
  assign \new_[12348]_  = A167 & A170;
  assign \new_[12352]_  = ~A200 & ~A199;
  assign \new_[12353]_  = ~A166 & \new_[12352]_ ;
  assign \new_[12354]_  = \new_[12353]_  & \new_[12348]_ ;
  assign \new_[12358]_  = A234 & A233;
  assign \new_[12359]_  = ~A202 & \new_[12358]_ ;
  assign \new_[12363]_  = A302 & A299;
  assign \new_[12364]_  = ~A298 & \new_[12363]_ ;
  assign \new_[12365]_  = \new_[12364]_  & \new_[12359]_ ;
  assign \new_[12368]_  = A167 & A170;
  assign \new_[12372]_  = ~A200 & ~A199;
  assign \new_[12373]_  = ~A166 & \new_[12372]_ ;
  assign \new_[12374]_  = \new_[12373]_  & \new_[12368]_ ;
  assign \new_[12378]_  = A234 & A233;
  assign \new_[12379]_  = ~A202 & \new_[12378]_ ;
  assign \new_[12383]_  = A269 & A266;
  assign \new_[12384]_  = ~A265 & \new_[12383]_ ;
  assign \new_[12385]_  = \new_[12384]_  & \new_[12379]_ ;
  assign \new_[12388]_  = A167 & A170;
  assign \new_[12392]_  = ~A200 & ~A199;
  assign \new_[12393]_  = ~A166 & \new_[12392]_ ;
  assign \new_[12394]_  = \new_[12393]_  & \new_[12388]_ ;
  assign \new_[12398]_  = A234 & A233;
  assign \new_[12399]_  = ~A202 & \new_[12398]_ ;
  assign \new_[12403]_  = A269 & ~A266;
  assign \new_[12404]_  = A265 & \new_[12403]_ ;
  assign \new_[12405]_  = \new_[12404]_  & \new_[12399]_ ;
  assign \new_[12408]_  = A167 & A170;
  assign \new_[12412]_  = ~A200 & ~A199;
  assign \new_[12413]_  = ~A166 & \new_[12412]_ ;
  assign \new_[12414]_  = \new_[12413]_  & \new_[12408]_ ;
  assign \new_[12418]_  = A233 & ~A232;
  assign \new_[12419]_  = ~A202 & \new_[12418]_ ;
  assign \new_[12423]_  = A300 & A299;
  assign \new_[12424]_  = A236 & \new_[12423]_ ;
  assign \new_[12425]_  = \new_[12424]_  & \new_[12419]_ ;
  assign \new_[12428]_  = A167 & A170;
  assign \new_[12432]_  = ~A200 & ~A199;
  assign \new_[12433]_  = ~A166 & \new_[12432]_ ;
  assign \new_[12434]_  = \new_[12433]_  & \new_[12428]_ ;
  assign \new_[12438]_  = A233 & ~A232;
  assign \new_[12439]_  = ~A202 & \new_[12438]_ ;
  assign \new_[12443]_  = A300 & A298;
  assign \new_[12444]_  = A236 & \new_[12443]_ ;
  assign \new_[12445]_  = \new_[12444]_  & \new_[12439]_ ;
  assign \new_[12448]_  = A167 & A170;
  assign \new_[12452]_  = ~A200 & ~A199;
  assign \new_[12453]_  = ~A166 & \new_[12452]_ ;
  assign \new_[12454]_  = \new_[12453]_  & \new_[12448]_ ;
  assign \new_[12458]_  = A233 & ~A232;
  assign \new_[12459]_  = ~A202 & \new_[12458]_ ;
  assign \new_[12463]_  = A267 & A265;
  assign \new_[12464]_  = A236 & \new_[12463]_ ;
  assign \new_[12465]_  = \new_[12464]_  & \new_[12459]_ ;
  assign \new_[12468]_  = A167 & A170;
  assign \new_[12472]_  = ~A200 & ~A199;
  assign \new_[12473]_  = ~A166 & \new_[12472]_ ;
  assign \new_[12474]_  = \new_[12473]_  & \new_[12468]_ ;
  assign \new_[12478]_  = A233 & ~A232;
  assign \new_[12479]_  = ~A202 & \new_[12478]_ ;
  assign \new_[12483]_  = A267 & A266;
  assign \new_[12484]_  = A236 & \new_[12483]_ ;
  assign \new_[12485]_  = \new_[12484]_  & \new_[12479]_ ;
  assign \new_[12488]_  = A167 & A170;
  assign \new_[12492]_  = ~A200 & ~A199;
  assign \new_[12493]_  = ~A166 & \new_[12492]_ ;
  assign \new_[12494]_  = \new_[12493]_  & \new_[12488]_ ;
  assign \new_[12498]_  = ~A233 & A232;
  assign \new_[12499]_  = ~A202 & \new_[12498]_ ;
  assign \new_[12503]_  = A300 & A299;
  assign \new_[12504]_  = A236 & \new_[12503]_ ;
  assign \new_[12505]_  = \new_[12504]_  & \new_[12499]_ ;
  assign \new_[12508]_  = A167 & A170;
  assign \new_[12512]_  = ~A200 & ~A199;
  assign \new_[12513]_  = ~A166 & \new_[12512]_ ;
  assign \new_[12514]_  = \new_[12513]_  & \new_[12508]_ ;
  assign \new_[12518]_  = ~A233 & A232;
  assign \new_[12519]_  = ~A202 & \new_[12518]_ ;
  assign \new_[12523]_  = A300 & A298;
  assign \new_[12524]_  = A236 & \new_[12523]_ ;
  assign \new_[12525]_  = \new_[12524]_  & \new_[12519]_ ;
  assign \new_[12528]_  = A167 & A170;
  assign \new_[12532]_  = ~A200 & ~A199;
  assign \new_[12533]_  = ~A166 & \new_[12532]_ ;
  assign \new_[12534]_  = \new_[12533]_  & \new_[12528]_ ;
  assign \new_[12538]_  = ~A233 & A232;
  assign \new_[12539]_  = ~A202 & \new_[12538]_ ;
  assign \new_[12543]_  = A267 & A265;
  assign \new_[12544]_  = A236 & \new_[12543]_ ;
  assign \new_[12545]_  = \new_[12544]_  & \new_[12539]_ ;
  assign \new_[12548]_  = A167 & A170;
  assign \new_[12552]_  = ~A200 & ~A199;
  assign \new_[12553]_  = ~A166 & \new_[12552]_ ;
  assign \new_[12554]_  = \new_[12553]_  & \new_[12548]_ ;
  assign \new_[12558]_  = ~A233 & A232;
  assign \new_[12559]_  = ~A202 & \new_[12558]_ ;
  assign \new_[12563]_  = A267 & A266;
  assign \new_[12564]_  = A236 & \new_[12563]_ ;
  assign \new_[12565]_  = \new_[12564]_  & \new_[12559]_ ;
  assign \new_[12568]_  = ~A167 & A170;
  assign \new_[12572]_  = ~A202 & ~A201;
  assign \new_[12573]_  = A166 & \new_[12572]_ ;
  assign \new_[12574]_  = \new_[12573]_  & \new_[12568]_ ;
  assign \new_[12578]_  = A234 & A232;
  assign \new_[12579]_  = ~A203 & \new_[12578]_ ;
  assign \new_[12583]_  = A302 & ~A299;
  assign \new_[12584]_  = A298 & \new_[12583]_ ;
  assign \new_[12585]_  = \new_[12584]_  & \new_[12579]_ ;
  assign \new_[12588]_  = ~A167 & A170;
  assign \new_[12592]_  = ~A202 & ~A201;
  assign \new_[12593]_  = A166 & \new_[12592]_ ;
  assign \new_[12594]_  = \new_[12593]_  & \new_[12588]_ ;
  assign \new_[12598]_  = A234 & A232;
  assign \new_[12599]_  = ~A203 & \new_[12598]_ ;
  assign \new_[12603]_  = A302 & A299;
  assign \new_[12604]_  = ~A298 & \new_[12603]_ ;
  assign \new_[12605]_  = \new_[12604]_  & \new_[12599]_ ;
  assign \new_[12608]_  = ~A167 & A170;
  assign \new_[12612]_  = ~A202 & ~A201;
  assign \new_[12613]_  = A166 & \new_[12612]_ ;
  assign \new_[12614]_  = \new_[12613]_  & \new_[12608]_ ;
  assign \new_[12618]_  = A234 & A232;
  assign \new_[12619]_  = ~A203 & \new_[12618]_ ;
  assign \new_[12623]_  = A269 & A266;
  assign \new_[12624]_  = ~A265 & \new_[12623]_ ;
  assign \new_[12625]_  = \new_[12624]_  & \new_[12619]_ ;
  assign \new_[12628]_  = ~A167 & A170;
  assign \new_[12632]_  = ~A202 & ~A201;
  assign \new_[12633]_  = A166 & \new_[12632]_ ;
  assign \new_[12634]_  = \new_[12633]_  & \new_[12628]_ ;
  assign \new_[12638]_  = A234 & A232;
  assign \new_[12639]_  = ~A203 & \new_[12638]_ ;
  assign \new_[12643]_  = A269 & ~A266;
  assign \new_[12644]_  = A265 & \new_[12643]_ ;
  assign \new_[12645]_  = \new_[12644]_  & \new_[12639]_ ;
  assign \new_[12648]_  = ~A167 & A170;
  assign \new_[12652]_  = ~A202 & ~A201;
  assign \new_[12653]_  = A166 & \new_[12652]_ ;
  assign \new_[12654]_  = \new_[12653]_  & \new_[12648]_ ;
  assign \new_[12658]_  = A234 & A233;
  assign \new_[12659]_  = ~A203 & \new_[12658]_ ;
  assign \new_[12663]_  = A302 & ~A299;
  assign \new_[12664]_  = A298 & \new_[12663]_ ;
  assign \new_[12665]_  = \new_[12664]_  & \new_[12659]_ ;
  assign \new_[12668]_  = ~A167 & A170;
  assign \new_[12672]_  = ~A202 & ~A201;
  assign \new_[12673]_  = A166 & \new_[12672]_ ;
  assign \new_[12674]_  = \new_[12673]_  & \new_[12668]_ ;
  assign \new_[12678]_  = A234 & A233;
  assign \new_[12679]_  = ~A203 & \new_[12678]_ ;
  assign \new_[12683]_  = A302 & A299;
  assign \new_[12684]_  = ~A298 & \new_[12683]_ ;
  assign \new_[12685]_  = \new_[12684]_  & \new_[12679]_ ;
  assign \new_[12688]_  = ~A167 & A170;
  assign \new_[12692]_  = ~A202 & ~A201;
  assign \new_[12693]_  = A166 & \new_[12692]_ ;
  assign \new_[12694]_  = \new_[12693]_  & \new_[12688]_ ;
  assign \new_[12698]_  = A234 & A233;
  assign \new_[12699]_  = ~A203 & \new_[12698]_ ;
  assign \new_[12703]_  = A269 & A266;
  assign \new_[12704]_  = ~A265 & \new_[12703]_ ;
  assign \new_[12705]_  = \new_[12704]_  & \new_[12699]_ ;
  assign \new_[12708]_  = ~A167 & A170;
  assign \new_[12712]_  = ~A202 & ~A201;
  assign \new_[12713]_  = A166 & \new_[12712]_ ;
  assign \new_[12714]_  = \new_[12713]_  & \new_[12708]_ ;
  assign \new_[12718]_  = A234 & A233;
  assign \new_[12719]_  = ~A203 & \new_[12718]_ ;
  assign \new_[12723]_  = A269 & ~A266;
  assign \new_[12724]_  = A265 & \new_[12723]_ ;
  assign \new_[12725]_  = \new_[12724]_  & \new_[12719]_ ;
  assign \new_[12728]_  = ~A167 & A170;
  assign \new_[12732]_  = ~A202 & ~A201;
  assign \new_[12733]_  = A166 & \new_[12732]_ ;
  assign \new_[12734]_  = \new_[12733]_  & \new_[12728]_ ;
  assign \new_[12738]_  = A233 & ~A232;
  assign \new_[12739]_  = ~A203 & \new_[12738]_ ;
  assign \new_[12743]_  = A300 & A299;
  assign \new_[12744]_  = A236 & \new_[12743]_ ;
  assign \new_[12745]_  = \new_[12744]_  & \new_[12739]_ ;
  assign \new_[12748]_  = ~A167 & A170;
  assign \new_[12752]_  = ~A202 & ~A201;
  assign \new_[12753]_  = A166 & \new_[12752]_ ;
  assign \new_[12754]_  = \new_[12753]_  & \new_[12748]_ ;
  assign \new_[12758]_  = A233 & ~A232;
  assign \new_[12759]_  = ~A203 & \new_[12758]_ ;
  assign \new_[12763]_  = A300 & A298;
  assign \new_[12764]_  = A236 & \new_[12763]_ ;
  assign \new_[12765]_  = \new_[12764]_  & \new_[12759]_ ;
  assign \new_[12768]_  = ~A167 & A170;
  assign \new_[12772]_  = ~A202 & ~A201;
  assign \new_[12773]_  = A166 & \new_[12772]_ ;
  assign \new_[12774]_  = \new_[12773]_  & \new_[12768]_ ;
  assign \new_[12778]_  = A233 & ~A232;
  assign \new_[12779]_  = ~A203 & \new_[12778]_ ;
  assign \new_[12783]_  = A267 & A265;
  assign \new_[12784]_  = A236 & \new_[12783]_ ;
  assign \new_[12785]_  = \new_[12784]_  & \new_[12779]_ ;
  assign \new_[12788]_  = ~A167 & A170;
  assign \new_[12792]_  = ~A202 & ~A201;
  assign \new_[12793]_  = A166 & \new_[12792]_ ;
  assign \new_[12794]_  = \new_[12793]_  & \new_[12788]_ ;
  assign \new_[12798]_  = A233 & ~A232;
  assign \new_[12799]_  = ~A203 & \new_[12798]_ ;
  assign \new_[12803]_  = A267 & A266;
  assign \new_[12804]_  = A236 & \new_[12803]_ ;
  assign \new_[12805]_  = \new_[12804]_  & \new_[12799]_ ;
  assign \new_[12808]_  = ~A167 & A170;
  assign \new_[12812]_  = ~A202 & ~A201;
  assign \new_[12813]_  = A166 & \new_[12812]_ ;
  assign \new_[12814]_  = \new_[12813]_  & \new_[12808]_ ;
  assign \new_[12818]_  = ~A233 & A232;
  assign \new_[12819]_  = ~A203 & \new_[12818]_ ;
  assign \new_[12823]_  = A300 & A299;
  assign \new_[12824]_  = A236 & \new_[12823]_ ;
  assign \new_[12825]_  = \new_[12824]_  & \new_[12819]_ ;
  assign \new_[12828]_  = ~A167 & A170;
  assign \new_[12832]_  = ~A202 & ~A201;
  assign \new_[12833]_  = A166 & \new_[12832]_ ;
  assign \new_[12834]_  = \new_[12833]_  & \new_[12828]_ ;
  assign \new_[12838]_  = ~A233 & A232;
  assign \new_[12839]_  = ~A203 & \new_[12838]_ ;
  assign \new_[12843]_  = A300 & A298;
  assign \new_[12844]_  = A236 & \new_[12843]_ ;
  assign \new_[12845]_  = \new_[12844]_  & \new_[12839]_ ;
  assign \new_[12848]_  = ~A167 & A170;
  assign \new_[12852]_  = ~A202 & ~A201;
  assign \new_[12853]_  = A166 & \new_[12852]_ ;
  assign \new_[12854]_  = \new_[12853]_  & \new_[12848]_ ;
  assign \new_[12858]_  = ~A233 & A232;
  assign \new_[12859]_  = ~A203 & \new_[12858]_ ;
  assign \new_[12863]_  = A267 & A265;
  assign \new_[12864]_  = A236 & \new_[12863]_ ;
  assign \new_[12865]_  = \new_[12864]_  & \new_[12859]_ ;
  assign \new_[12868]_  = ~A167 & A170;
  assign \new_[12872]_  = ~A202 & ~A201;
  assign \new_[12873]_  = A166 & \new_[12872]_ ;
  assign \new_[12874]_  = \new_[12873]_  & \new_[12868]_ ;
  assign \new_[12878]_  = ~A233 & A232;
  assign \new_[12879]_  = ~A203 & \new_[12878]_ ;
  assign \new_[12883]_  = A267 & A266;
  assign \new_[12884]_  = A236 & \new_[12883]_ ;
  assign \new_[12885]_  = \new_[12884]_  & \new_[12879]_ ;
  assign \new_[12888]_  = ~A167 & A170;
  assign \new_[12892]_  = A200 & A199;
  assign \new_[12893]_  = A166 & \new_[12892]_ ;
  assign \new_[12894]_  = \new_[12893]_  & \new_[12888]_ ;
  assign \new_[12898]_  = A235 & ~A202;
  assign \new_[12899]_  = ~A201 & \new_[12898]_ ;
  assign \new_[12903]_  = A302 & ~A299;
  assign \new_[12904]_  = A298 & \new_[12903]_ ;
  assign \new_[12905]_  = \new_[12904]_  & \new_[12899]_ ;
  assign \new_[12908]_  = ~A167 & A170;
  assign \new_[12912]_  = A200 & A199;
  assign \new_[12913]_  = A166 & \new_[12912]_ ;
  assign \new_[12914]_  = \new_[12913]_  & \new_[12908]_ ;
  assign \new_[12918]_  = A235 & ~A202;
  assign \new_[12919]_  = ~A201 & \new_[12918]_ ;
  assign \new_[12923]_  = A302 & A299;
  assign \new_[12924]_  = ~A298 & \new_[12923]_ ;
  assign \new_[12925]_  = \new_[12924]_  & \new_[12919]_ ;
  assign \new_[12928]_  = ~A167 & A170;
  assign \new_[12932]_  = A200 & A199;
  assign \new_[12933]_  = A166 & \new_[12932]_ ;
  assign \new_[12934]_  = \new_[12933]_  & \new_[12928]_ ;
  assign \new_[12938]_  = A235 & ~A202;
  assign \new_[12939]_  = ~A201 & \new_[12938]_ ;
  assign \new_[12943]_  = A269 & A266;
  assign \new_[12944]_  = ~A265 & \new_[12943]_ ;
  assign \new_[12945]_  = \new_[12944]_  & \new_[12939]_ ;
  assign \new_[12948]_  = ~A167 & A170;
  assign \new_[12952]_  = A200 & A199;
  assign \new_[12953]_  = A166 & \new_[12952]_ ;
  assign \new_[12954]_  = \new_[12953]_  & \new_[12948]_ ;
  assign \new_[12958]_  = A235 & ~A202;
  assign \new_[12959]_  = ~A201 & \new_[12958]_ ;
  assign \new_[12963]_  = A269 & ~A266;
  assign \new_[12964]_  = A265 & \new_[12963]_ ;
  assign \new_[12965]_  = \new_[12964]_  & \new_[12959]_ ;
  assign \new_[12968]_  = ~A167 & A170;
  assign \new_[12972]_  = A200 & A199;
  assign \new_[12973]_  = A166 & \new_[12972]_ ;
  assign \new_[12974]_  = \new_[12973]_  & \new_[12968]_ ;
  assign \new_[12978]_  = A232 & ~A202;
  assign \new_[12979]_  = ~A201 & \new_[12978]_ ;
  assign \new_[12983]_  = A300 & A299;
  assign \new_[12984]_  = A234 & \new_[12983]_ ;
  assign \new_[12985]_  = \new_[12984]_  & \new_[12979]_ ;
  assign \new_[12988]_  = ~A167 & A170;
  assign \new_[12992]_  = A200 & A199;
  assign \new_[12993]_  = A166 & \new_[12992]_ ;
  assign \new_[12994]_  = \new_[12993]_  & \new_[12988]_ ;
  assign \new_[12998]_  = A232 & ~A202;
  assign \new_[12999]_  = ~A201 & \new_[12998]_ ;
  assign \new_[13003]_  = A300 & A298;
  assign \new_[13004]_  = A234 & \new_[13003]_ ;
  assign \new_[13005]_  = \new_[13004]_  & \new_[12999]_ ;
  assign \new_[13008]_  = ~A167 & A170;
  assign \new_[13012]_  = A200 & A199;
  assign \new_[13013]_  = A166 & \new_[13012]_ ;
  assign \new_[13014]_  = \new_[13013]_  & \new_[13008]_ ;
  assign \new_[13018]_  = A232 & ~A202;
  assign \new_[13019]_  = ~A201 & \new_[13018]_ ;
  assign \new_[13023]_  = A267 & A265;
  assign \new_[13024]_  = A234 & \new_[13023]_ ;
  assign \new_[13025]_  = \new_[13024]_  & \new_[13019]_ ;
  assign \new_[13028]_  = ~A167 & A170;
  assign \new_[13032]_  = A200 & A199;
  assign \new_[13033]_  = A166 & \new_[13032]_ ;
  assign \new_[13034]_  = \new_[13033]_  & \new_[13028]_ ;
  assign \new_[13038]_  = A232 & ~A202;
  assign \new_[13039]_  = ~A201 & \new_[13038]_ ;
  assign \new_[13043]_  = A267 & A266;
  assign \new_[13044]_  = A234 & \new_[13043]_ ;
  assign \new_[13045]_  = \new_[13044]_  & \new_[13039]_ ;
  assign \new_[13048]_  = ~A167 & A170;
  assign \new_[13052]_  = A200 & A199;
  assign \new_[13053]_  = A166 & \new_[13052]_ ;
  assign \new_[13054]_  = \new_[13053]_  & \new_[13048]_ ;
  assign \new_[13058]_  = A233 & ~A202;
  assign \new_[13059]_  = ~A201 & \new_[13058]_ ;
  assign \new_[13063]_  = A300 & A299;
  assign \new_[13064]_  = A234 & \new_[13063]_ ;
  assign \new_[13065]_  = \new_[13064]_  & \new_[13059]_ ;
  assign \new_[13068]_  = ~A167 & A170;
  assign \new_[13072]_  = A200 & A199;
  assign \new_[13073]_  = A166 & \new_[13072]_ ;
  assign \new_[13074]_  = \new_[13073]_  & \new_[13068]_ ;
  assign \new_[13078]_  = A233 & ~A202;
  assign \new_[13079]_  = ~A201 & \new_[13078]_ ;
  assign \new_[13083]_  = A300 & A298;
  assign \new_[13084]_  = A234 & \new_[13083]_ ;
  assign \new_[13085]_  = \new_[13084]_  & \new_[13079]_ ;
  assign \new_[13088]_  = ~A167 & A170;
  assign \new_[13092]_  = A200 & A199;
  assign \new_[13093]_  = A166 & \new_[13092]_ ;
  assign \new_[13094]_  = \new_[13093]_  & \new_[13088]_ ;
  assign \new_[13098]_  = A233 & ~A202;
  assign \new_[13099]_  = ~A201 & \new_[13098]_ ;
  assign \new_[13103]_  = A267 & A265;
  assign \new_[13104]_  = A234 & \new_[13103]_ ;
  assign \new_[13105]_  = \new_[13104]_  & \new_[13099]_ ;
  assign \new_[13108]_  = ~A167 & A170;
  assign \new_[13112]_  = A200 & A199;
  assign \new_[13113]_  = A166 & \new_[13112]_ ;
  assign \new_[13114]_  = \new_[13113]_  & \new_[13108]_ ;
  assign \new_[13118]_  = A233 & ~A202;
  assign \new_[13119]_  = ~A201 & \new_[13118]_ ;
  assign \new_[13123]_  = A267 & A266;
  assign \new_[13124]_  = A234 & \new_[13123]_ ;
  assign \new_[13125]_  = \new_[13124]_  & \new_[13119]_ ;
  assign \new_[13128]_  = ~A167 & A170;
  assign \new_[13132]_  = A200 & A199;
  assign \new_[13133]_  = A166 & \new_[13132]_ ;
  assign \new_[13134]_  = \new_[13133]_  & \new_[13128]_ ;
  assign \new_[13138]_  = ~A232 & ~A202;
  assign \new_[13139]_  = ~A201 & \new_[13138]_ ;
  assign \new_[13143]_  = A301 & A236;
  assign \new_[13144]_  = A233 & \new_[13143]_ ;
  assign \new_[13145]_  = \new_[13144]_  & \new_[13139]_ ;
  assign \new_[13148]_  = ~A167 & A170;
  assign \new_[13152]_  = A200 & A199;
  assign \new_[13153]_  = A166 & \new_[13152]_ ;
  assign \new_[13154]_  = \new_[13153]_  & \new_[13148]_ ;
  assign \new_[13158]_  = ~A232 & ~A202;
  assign \new_[13159]_  = ~A201 & \new_[13158]_ ;
  assign \new_[13163]_  = A268 & A236;
  assign \new_[13164]_  = A233 & \new_[13163]_ ;
  assign \new_[13165]_  = \new_[13164]_  & \new_[13159]_ ;
  assign \new_[13168]_  = ~A167 & A170;
  assign \new_[13172]_  = A200 & A199;
  assign \new_[13173]_  = A166 & \new_[13172]_ ;
  assign \new_[13174]_  = \new_[13173]_  & \new_[13168]_ ;
  assign \new_[13178]_  = A232 & ~A202;
  assign \new_[13179]_  = ~A201 & \new_[13178]_ ;
  assign \new_[13183]_  = A301 & A236;
  assign \new_[13184]_  = ~A233 & \new_[13183]_ ;
  assign \new_[13185]_  = \new_[13184]_  & \new_[13179]_ ;
  assign \new_[13188]_  = ~A167 & A170;
  assign \new_[13192]_  = A200 & A199;
  assign \new_[13193]_  = A166 & \new_[13192]_ ;
  assign \new_[13194]_  = \new_[13193]_  & \new_[13188]_ ;
  assign \new_[13198]_  = A232 & ~A202;
  assign \new_[13199]_  = ~A201 & \new_[13198]_ ;
  assign \new_[13203]_  = A268 & A236;
  assign \new_[13204]_  = ~A233 & \new_[13203]_ ;
  assign \new_[13205]_  = \new_[13204]_  & \new_[13199]_ ;
  assign \new_[13208]_  = ~A167 & A170;
  assign \new_[13212]_  = ~A200 & ~A199;
  assign \new_[13213]_  = A166 & \new_[13212]_ ;
  assign \new_[13214]_  = \new_[13213]_  & \new_[13208]_ ;
  assign \new_[13218]_  = A234 & A232;
  assign \new_[13219]_  = ~A202 & \new_[13218]_ ;
  assign \new_[13223]_  = A302 & ~A299;
  assign \new_[13224]_  = A298 & \new_[13223]_ ;
  assign \new_[13225]_  = \new_[13224]_  & \new_[13219]_ ;
  assign \new_[13228]_  = ~A167 & A170;
  assign \new_[13232]_  = ~A200 & ~A199;
  assign \new_[13233]_  = A166 & \new_[13232]_ ;
  assign \new_[13234]_  = \new_[13233]_  & \new_[13228]_ ;
  assign \new_[13238]_  = A234 & A232;
  assign \new_[13239]_  = ~A202 & \new_[13238]_ ;
  assign \new_[13243]_  = A302 & A299;
  assign \new_[13244]_  = ~A298 & \new_[13243]_ ;
  assign \new_[13245]_  = \new_[13244]_  & \new_[13239]_ ;
  assign \new_[13248]_  = ~A167 & A170;
  assign \new_[13252]_  = ~A200 & ~A199;
  assign \new_[13253]_  = A166 & \new_[13252]_ ;
  assign \new_[13254]_  = \new_[13253]_  & \new_[13248]_ ;
  assign \new_[13258]_  = A234 & A232;
  assign \new_[13259]_  = ~A202 & \new_[13258]_ ;
  assign \new_[13263]_  = A269 & A266;
  assign \new_[13264]_  = ~A265 & \new_[13263]_ ;
  assign \new_[13265]_  = \new_[13264]_  & \new_[13259]_ ;
  assign \new_[13268]_  = ~A167 & A170;
  assign \new_[13272]_  = ~A200 & ~A199;
  assign \new_[13273]_  = A166 & \new_[13272]_ ;
  assign \new_[13274]_  = \new_[13273]_  & \new_[13268]_ ;
  assign \new_[13278]_  = A234 & A232;
  assign \new_[13279]_  = ~A202 & \new_[13278]_ ;
  assign \new_[13283]_  = A269 & ~A266;
  assign \new_[13284]_  = A265 & \new_[13283]_ ;
  assign \new_[13285]_  = \new_[13284]_  & \new_[13279]_ ;
  assign \new_[13288]_  = ~A167 & A170;
  assign \new_[13292]_  = ~A200 & ~A199;
  assign \new_[13293]_  = A166 & \new_[13292]_ ;
  assign \new_[13294]_  = \new_[13293]_  & \new_[13288]_ ;
  assign \new_[13298]_  = A234 & A233;
  assign \new_[13299]_  = ~A202 & \new_[13298]_ ;
  assign \new_[13303]_  = A302 & ~A299;
  assign \new_[13304]_  = A298 & \new_[13303]_ ;
  assign \new_[13305]_  = \new_[13304]_  & \new_[13299]_ ;
  assign \new_[13308]_  = ~A167 & A170;
  assign \new_[13312]_  = ~A200 & ~A199;
  assign \new_[13313]_  = A166 & \new_[13312]_ ;
  assign \new_[13314]_  = \new_[13313]_  & \new_[13308]_ ;
  assign \new_[13318]_  = A234 & A233;
  assign \new_[13319]_  = ~A202 & \new_[13318]_ ;
  assign \new_[13323]_  = A302 & A299;
  assign \new_[13324]_  = ~A298 & \new_[13323]_ ;
  assign \new_[13325]_  = \new_[13324]_  & \new_[13319]_ ;
  assign \new_[13328]_  = ~A167 & A170;
  assign \new_[13332]_  = ~A200 & ~A199;
  assign \new_[13333]_  = A166 & \new_[13332]_ ;
  assign \new_[13334]_  = \new_[13333]_  & \new_[13328]_ ;
  assign \new_[13338]_  = A234 & A233;
  assign \new_[13339]_  = ~A202 & \new_[13338]_ ;
  assign \new_[13343]_  = A269 & A266;
  assign \new_[13344]_  = ~A265 & \new_[13343]_ ;
  assign \new_[13345]_  = \new_[13344]_  & \new_[13339]_ ;
  assign \new_[13348]_  = ~A167 & A170;
  assign \new_[13352]_  = ~A200 & ~A199;
  assign \new_[13353]_  = A166 & \new_[13352]_ ;
  assign \new_[13354]_  = \new_[13353]_  & \new_[13348]_ ;
  assign \new_[13358]_  = A234 & A233;
  assign \new_[13359]_  = ~A202 & \new_[13358]_ ;
  assign \new_[13363]_  = A269 & ~A266;
  assign \new_[13364]_  = A265 & \new_[13363]_ ;
  assign \new_[13365]_  = \new_[13364]_  & \new_[13359]_ ;
  assign \new_[13368]_  = ~A167 & A170;
  assign \new_[13372]_  = ~A200 & ~A199;
  assign \new_[13373]_  = A166 & \new_[13372]_ ;
  assign \new_[13374]_  = \new_[13373]_  & \new_[13368]_ ;
  assign \new_[13378]_  = A233 & ~A232;
  assign \new_[13379]_  = ~A202 & \new_[13378]_ ;
  assign \new_[13383]_  = A300 & A299;
  assign \new_[13384]_  = A236 & \new_[13383]_ ;
  assign \new_[13385]_  = \new_[13384]_  & \new_[13379]_ ;
  assign \new_[13388]_  = ~A167 & A170;
  assign \new_[13392]_  = ~A200 & ~A199;
  assign \new_[13393]_  = A166 & \new_[13392]_ ;
  assign \new_[13394]_  = \new_[13393]_  & \new_[13388]_ ;
  assign \new_[13398]_  = A233 & ~A232;
  assign \new_[13399]_  = ~A202 & \new_[13398]_ ;
  assign \new_[13403]_  = A300 & A298;
  assign \new_[13404]_  = A236 & \new_[13403]_ ;
  assign \new_[13405]_  = \new_[13404]_  & \new_[13399]_ ;
  assign \new_[13408]_  = ~A167 & A170;
  assign \new_[13412]_  = ~A200 & ~A199;
  assign \new_[13413]_  = A166 & \new_[13412]_ ;
  assign \new_[13414]_  = \new_[13413]_  & \new_[13408]_ ;
  assign \new_[13418]_  = A233 & ~A232;
  assign \new_[13419]_  = ~A202 & \new_[13418]_ ;
  assign \new_[13423]_  = A267 & A265;
  assign \new_[13424]_  = A236 & \new_[13423]_ ;
  assign \new_[13425]_  = \new_[13424]_  & \new_[13419]_ ;
  assign \new_[13428]_  = ~A167 & A170;
  assign \new_[13432]_  = ~A200 & ~A199;
  assign \new_[13433]_  = A166 & \new_[13432]_ ;
  assign \new_[13434]_  = \new_[13433]_  & \new_[13428]_ ;
  assign \new_[13438]_  = A233 & ~A232;
  assign \new_[13439]_  = ~A202 & \new_[13438]_ ;
  assign \new_[13443]_  = A267 & A266;
  assign \new_[13444]_  = A236 & \new_[13443]_ ;
  assign \new_[13445]_  = \new_[13444]_  & \new_[13439]_ ;
  assign \new_[13448]_  = ~A167 & A170;
  assign \new_[13452]_  = ~A200 & ~A199;
  assign \new_[13453]_  = A166 & \new_[13452]_ ;
  assign \new_[13454]_  = \new_[13453]_  & \new_[13448]_ ;
  assign \new_[13458]_  = ~A233 & A232;
  assign \new_[13459]_  = ~A202 & \new_[13458]_ ;
  assign \new_[13463]_  = A300 & A299;
  assign \new_[13464]_  = A236 & \new_[13463]_ ;
  assign \new_[13465]_  = \new_[13464]_  & \new_[13459]_ ;
  assign \new_[13468]_  = ~A167 & A170;
  assign \new_[13472]_  = ~A200 & ~A199;
  assign \new_[13473]_  = A166 & \new_[13472]_ ;
  assign \new_[13474]_  = \new_[13473]_  & \new_[13468]_ ;
  assign \new_[13478]_  = ~A233 & A232;
  assign \new_[13479]_  = ~A202 & \new_[13478]_ ;
  assign \new_[13483]_  = A300 & A298;
  assign \new_[13484]_  = A236 & \new_[13483]_ ;
  assign \new_[13485]_  = \new_[13484]_  & \new_[13479]_ ;
  assign \new_[13488]_  = ~A167 & A170;
  assign \new_[13492]_  = ~A200 & ~A199;
  assign \new_[13493]_  = A166 & \new_[13492]_ ;
  assign \new_[13494]_  = \new_[13493]_  & \new_[13488]_ ;
  assign \new_[13498]_  = ~A233 & A232;
  assign \new_[13499]_  = ~A202 & \new_[13498]_ ;
  assign \new_[13503]_  = A267 & A265;
  assign \new_[13504]_  = A236 & \new_[13503]_ ;
  assign \new_[13505]_  = \new_[13504]_  & \new_[13499]_ ;
  assign \new_[13508]_  = ~A167 & A170;
  assign \new_[13512]_  = ~A200 & ~A199;
  assign \new_[13513]_  = A166 & \new_[13512]_ ;
  assign \new_[13514]_  = \new_[13513]_  & \new_[13508]_ ;
  assign \new_[13518]_  = ~A233 & A232;
  assign \new_[13519]_  = ~A202 & \new_[13518]_ ;
  assign \new_[13523]_  = A267 & A266;
  assign \new_[13524]_  = A236 & \new_[13523]_ ;
  assign \new_[13525]_  = \new_[13524]_  & \new_[13519]_ ;
  assign \new_[13528]_  = A199 & A169;
  assign \new_[13532]_  = ~A202 & ~A201;
  assign \new_[13533]_  = A200 & \new_[13532]_ ;
  assign \new_[13534]_  = \new_[13533]_  & \new_[13528]_ ;
  assign \new_[13538]_  = A236 & A233;
  assign \new_[13539]_  = ~A232 & \new_[13538]_ ;
  assign \new_[13543]_  = A302 & ~A299;
  assign \new_[13544]_  = A298 & \new_[13543]_ ;
  assign \new_[13545]_  = \new_[13544]_  & \new_[13539]_ ;
  assign \new_[13548]_  = A199 & A169;
  assign \new_[13552]_  = ~A202 & ~A201;
  assign \new_[13553]_  = A200 & \new_[13552]_ ;
  assign \new_[13554]_  = \new_[13553]_  & \new_[13548]_ ;
  assign \new_[13558]_  = A236 & A233;
  assign \new_[13559]_  = ~A232 & \new_[13558]_ ;
  assign \new_[13563]_  = A302 & A299;
  assign \new_[13564]_  = ~A298 & \new_[13563]_ ;
  assign \new_[13565]_  = \new_[13564]_  & \new_[13559]_ ;
  assign \new_[13568]_  = A199 & A169;
  assign \new_[13572]_  = ~A202 & ~A201;
  assign \new_[13573]_  = A200 & \new_[13572]_ ;
  assign \new_[13574]_  = \new_[13573]_  & \new_[13568]_ ;
  assign \new_[13578]_  = A236 & A233;
  assign \new_[13579]_  = ~A232 & \new_[13578]_ ;
  assign \new_[13583]_  = A269 & A266;
  assign \new_[13584]_  = ~A265 & \new_[13583]_ ;
  assign \new_[13585]_  = \new_[13584]_  & \new_[13579]_ ;
  assign \new_[13588]_  = A199 & A169;
  assign \new_[13592]_  = ~A202 & ~A201;
  assign \new_[13593]_  = A200 & \new_[13592]_ ;
  assign \new_[13594]_  = \new_[13593]_  & \new_[13588]_ ;
  assign \new_[13598]_  = A236 & A233;
  assign \new_[13599]_  = ~A232 & \new_[13598]_ ;
  assign \new_[13603]_  = A269 & ~A266;
  assign \new_[13604]_  = A265 & \new_[13603]_ ;
  assign \new_[13605]_  = \new_[13604]_  & \new_[13599]_ ;
  assign \new_[13608]_  = A199 & A169;
  assign \new_[13612]_  = ~A202 & ~A201;
  assign \new_[13613]_  = A200 & \new_[13612]_ ;
  assign \new_[13614]_  = \new_[13613]_  & \new_[13608]_ ;
  assign \new_[13618]_  = A236 & ~A233;
  assign \new_[13619]_  = A232 & \new_[13618]_ ;
  assign \new_[13623]_  = A302 & ~A299;
  assign \new_[13624]_  = A298 & \new_[13623]_ ;
  assign \new_[13625]_  = \new_[13624]_  & \new_[13619]_ ;
  assign \new_[13628]_  = A199 & A169;
  assign \new_[13632]_  = ~A202 & ~A201;
  assign \new_[13633]_  = A200 & \new_[13632]_ ;
  assign \new_[13634]_  = \new_[13633]_  & \new_[13628]_ ;
  assign \new_[13638]_  = A236 & ~A233;
  assign \new_[13639]_  = A232 & \new_[13638]_ ;
  assign \new_[13643]_  = A302 & A299;
  assign \new_[13644]_  = ~A298 & \new_[13643]_ ;
  assign \new_[13645]_  = \new_[13644]_  & \new_[13639]_ ;
  assign \new_[13648]_  = A199 & A169;
  assign \new_[13652]_  = ~A202 & ~A201;
  assign \new_[13653]_  = A200 & \new_[13652]_ ;
  assign \new_[13654]_  = \new_[13653]_  & \new_[13648]_ ;
  assign \new_[13658]_  = A236 & ~A233;
  assign \new_[13659]_  = A232 & \new_[13658]_ ;
  assign \new_[13663]_  = A269 & A266;
  assign \new_[13664]_  = ~A265 & \new_[13663]_ ;
  assign \new_[13665]_  = \new_[13664]_  & \new_[13659]_ ;
  assign \new_[13668]_  = A199 & A169;
  assign \new_[13672]_  = ~A202 & ~A201;
  assign \new_[13673]_  = A200 & \new_[13672]_ ;
  assign \new_[13674]_  = \new_[13673]_  & \new_[13668]_ ;
  assign \new_[13678]_  = A236 & ~A233;
  assign \new_[13679]_  = A232 & \new_[13678]_ ;
  assign \new_[13683]_  = A269 & ~A266;
  assign \new_[13684]_  = A265 & \new_[13683]_ ;
  assign \new_[13685]_  = \new_[13684]_  & \new_[13679]_ ;
  assign \new_[13689]_  = A199 & A166;
  assign \new_[13690]_  = A168 & \new_[13689]_ ;
  assign \new_[13694]_  = ~A202 & ~A201;
  assign \new_[13695]_  = A200 & \new_[13694]_ ;
  assign \new_[13696]_  = \new_[13695]_  & \new_[13690]_ ;
  assign \new_[13700]_  = A236 & A233;
  assign \new_[13701]_  = ~A232 & \new_[13700]_ ;
  assign \new_[13705]_  = A302 & ~A299;
  assign \new_[13706]_  = A298 & \new_[13705]_ ;
  assign \new_[13707]_  = \new_[13706]_  & \new_[13701]_ ;
  assign \new_[13711]_  = A199 & A166;
  assign \new_[13712]_  = A168 & \new_[13711]_ ;
  assign \new_[13716]_  = ~A202 & ~A201;
  assign \new_[13717]_  = A200 & \new_[13716]_ ;
  assign \new_[13718]_  = \new_[13717]_  & \new_[13712]_ ;
  assign \new_[13722]_  = A236 & A233;
  assign \new_[13723]_  = ~A232 & \new_[13722]_ ;
  assign \new_[13727]_  = A302 & A299;
  assign \new_[13728]_  = ~A298 & \new_[13727]_ ;
  assign \new_[13729]_  = \new_[13728]_  & \new_[13723]_ ;
  assign \new_[13733]_  = A199 & A166;
  assign \new_[13734]_  = A168 & \new_[13733]_ ;
  assign \new_[13738]_  = ~A202 & ~A201;
  assign \new_[13739]_  = A200 & \new_[13738]_ ;
  assign \new_[13740]_  = \new_[13739]_  & \new_[13734]_ ;
  assign \new_[13744]_  = A236 & A233;
  assign \new_[13745]_  = ~A232 & \new_[13744]_ ;
  assign \new_[13749]_  = A269 & A266;
  assign \new_[13750]_  = ~A265 & \new_[13749]_ ;
  assign \new_[13751]_  = \new_[13750]_  & \new_[13745]_ ;
  assign \new_[13755]_  = A199 & A166;
  assign \new_[13756]_  = A168 & \new_[13755]_ ;
  assign \new_[13760]_  = ~A202 & ~A201;
  assign \new_[13761]_  = A200 & \new_[13760]_ ;
  assign \new_[13762]_  = \new_[13761]_  & \new_[13756]_ ;
  assign \new_[13766]_  = A236 & A233;
  assign \new_[13767]_  = ~A232 & \new_[13766]_ ;
  assign \new_[13771]_  = A269 & ~A266;
  assign \new_[13772]_  = A265 & \new_[13771]_ ;
  assign \new_[13773]_  = \new_[13772]_  & \new_[13767]_ ;
  assign \new_[13777]_  = A199 & A166;
  assign \new_[13778]_  = A168 & \new_[13777]_ ;
  assign \new_[13782]_  = ~A202 & ~A201;
  assign \new_[13783]_  = A200 & \new_[13782]_ ;
  assign \new_[13784]_  = \new_[13783]_  & \new_[13778]_ ;
  assign \new_[13788]_  = A236 & ~A233;
  assign \new_[13789]_  = A232 & \new_[13788]_ ;
  assign \new_[13793]_  = A302 & ~A299;
  assign \new_[13794]_  = A298 & \new_[13793]_ ;
  assign \new_[13795]_  = \new_[13794]_  & \new_[13789]_ ;
  assign \new_[13799]_  = A199 & A166;
  assign \new_[13800]_  = A168 & \new_[13799]_ ;
  assign \new_[13804]_  = ~A202 & ~A201;
  assign \new_[13805]_  = A200 & \new_[13804]_ ;
  assign \new_[13806]_  = \new_[13805]_  & \new_[13800]_ ;
  assign \new_[13810]_  = A236 & ~A233;
  assign \new_[13811]_  = A232 & \new_[13810]_ ;
  assign \new_[13815]_  = A302 & A299;
  assign \new_[13816]_  = ~A298 & \new_[13815]_ ;
  assign \new_[13817]_  = \new_[13816]_  & \new_[13811]_ ;
  assign \new_[13821]_  = A199 & A166;
  assign \new_[13822]_  = A168 & \new_[13821]_ ;
  assign \new_[13826]_  = ~A202 & ~A201;
  assign \new_[13827]_  = A200 & \new_[13826]_ ;
  assign \new_[13828]_  = \new_[13827]_  & \new_[13822]_ ;
  assign \new_[13832]_  = A236 & ~A233;
  assign \new_[13833]_  = A232 & \new_[13832]_ ;
  assign \new_[13837]_  = A269 & A266;
  assign \new_[13838]_  = ~A265 & \new_[13837]_ ;
  assign \new_[13839]_  = \new_[13838]_  & \new_[13833]_ ;
  assign \new_[13843]_  = A199 & A166;
  assign \new_[13844]_  = A168 & \new_[13843]_ ;
  assign \new_[13848]_  = ~A202 & ~A201;
  assign \new_[13849]_  = A200 & \new_[13848]_ ;
  assign \new_[13850]_  = \new_[13849]_  & \new_[13844]_ ;
  assign \new_[13854]_  = A236 & ~A233;
  assign \new_[13855]_  = A232 & \new_[13854]_ ;
  assign \new_[13859]_  = A269 & ~A266;
  assign \new_[13860]_  = A265 & \new_[13859]_ ;
  assign \new_[13861]_  = \new_[13860]_  & \new_[13855]_ ;
  assign \new_[13865]_  = A199 & A167;
  assign \new_[13866]_  = A168 & \new_[13865]_ ;
  assign \new_[13870]_  = ~A202 & ~A201;
  assign \new_[13871]_  = A200 & \new_[13870]_ ;
  assign \new_[13872]_  = \new_[13871]_  & \new_[13866]_ ;
  assign \new_[13876]_  = A236 & A233;
  assign \new_[13877]_  = ~A232 & \new_[13876]_ ;
  assign \new_[13881]_  = A302 & ~A299;
  assign \new_[13882]_  = A298 & \new_[13881]_ ;
  assign \new_[13883]_  = \new_[13882]_  & \new_[13877]_ ;
  assign \new_[13887]_  = A199 & A167;
  assign \new_[13888]_  = A168 & \new_[13887]_ ;
  assign \new_[13892]_  = ~A202 & ~A201;
  assign \new_[13893]_  = A200 & \new_[13892]_ ;
  assign \new_[13894]_  = \new_[13893]_  & \new_[13888]_ ;
  assign \new_[13898]_  = A236 & A233;
  assign \new_[13899]_  = ~A232 & \new_[13898]_ ;
  assign \new_[13903]_  = A302 & A299;
  assign \new_[13904]_  = ~A298 & \new_[13903]_ ;
  assign \new_[13905]_  = \new_[13904]_  & \new_[13899]_ ;
  assign \new_[13909]_  = A199 & A167;
  assign \new_[13910]_  = A168 & \new_[13909]_ ;
  assign \new_[13914]_  = ~A202 & ~A201;
  assign \new_[13915]_  = A200 & \new_[13914]_ ;
  assign \new_[13916]_  = \new_[13915]_  & \new_[13910]_ ;
  assign \new_[13920]_  = A236 & A233;
  assign \new_[13921]_  = ~A232 & \new_[13920]_ ;
  assign \new_[13925]_  = A269 & A266;
  assign \new_[13926]_  = ~A265 & \new_[13925]_ ;
  assign \new_[13927]_  = \new_[13926]_  & \new_[13921]_ ;
  assign \new_[13931]_  = A199 & A167;
  assign \new_[13932]_  = A168 & \new_[13931]_ ;
  assign \new_[13936]_  = ~A202 & ~A201;
  assign \new_[13937]_  = A200 & \new_[13936]_ ;
  assign \new_[13938]_  = \new_[13937]_  & \new_[13932]_ ;
  assign \new_[13942]_  = A236 & A233;
  assign \new_[13943]_  = ~A232 & \new_[13942]_ ;
  assign \new_[13947]_  = A269 & ~A266;
  assign \new_[13948]_  = A265 & \new_[13947]_ ;
  assign \new_[13949]_  = \new_[13948]_  & \new_[13943]_ ;
  assign \new_[13953]_  = A199 & A167;
  assign \new_[13954]_  = A168 & \new_[13953]_ ;
  assign \new_[13958]_  = ~A202 & ~A201;
  assign \new_[13959]_  = A200 & \new_[13958]_ ;
  assign \new_[13960]_  = \new_[13959]_  & \new_[13954]_ ;
  assign \new_[13964]_  = A236 & ~A233;
  assign \new_[13965]_  = A232 & \new_[13964]_ ;
  assign \new_[13969]_  = A302 & ~A299;
  assign \new_[13970]_  = A298 & \new_[13969]_ ;
  assign \new_[13971]_  = \new_[13970]_  & \new_[13965]_ ;
  assign \new_[13975]_  = A199 & A167;
  assign \new_[13976]_  = A168 & \new_[13975]_ ;
  assign \new_[13980]_  = ~A202 & ~A201;
  assign \new_[13981]_  = A200 & \new_[13980]_ ;
  assign \new_[13982]_  = \new_[13981]_  & \new_[13976]_ ;
  assign \new_[13986]_  = A236 & ~A233;
  assign \new_[13987]_  = A232 & \new_[13986]_ ;
  assign \new_[13991]_  = A302 & A299;
  assign \new_[13992]_  = ~A298 & \new_[13991]_ ;
  assign \new_[13993]_  = \new_[13992]_  & \new_[13987]_ ;
  assign \new_[13997]_  = A199 & A167;
  assign \new_[13998]_  = A168 & \new_[13997]_ ;
  assign \new_[14002]_  = ~A202 & ~A201;
  assign \new_[14003]_  = A200 & \new_[14002]_ ;
  assign \new_[14004]_  = \new_[14003]_  & \new_[13998]_ ;
  assign \new_[14008]_  = A236 & ~A233;
  assign \new_[14009]_  = A232 & \new_[14008]_ ;
  assign \new_[14013]_  = A269 & A266;
  assign \new_[14014]_  = ~A265 & \new_[14013]_ ;
  assign \new_[14015]_  = \new_[14014]_  & \new_[14009]_ ;
  assign \new_[14019]_  = A199 & A167;
  assign \new_[14020]_  = A168 & \new_[14019]_ ;
  assign \new_[14024]_  = ~A202 & ~A201;
  assign \new_[14025]_  = A200 & \new_[14024]_ ;
  assign \new_[14026]_  = \new_[14025]_  & \new_[14020]_ ;
  assign \new_[14030]_  = A236 & ~A233;
  assign \new_[14031]_  = A232 & \new_[14030]_ ;
  assign \new_[14035]_  = A269 & ~A266;
  assign \new_[14036]_  = A265 & \new_[14035]_ ;
  assign \new_[14037]_  = \new_[14036]_  & \new_[14031]_ ;
  assign \new_[14041]_  = ~A166 & A167;
  assign \new_[14042]_  = A170 & \new_[14041]_ ;
  assign \new_[14046]_  = ~A203 & ~A202;
  assign \new_[14047]_  = ~A201 & \new_[14046]_ ;
  assign \new_[14048]_  = \new_[14047]_  & \new_[14042]_ ;
  assign \new_[14052]_  = A236 & A233;
  assign \new_[14053]_  = ~A232 & \new_[14052]_ ;
  assign \new_[14057]_  = A302 & ~A299;
  assign \new_[14058]_  = A298 & \new_[14057]_ ;
  assign \new_[14059]_  = \new_[14058]_  & \new_[14053]_ ;
  assign \new_[14063]_  = ~A166 & A167;
  assign \new_[14064]_  = A170 & \new_[14063]_ ;
  assign \new_[14068]_  = ~A203 & ~A202;
  assign \new_[14069]_  = ~A201 & \new_[14068]_ ;
  assign \new_[14070]_  = \new_[14069]_  & \new_[14064]_ ;
  assign \new_[14074]_  = A236 & A233;
  assign \new_[14075]_  = ~A232 & \new_[14074]_ ;
  assign \new_[14079]_  = A302 & A299;
  assign \new_[14080]_  = ~A298 & \new_[14079]_ ;
  assign \new_[14081]_  = \new_[14080]_  & \new_[14075]_ ;
  assign \new_[14085]_  = ~A166 & A167;
  assign \new_[14086]_  = A170 & \new_[14085]_ ;
  assign \new_[14090]_  = ~A203 & ~A202;
  assign \new_[14091]_  = ~A201 & \new_[14090]_ ;
  assign \new_[14092]_  = \new_[14091]_  & \new_[14086]_ ;
  assign \new_[14096]_  = A236 & A233;
  assign \new_[14097]_  = ~A232 & \new_[14096]_ ;
  assign \new_[14101]_  = A269 & A266;
  assign \new_[14102]_  = ~A265 & \new_[14101]_ ;
  assign \new_[14103]_  = \new_[14102]_  & \new_[14097]_ ;
  assign \new_[14107]_  = ~A166 & A167;
  assign \new_[14108]_  = A170 & \new_[14107]_ ;
  assign \new_[14112]_  = ~A203 & ~A202;
  assign \new_[14113]_  = ~A201 & \new_[14112]_ ;
  assign \new_[14114]_  = \new_[14113]_  & \new_[14108]_ ;
  assign \new_[14118]_  = A236 & A233;
  assign \new_[14119]_  = ~A232 & \new_[14118]_ ;
  assign \new_[14123]_  = A269 & ~A266;
  assign \new_[14124]_  = A265 & \new_[14123]_ ;
  assign \new_[14125]_  = \new_[14124]_  & \new_[14119]_ ;
  assign \new_[14129]_  = ~A166 & A167;
  assign \new_[14130]_  = A170 & \new_[14129]_ ;
  assign \new_[14134]_  = ~A203 & ~A202;
  assign \new_[14135]_  = ~A201 & \new_[14134]_ ;
  assign \new_[14136]_  = \new_[14135]_  & \new_[14130]_ ;
  assign \new_[14140]_  = A236 & ~A233;
  assign \new_[14141]_  = A232 & \new_[14140]_ ;
  assign \new_[14145]_  = A302 & ~A299;
  assign \new_[14146]_  = A298 & \new_[14145]_ ;
  assign \new_[14147]_  = \new_[14146]_  & \new_[14141]_ ;
  assign \new_[14151]_  = ~A166 & A167;
  assign \new_[14152]_  = A170 & \new_[14151]_ ;
  assign \new_[14156]_  = ~A203 & ~A202;
  assign \new_[14157]_  = ~A201 & \new_[14156]_ ;
  assign \new_[14158]_  = \new_[14157]_  & \new_[14152]_ ;
  assign \new_[14162]_  = A236 & ~A233;
  assign \new_[14163]_  = A232 & \new_[14162]_ ;
  assign \new_[14167]_  = A302 & A299;
  assign \new_[14168]_  = ~A298 & \new_[14167]_ ;
  assign \new_[14169]_  = \new_[14168]_  & \new_[14163]_ ;
  assign \new_[14173]_  = ~A166 & A167;
  assign \new_[14174]_  = A170 & \new_[14173]_ ;
  assign \new_[14178]_  = ~A203 & ~A202;
  assign \new_[14179]_  = ~A201 & \new_[14178]_ ;
  assign \new_[14180]_  = \new_[14179]_  & \new_[14174]_ ;
  assign \new_[14184]_  = A236 & ~A233;
  assign \new_[14185]_  = A232 & \new_[14184]_ ;
  assign \new_[14189]_  = A269 & A266;
  assign \new_[14190]_  = ~A265 & \new_[14189]_ ;
  assign \new_[14191]_  = \new_[14190]_  & \new_[14185]_ ;
  assign \new_[14195]_  = ~A166 & A167;
  assign \new_[14196]_  = A170 & \new_[14195]_ ;
  assign \new_[14200]_  = ~A203 & ~A202;
  assign \new_[14201]_  = ~A201 & \new_[14200]_ ;
  assign \new_[14202]_  = \new_[14201]_  & \new_[14196]_ ;
  assign \new_[14206]_  = A236 & ~A233;
  assign \new_[14207]_  = A232 & \new_[14206]_ ;
  assign \new_[14211]_  = A269 & ~A266;
  assign \new_[14212]_  = A265 & \new_[14211]_ ;
  assign \new_[14213]_  = \new_[14212]_  & \new_[14207]_ ;
  assign \new_[14217]_  = ~A166 & A167;
  assign \new_[14218]_  = A170 & \new_[14217]_ ;
  assign \new_[14222]_  = ~A201 & A200;
  assign \new_[14223]_  = A199 & \new_[14222]_ ;
  assign \new_[14224]_  = \new_[14223]_  & \new_[14218]_ ;
  assign \new_[14228]_  = A234 & A232;
  assign \new_[14229]_  = ~A202 & \new_[14228]_ ;
  assign \new_[14233]_  = A302 & ~A299;
  assign \new_[14234]_  = A298 & \new_[14233]_ ;
  assign \new_[14235]_  = \new_[14234]_  & \new_[14229]_ ;
  assign \new_[14239]_  = ~A166 & A167;
  assign \new_[14240]_  = A170 & \new_[14239]_ ;
  assign \new_[14244]_  = ~A201 & A200;
  assign \new_[14245]_  = A199 & \new_[14244]_ ;
  assign \new_[14246]_  = \new_[14245]_  & \new_[14240]_ ;
  assign \new_[14250]_  = A234 & A232;
  assign \new_[14251]_  = ~A202 & \new_[14250]_ ;
  assign \new_[14255]_  = A302 & A299;
  assign \new_[14256]_  = ~A298 & \new_[14255]_ ;
  assign \new_[14257]_  = \new_[14256]_  & \new_[14251]_ ;
  assign \new_[14261]_  = ~A166 & A167;
  assign \new_[14262]_  = A170 & \new_[14261]_ ;
  assign \new_[14266]_  = ~A201 & A200;
  assign \new_[14267]_  = A199 & \new_[14266]_ ;
  assign \new_[14268]_  = \new_[14267]_  & \new_[14262]_ ;
  assign \new_[14272]_  = A234 & A232;
  assign \new_[14273]_  = ~A202 & \new_[14272]_ ;
  assign \new_[14277]_  = A269 & A266;
  assign \new_[14278]_  = ~A265 & \new_[14277]_ ;
  assign \new_[14279]_  = \new_[14278]_  & \new_[14273]_ ;
  assign \new_[14283]_  = ~A166 & A167;
  assign \new_[14284]_  = A170 & \new_[14283]_ ;
  assign \new_[14288]_  = ~A201 & A200;
  assign \new_[14289]_  = A199 & \new_[14288]_ ;
  assign \new_[14290]_  = \new_[14289]_  & \new_[14284]_ ;
  assign \new_[14294]_  = A234 & A232;
  assign \new_[14295]_  = ~A202 & \new_[14294]_ ;
  assign \new_[14299]_  = A269 & ~A266;
  assign \new_[14300]_  = A265 & \new_[14299]_ ;
  assign \new_[14301]_  = \new_[14300]_  & \new_[14295]_ ;
  assign \new_[14305]_  = ~A166 & A167;
  assign \new_[14306]_  = A170 & \new_[14305]_ ;
  assign \new_[14310]_  = ~A201 & A200;
  assign \new_[14311]_  = A199 & \new_[14310]_ ;
  assign \new_[14312]_  = \new_[14311]_  & \new_[14306]_ ;
  assign \new_[14316]_  = A234 & A233;
  assign \new_[14317]_  = ~A202 & \new_[14316]_ ;
  assign \new_[14321]_  = A302 & ~A299;
  assign \new_[14322]_  = A298 & \new_[14321]_ ;
  assign \new_[14323]_  = \new_[14322]_  & \new_[14317]_ ;
  assign \new_[14327]_  = ~A166 & A167;
  assign \new_[14328]_  = A170 & \new_[14327]_ ;
  assign \new_[14332]_  = ~A201 & A200;
  assign \new_[14333]_  = A199 & \new_[14332]_ ;
  assign \new_[14334]_  = \new_[14333]_  & \new_[14328]_ ;
  assign \new_[14338]_  = A234 & A233;
  assign \new_[14339]_  = ~A202 & \new_[14338]_ ;
  assign \new_[14343]_  = A302 & A299;
  assign \new_[14344]_  = ~A298 & \new_[14343]_ ;
  assign \new_[14345]_  = \new_[14344]_  & \new_[14339]_ ;
  assign \new_[14349]_  = ~A166 & A167;
  assign \new_[14350]_  = A170 & \new_[14349]_ ;
  assign \new_[14354]_  = ~A201 & A200;
  assign \new_[14355]_  = A199 & \new_[14354]_ ;
  assign \new_[14356]_  = \new_[14355]_  & \new_[14350]_ ;
  assign \new_[14360]_  = A234 & A233;
  assign \new_[14361]_  = ~A202 & \new_[14360]_ ;
  assign \new_[14365]_  = A269 & A266;
  assign \new_[14366]_  = ~A265 & \new_[14365]_ ;
  assign \new_[14367]_  = \new_[14366]_  & \new_[14361]_ ;
  assign \new_[14371]_  = ~A166 & A167;
  assign \new_[14372]_  = A170 & \new_[14371]_ ;
  assign \new_[14376]_  = ~A201 & A200;
  assign \new_[14377]_  = A199 & \new_[14376]_ ;
  assign \new_[14378]_  = \new_[14377]_  & \new_[14372]_ ;
  assign \new_[14382]_  = A234 & A233;
  assign \new_[14383]_  = ~A202 & \new_[14382]_ ;
  assign \new_[14387]_  = A269 & ~A266;
  assign \new_[14388]_  = A265 & \new_[14387]_ ;
  assign \new_[14389]_  = \new_[14388]_  & \new_[14383]_ ;
  assign \new_[14393]_  = ~A166 & A167;
  assign \new_[14394]_  = A170 & \new_[14393]_ ;
  assign \new_[14398]_  = ~A201 & A200;
  assign \new_[14399]_  = A199 & \new_[14398]_ ;
  assign \new_[14400]_  = \new_[14399]_  & \new_[14394]_ ;
  assign \new_[14404]_  = A233 & ~A232;
  assign \new_[14405]_  = ~A202 & \new_[14404]_ ;
  assign \new_[14409]_  = A300 & A299;
  assign \new_[14410]_  = A236 & \new_[14409]_ ;
  assign \new_[14411]_  = \new_[14410]_  & \new_[14405]_ ;
  assign \new_[14415]_  = ~A166 & A167;
  assign \new_[14416]_  = A170 & \new_[14415]_ ;
  assign \new_[14420]_  = ~A201 & A200;
  assign \new_[14421]_  = A199 & \new_[14420]_ ;
  assign \new_[14422]_  = \new_[14421]_  & \new_[14416]_ ;
  assign \new_[14426]_  = A233 & ~A232;
  assign \new_[14427]_  = ~A202 & \new_[14426]_ ;
  assign \new_[14431]_  = A300 & A298;
  assign \new_[14432]_  = A236 & \new_[14431]_ ;
  assign \new_[14433]_  = \new_[14432]_  & \new_[14427]_ ;
  assign \new_[14437]_  = ~A166 & A167;
  assign \new_[14438]_  = A170 & \new_[14437]_ ;
  assign \new_[14442]_  = ~A201 & A200;
  assign \new_[14443]_  = A199 & \new_[14442]_ ;
  assign \new_[14444]_  = \new_[14443]_  & \new_[14438]_ ;
  assign \new_[14448]_  = A233 & ~A232;
  assign \new_[14449]_  = ~A202 & \new_[14448]_ ;
  assign \new_[14453]_  = A267 & A265;
  assign \new_[14454]_  = A236 & \new_[14453]_ ;
  assign \new_[14455]_  = \new_[14454]_  & \new_[14449]_ ;
  assign \new_[14459]_  = ~A166 & A167;
  assign \new_[14460]_  = A170 & \new_[14459]_ ;
  assign \new_[14464]_  = ~A201 & A200;
  assign \new_[14465]_  = A199 & \new_[14464]_ ;
  assign \new_[14466]_  = \new_[14465]_  & \new_[14460]_ ;
  assign \new_[14470]_  = A233 & ~A232;
  assign \new_[14471]_  = ~A202 & \new_[14470]_ ;
  assign \new_[14475]_  = A267 & A266;
  assign \new_[14476]_  = A236 & \new_[14475]_ ;
  assign \new_[14477]_  = \new_[14476]_  & \new_[14471]_ ;
  assign \new_[14481]_  = ~A166 & A167;
  assign \new_[14482]_  = A170 & \new_[14481]_ ;
  assign \new_[14486]_  = ~A201 & A200;
  assign \new_[14487]_  = A199 & \new_[14486]_ ;
  assign \new_[14488]_  = \new_[14487]_  & \new_[14482]_ ;
  assign \new_[14492]_  = ~A233 & A232;
  assign \new_[14493]_  = ~A202 & \new_[14492]_ ;
  assign \new_[14497]_  = A300 & A299;
  assign \new_[14498]_  = A236 & \new_[14497]_ ;
  assign \new_[14499]_  = \new_[14498]_  & \new_[14493]_ ;
  assign \new_[14503]_  = ~A166 & A167;
  assign \new_[14504]_  = A170 & \new_[14503]_ ;
  assign \new_[14508]_  = ~A201 & A200;
  assign \new_[14509]_  = A199 & \new_[14508]_ ;
  assign \new_[14510]_  = \new_[14509]_  & \new_[14504]_ ;
  assign \new_[14514]_  = ~A233 & A232;
  assign \new_[14515]_  = ~A202 & \new_[14514]_ ;
  assign \new_[14519]_  = A300 & A298;
  assign \new_[14520]_  = A236 & \new_[14519]_ ;
  assign \new_[14521]_  = \new_[14520]_  & \new_[14515]_ ;
  assign \new_[14525]_  = ~A166 & A167;
  assign \new_[14526]_  = A170 & \new_[14525]_ ;
  assign \new_[14530]_  = ~A201 & A200;
  assign \new_[14531]_  = A199 & \new_[14530]_ ;
  assign \new_[14532]_  = \new_[14531]_  & \new_[14526]_ ;
  assign \new_[14536]_  = ~A233 & A232;
  assign \new_[14537]_  = ~A202 & \new_[14536]_ ;
  assign \new_[14541]_  = A267 & A265;
  assign \new_[14542]_  = A236 & \new_[14541]_ ;
  assign \new_[14543]_  = \new_[14542]_  & \new_[14537]_ ;
  assign \new_[14547]_  = ~A166 & A167;
  assign \new_[14548]_  = A170 & \new_[14547]_ ;
  assign \new_[14552]_  = ~A201 & A200;
  assign \new_[14553]_  = A199 & \new_[14552]_ ;
  assign \new_[14554]_  = \new_[14553]_  & \new_[14548]_ ;
  assign \new_[14558]_  = ~A233 & A232;
  assign \new_[14559]_  = ~A202 & \new_[14558]_ ;
  assign \new_[14563]_  = A267 & A266;
  assign \new_[14564]_  = A236 & \new_[14563]_ ;
  assign \new_[14565]_  = \new_[14564]_  & \new_[14559]_ ;
  assign \new_[14569]_  = ~A166 & A167;
  assign \new_[14570]_  = A170 & \new_[14569]_ ;
  assign \new_[14574]_  = ~A202 & ~A200;
  assign \new_[14575]_  = ~A199 & \new_[14574]_ ;
  assign \new_[14576]_  = \new_[14575]_  & \new_[14570]_ ;
  assign \new_[14580]_  = A236 & A233;
  assign \new_[14581]_  = ~A232 & \new_[14580]_ ;
  assign \new_[14585]_  = A302 & ~A299;
  assign \new_[14586]_  = A298 & \new_[14585]_ ;
  assign \new_[14587]_  = \new_[14586]_  & \new_[14581]_ ;
  assign \new_[14591]_  = ~A166 & A167;
  assign \new_[14592]_  = A170 & \new_[14591]_ ;
  assign \new_[14596]_  = ~A202 & ~A200;
  assign \new_[14597]_  = ~A199 & \new_[14596]_ ;
  assign \new_[14598]_  = \new_[14597]_  & \new_[14592]_ ;
  assign \new_[14602]_  = A236 & A233;
  assign \new_[14603]_  = ~A232 & \new_[14602]_ ;
  assign \new_[14607]_  = A302 & A299;
  assign \new_[14608]_  = ~A298 & \new_[14607]_ ;
  assign \new_[14609]_  = \new_[14608]_  & \new_[14603]_ ;
  assign \new_[14613]_  = ~A166 & A167;
  assign \new_[14614]_  = A170 & \new_[14613]_ ;
  assign \new_[14618]_  = ~A202 & ~A200;
  assign \new_[14619]_  = ~A199 & \new_[14618]_ ;
  assign \new_[14620]_  = \new_[14619]_  & \new_[14614]_ ;
  assign \new_[14624]_  = A236 & A233;
  assign \new_[14625]_  = ~A232 & \new_[14624]_ ;
  assign \new_[14629]_  = A269 & A266;
  assign \new_[14630]_  = ~A265 & \new_[14629]_ ;
  assign \new_[14631]_  = \new_[14630]_  & \new_[14625]_ ;
  assign \new_[14635]_  = ~A166 & A167;
  assign \new_[14636]_  = A170 & \new_[14635]_ ;
  assign \new_[14640]_  = ~A202 & ~A200;
  assign \new_[14641]_  = ~A199 & \new_[14640]_ ;
  assign \new_[14642]_  = \new_[14641]_  & \new_[14636]_ ;
  assign \new_[14646]_  = A236 & A233;
  assign \new_[14647]_  = ~A232 & \new_[14646]_ ;
  assign \new_[14651]_  = A269 & ~A266;
  assign \new_[14652]_  = A265 & \new_[14651]_ ;
  assign \new_[14653]_  = \new_[14652]_  & \new_[14647]_ ;
  assign \new_[14657]_  = ~A166 & A167;
  assign \new_[14658]_  = A170 & \new_[14657]_ ;
  assign \new_[14662]_  = ~A202 & ~A200;
  assign \new_[14663]_  = ~A199 & \new_[14662]_ ;
  assign \new_[14664]_  = \new_[14663]_  & \new_[14658]_ ;
  assign \new_[14668]_  = A236 & ~A233;
  assign \new_[14669]_  = A232 & \new_[14668]_ ;
  assign \new_[14673]_  = A302 & ~A299;
  assign \new_[14674]_  = A298 & \new_[14673]_ ;
  assign \new_[14675]_  = \new_[14674]_  & \new_[14669]_ ;
  assign \new_[14679]_  = ~A166 & A167;
  assign \new_[14680]_  = A170 & \new_[14679]_ ;
  assign \new_[14684]_  = ~A202 & ~A200;
  assign \new_[14685]_  = ~A199 & \new_[14684]_ ;
  assign \new_[14686]_  = \new_[14685]_  & \new_[14680]_ ;
  assign \new_[14690]_  = A236 & ~A233;
  assign \new_[14691]_  = A232 & \new_[14690]_ ;
  assign \new_[14695]_  = A302 & A299;
  assign \new_[14696]_  = ~A298 & \new_[14695]_ ;
  assign \new_[14697]_  = \new_[14696]_  & \new_[14691]_ ;
  assign \new_[14701]_  = ~A166 & A167;
  assign \new_[14702]_  = A170 & \new_[14701]_ ;
  assign \new_[14706]_  = ~A202 & ~A200;
  assign \new_[14707]_  = ~A199 & \new_[14706]_ ;
  assign \new_[14708]_  = \new_[14707]_  & \new_[14702]_ ;
  assign \new_[14712]_  = A236 & ~A233;
  assign \new_[14713]_  = A232 & \new_[14712]_ ;
  assign \new_[14717]_  = A269 & A266;
  assign \new_[14718]_  = ~A265 & \new_[14717]_ ;
  assign \new_[14719]_  = \new_[14718]_  & \new_[14713]_ ;
  assign \new_[14723]_  = ~A166 & A167;
  assign \new_[14724]_  = A170 & \new_[14723]_ ;
  assign \new_[14728]_  = ~A202 & ~A200;
  assign \new_[14729]_  = ~A199 & \new_[14728]_ ;
  assign \new_[14730]_  = \new_[14729]_  & \new_[14724]_ ;
  assign \new_[14734]_  = A236 & ~A233;
  assign \new_[14735]_  = A232 & \new_[14734]_ ;
  assign \new_[14739]_  = A269 & ~A266;
  assign \new_[14740]_  = A265 & \new_[14739]_ ;
  assign \new_[14741]_  = \new_[14740]_  & \new_[14735]_ ;
  assign \new_[14745]_  = A166 & ~A167;
  assign \new_[14746]_  = A170 & \new_[14745]_ ;
  assign \new_[14750]_  = ~A203 & ~A202;
  assign \new_[14751]_  = ~A201 & \new_[14750]_ ;
  assign \new_[14752]_  = \new_[14751]_  & \new_[14746]_ ;
  assign \new_[14756]_  = A236 & A233;
  assign \new_[14757]_  = ~A232 & \new_[14756]_ ;
  assign \new_[14761]_  = A302 & ~A299;
  assign \new_[14762]_  = A298 & \new_[14761]_ ;
  assign \new_[14763]_  = \new_[14762]_  & \new_[14757]_ ;
  assign \new_[14767]_  = A166 & ~A167;
  assign \new_[14768]_  = A170 & \new_[14767]_ ;
  assign \new_[14772]_  = ~A203 & ~A202;
  assign \new_[14773]_  = ~A201 & \new_[14772]_ ;
  assign \new_[14774]_  = \new_[14773]_  & \new_[14768]_ ;
  assign \new_[14778]_  = A236 & A233;
  assign \new_[14779]_  = ~A232 & \new_[14778]_ ;
  assign \new_[14783]_  = A302 & A299;
  assign \new_[14784]_  = ~A298 & \new_[14783]_ ;
  assign \new_[14785]_  = \new_[14784]_  & \new_[14779]_ ;
  assign \new_[14789]_  = A166 & ~A167;
  assign \new_[14790]_  = A170 & \new_[14789]_ ;
  assign \new_[14794]_  = ~A203 & ~A202;
  assign \new_[14795]_  = ~A201 & \new_[14794]_ ;
  assign \new_[14796]_  = \new_[14795]_  & \new_[14790]_ ;
  assign \new_[14800]_  = A236 & A233;
  assign \new_[14801]_  = ~A232 & \new_[14800]_ ;
  assign \new_[14805]_  = A269 & A266;
  assign \new_[14806]_  = ~A265 & \new_[14805]_ ;
  assign \new_[14807]_  = \new_[14806]_  & \new_[14801]_ ;
  assign \new_[14811]_  = A166 & ~A167;
  assign \new_[14812]_  = A170 & \new_[14811]_ ;
  assign \new_[14816]_  = ~A203 & ~A202;
  assign \new_[14817]_  = ~A201 & \new_[14816]_ ;
  assign \new_[14818]_  = \new_[14817]_  & \new_[14812]_ ;
  assign \new_[14822]_  = A236 & A233;
  assign \new_[14823]_  = ~A232 & \new_[14822]_ ;
  assign \new_[14827]_  = A269 & ~A266;
  assign \new_[14828]_  = A265 & \new_[14827]_ ;
  assign \new_[14829]_  = \new_[14828]_  & \new_[14823]_ ;
  assign \new_[14833]_  = A166 & ~A167;
  assign \new_[14834]_  = A170 & \new_[14833]_ ;
  assign \new_[14838]_  = ~A203 & ~A202;
  assign \new_[14839]_  = ~A201 & \new_[14838]_ ;
  assign \new_[14840]_  = \new_[14839]_  & \new_[14834]_ ;
  assign \new_[14844]_  = A236 & ~A233;
  assign \new_[14845]_  = A232 & \new_[14844]_ ;
  assign \new_[14849]_  = A302 & ~A299;
  assign \new_[14850]_  = A298 & \new_[14849]_ ;
  assign \new_[14851]_  = \new_[14850]_  & \new_[14845]_ ;
  assign \new_[14855]_  = A166 & ~A167;
  assign \new_[14856]_  = A170 & \new_[14855]_ ;
  assign \new_[14860]_  = ~A203 & ~A202;
  assign \new_[14861]_  = ~A201 & \new_[14860]_ ;
  assign \new_[14862]_  = \new_[14861]_  & \new_[14856]_ ;
  assign \new_[14866]_  = A236 & ~A233;
  assign \new_[14867]_  = A232 & \new_[14866]_ ;
  assign \new_[14871]_  = A302 & A299;
  assign \new_[14872]_  = ~A298 & \new_[14871]_ ;
  assign \new_[14873]_  = \new_[14872]_  & \new_[14867]_ ;
  assign \new_[14877]_  = A166 & ~A167;
  assign \new_[14878]_  = A170 & \new_[14877]_ ;
  assign \new_[14882]_  = ~A203 & ~A202;
  assign \new_[14883]_  = ~A201 & \new_[14882]_ ;
  assign \new_[14884]_  = \new_[14883]_  & \new_[14878]_ ;
  assign \new_[14888]_  = A236 & ~A233;
  assign \new_[14889]_  = A232 & \new_[14888]_ ;
  assign \new_[14893]_  = A269 & A266;
  assign \new_[14894]_  = ~A265 & \new_[14893]_ ;
  assign \new_[14895]_  = \new_[14894]_  & \new_[14889]_ ;
  assign \new_[14899]_  = A166 & ~A167;
  assign \new_[14900]_  = A170 & \new_[14899]_ ;
  assign \new_[14904]_  = ~A203 & ~A202;
  assign \new_[14905]_  = ~A201 & \new_[14904]_ ;
  assign \new_[14906]_  = \new_[14905]_  & \new_[14900]_ ;
  assign \new_[14910]_  = A236 & ~A233;
  assign \new_[14911]_  = A232 & \new_[14910]_ ;
  assign \new_[14915]_  = A269 & ~A266;
  assign \new_[14916]_  = A265 & \new_[14915]_ ;
  assign \new_[14917]_  = \new_[14916]_  & \new_[14911]_ ;
  assign \new_[14921]_  = A166 & ~A167;
  assign \new_[14922]_  = A170 & \new_[14921]_ ;
  assign \new_[14926]_  = ~A201 & A200;
  assign \new_[14927]_  = A199 & \new_[14926]_ ;
  assign \new_[14928]_  = \new_[14927]_  & \new_[14922]_ ;
  assign \new_[14932]_  = A234 & A232;
  assign \new_[14933]_  = ~A202 & \new_[14932]_ ;
  assign \new_[14937]_  = A302 & ~A299;
  assign \new_[14938]_  = A298 & \new_[14937]_ ;
  assign \new_[14939]_  = \new_[14938]_  & \new_[14933]_ ;
  assign \new_[14943]_  = A166 & ~A167;
  assign \new_[14944]_  = A170 & \new_[14943]_ ;
  assign \new_[14948]_  = ~A201 & A200;
  assign \new_[14949]_  = A199 & \new_[14948]_ ;
  assign \new_[14950]_  = \new_[14949]_  & \new_[14944]_ ;
  assign \new_[14954]_  = A234 & A232;
  assign \new_[14955]_  = ~A202 & \new_[14954]_ ;
  assign \new_[14959]_  = A302 & A299;
  assign \new_[14960]_  = ~A298 & \new_[14959]_ ;
  assign \new_[14961]_  = \new_[14960]_  & \new_[14955]_ ;
  assign \new_[14965]_  = A166 & ~A167;
  assign \new_[14966]_  = A170 & \new_[14965]_ ;
  assign \new_[14970]_  = ~A201 & A200;
  assign \new_[14971]_  = A199 & \new_[14970]_ ;
  assign \new_[14972]_  = \new_[14971]_  & \new_[14966]_ ;
  assign \new_[14976]_  = A234 & A232;
  assign \new_[14977]_  = ~A202 & \new_[14976]_ ;
  assign \new_[14981]_  = A269 & A266;
  assign \new_[14982]_  = ~A265 & \new_[14981]_ ;
  assign \new_[14983]_  = \new_[14982]_  & \new_[14977]_ ;
  assign \new_[14987]_  = A166 & ~A167;
  assign \new_[14988]_  = A170 & \new_[14987]_ ;
  assign \new_[14992]_  = ~A201 & A200;
  assign \new_[14993]_  = A199 & \new_[14992]_ ;
  assign \new_[14994]_  = \new_[14993]_  & \new_[14988]_ ;
  assign \new_[14998]_  = A234 & A232;
  assign \new_[14999]_  = ~A202 & \new_[14998]_ ;
  assign \new_[15003]_  = A269 & ~A266;
  assign \new_[15004]_  = A265 & \new_[15003]_ ;
  assign \new_[15005]_  = \new_[15004]_  & \new_[14999]_ ;
  assign \new_[15009]_  = A166 & ~A167;
  assign \new_[15010]_  = A170 & \new_[15009]_ ;
  assign \new_[15014]_  = ~A201 & A200;
  assign \new_[15015]_  = A199 & \new_[15014]_ ;
  assign \new_[15016]_  = \new_[15015]_  & \new_[15010]_ ;
  assign \new_[15020]_  = A234 & A233;
  assign \new_[15021]_  = ~A202 & \new_[15020]_ ;
  assign \new_[15025]_  = A302 & ~A299;
  assign \new_[15026]_  = A298 & \new_[15025]_ ;
  assign \new_[15027]_  = \new_[15026]_  & \new_[15021]_ ;
  assign \new_[15031]_  = A166 & ~A167;
  assign \new_[15032]_  = A170 & \new_[15031]_ ;
  assign \new_[15036]_  = ~A201 & A200;
  assign \new_[15037]_  = A199 & \new_[15036]_ ;
  assign \new_[15038]_  = \new_[15037]_  & \new_[15032]_ ;
  assign \new_[15042]_  = A234 & A233;
  assign \new_[15043]_  = ~A202 & \new_[15042]_ ;
  assign \new_[15047]_  = A302 & A299;
  assign \new_[15048]_  = ~A298 & \new_[15047]_ ;
  assign \new_[15049]_  = \new_[15048]_  & \new_[15043]_ ;
  assign \new_[15053]_  = A166 & ~A167;
  assign \new_[15054]_  = A170 & \new_[15053]_ ;
  assign \new_[15058]_  = ~A201 & A200;
  assign \new_[15059]_  = A199 & \new_[15058]_ ;
  assign \new_[15060]_  = \new_[15059]_  & \new_[15054]_ ;
  assign \new_[15064]_  = A234 & A233;
  assign \new_[15065]_  = ~A202 & \new_[15064]_ ;
  assign \new_[15069]_  = A269 & A266;
  assign \new_[15070]_  = ~A265 & \new_[15069]_ ;
  assign \new_[15071]_  = \new_[15070]_  & \new_[15065]_ ;
  assign \new_[15075]_  = A166 & ~A167;
  assign \new_[15076]_  = A170 & \new_[15075]_ ;
  assign \new_[15080]_  = ~A201 & A200;
  assign \new_[15081]_  = A199 & \new_[15080]_ ;
  assign \new_[15082]_  = \new_[15081]_  & \new_[15076]_ ;
  assign \new_[15086]_  = A234 & A233;
  assign \new_[15087]_  = ~A202 & \new_[15086]_ ;
  assign \new_[15091]_  = A269 & ~A266;
  assign \new_[15092]_  = A265 & \new_[15091]_ ;
  assign \new_[15093]_  = \new_[15092]_  & \new_[15087]_ ;
  assign \new_[15097]_  = A166 & ~A167;
  assign \new_[15098]_  = A170 & \new_[15097]_ ;
  assign \new_[15102]_  = ~A201 & A200;
  assign \new_[15103]_  = A199 & \new_[15102]_ ;
  assign \new_[15104]_  = \new_[15103]_  & \new_[15098]_ ;
  assign \new_[15108]_  = A233 & ~A232;
  assign \new_[15109]_  = ~A202 & \new_[15108]_ ;
  assign \new_[15113]_  = A300 & A299;
  assign \new_[15114]_  = A236 & \new_[15113]_ ;
  assign \new_[15115]_  = \new_[15114]_  & \new_[15109]_ ;
  assign \new_[15119]_  = A166 & ~A167;
  assign \new_[15120]_  = A170 & \new_[15119]_ ;
  assign \new_[15124]_  = ~A201 & A200;
  assign \new_[15125]_  = A199 & \new_[15124]_ ;
  assign \new_[15126]_  = \new_[15125]_  & \new_[15120]_ ;
  assign \new_[15130]_  = A233 & ~A232;
  assign \new_[15131]_  = ~A202 & \new_[15130]_ ;
  assign \new_[15135]_  = A300 & A298;
  assign \new_[15136]_  = A236 & \new_[15135]_ ;
  assign \new_[15137]_  = \new_[15136]_  & \new_[15131]_ ;
  assign \new_[15141]_  = A166 & ~A167;
  assign \new_[15142]_  = A170 & \new_[15141]_ ;
  assign \new_[15146]_  = ~A201 & A200;
  assign \new_[15147]_  = A199 & \new_[15146]_ ;
  assign \new_[15148]_  = \new_[15147]_  & \new_[15142]_ ;
  assign \new_[15152]_  = A233 & ~A232;
  assign \new_[15153]_  = ~A202 & \new_[15152]_ ;
  assign \new_[15157]_  = A267 & A265;
  assign \new_[15158]_  = A236 & \new_[15157]_ ;
  assign \new_[15159]_  = \new_[15158]_  & \new_[15153]_ ;
  assign \new_[15163]_  = A166 & ~A167;
  assign \new_[15164]_  = A170 & \new_[15163]_ ;
  assign \new_[15168]_  = ~A201 & A200;
  assign \new_[15169]_  = A199 & \new_[15168]_ ;
  assign \new_[15170]_  = \new_[15169]_  & \new_[15164]_ ;
  assign \new_[15174]_  = A233 & ~A232;
  assign \new_[15175]_  = ~A202 & \new_[15174]_ ;
  assign \new_[15179]_  = A267 & A266;
  assign \new_[15180]_  = A236 & \new_[15179]_ ;
  assign \new_[15181]_  = \new_[15180]_  & \new_[15175]_ ;
  assign \new_[15185]_  = A166 & ~A167;
  assign \new_[15186]_  = A170 & \new_[15185]_ ;
  assign \new_[15190]_  = ~A201 & A200;
  assign \new_[15191]_  = A199 & \new_[15190]_ ;
  assign \new_[15192]_  = \new_[15191]_  & \new_[15186]_ ;
  assign \new_[15196]_  = ~A233 & A232;
  assign \new_[15197]_  = ~A202 & \new_[15196]_ ;
  assign \new_[15201]_  = A300 & A299;
  assign \new_[15202]_  = A236 & \new_[15201]_ ;
  assign \new_[15203]_  = \new_[15202]_  & \new_[15197]_ ;
  assign \new_[15207]_  = A166 & ~A167;
  assign \new_[15208]_  = A170 & \new_[15207]_ ;
  assign \new_[15212]_  = ~A201 & A200;
  assign \new_[15213]_  = A199 & \new_[15212]_ ;
  assign \new_[15214]_  = \new_[15213]_  & \new_[15208]_ ;
  assign \new_[15218]_  = ~A233 & A232;
  assign \new_[15219]_  = ~A202 & \new_[15218]_ ;
  assign \new_[15223]_  = A300 & A298;
  assign \new_[15224]_  = A236 & \new_[15223]_ ;
  assign \new_[15225]_  = \new_[15224]_  & \new_[15219]_ ;
  assign \new_[15229]_  = A166 & ~A167;
  assign \new_[15230]_  = A170 & \new_[15229]_ ;
  assign \new_[15234]_  = ~A201 & A200;
  assign \new_[15235]_  = A199 & \new_[15234]_ ;
  assign \new_[15236]_  = \new_[15235]_  & \new_[15230]_ ;
  assign \new_[15240]_  = ~A233 & A232;
  assign \new_[15241]_  = ~A202 & \new_[15240]_ ;
  assign \new_[15245]_  = A267 & A265;
  assign \new_[15246]_  = A236 & \new_[15245]_ ;
  assign \new_[15247]_  = \new_[15246]_  & \new_[15241]_ ;
  assign \new_[15251]_  = A166 & ~A167;
  assign \new_[15252]_  = A170 & \new_[15251]_ ;
  assign \new_[15256]_  = ~A201 & A200;
  assign \new_[15257]_  = A199 & \new_[15256]_ ;
  assign \new_[15258]_  = \new_[15257]_  & \new_[15252]_ ;
  assign \new_[15262]_  = ~A233 & A232;
  assign \new_[15263]_  = ~A202 & \new_[15262]_ ;
  assign \new_[15267]_  = A267 & A266;
  assign \new_[15268]_  = A236 & \new_[15267]_ ;
  assign \new_[15269]_  = \new_[15268]_  & \new_[15263]_ ;
  assign \new_[15273]_  = A166 & ~A167;
  assign \new_[15274]_  = A170 & \new_[15273]_ ;
  assign \new_[15278]_  = ~A202 & ~A200;
  assign \new_[15279]_  = ~A199 & \new_[15278]_ ;
  assign \new_[15280]_  = \new_[15279]_  & \new_[15274]_ ;
  assign \new_[15284]_  = A236 & A233;
  assign \new_[15285]_  = ~A232 & \new_[15284]_ ;
  assign \new_[15289]_  = A302 & ~A299;
  assign \new_[15290]_  = A298 & \new_[15289]_ ;
  assign \new_[15291]_  = \new_[15290]_  & \new_[15285]_ ;
  assign \new_[15295]_  = A166 & ~A167;
  assign \new_[15296]_  = A170 & \new_[15295]_ ;
  assign \new_[15300]_  = ~A202 & ~A200;
  assign \new_[15301]_  = ~A199 & \new_[15300]_ ;
  assign \new_[15302]_  = \new_[15301]_  & \new_[15296]_ ;
  assign \new_[15306]_  = A236 & A233;
  assign \new_[15307]_  = ~A232 & \new_[15306]_ ;
  assign \new_[15311]_  = A302 & A299;
  assign \new_[15312]_  = ~A298 & \new_[15311]_ ;
  assign \new_[15313]_  = \new_[15312]_  & \new_[15307]_ ;
  assign \new_[15317]_  = A166 & ~A167;
  assign \new_[15318]_  = A170 & \new_[15317]_ ;
  assign \new_[15322]_  = ~A202 & ~A200;
  assign \new_[15323]_  = ~A199 & \new_[15322]_ ;
  assign \new_[15324]_  = \new_[15323]_  & \new_[15318]_ ;
  assign \new_[15328]_  = A236 & A233;
  assign \new_[15329]_  = ~A232 & \new_[15328]_ ;
  assign \new_[15333]_  = A269 & A266;
  assign \new_[15334]_  = ~A265 & \new_[15333]_ ;
  assign \new_[15335]_  = \new_[15334]_  & \new_[15329]_ ;
  assign \new_[15339]_  = A166 & ~A167;
  assign \new_[15340]_  = A170 & \new_[15339]_ ;
  assign \new_[15344]_  = ~A202 & ~A200;
  assign \new_[15345]_  = ~A199 & \new_[15344]_ ;
  assign \new_[15346]_  = \new_[15345]_  & \new_[15340]_ ;
  assign \new_[15350]_  = A236 & A233;
  assign \new_[15351]_  = ~A232 & \new_[15350]_ ;
  assign \new_[15355]_  = A269 & ~A266;
  assign \new_[15356]_  = A265 & \new_[15355]_ ;
  assign \new_[15357]_  = \new_[15356]_  & \new_[15351]_ ;
  assign \new_[15361]_  = A166 & ~A167;
  assign \new_[15362]_  = A170 & \new_[15361]_ ;
  assign \new_[15366]_  = ~A202 & ~A200;
  assign \new_[15367]_  = ~A199 & \new_[15366]_ ;
  assign \new_[15368]_  = \new_[15367]_  & \new_[15362]_ ;
  assign \new_[15372]_  = A236 & ~A233;
  assign \new_[15373]_  = A232 & \new_[15372]_ ;
  assign \new_[15377]_  = A302 & ~A299;
  assign \new_[15378]_  = A298 & \new_[15377]_ ;
  assign \new_[15379]_  = \new_[15378]_  & \new_[15373]_ ;
  assign \new_[15383]_  = A166 & ~A167;
  assign \new_[15384]_  = A170 & \new_[15383]_ ;
  assign \new_[15388]_  = ~A202 & ~A200;
  assign \new_[15389]_  = ~A199 & \new_[15388]_ ;
  assign \new_[15390]_  = \new_[15389]_  & \new_[15384]_ ;
  assign \new_[15394]_  = A236 & ~A233;
  assign \new_[15395]_  = A232 & \new_[15394]_ ;
  assign \new_[15399]_  = A302 & A299;
  assign \new_[15400]_  = ~A298 & \new_[15399]_ ;
  assign \new_[15401]_  = \new_[15400]_  & \new_[15395]_ ;
  assign \new_[15405]_  = A166 & ~A167;
  assign \new_[15406]_  = A170 & \new_[15405]_ ;
  assign \new_[15410]_  = ~A202 & ~A200;
  assign \new_[15411]_  = ~A199 & \new_[15410]_ ;
  assign \new_[15412]_  = \new_[15411]_  & \new_[15406]_ ;
  assign \new_[15416]_  = A236 & ~A233;
  assign \new_[15417]_  = A232 & \new_[15416]_ ;
  assign \new_[15421]_  = A269 & A266;
  assign \new_[15422]_  = ~A265 & \new_[15421]_ ;
  assign \new_[15423]_  = \new_[15422]_  & \new_[15417]_ ;
  assign \new_[15427]_  = A166 & ~A167;
  assign \new_[15428]_  = A170 & \new_[15427]_ ;
  assign \new_[15432]_  = ~A202 & ~A200;
  assign \new_[15433]_  = ~A199 & \new_[15432]_ ;
  assign \new_[15434]_  = \new_[15433]_  & \new_[15428]_ ;
  assign \new_[15438]_  = A236 & ~A233;
  assign \new_[15439]_  = A232 & \new_[15438]_ ;
  assign \new_[15443]_  = A269 & ~A266;
  assign \new_[15444]_  = A265 & \new_[15443]_ ;
  assign \new_[15445]_  = \new_[15444]_  & \new_[15439]_ ;
  assign \new_[15449]_  = ~A166 & A167;
  assign \new_[15450]_  = A170 & \new_[15449]_ ;
  assign \new_[15454]_  = ~A201 & A200;
  assign \new_[15455]_  = A199 & \new_[15454]_ ;
  assign \new_[15456]_  = \new_[15455]_  & \new_[15450]_ ;
  assign \new_[15460]_  = A233 & ~A232;
  assign \new_[15461]_  = ~A202 & \new_[15460]_ ;
  assign \new_[15464]_  = A298 & A236;
  assign \new_[15467]_  = A302 & ~A299;
  assign \new_[15468]_  = \new_[15467]_  & \new_[15464]_ ;
  assign \new_[15469]_  = \new_[15468]_  & \new_[15461]_ ;
  assign \new_[15473]_  = ~A166 & A167;
  assign \new_[15474]_  = A170 & \new_[15473]_ ;
  assign \new_[15478]_  = ~A201 & A200;
  assign \new_[15479]_  = A199 & \new_[15478]_ ;
  assign \new_[15480]_  = \new_[15479]_  & \new_[15474]_ ;
  assign \new_[15484]_  = A233 & ~A232;
  assign \new_[15485]_  = ~A202 & \new_[15484]_ ;
  assign \new_[15488]_  = ~A298 & A236;
  assign \new_[15491]_  = A302 & A299;
  assign \new_[15492]_  = \new_[15491]_  & \new_[15488]_ ;
  assign \new_[15493]_  = \new_[15492]_  & \new_[15485]_ ;
  assign \new_[15497]_  = ~A166 & A167;
  assign \new_[15498]_  = A170 & \new_[15497]_ ;
  assign \new_[15502]_  = ~A201 & A200;
  assign \new_[15503]_  = A199 & \new_[15502]_ ;
  assign \new_[15504]_  = \new_[15503]_  & \new_[15498]_ ;
  assign \new_[15508]_  = A233 & ~A232;
  assign \new_[15509]_  = ~A202 & \new_[15508]_ ;
  assign \new_[15512]_  = ~A265 & A236;
  assign \new_[15515]_  = A269 & A266;
  assign \new_[15516]_  = \new_[15515]_  & \new_[15512]_ ;
  assign \new_[15517]_  = \new_[15516]_  & \new_[15509]_ ;
  assign \new_[15521]_  = ~A166 & A167;
  assign \new_[15522]_  = A170 & \new_[15521]_ ;
  assign \new_[15526]_  = ~A201 & A200;
  assign \new_[15527]_  = A199 & \new_[15526]_ ;
  assign \new_[15528]_  = \new_[15527]_  & \new_[15522]_ ;
  assign \new_[15532]_  = A233 & ~A232;
  assign \new_[15533]_  = ~A202 & \new_[15532]_ ;
  assign \new_[15536]_  = A265 & A236;
  assign \new_[15539]_  = A269 & ~A266;
  assign \new_[15540]_  = \new_[15539]_  & \new_[15536]_ ;
  assign \new_[15541]_  = \new_[15540]_  & \new_[15533]_ ;
  assign \new_[15545]_  = ~A166 & A167;
  assign \new_[15546]_  = A170 & \new_[15545]_ ;
  assign \new_[15550]_  = ~A201 & A200;
  assign \new_[15551]_  = A199 & \new_[15550]_ ;
  assign \new_[15552]_  = \new_[15551]_  & \new_[15546]_ ;
  assign \new_[15556]_  = ~A233 & A232;
  assign \new_[15557]_  = ~A202 & \new_[15556]_ ;
  assign \new_[15560]_  = A298 & A236;
  assign \new_[15563]_  = A302 & ~A299;
  assign \new_[15564]_  = \new_[15563]_  & \new_[15560]_ ;
  assign \new_[15565]_  = \new_[15564]_  & \new_[15557]_ ;
  assign \new_[15569]_  = ~A166 & A167;
  assign \new_[15570]_  = A170 & \new_[15569]_ ;
  assign \new_[15574]_  = ~A201 & A200;
  assign \new_[15575]_  = A199 & \new_[15574]_ ;
  assign \new_[15576]_  = \new_[15575]_  & \new_[15570]_ ;
  assign \new_[15580]_  = ~A233 & A232;
  assign \new_[15581]_  = ~A202 & \new_[15580]_ ;
  assign \new_[15584]_  = ~A298 & A236;
  assign \new_[15587]_  = A302 & A299;
  assign \new_[15588]_  = \new_[15587]_  & \new_[15584]_ ;
  assign \new_[15589]_  = \new_[15588]_  & \new_[15581]_ ;
  assign \new_[15593]_  = ~A166 & A167;
  assign \new_[15594]_  = A170 & \new_[15593]_ ;
  assign \new_[15598]_  = ~A201 & A200;
  assign \new_[15599]_  = A199 & \new_[15598]_ ;
  assign \new_[15600]_  = \new_[15599]_  & \new_[15594]_ ;
  assign \new_[15604]_  = ~A233 & A232;
  assign \new_[15605]_  = ~A202 & \new_[15604]_ ;
  assign \new_[15608]_  = ~A265 & A236;
  assign \new_[15611]_  = A269 & A266;
  assign \new_[15612]_  = \new_[15611]_  & \new_[15608]_ ;
  assign \new_[15613]_  = \new_[15612]_  & \new_[15605]_ ;
  assign \new_[15617]_  = ~A166 & A167;
  assign \new_[15618]_  = A170 & \new_[15617]_ ;
  assign \new_[15622]_  = ~A201 & A200;
  assign \new_[15623]_  = A199 & \new_[15622]_ ;
  assign \new_[15624]_  = \new_[15623]_  & \new_[15618]_ ;
  assign \new_[15628]_  = ~A233 & A232;
  assign \new_[15629]_  = ~A202 & \new_[15628]_ ;
  assign \new_[15632]_  = A265 & A236;
  assign \new_[15635]_  = A269 & ~A266;
  assign \new_[15636]_  = \new_[15635]_  & \new_[15632]_ ;
  assign \new_[15637]_  = \new_[15636]_  & \new_[15629]_ ;
  assign \new_[15641]_  = A166 & ~A167;
  assign \new_[15642]_  = A170 & \new_[15641]_ ;
  assign \new_[15646]_  = ~A201 & A200;
  assign \new_[15647]_  = A199 & \new_[15646]_ ;
  assign \new_[15648]_  = \new_[15647]_  & \new_[15642]_ ;
  assign \new_[15652]_  = A233 & ~A232;
  assign \new_[15653]_  = ~A202 & \new_[15652]_ ;
  assign \new_[15656]_  = A298 & A236;
  assign \new_[15659]_  = A302 & ~A299;
  assign \new_[15660]_  = \new_[15659]_  & \new_[15656]_ ;
  assign \new_[15661]_  = \new_[15660]_  & \new_[15653]_ ;
  assign \new_[15665]_  = A166 & ~A167;
  assign \new_[15666]_  = A170 & \new_[15665]_ ;
  assign \new_[15670]_  = ~A201 & A200;
  assign \new_[15671]_  = A199 & \new_[15670]_ ;
  assign \new_[15672]_  = \new_[15671]_  & \new_[15666]_ ;
  assign \new_[15676]_  = A233 & ~A232;
  assign \new_[15677]_  = ~A202 & \new_[15676]_ ;
  assign \new_[15680]_  = ~A298 & A236;
  assign \new_[15683]_  = A302 & A299;
  assign \new_[15684]_  = \new_[15683]_  & \new_[15680]_ ;
  assign \new_[15685]_  = \new_[15684]_  & \new_[15677]_ ;
  assign \new_[15689]_  = A166 & ~A167;
  assign \new_[15690]_  = A170 & \new_[15689]_ ;
  assign \new_[15694]_  = ~A201 & A200;
  assign \new_[15695]_  = A199 & \new_[15694]_ ;
  assign \new_[15696]_  = \new_[15695]_  & \new_[15690]_ ;
  assign \new_[15700]_  = A233 & ~A232;
  assign \new_[15701]_  = ~A202 & \new_[15700]_ ;
  assign \new_[15704]_  = ~A265 & A236;
  assign \new_[15707]_  = A269 & A266;
  assign \new_[15708]_  = \new_[15707]_  & \new_[15704]_ ;
  assign \new_[15709]_  = \new_[15708]_  & \new_[15701]_ ;
  assign \new_[15713]_  = A166 & ~A167;
  assign \new_[15714]_  = A170 & \new_[15713]_ ;
  assign \new_[15718]_  = ~A201 & A200;
  assign \new_[15719]_  = A199 & \new_[15718]_ ;
  assign \new_[15720]_  = \new_[15719]_  & \new_[15714]_ ;
  assign \new_[15724]_  = A233 & ~A232;
  assign \new_[15725]_  = ~A202 & \new_[15724]_ ;
  assign \new_[15728]_  = A265 & A236;
  assign \new_[15731]_  = A269 & ~A266;
  assign \new_[15732]_  = \new_[15731]_  & \new_[15728]_ ;
  assign \new_[15733]_  = \new_[15732]_  & \new_[15725]_ ;
  assign \new_[15737]_  = A166 & ~A167;
  assign \new_[15738]_  = A170 & \new_[15737]_ ;
  assign \new_[15742]_  = ~A201 & A200;
  assign \new_[15743]_  = A199 & \new_[15742]_ ;
  assign \new_[15744]_  = \new_[15743]_  & \new_[15738]_ ;
  assign \new_[15748]_  = ~A233 & A232;
  assign \new_[15749]_  = ~A202 & \new_[15748]_ ;
  assign \new_[15752]_  = A298 & A236;
  assign \new_[15755]_  = A302 & ~A299;
  assign \new_[15756]_  = \new_[15755]_  & \new_[15752]_ ;
  assign \new_[15757]_  = \new_[15756]_  & \new_[15749]_ ;
  assign \new_[15761]_  = A166 & ~A167;
  assign \new_[15762]_  = A170 & \new_[15761]_ ;
  assign \new_[15766]_  = ~A201 & A200;
  assign \new_[15767]_  = A199 & \new_[15766]_ ;
  assign \new_[15768]_  = \new_[15767]_  & \new_[15762]_ ;
  assign \new_[15772]_  = ~A233 & A232;
  assign \new_[15773]_  = ~A202 & \new_[15772]_ ;
  assign \new_[15776]_  = ~A298 & A236;
  assign \new_[15779]_  = A302 & A299;
  assign \new_[15780]_  = \new_[15779]_  & \new_[15776]_ ;
  assign \new_[15781]_  = \new_[15780]_  & \new_[15773]_ ;
  assign \new_[15785]_  = A166 & ~A167;
  assign \new_[15786]_  = A170 & \new_[15785]_ ;
  assign \new_[15790]_  = ~A201 & A200;
  assign \new_[15791]_  = A199 & \new_[15790]_ ;
  assign \new_[15792]_  = \new_[15791]_  & \new_[15786]_ ;
  assign \new_[15796]_  = ~A233 & A232;
  assign \new_[15797]_  = ~A202 & \new_[15796]_ ;
  assign \new_[15800]_  = ~A265 & A236;
  assign \new_[15803]_  = A269 & A266;
  assign \new_[15804]_  = \new_[15803]_  & \new_[15800]_ ;
  assign \new_[15805]_  = \new_[15804]_  & \new_[15797]_ ;
  assign \new_[15809]_  = A166 & ~A167;
  assign \new_[15810]_  = A170 & \new_[15809]_ ;
  assign \new_[15814]_  = ~A201 & A200;
  assign \new_[15815]_  = A199 & \new_[15814]_ ;
  assign \new_[15816]_  = \new_[15815]_  & \new_[15810]_ ;
  assign \new_[15820]_  = ~A233 & A232;
  assign \new_[15821]_  = ~A202 & \new_[15820]_ ;
  assign \new_[15824]_  = A265 & A236;
  assign \new_[15827]_  = A269 & ~A266;
  assign \new_[15828]_  = \new_[15827]_  & \new_[15824]_ ;
  assign \new_[15829]_  = \new_[15828]_  & \new_[15821]_ ;
endmodule


