module top ( 
    i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_, i_10_,
    i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_, i_4_,
    i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_, i_24_,
    i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_, i_32_,
    i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_, i_19_,
    i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_, i_38_,
    i_29_, i_51_, i_44_, i_37_,
    o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_  );
  input  i_63_, i_50_, i_64_, i_61_, i_62_, i_40_, i_30_, i_20_, i_9_,
    i_10_, i_7_, i_8_, i_5_, i_6_, i_27_, i_14_, i_3_, i_39_, i_28_, i_13_,
    i_4_, i_25_, i_12_, i_1_, i_26_, i_11_, i_2_, i_49_, i_23_, i_18_,
    i_24_, i_17_, i_0_, i_21_, i_16_, i_59_, i_22_, i_15_, i_58_, i_45_,
    i_32_, i_57_, i_46_, i_31_, i_56_, i_47_, i_34_, i_55_, i_48_, i_33_,
    i_19_, i_54_, i_41_, i_36_, i_60_, i_53_, i_42_, i_35_, i_52_, i_43_,
    i_38_, i_29_, i_51_, i_44_, i_37_;
  output o_1_, o_19_, o_2_, o_0_, o_29_, o_60_, o_39_, o_38_, o_25_, o_12_,
    o_37_, o_26_, o_11_, o_50_, o_36_, o_27_, o_14_, o_35_, o_28_, o_13_,
    o_34_, o_21_, o_16_, o_40_, o_33_, o_22_, o_15_, o_32_, o_23_, o_18_,
    o_31_, o_24_, o_17_, o_56_, o_43_, o_30_, o_55_, o_44_, o_58_, o_41_,
    o_57_, o_42_, o_20_, o_52_, o_47_, o_51_, o_48_, o_54_, o_45_, o_10_,
    o_53_, o_46_, o_61_, o_9_, o_62_, o_63_, o_49_, o_7_, o_64_, o_8_,
    o_5_, o_59_, o_6_, o_3_, o_4_;
  wire new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n424_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n473_, new_n474_, new_n475_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_,
    new_n578_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_;
  assign new_n131_ = ~i_59_ & ~i_60_;
  assign new_n132_ = ~i_58_ & new_n131_;
  assign new_n133_ = ~i_61_ & ~i_62_;
  assign new_n134_ = ~i_56_ & ~i_55_;
  assign new_n135_ = ~i_54_ & new_n134_;
  assign new_n136_ = new_n132_ & new_n133_;
  assign new_n137_ = new_n135_ & new_n136_;
  assign new_n138_ = ~i_46_ & ~i_47_;
  assign new_n139_ = ~i_43_ & new_n138_;
  assign new_n140_ = ~i_53_ & ~i_51_;
  assign new_n141_ = ~i_50_ & new_n140_;
  assign new_n142_ = ~i_41_ & ~i_42_;
  assign new_n143_ = ~i_40_ & new_n142_;
  assign new_n144_ = new_n139_ & new_n141_;
  assign new_n145_ = new_n143_ & new_n144_;
  assign new_n146_ = new_n137_ & new_n145_;
  assign new_n147_ = ~i_18_ & ~i_22_;
  assign new_n148_ = ~i_17_ & new_n147_;
  assign new_n149_ = ~i_25_ & ~i_26_;
  assign new_n150_ = ~i_24_ & new_n149_;
  assign new_n151_ = ~i_14_ & ~i_15_;
  assign new_n152_ = ~i_11_ & new_n151_;
  assign new_n153_ = new_n148_ & new_n150_;
  assign new_n154_ = new_n152_ & new_n153_;
  assign new_n155_ = ~i_34_ & ~i_33_;
  assign new_n156_ = ~i_31_ & new_n155_;
  assign new_n157_ = ~i_39_ & ~i_37_;
  assign new_n158_ = ~i_35_ & new_n157_;
  assign new_n159_ = ~i_30_ & i_29_;
  assign new_n160_ = ~i_28_ & new_n159_;
  assign new_n161_ = new_n156_ & new_n158_;
  assign new_n162_ = new_n160_ & new_n161_;
  assign new_n163_ = ~i_7_ & ~i_6_;
  assign new_n164_ = i_5_ & new_n163_;
  assign new_n165_ = ~i_9_ & ~i_10_;
  assign new_n166_ = ~i_8_ & new_n165_;
  assign new_n167_ = ~i_3_ & ~i_4_;
  assign new_n168_ = ~i_0_ & new_n167_;
  assign new_n169_ = new_n164_ & new_n166_;
  assign new_n170_ = new_n168_ & new_n169_;
  assign new_n171_ = new_n154_ & new_n162_;
  assign new_n172_ = new_n170_ & new_n171_;
  assign o_1_ = new_n146_ & new_n172_;
  assign new_n174_ = ~i_54_ & ~i_53_;
  assign new_n175_ = ~i_51_ & new_n174_;
  assign new_n176_ = ~i_57_ & ~i_56_;
  assign new_n177_ = ~i_55_ & new_n176_;
  assign new_n178_ = ~i_50_ & ~i_49_;
  assign new_n179_ = ~i_48_ & new_n178_;
  assign new_n180_ = new_n175_ & new_n177_;
  assign new_n181_ = new_n179_ & new_n180_;
  assign new_n182_ = i_64_ & ~i_62_;
  assign new_n183_ = ~i_61_ & new_n182_;
  assign new_n184_ = new_n132_ & new_n183_;
  assign new_n185_ = ~i_42_ & ~i_43_;
  assign new_n186_ = ~i_41_ & new_n185_;
  assign new_n187_ = ~i_45_ & new_n138_;
  assign new_n188_ = ~i_40_ & ~i_39_;
  assign new_n189_ = ~i_37_ & new_n188_;
  assign new_n190_ = new_n186_ & new_n187_;
  assign new_n191_ = new_n189_ & new_n190_;
  assign new_n192_ = new_n181_ & new_n184_;
  assign new_n193_ = new_n191_ & new_n192_;
  assign new_n194_ = ~i_17_ & ~i_15_;
  assign new_n195_ = ~i_14_ & new_n194_;
  assign new_n196_ = ~i_24_ & ~i_22_;
  assign new_n197_ = ~i_18_ & new_n196_;
  assign new_n198_ = ~i_10_ & ~i_11_;
  assign new_n199_ = ~i_9_ & new_n198_;
  assign new_n200_ = new_n195_ & new_n197_;
  assign new_n201_ = new_n199_ & new_n200_;
  assign new_n202_ = ~i_30_ & ~i_31_;
  assign new_n203_ = i_29_ & new_n202_;
  assign new_n204_ = ~i_34_ & ~i_35_;
  assign new_n205_ = ~i_33_ & new_n204_;
  assign new_n206_ = ~i_28_ & ~i_26_;
  assign new_n207_ = ~i_25_ & new_n206_;
  assign new_n208_ = new_n203_ & new_n205_;
  assign new_n209_ = new_n207_ & new_n208_;
  assign new_n210_ = ~i_5_ & ~i_4_;
  assign new_n211_ = ~i_3_ & new_n210_;
  assign new_n212_ = ~i_7_ & ~i_8_;
  assign new_n213_ = ~i_6_ & new_n212_;
  assign new_n214_ = ~i_1_ & ~i_2_;
  assign new_n215_ = ~i_0_ & new_n214_;
  assign new_n216_ = new_n211_ & new_n213_;
  assign new_n217_ = new_n215_ & new_n216_;
  assign new_n218_ = new_n201_ & new_n209_;
  assign new_n219_ = new_n217_ & new_n218_;
  assign o_19_ = new_n193_ & new_n219_;
  assign new_n221_ = ~i_40_ & ~i_41_;
  assign new_n222_ = ~i_39_ & new_n221_;
  assign new_n223_ = ~i_43_ & ~i_44_;
  assign new_n224_ = ~i_42_ & new_n223_;
  assign new_n225_ = ~i_38_ & ~i_37_;
  assign new_n226_ = ~i_36_ & new_n225_;
  assign new_n227_ = new_n222_ & new_n224_;
  assign new_n228_ = new_n226_ & new_n227_;
  assign new_n229_ = ~i_53_ & ~i_52_;
  assign new_n230_ = ~i_51_ & new_n229_;
  assign new_n231_ = new_n179_ & new_n230_;
  assign new_n232_ = new_n187_ & new_n231_;
  assign new_n233_ = ~i_32_ & ~i_31_;
  assign new_n234_ = ~i_30_ & new_n233_;
  assign new_n235_ = ~i_28_ & i_29_;
  assign new_n236_ = i_27_ & new_n235_;
  assign new_n237_ = new_n205_ & new_n234_;
  assign new_n238_ = new_n236_ & new_n237_;
  assign new_n239_ = new_n228_ & new_n232_;
  assign new_n240_ = new_n238_ & new_n239_;
  assign new_n241_ = ~i_63_ & ~i_64_;
  assign new_n242_ = ~i_59_ & ~i_58_;
  assign new_n243_ = ~i_57_ & new_n242_;
  assign new_n244_ = ~i_60_ & new_n133_;
  assign new_n245_ = new_n243_ & new_n244_;
  assign new_n246_ = new_n135_ & new_n245_;
  assign new_n247_ = new_n241_ & new_n246_;
  assign new_n248_ = ~i_14_ & ~i_13_;
  assign new_n249_ = ~i_12_ & new_n248_;
  assign new_n250_ = ~i_17_ & ~i_16_;
  assign new_n251_ = ~i_15_ & new_n250_;
  assign new_n252_ = new_n249_ & new_n251_;
  assign new_n253_ = new_n199_ & new_n252_;
  assign new_n254_ = ~i_23_ & ~i_22_;
  assign new_n255_ = ~i_21_ & new_n254_;
  assign new_n256_ = ~i_20_ & ~i_19_;
  assign new_n257_ = ~i_18_ & new_n256_;
  assign new_n258_ = new_n150_ & new_n255_;
  assign new_n259_ = new_n257_ & new_n258_;
  assign new_n260_ = new_n253_ & new_n259_;
  assign new_n261_ = new_n217_ & new_n260_;
  assign new_n262_ = new_n240_ & new_n247_;
  assign o_2_ = new_n261_ & new_n262_;
  assign new_n264_ = ~i_56_ & new_n242_;
  assign new_n265_ = ~i_55_ & ~i_54_;
  assign new_n266_ = ~i_53_ & new_n265_;
  assign new_n267_ = new_n244_ & new_n264_;
  assign new_n268_ = new_n266_ & new_n267_;
  assign new_n269_ = i_45_ & ~i_46_;
  assign new_n270_ = ~i_43_ & new_n269_;
  assign new_n271_ = ~i_50_ & ~i_51_;
  assign new_n272_ = ~i_47_ & new_n271_;
  assign new_n273_ = new_n270_ & new_n272_;
  assign new_n274_ = new_n143_ & new_n273_;
  assign new_n275_ = new_n268_ & new_n274_;
  assign new_n276_ = ~i_5_ & new_n163_;
  assign new_n277_ = new_n166_ & new_n276_;
  assign new_n278_ = new_n168_ & new_n277_;
  assign new_n279_ = new_n171_ & new_n278_;
  assign o_0_ = new_n275_ & new_n279_;
  assign new_n281_ = ~i_50_ & ~i_58_;
  assign new_n282_ = ~i_46_ & new_n281_;
  assign new_n283_ = i_60_ & new_n282_;
  assign new_n284_ = i_29_ & ~i_37_;
  assign new_n285_ = ~i_28_ & new_n284_;
  assign new_n286_ = ~i_40_ & ~i_43_;
  assign new_n287_ = ~i_39_ & new_n286_;
  assign new_n288_ = ~i_10_ & new_n151_;
  assign new_n289_ = new_n285_ & new_n287_;
  assign new_n290_ = new_n288_ & new_n289_;
  assign o_29_ = new_n283_ & new_n290_;
  assign new_n292_ = ~i_50_ & ~i_47_;
  assign new_n293_ = ~i_46_ & new_n292_;
  assign new_n294_ = ~i_30_ & ~i_37_;
  assign new_n295_ = i_29_ & new_n294_;
  assign new_n296_ = new_n287_ & new_n293_;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = ~i_58_ & ~i_60_;
  assign new_n299_ = ~i_56_ & new_n298_;
  assign new_n300_ = ~i_28_ & ~i_25_;
  assign new_n301_ = ~i_24_ & new_n300_;
  assign new_n302_ = ~i_10_ & ~i_8_;
  assign new_n303_ = i_7_ & new_n302_;
  assign new_n304_ = new_n152_ & new_n301_;
  assign new_n305_ = new_n303_ & new_n304_;
  assign new_n306_ = new_n297_ & new_n299_;
  assign o_60_ = new_n305_ & new_n306_;
  assign new_n308_ = ~i_55_ & ~i_51_;
  assign new_n309_ = ~i_50_ & new_n308_;
  assign new_n310_ = new_n133_ & new_n299_;
  assign new_n311_ = new_n309_ & new_n310_;
  assign new_n312_ = ~i_15_ & new_n147_;
  assign new_n313_ = new_n150_ & new_n160_;
  assign new_n314_ = new_n312_ & new_n313_;
  assign new_n315_ = ~i_41_ & i_42_;
  assign new_n316_ = ~i_40_ & new_n315_;
  assign new_n317_ = new_n139_ & new_n316_;
  assign new_n318_ = new_n158_ & new_n317_;
  assign new_n319_ = ~i_14_ & ~i_11_;
  assign new_n320_ = ~i_10_ & new_n319_;
  assign new_n321_ = new_n213_ & new_n320_;
  assign new_n322_ = new_n168_ & new_n321_;
  assign new_n323_ = new_n314_ & new_n318_;
  assign new_n324_ = new_n322_ & new_n323_;
  assign o_39_ = new_n311_ & new_n324_;
  assign new_n326_ = i_59_ & ~i_58_;
  assign new_n327_ = ~i_56_ & new_n326_;
  assign new_n328_ = new_n244_ & new_n327_;
  assign new_n329_ = new_n309_ & new_n328_;
  assign new_n330_ = new_n139_ & new_n143_;
  assign new_n331_ = new_n158_ & new_n330_;
  assign new_n332_ = new_n314_ & new_n331_;
  assign new_n333_ = new_n322_ & new_n332_;
  assign o_38_ = new_n329_ & new_n333_;
  assign new_n335_ = ~i_50_ & new_n298_;
  assign new_n336_ = ~i_46_ & ~i_43_;
  assign new_n337_ = ~i_40_ & new_n336_;
  assign new_n338_ = new_n335_ & new_n337_;
  assign new_n339_ = i_24_ & new_n300_;
  assign new_n340_ = i_29_ & new_n157_;
  assign new_n341_ = new_n339_ & new_n340_;
  assign new_n342_ = new_n288_ & new_n341_;
  assign o_25_ = new_n338_ & new_n342_;
  assign new_n344_ = new_n222_ & new_n295_;
  assign new_n345_ = new_n207_ & new_n344_;
  assign new_n346_ = ~i_58_ & ~i_56_;
  assign new_n347_ = ~i_50_ & new_n346_;
  assign new_n348_ = ~i_62_ & ~i_60_;
  assign new_n349_ = new_n347_ & new_n348_;
  assign new_n350_ = new_n139_ & new_n349_;
  assign new_n351_ = ~i_8_ & new_n198_;
  assign new_n352_ = ~i_24_ & ~i_15_;
  assign new_n353_ = ~i_14_ & new_n352_;
  assign new_n354_ = ~i_7_ & i_6_;
  assign new_n355_ = ~i_3_ & new_n354_;
  assign new_n356_ = new_n351_ & new_n353_;
  assign new_n357_ = new_n355_ & new_n356_;
  assign new_n358_ = new_n345_ & new_n350_;
  assign o_12_ = new_n357_ & new_n358_;
  assign new_n360_ = ~i_45_ & ~i_43_;
  assign new_n361_ = ~i_42_ & new_n360_;
  assign new_n362_ = ~i_47_ & ~i_48_;
  assign new_n363_ = ~i_46_ & new_n362_;
  assign new_n364_ = new_n361_ & new_n363_;
  assign new_n365_ = new_n222_ & new_n364_;
  assign new_n366_ = ~i_52_ & new_n174_;
  assign new_n367_ = ~i_49_ & new_n271_;
  assign new_n368_ = new_n177_ & new_n366_;
  assign new_n369_ = new_n367_ & new_n368_;
  assign new_n370_ = ~i_32_ & new_n155_;
  assign new_n371_ = ~i_36_ & ~i_37_;
  assign new_n372_ = ~i_35_ & new_n371_;
  assign new_n373_ = new_n370_ & new_n372_;
  assign new_n374_ = new_n203_ & new_n373_;
  assign new_n375_ = new_n365_ & new_n369_;
  assign new_n376_ = new_n374_ & new_n375_;
  assign new_n377_ = ~i_63_ & ~i_62_;
  assign new_n378_ = ~i_61_ & new_n377_;
  assign new_n379_ = ~i_64_ & new_n378_;
  assign new_n380_ = new_n132_ & new_n379_;
  assign new_n381_ = ~i_21_ & new_n196_;
  assign new_n382_ = ~i_20_ & i_19_;
  assign new_n383_ = ~i_18_ & new_n382_;
  assign new_n384_ = new_n207_ & new_n381_;
  assign new_n385_ = new_n383_ & new_n384_;
  assign new_n386_ = new_n253_ & new_n385_;
  assign new_n387_ = new_n217_ & new_n386_;
  assign new_n388_ = new_n376_ & new_n380_;
  assign o_37_ = new_n387_ & new_n388_;
  assign new_n390_ = ~i_45_ & ~i_46_;
  assign new_n391_ = ~i_43_ & new_n390_;
  assign new_n392_ = ~i_49_ & ~i_48_;
  assign new_n393_ = ~i_47_ & new_n392_;
  assign new_n394_ = new_n391_ & new_n393_;
  assign new_n395_ = new_n143_ & new_n394_;
  assign new_n396_ = ~i_58_ & ~i_57_;
  assign new_n397_ = ~i_56_ & new_n396_;
  assign new_n398_ = ~i_52_ & ~i_51_;
  assign new_n399_ = ~i_50_ & new_n398_;
  assign new_n400_ = new_n266_ & new_n397_;
  assign new_n401_ = new_n399_ & new_n400_;
  assign new_n402_ = ~i_36_ & new_n157_;
  assign new_n403_ = i_32_ & ~i_31_;
  assign new_n404_ = ~i_30_ & new_n403_;
  assign new_n405_ = new_n205_ & new_n402_;
  assign new_n406_ = new_n404_ & new_n405_;
  assign new_n407_ = new_n395_ & new_n401_;
  assign new_n408_ = new_n406_ & new_n407_;
  assign new_n409_ = ~i_62_ & new_n241_;
  assign new_n410_ = ~i_61_ & ~i_60_;
  assign new_n411_ = ~i_59_ & new_n410_;
  assign new_n412_ = new_n409_ & new_n411_;
  assign new_n413_ = ~i_25_ & ~i_24_;
  assign new_n414_ = ~i_22_ & new_n413_;
  assign new_n415_ = ~i_26_ & new_n235_;
  assign new_n416_ = ~i_20_ & ~i_21_;
  assign new_n417_ = ~i_18_ & new_n416_;
  assign new_n418_ = new_n414_ & new_n415_;
  assign new_n419_ = new_n417_ & new_n418_;
  assign new_n420_ = new_n253_ & new_n419_;
  assign new_n421_ = new_n217_ & new_n420_;
  assign new_n422_ = new_n408_ & new_n412_;
  assign o_26_ = new_n421_ & new_n422_;
  assign new_n424_ = i_29_ & i_37_;
  assign o_11_ = ~i_15_ & new_n424_;
  assign new_n426_ = i_57_ & ~i_56_;
  assign new_n427_ = ~i_55_ & new_n426_;
  assign new_n428_ = new_n175_ & new_n427_;
  assign new_n429_ = new_n179_ & new_n428_;
  assign new_n430_ = new_n136_ & new_n429_;
  assign new_n431_ = new_n191_ & new_n430_;
  assign o_50_ = new_n219_ & new_n431_;
  assign new_n433_ = i_61_ & ~i_62_;
  assign new_n434_ = ~i_60_ & new_n433_;
  assign new_n435_ = ~i_55_ & new_n346_;
  assign new_n436_ = new_n434_ & new_n435_;
  assign new_n437_ = ~i_30_ & ~i_35_;
  assign new_n438_ = i_29_ & new_n437_;
  assign new_n439_ = new_n207_ & new_n438_;
  assign new_n440_ = new_n197_ & new_n439_;
  assign new_n441_ = ~i_41_ & new_n336_;
  assign new_n442_ = new_n272_ & new_n441_;
  assign new_n443_ = new_n189_ & new_n442_;
  assign new_n444_ = ~i_7_ & new_n302_;
  assign new_n445_ = ~i_6_ & ~i_3_;
  assign new_n446_ = ~i_0_ & new_n445_;
  assign new_n447_ = new_n152_ & new_n444_;
  assign new_n448_ = new_n446_ & new_n447_;
  assign new_n449_ = new_n440_ & new_n443_;
  assign new_n450_ = new_n448_ & new_n449_;
  assign o_36_ = new_n436_ & new_n450_;
  assign new_n452_ = new_n179_ & new_n187_;
  assign new_n453_ = new_n186_ & new_n452_;
  assign new_n454_ = new_n135_ & new_n243_;
  assign new_n455_ = new_n230_ & new_n454_;
  assign new_n456_ = ~i_36_ & ~i_35_;
  assign new_n457_ = ~i_34_ & new_n456_;
  assign new_n458_ = ~i_31_ & ~i_33_;
  assign new_n459_ = ~i_30_ & new_n458_;
  assign new_n460_ = new_n189_ & new_n457_;
  assign new_n461_ = new_n459_ & new_n460_;
  assign new_n462_ = new_n453_ & new_n455_;
  assign new_n463_ = new_n461_ & new_n462_;
  assign new_n464_ = new_n241_ & new_n244_;
  assign new_n465_ = ~i_14_ & i_13_;
  assign new_n466_ = ~i_12_ & new_n465_;
  assign new_n467_ = new_n251_ & new_n466_;
  assign new_n468_ = new_n199_ & new_n467_;
  assign new_n469_ = new_n419_ & new_n468_;
  assign new_n470_ = new_n217_ & new_n469_;
  assign new_n471_ = new_n463_ & new_n464_;
  assign o_27_ = new_n470_ & new_n471_;
  assign new_n473_ = i_50_ & ~i_58_;
  assign new_n474_ = ~i_43_ & new_n473_;
  assign new_n475_ = new_n285_ & new_n474_;
  assign o_14_ = new_n288_ & new_n475_;
  assign new_n477_ = ~i_58_ & new_n410_;
  assign new_n478_ = ~i_51_ & new_n134_;
  assign new_n479_ = ~i_62_ & new_n477_;
  assign new_n480_ = new_n478_ & new_n479_;
  assign new_n481_ = ~i_41_ & ~i_43_;
  assign new_n482_ = ~i_40_ & new_n481_;
  assign new_n483_ = new_n293_ & new_n482_;
  assign new_n484_ = new_n158_ & new_n483_;
  assign new_n485_ = ~i_3_ & i_4_;
  assign new_n486_ = ~i_0_ & new_n485_;
  assign new_n487_ = new_n321_ & new_n486_;
  assign new_n488_ = new_n314_ & new_n484_;
  assign new_n489_ = new_n487_ & new_n488_;
  assign o_35_ = new_n480_ & new_n489_;
  assign new_n491_ = ~i_50_ & ~i_46_;
  assign new_n492_ = ~i_43_ & new_n491_;
  assign new_n493_ = new_n298_ & new_n492_;
  assign new_n494_ = i_25_ & new_n235_;
  assign new_n495_ = new_n189_ & new_n494_;
  assign new_n496_ = new_n288_ & new_n495_;
  assign o_28_ = new_n493_ & new_n496_;
  assign new_n498_ = ~i_30_ & new_n157_;
  assign new_n499_ = i_41_ & ~i_43_;
  assign new_n500_ = ~i_40_ & new_n499_;
  assign new_n501_ = new_n498_ & new_n500_;
  assign new_n502_ = new_n415_ & new_n501_;
  assign new_n503_ = ~i_62_ & new_n299_;
  assign new_n504_ = new_n293_ & new_n503_;
  assign new_n505_ = ~i_15_ & new_n413_;
  assign new_n506_ = ~i_3_ & new_n212_;
  assign new_n507_ = new_n320_ & new_n505_;
  assign new_n508_ = new_n506_ & new_n507_;
  assign new_n509_ = new_n502_ & new_n504_;
  assign o_13_ = new_n508_ & new_n509_;
  assign new_n511_ = ~i_43_ & ~i_37_;
  assign new_n512_ = i_29_ & new_n511_;
  assign new_n513_ = ~i_28_ & ~i_15_;
  assign new_n514_ = ~i_14_ & new_n513_;
  assign new_n515_ = i_58_ & new_n512_;
  assign o_34_ = new_n514_ & new_n515_;
  assign new_n517_ = new_n207_ & new_n295_;
  assign new_n518_ = new_n197_ & new_n517_;
  assign new_n519_ = new_n139_ & new_n347_;
  assign new_n520_ = new_n222_ & new_n519_;
  assign new_n521_ = i_0_ & new_n445_;
  assign new_n522_ = new_n447_ & new_n521_;
  assign new_n523_ = new_n518_ & new_n520_;
  assign new_n524_ = new_n522_ & new_n523_;
  assign o_21_ = new_n348_ & new_n524_;
  assign new_n526_ = i_26_ & new_n235_;
  assign new_n527_ = new_n337_ & new_n498_;
  assign new_n528_ = new_n526_ & new_n527_;
  assign new_n529_ = ~i_58_ & new_n348_;
  assign new_n530_ = ~i_50_ & ~i_56_;
  assign new_n531_ = ~i_47_ & new_n530_;
  assign new_n532_ = new_n529_ & new_n531_;
  assign new_n533_ = new_n528_ & new_n532_;
  assign o_16_ = new_n508_ & new_n533_;
  assign new_n535_ = i_54_ & new_n134_;
  assign new_n536_ = ~i_42_ & new_n336_;
  assign new_n537_ = new_n272_ & new_n535_;
  assign new_n538_ = new_n536_ & new_n537_;
  assign new_n539_ = new_n136_ & new_n538_;
  assign new_n540_ = new_n197_ & new_n207_;
  assign new_n541_ = new_n195_ & new_n540_;
  assign new_n542_ = ~i_35_ & ~i_37_;
  assign new_n543_ = ~i_34_ & new_n542_;
  assign new_n544_ = ~i_30_ & ~i_33_;
  assign new_n545_ = i_29_ & new_n544_;
  assign new_n546_ = new_n222_ & new_n543_;
  assign new_n547_ = new_n545_ & new_n546_;
  assign new_n548_ = new_n199_ & new_n213_;
  assign new_n549_ = new_n168_ & new_n548_;
  assign new_n550_ = new_n541_ & new_n547_;
  assign new_n551_ = new_n549_ & new_n550_;
  assign o_40_ = new_n539_ & new_n551_;
  assign new_n553_ = i_39_ & new_n286_;
  assign new_n554_ = new_n285_ & new_n553_;
  assign new_n555_ = new_n288_ & new_n554_;
  assign o_33_ = new_n281_ & new_n555_;
  assign new_n557_ = new_n266_ & new_n367_;
  assign new_n558_ = new_n363_ & new_n557_;
  assign new_n559_ = new_n397_ & new_n412_;
  assign new_n560_ = i_36_ & ~i_37_;
  assign new_n561_ = ~i_35_ & new_n560_;
  assign new_n562_ = new_n222_ & new_n361_;
  assign new_n563_ = new_n561_ & new_n562_;
  assign new_n564_ = new_n558_ & new_n559_;
  assign new_n565_ = new_n563_ & new_n564_;
  assign new_n566_ = ~i_12_ & new_n151_;
  assign new_n567_ = new_n148_ & new_n566_;
  assign new_n568_ = new_n199_ & new_n567_;
  assign new_n569_ = new_n156_ & new_n160_;
  assign new_n570_ = new_n150_ & new_n569_;
  assign new_n571_ = new_n568_ & new_n570_;
  assign new_n572_ = new_n217_ & new_n571_;
  assign o_22_ = new_n565_ & new_n572_;
  assign new_n574_ = ~i_58_ & ~i_43_;
  assign new_n575_ = i_10_ & new_n151_;
  assign new_n576_ = new_n285_ & new_n574_;
  assign o_15_ = new_n575_ & new_n576_;
  assign new_n578_ = i_46_ & new_n281_;
  assign o_32_ = new_n290_ & new_n578_;
  assign new_n580_ = new_n393_ & new_n399_;
  assign new_n581_ = new_n391_ & new_n580_;
  assign new_n582_ = new_n397_ & new_n411_;
  assign new_n583_ = new_n266_ & new_n582_;
  assign new_n584_ = new_n143_ & new_n402_;
  assign new_n585_ = new_n205_ & new_n584_;
  assign new_n586_ = new_n581_ & new_n583_;
  assign new_n587_ = new_n585_ & new_n586_;
  assign new_n588_ = ~i_18_ & ~i_17_;
  assign new_n589_ = i_16_ & new_n588_;
  assign new_n590_ = new_n566_ & new_n589_;
  assign new_n591_ = new_n199_ & new_n590_;
  assign new_n592_ = new_n203_ & new_n207_;
  assign new_n593_ = new_n381_ & new_n592_;
  assign new_n594_ = new_n591_ & new_n593_;
  assign new_n595_ = new_n217_ & new_n594_;
  assign new_n596_ = new_n409_ & new_n587_;
  assign o_23_ = new_n595_ & new_n596_;
  assign new_n598_ = i_62_ & new_n299_;
  assign new_n599_ = new_n304_ & new_n444_;
  assign new_n600_ = new_n297_ & new_n598_;
  assign o_18_ = new_n599_ & new_n600_;
  assign new_n602_ = new_n175_ & new_n179_;
  assign new_n603_ = new_n187_ & new_n602_;
  assign new_n604_ = new_n132_ & new_n378_;
  assign new_n605_ = new_n177_ & new_n604_;
  assign new_n606_ = new_n186_ & new_n189_;
  assign new_n607_ = new_n457_ & new_n606_;
  assign new_n608_ = new_n603_ & new_n605_;
  assign new_n609_ = new_n607_ & new_n608_;
  assign new_n610_ = ~i_18_ & i_21_;
  assign new_n611_ = ~i_17_ & new_n610_;
  assign new_n612_ = new_n566_ & new_n611_;
  assign new_n613_ = new_n199_ & new_n612_;
  assign new_n614_ = new_n415_ & new_n459_;
  assign new_n615_ = new_n414_ & new_n614_;
  assign new_n616_ = new_n613_ & new_n615_;
  assign new_n617_ = new_n217_ & new_n616_;
  assign new_n618_ = ~i_64_ & new_n609_;
  assign o_31_ = new_n617_ & new_n618_;
  assign new_n620_ = ~i_60_ & new_n282_;
  assign new_n621_ = new_n287_ & new_n620_;
  assign new_n622_ = ~i_14_ & i_11_;
  assign new_n623_ = ~i_10_ & new_n622_;
  assign new_n624_ = new_n285_ & new_n505_;
  assign new_n625_ = new_n623_ & new_n624_;
  assign o_24_ = new_n621_ & new_n625_;
  assign new_n627_ = new_n139_ & new_n189_;
  assign new_n628_ = new_n160_ & new_n627_;
  assign new_n629_ = i_3_ & new_n212_;
  assign new_n630_ = new_n507_ & new_n629_;
  assign new_n631_ = new_n349_ & new_n628_;
  assign o_17_ = new_n630_ & new_n631_;
  assign new_n633_ = new_n363_ & new_n367_;
  assign new_n634_ = new_n361_ & new_n633_;
  assign new_n635_ = new_n132_ & new_n177_;
  assign new_n636_ = new_n366_ & new_n635_;
  assign new_n637_ = new_n222_ & new_n372_;
  assign new_n638_ = new_n156_ & new_n637_;
  assign new_n639_ = new_n634_ & new_n636_;
  assign new_n640_ = new_n638_ & new_n639_;
  assign new_n641_ = ~i_16_ & new_n588_;
  assign new_n642_ = new_n566_ & new_n641_;
  assign new_n643_ = new_n199_ & new_n642_;
  assign new_n644_ = ~i_21_ & ~i_22_;
  assign new_n645_ = i_20_ & new_n644_;
  assign new_n646_ = new_n313_ & new_n645_;
  assign new_n647_ = new_n643_ & new_n646_;
  assign new_n648_ = new_n217_ & new_n647_;
  assign new_n649_ = new_n379_ & new_n640_;
  assign o_56_ = new_n648_ & new_n649_;
  assign new_n651_ = new_n132_ & new_n135_;
  assign new_n652_ = new_n141_ & new_n651_;
  assign new_n653_ = new_n133_ & new_n652_;
  assign new_n654_ = new_n191_ & new_n653_;
  assign new_n655_ = i_1_ & ~i_2_;
  assign new_n656_ = ~i_0_ & new_n655_;
  assign new_n657_ = new_n216_ & new_n656_;
  assign new_n658_ = new_n218_ & new_n657_;
  assign o_43_ = new_n654_ & new_n658_;
  assign new_n660_ = ~i_53_ & i_52_;
  assign new_n661_ = ~i_51_ & new_n660_;
  assign new_n662_ = new_n179_ & new_n661_;
  assign new_n663_ = new_n187_ & new_n662_;
  assign new_n664_ = new_n246_ & new_n663_;
  assign new_n665_ = new_n607_ & new_n664_;
  assign new_n666_ = ~i_18_ & ~i_21_;
  assign new_n667_ = ~i_17_ & new_n666_;
  assign new_n668_ = new_n566_ & new_n667_;
  assign new_n669_ = new_n199_ & new_n668_;
  assign new_n670_ = new_n615_ & new_n669_;
  assign new_n671_ = new_n217_ & new_n670_;
  assign new_n672_ = new_n241_ & new_n665_;
  assign o_30_ = new_n671_ & new_n672_;
  assign new_n674_ = ~i_30_ & i_35_;
  assign new_n675_ = i_29_ & new_n674_;
  assign new_n676_ = new_n207_ & new_n675_;
  assign new_n677_ = new_n197_ & new_n676_;
  assign new_n678_ = new_n443_ & new_n677_;
  assign new_n679_ = new_n448_ & new_n678_;
  assign o_55_ = new_n503_ & new_n679_;
  assign new_n681_ = new_n411_ & new_n435_;
  assign new_n682_ = new_n175_ & new_n681_;
  assign new_n683_ = new_n293_ & new_n361_;
  assign new_n684_ = new_n222_ & new_n683_;
  assign new_n685_ = ~i_62_ & new_n682_;
  assign new_n686_ = new_n684_ & new_n685_;
  assign new_n687_ = ~i_15_ & new_n588_;
  assign new_n688_ = new_n414_ & new_n687_;
  assign new_n689_ = new_n320_ & new_n688_;
  assign new_n690_ = new_n459_ & new_n543_;
  assign new_n691_ = new_n415_ & new_n690_;
  assign new_n692_ = ~i_5_ & ~i_6_;
  assign new_n693_ = ~i_4_ & new_n692_;
  assign new_n694_ = ~i_9_ & ~i_8_;
  assign new_n695_ = ~i_7_ & new_n694_;
  assign new_n696_ = ~i_3_ & i_2_;
  assign new_n697_ = ~i_0_ & new_n696_;
  assign new_n698_ = new_n693_ & new_n695_;
  assign new_n699_ = new_n697_ & new_n698_;
  assign new_n700_ = new_n689_ & new_n691_;
  assign new_n701_ = new_n699_ & new_n700_;
  assign o_44_ = new_n686_ & new_n701_;
  assign new_n703_ = new_n160_ & new_n189_;
  assign new_n704_ = new_n150_ & new_n703_;
  assign new_n705_ = new_n441_ & new_n532_;
  assign new_n706_ = i_22_ & ~i_15_;
  assign new_n707_ = ~i_14_ & new_n706_;
  assign new_n708_ = ~i_3_ & new_n163_;
  assign new_n709_ = new_n351_ & new_n707_;
  assign new_n710_ = new_n708_ & new_n709_;
  assign new_n711_ = new_n704_ & new_n705_;
  assign o_58_ = new_n710_ & new_n711_;
  assign new_n713_ = ~i_62_ & new_n411_;
  assign new_n714_ = new_n272_ & new_n435_;
  assign new_n715_ = new_n536_ & new_n714_;
  assign new_n716_ = new_n713_ & new_n715_;
  assign new_n717_ = ~i_30_ & i_33_;
  assign new_n718_ = i_29_ & new_n717_;
  assign new_n719_ = new_n546_ & new_n718_;
  assign new_n720_ = new_n541_ & new_n719_;
  assign new_n721_ = new_n549_ & new_n720_;
  assign o_41_ = new_n716_ & new_n721_;
  assign new_n723_ = new_n415_ & new_n498_;
  assign new_n724_ = new_n414_ & new_n723_;
  assign new_n725_ = new_n293_ & new_n299_;
  assign new_n726_ = new_n482_ & new_n725_;
  assign new_n727_ = i_18_ & ~i_15_;
  assign new_n728_ = ~i_14_ & new_n727_;
  assign new_n729_ = new_n351_ & new_n728_;
  assign new_n730_ = new_n708_ & new_n729_;
  assign new_n731_ = new_n724_ & new_n726_;
  assign new_n732_ = new_n730_ & new_n731_;
  assign o_57_ = ~i_62_ & new_n732_;
  assign new_n734_ = i_49_ & new_n271_;
  assign new_n735_ = new_n264_ & new_n266_;
  assign new_n736_ = new_n734_ & new_n735_;
  assign new_n737_ = new_n244_ & new_n736_;
  assign new_n738_ = new_n191_ & new_n737_;
  assign o_42_ = new_n219_ & new_n738_;
  assign new_n740_ = ~i_56_ & i_51_;
  assign new_n741_ = ~i_50_ & new_n740_;
  assign new_n742_ = new_n139_ & new_n741_;
  assign new_n743_ = new_n222_ & new_n742_;
  assign new_n744_ = new_n518_ & new_n743_;
  assign new_n745_ = new_n448_ & new_n744_;
  assign o_20_ = new_n529_ & new_n745_;
  assign new_n747_ = new_n135_ & new_n141_;
  assign new_n748_ = new_n393_ & new_n747_;
  assign new_n749_ = new_n243_ & new_n464_;
  assign new_n750_ = new_n143_ & new_n391_;
  assign new_n751_ = new_n158_ & new_n750_;
  assign new_n752_ = new_n748_ & new_n749_;
  assign new_n753_ = new_n751_ & new_n752_;
  assign new_n754_ = i_12_ & new_n151_;
  assign new_n755_ = new_n148_ & new_n754_;
  assign new_n756_ = new_n199_ & new_n755_;
  assign new_n757_ = new_n570_ & new_n756_;
  assign new_n758_ = new_n217_ & new_n757_;
  assign o_52_ = new_n753_ & new_n758_;
  assign new_n760_ = new_n272_ & new_n681_;
  assign new_n761_ = ~i_62_ & new_n760_;
  assign new_n762_ = ~i_18_ & i_17_;
  assign new_n763_ = ~i_15_ & new_n762_;
  assign new_n764_ = new_n418_ & new_n763_;
  assign new_n765_ = ~i_30_ & new_n542_;
  assign new_n766_ = new_n222_ & new_n536_;
  assign new_n767_ = new_n765_ & new_n766_;
  assign new_n768_ = new_n764_ & new_n767_;
  assign new_n769_ = new_n322_ & new_n768_;
  assign o_47_ = new_n761_ & new_n769_;
  assign new_n771_ = i_48_ & new_n178_;
  assign new_n772_ = new_n175_ & new_n435_;
  assign new_n773_ = new_n771_ & new_n772_;
  assign new_n774_ = new_n713_ & new_n773_;
  assign new_n775_ = new_n191_ & new_n774_;
  assign o_51_ = new_n219_ & new_n775_;
  assign new_n777_ = new_n435_ & new_n713_;
  assign new_n778_ = new_n175_ & new_n293_;
  assign new_n779_ = new_n186_ & new_n778_;
  assign new_n780_ = new_n777_ & new_n779_;
  assign new_n781_ = ~i_30_ & i_31_;
  assign new_n782_ = i_29_ & new_n781_;
  assign new_n783_ = new_n189_ & new_n205_;
  assign new_n784_ = new_n782_ & new_n783_;
  assign new_n785_ = new_n541_ & new_n784_;
  assign new_n786_ = new_n549_ & new_n785_;
  assign o_48_ = new_n780_ & new_n786_;
  assign new_n788_ = i_55_ & new_n346_;
  assign new_n789_ = new_n348_ & new_n788_;
  assign o_54_ = new_n450_ & new_n789_;
  assign new_n791_ = new_n264_ & new_n309_;
  assign new_n792_ = new_n139_ & new_n791_;
  assign new_n793_ = new_n244_ & new_n792_;
  assign new_n794_ = ~i_30_ & i_34_;
  assign new_n795_ = i_29_ & new_n794_;
  assign new_n796_ = new_n143_ & new_n158_;
  assign new_n797_ = new_n795_ & new_n796_;
  assign new_n798_ = new_n541_ & new_n797_;
  assign new_n799_ = new_n549_ & new_n798_;
  assign o_45_ = new_n793_ & new_n799_;
  assign new_n801_ = i_28_ & i_29_;
  assign new_n802_ = ~i_15_ & new_n801_;
  assign o_10_ = ~i_37_ & new_n802_;
  assign new_n804_ = i_63_ & ~i_62_;
  assign new_n805_ = ~i_61_ & new_n804_;
  assign new_n806_ = ~i_64_ & new_n805_;
  assign new_n807_ = new_n132_ & new_n806_;
  assign new_n808_ = new_n181_ & new_n807_;
  assign new_n809_ = new_n191_ & new_n808_;
  assign o_53_ = new_n219_ & new_n809_;
  assign new_n811_ = new_n132_ & new_n478_;
  assign new_n812_ = new_n293_ & new_n811_;
  assign new_n813_ = new_n133_ & new_n812_;
  assign new_n814_ = new_n438_ & new_n606_;
  assign new_n815_ = i_9_ & new_n198_;
  assign new_n816_ = new_n213_ & new_n815_;
  assign new_n817_ = new_n168_ & new_n816_;
  assign new_n818_ = new_n541_ & new_n814_;
  assign new_n819_ = new_n817_ & new_n818_;
  assign o_46_ = new_n813_ & new_n819_;
  assign new_n821_ = new_n337_ & new_n531_;
  assign new_n822_ = new_n498_ & new_n821_;
  assign new_n823_ = ~i_25_ & new_n235_;
  assign new_n824_ = i_8_ & new_n198_;
  assign new_n825_ = new_n353_ & new_n823_;
  assign new_n826_ = new_n824_ & new_n825_;
  assign new_n827_ = new_n298_ & new_n822_;
  assign o_61_ = new_n826_ & new_n827_;
  assign new_n829_ = new_n135_ & new_n230_;
  assign new_n830_ = new_n179_ & new_n829_;
  assign new_n831_ = ~i_32_ & ~i_33_;
  assign new_n832_ = ~i_31_ & new_n831_;
  assign new_n833_ = new_n457_ & new_n832_;
  assign new_n834_ = new_n160_ & new_n833_;
  assign new_n835_ = new_n191_ & new_n830_;
  assign new_n836_ = new_n834_ & new_n835_;
  assign new_n837_ = i_23_ & ~i_22_;
  assign new_n838_ = ~i_21_ & new_n837_;
  assign new_n839_ = new_n150_ & new_n838_;
  assign new_n840_ = new_n257_ & new_n839_;
  assign new_n841_ = new_n253_ & new_n840_;
  assign new_n842_ = new_n217_ & new_n841_;
  assign new_n843_ = new_n749_ & new_n836_;
  assign o_9_ = new_n842_ & new_n843_;
  assign new_n845_ = ~i_46_ & i_47_;
  assign new_n846_ = ~i_43_ & new_n845_;
  assign new_n847_ = new_n347_ & new_n846_;
  assign new_n848_ = new_n189_ & new_n847_;
  assign new_n849_ = new_n160_ & new_n505_;
  assign new_n850_ = new_n320_ & new_n849_;
  assign new_n851_ = ~i_60_ & new_n848_;
  assign o_62_ = new_n850_ & new_n851_;
  assign new_n853_ = i_56_ & new_n298_;
  assign new_n854_ = new_n492_ & new_n853_;
  assign new_n855_ = new_n189_ & new_n854_;
  assign o_63_ = new_n850_ & new_n855_;
  assign new_n857_ = i_53_ & new_n265_;
  assign new_n858_ = new_n272_ & new_n857_;
  assign new_n859_ = new_n536_ & new_n858_;
  assign new_n860_ = new_n267_ & new_n859_;
  assign o_49_ = new_n551_ & new_n860_;
  assign new_n862_ = i_43_ & ~i_37_;
  assign new_n863_ = ~i_15_ & new_n235_;
  assign o_7_ = new_n862_ & new_n863_;
  assign new_n865_ = new_n189_ & new_n493_;
  assign new_n866_ = i_30_ & i_29_;
  assign new_n867_ = ~i_28_ & new_n866_;
  assign new_n868_ = new_n505_ & new_n867_;
  assign new_n869_ = new_n320_ & new_n868_;
  assign o_64_ = new_n865_ & new_n869_;
  assign new_n871_ = ~i_39_ & i_38_;
  assign new_n872_ = ~i_37_ & new_n871_;
  assign new_n873_ = new_n750_ & new_n872_;
  assign new_n874_ = new_n266_ & new_n399_;
  assign new_n875_ = new_n393_ & new_n874_;
  assign new_n876_ = new_n873_ & new_n875_;
  assign new_n877_ = new_n834_ & new_n876_;
  assign new_n878_ = new_n559_ & new_n877_;
  assign o_8_ = new_n261_ & new_n878_;
  assign new_n880_ = ~i_50_ & ~i_43_;
  assign new_n881_ = i_40_ & new_n880_;
  assign new_n882_ = new_n285_ & new_n881_;
  assign new_n883_ = new_n288_ & new_n882_;
  assign o_59_ = ~i_58_ & new_n883_;
  assign new_n885_ = i_14_ & new_n513_;
  assign o_6_ = new_n512_ & new_n885_;
  assign new_n887_ = ~i_45_ & i_44_;
  assign new_n888_ = ~i_43_ & new_n887_;
  assign new_n889_ = ~i_39_ & ~i_38_;
  assign new_n890_ = ~i_37_ & new_n889_;
  assign new_n891_ = new_n143_ & new_n888_;
  assign new_n892_ = new_n890_ & new_n891_;
  assign new_n893_ = new_n366_ & new_n367_;
  assign new_n894_ = new_n363_ & new_n893_;
  assign new_n895_ = new_n892_ & new_n894_;
  assign new_n896_ = new_n834_ & new_n895_;
  assign new_n897_ = ~i_64_ & new_n605_;
  assign new_n898_ = new_n896_ & new_n897_;
  assign o_3_ = new_n261_ & new_n898_;
  assign o_4_ = i_15_ & i_29_;
  assign o_5_ = i_29_;
endmodule

