module pcler8_cl ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0,
    b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0;
  output b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0;
  wire new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n63_, new_n64_, new_n65_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_;
  assign new_n45_ = t & u;
  assign new_n46_ = v & new_n45_;
  assign new_n47_ = w & new_n46_;
  assign new_n48_ = x & new_n47_;
  assign new_n49_ = y & new_n48_;
  assign new_n50_ = z & new_n49_;
  assign new_n51_ = ~i & j;
  assign new_n52_ = ~k & new_n51_;
  assign new_n53_ = a0 & new_n50_;
  assign b0 = new_n52_ & new_n53_;
  assign c0 = a & i;
  assign d0 = b & i;
  assign e0 = c & i;
  assign f0 = d & i;
  assign g0 = e & i;
  assign h0 = f & i;
  assign i0 = g & i;
  assign j0 = h & i;
  assign new_n63_ = l & b0;
  assign new_n64_ = ~t & new_n52_;
  assign new_n65_ = ~new_n63_ & ~new_n64_;
  assign k0 = c0 | ~new_n65_;
  assign new_n67_ = ~t & u;
  assign new_n68_ = t & ~u;
  assign new_n69_ = ~new_n67_ & ~new_n68_;
  assign new_n70_ = new_n52_ & ~new_n69_;
  assign new_n71_ = m & b0;
  assign new_n72_ = ~d0 & ~new_n71_;
  assign l0 = new_n70_ | ~new_n72_;
  assign new_n74_ = ~v & new_n45_;
  assign new_n75_ = v & ~new_n45_;
  assign new_n76_ = ~new_n74_ & ~new_n75_;
  assign new_n77_ = new_n52_ & ~new_n76_;
  assign new_n78_ = n & b0;
  assign new_n79_ = ~e0 & ~new_n78_;
  assign m0 = new_n77_ | ~new_n79_;
  assign new_n81_ = ~w & new_n46_;
  assign new_n82_ = w & ~new_n46_;
  assign new_n83_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = new_n52_ & ~new_n83_;
  assign new_n85_ = o & b0;
  assign new_n86_ = ~f0 & ~new_n85_;
  assign n0 = new_n84_ | ~new_n86_;
  assign new_n88_ = ~x & new_n47_;
  assign new_n89_ = x & ~new_n47_;
  assign new_n90_ = ~new_n88_ & ~new_n89_;
  assign new_n91_ = new_n52_ & ~new_n90_;
  assign new_n92_ = p & b0;
  assign new_n93_ = ~g0 & ~new_n92_;
  assign o0 = new_n91_ | ~new_n93_;
  assign new_n95_ = ~y & new_n48_;
  assign new_n96_ = y & ~new_n48_;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign new_n98_ = new_n52_ & ~new_n97_;
  assign new_n99_ = q & b0;
  assign new_n100_ = ~h0 & ~new_n99_;
  assign p0 = new_n98_ | ~new_n100_;
  assign new_n102_ = ~z & new_n49_;
  assign new_n103_ = z & ~new_n49_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = new_n52_ & ~new_n104_;
  assign new_n106_ = r & b0;
  assign new_n107_ = ~i0 & ~new_n106_;
  assign q0 = new_n105_ | ~new_n107_;
  assign new_n109_ = ~a0 & new_n50_;
  assign new_n110_ = a0 & ~new_n50_;
  assign new_n111_ = ~new_n109_ & ~new_n110_;
  assign new_n112_ = new_n52_ & ~new_n111_;
  assign new_n113_ = s & b0;
  assign new_n114_ = ~j0 & ~new_n113_;
  assign r0 = new_n112_ | ~new_n114_;
endmodule

