module top ( 
    v_6_, v_7_, v_4_, v_5_, v_2_, v_3_, v_0_, v_1_,
    sqrt_3_, sqrt_2_, sqrt_1_, sqrt_0_  );
  input  v_6_, v_7_, v_4_, v_5_, v_2_, v_3_, v_0_, v_1_;
  output sqrt_3_, sqrt_2_, sqrt_1_, sqrt_0_;
  wire new_n14_, new_n15_, new_n16_, new_n17_, new_n19_, new_n20_, new_n21_,
    new_n22_, new_n23_, new_n24_, new_n25_, new_n26_, new_n27_, new_n28_,
    new_n29_, new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_,
    new_n36_, new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_,
    new_n43_, new_n44_, new_n45_, new_n46_, new_n48_, new_n49_, new_n50_,
    new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_,
    new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_,
    new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_;
  assign sqrt_3_ = v_6_ | v_7_;
  assign new_n14_ = ~v_6_ & v_5_;
  assign new_n15_ = ~v_6_ & v_4_;
  assign new_n16_ = v_6_ & v_7_;
  assign new_n17_ = ~new_n14_ & ~new_n15_;
  assign sqrt_2_ = new_n16_ | ~new_n17_;
  assign new_n19_ = v_5_ & v_2_;
  assign new_n20_ = ~v_7_ & new_n19_;
  assign new_n21_ = ~v_4_ & ~v_5_;
  assign new_n22_ = ~v_6_ & new_n21_;
  assign new_n23_ = v_3_ & new_n22_;
  assign new_n24_ = v_5_ & v_3_;
  assign new_n25_ = ~v_7_ & new_n24_;
  assign new_n26_ = v_7_ & new_n21_;
  assign new_n27_ = v_3_ & new_n26_;
  assign new_n28_ = ~new_n23_ & ~new_n25_;
  assign new_n29_ = ~new_n27_ & new_n28_;
  assign new_n30_ = v_2_ & new_n22_;
  assign new_n31_ = v_6_ & v_4_;
  assign new_n32_ = v_7_ & new_n31_;
  assign new_n33_ = v_2_ & new_n26_;
  assign new_n34_ = ~new_n30_ & ~new_n32_;
  assign new_n35_ = ~new_n33_ & new_n34_;
  assign new_n36_ = v_6_ & v_5_;
  assign new_n37_ = v_7_ & new_n36_;
  assign new_n38_ = v_4_ & v_5_;
  assign new_n39_ = ~v_7_ & new_n38_;
  assign new_n40_ = ~v_6_ & ~v_5_;
  assign new_n41_ = v_7_ & new_n40_;
  assign new_n42_ = ~v_4_ & new_n41_;
  assign new_n43_ = ~new_n37_ & ~new_n39_;
  assign new_n44_ = ~new_n42_ & new_n43_;
  assign new_n45_ = new_n29_ & new_n35_;
  assign new_n46_ = new_n44_ & new_n45_;
  assign sqrt_1_ = new_n20_ | ~new_n46_;
  assign new_n48_ = v_4_ & v_0_;
  assign new_n49_ = v_6_ & ~v_5_;
  assign new_n50_ = ~v_7_ & new_n49_;
  assign new_n51_ = new_n48_ & new_n50_;
  assign new_n52_ = ~v_2_ & v_0_;
  assign new_n53_ = ~v_3_ & new_n52_;
  assign new_n54_ = ~v_4_ & v_5_;
  assign new_n55_ = v_6_ & new_n54_;
  assign new_n56_ = new_n53_ & new_n55_;
  assign new_n57_ = ~new_n42_ & ~new_n51_;
  assign new_n58_ = ~new_n56_ & new_n57_;
  assign new_n59_ = v_4_ & v_3_;
  assign new_n60_ = ~v_7_ & new_n59_;
  assign new_n61_ = v_1_ & new_n60_;
  assign new_n62_ = new_n22_ & new_n52_;
  assign new_n63_ = v_2_ & new_n37_;
  assign new_n64_ = ~new_n61_ & ~new_n62_;
  assign new_n65_ = ~new_n63_ & new_n64_;
  assign new_n66_ = v_7_ & new_n24_;
  assign new_n67_ = v_1_ & new_n66_;
  assign new_n68_ = ~v_6_ & new_n38_;
  assign new_n69_ = v_1_ & new_n68_;
  assign new_n70_ = ~v_2_ & v_1_;
  assign new_n71_ = new_n22_ & new_n70_;
  assign new_n72_ = ~new_n67_ & ~new_n69_;
  assign new_n73_ = ~new_n71_ & new_n72_;
  assign new_n74_ = new_n58_ & new_n65_;
  assign new_n75_ = new_n73_ & new_n74_;
  assign new_n76_ = ~v_2_ & ~v_3_;
  assign new_n77_ = ~v_7_ & new_n54_;
  assign new_n78_ = new_n76_ & new_n77_;
  assign new_n79_ = v_2_ & v_3_;
  assign new_n80_ = new_n22_ & new_n79_;
  assign new_n81_ = new_n26_ & new_n76_;
  assign new_n82_ = ~new_n78_ & ~new_n80_;
  assign new_n83_ = ~new_n81_ & new_n82_;
  assign new_n84_ = v_0_ & new_n60_;
  assign new_n85_ = v_0_ & new_n68_;
  assign new_n86_ = v_7_ & new_n38_;
  assign new_n87_ = v_0_ & new_n66_;
  assign new_n88_ = ~new_n85_ & ~new_n86_;
  assign new_n89_ = ~new_n87_ & new_n88_;
  assign new_n90_ = new_n83_ & ~new_n84_;
  assign new_n91_ = new_n89_ & new_n90_;
  assign new_n92_ = v_2_ & new_n68_;
  assign new_n93_ = v_2_ & new_n66_;
  assign new_n94_ = v_3_ & new_n68_;
  assign new_n95_ = ~new_n92_ & ~new_n93_;
  assign new_n96_ = ~new_n94_ & new_n95_;
  assign new_n97_ = v_4_ & v_1_;
  assign new_n98_ = new_n50_ & new_n97_;
  assign new_n99_ = v_2_ & new_n60_;
  assign new_n100_ = ~v_3_ & new_n70_;
  assign new_n101_ = new_n55_ & new_n100_;
  assign new_n102_ = ~new_n98_ & ~new_n99_;
  assign new_n103_ = ~new_n101_ & new_n102_;
  assign new_n104_ = new_n50_ & new_n59_;
  assign new_n105_ = v_4_ & v_2_;
  assign new_n106_ = new_n50_ & new_n105_;
  assign new_n107_ = v_3_ & new_n37_;
  assign new_n108_ = ~new_n104_ & ~new_n106_;
  assign new_n109_ = ~new_n107_ & new_n108_;
  assign new_n110_ = new_n96_ & new_n103_;
  assign new_n111_ = new_n109_ & new_n110_;
  assign new_n112_ = new_n75_ & new_n91_;
  assign sqrt_0_ = ~new_n111_ | ~new_n112_;
endmodule

