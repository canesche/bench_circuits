module top ( clock, 
    pa, pclk, pb, pc, pd, pe, pf, pg,
    pt, pu, pv, pw  );
  input  clock;
  input  pa, pclk, pb, pc, pd, pe, pf, pg;
  output pt, pu, pv, pw;
  reg nq, nm, nn, no, np, ni, nj, nk, nl, nh, nr, ns;
  wire new_n49_, new_n50_, new_n51_1_, new_n52_, new_n53_, new_n55_,
    new_n56_1_, new_n57_, new_n58_, new_n60_, new_n61_1_, new_n62_,
    new_n63_, new_n64_, new_n65_, new_n66_1_, new_n68_, new_n69_, new_n70_,
    new_n71_1_, new_n73_, new_n74_, new_n75_, new_n76_1_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_1_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n234_, new_n235_, new_n236_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n274_, new_n275_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n300_,
    new_n302_, n26, n31, n36, n41, n46, n51, n56, n61, n66, n71, n76, n81;
  assign new_n49_ = ~pa & ~pb;
  assign new_n50_ = ~pa & pc;
  assign new_n51_1_ = ~new_n49_ & ~new_n50_;
  assign new_n52_ = ~pa & new_n51_1_;
  assign new_n53_ = ~pa & pb;
  assign n51 = pe & new_n53_;
  assign new_n55_ = new_n52_ & n51;
  assign new_n56_1_ = ~nr & new_n55_;
  assign new_n57_ = ~ns & new_n56_1_;
  assign new_n58_ = ~nq & new_n57_;
  assign n56 = pf & new_n53_;
  assign new_n60_ = new_n52_ & n56;
  assign new_n61_1_ = ~ns & new_n60_;
  assign new_n62_ = n51 & new_n61_1_;
  assign new_n63_ = ~nq & new_n62_;
  assign new_n64_ = ~ns & new_n52_;
  assign new_n65_ = n56 & new_n64_;
  assign new_n66_1_ = ~nr & new_n65_;
  assign n61 = pg & new_n53_;
  assign new_n68_ = new_n60_ & n61;
  assign new_n69_ = ~nr & new_n68_;
  assign new_n70_ = new_n52_ & n61;
  assign new_n71_1_ = ~ns & new_n70_;
  assign n71 = pd & new_n53_;
  assign new_n73_ = n51 & n61;
  assign new_n74_ = ~nr & new_n73_;
  assign new_n75_ = n71 & new_n74_;
  assign new_n76_1_ = ~np & new_n75_;
  assign new_n77_ = new_n52_ & new_n76_1_;
  assign new_n78_ = n56 & n61;
  assign new_n79_ = ~nq & new_n78_;
  assign new_n80_ = n71 & new_n79_;
  assign new_n81_1_ = ~np & new_n80_;
  assign new_n82_ = new_n52_ & new_n81_1_;
  assign new_n83_ = n71 & new_n78_;
  assign new_n84_ = n51 & new_n83_;
  assign new_n85_ = ~np & new_n84_;
  assign new_n86_ = new_n52_ & new_n85_;
  assign new_n87_ = n51 & n56;
  assign new_n88_ = ~ns & new_n87_;
  assign new_n89_ = n71 & new_n88_;
  assign new_n90_ = ~np & new_n89_;
  assign new_n91_ = new_n52_ & new_n90_;
  assign new_n92_ = n61 & n71;
  assign new_n93_ = ~nq & new_n92_;
  assign new_n94_ = ~nr & new_n93_;
  assign new_n95_ = ~np & new_n94_;
  assign new_n96_ = new_n52_ & new_n95_;
  assign new_n97_ = n56 & n71;
  assign new_n98_ = ~nq & new_n97_;
  assign new_n99_ = ~ns & new_n98_;
  assign new_n100_ = ~np & new_n99_;
  assign new_n101_ = new_n52_ & new_n100_;
  assign new_n102_ = ~ns & n71;
  assign new_n103_ = ~nq & new_n102_;
  assign new_n104_ = ~nr & new_n103_;
  assign new_n105_ = ~np & new_n104_;
  assign new_n106_ = new_n52_ & new_n105_;
  assign new_n107_ = n51 & n71;
  assign new_n108_ = ~nr & new_n107_;
  assign new_n109_ = ~ns & new_n108_;
  assign new_n110_ = ~np & new_n109_;
  assign new_n111_ = new_n52_ & new_n110_;
  assign new_n112_ = ~nr & new_n70_;
  assign new_n113_ = n51 & new_n112_;
  assign new_n114_ = ~nq & new_n113_;
  assign new_n115_ = n51 & new_n70_;
  assign new_n116_ = n56 & new_n115_;
  assign new_n117_ = ~nq & new_n116_;
  assign new_n118_ = ~new_n111_ & ~new_n114_;
  assign new_n119_ = ~new_n117_ & new_n118_;
  assign new_n120_ = ~new_n101_ & ~new_n106_;
  assign new_n121_ = ~new_n91_ & ~new_n96_;
  assign new_n122_ = new_n120_ & new_n121_;
  assign new_n123_ = new_n119_ & new_n122_;
  assign new_n124_ = ~new_n82_ & ~new_n86_;
  assign new_n125_ = ~new_n71_1_ & ~new_n77_;
  assign new_n126_ = new_n124_ & new_n125_;
  assign new_n127_ = ~new_n58_ & ~new_n63_;
  assign new_n128_ = ~new_n66_1_ & ~new_n69_;
  assign new_n129_ = new_n127_ & new_n128_;
  assign new_n130_ = new_n126_ & new_n129_;
  assign new_n131_ = new_n123_ & new_n130_;
  assign new_n132_ = new_n52_ & new_n131_;
  assign new_n133_ = nq & new_n132_;
  assign new_n134_ = ~pc & ~new_n131_;
  assign new_n135_ = n51 & new_n134_;
  assign new_n136_ = ~new_n133_ & ~new_n135_;
  assign n26 = new_n52_ & ~new_n136_;
  assign new_n138_ = np & new_n132_;
  assign new_n139_ = n71 & new_n134_;
  assign new_n140_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = ~nn & new_n55_;
  assign new_n142_ = ~no & new_n141_;
  assign new_n143_ = ~nm & new_n142_;
  assign new_n144_ = ~no & new_n60_;
  assign new_n145_ = n51 & new_n144_;
  assign new_n146_ = ~nm & new_n145_;
  assign new_n147_ = ~no & new_n52_;
  assign new_n148_ = n56 & new_n147_;
  assign new_n149_ = ~nn & new_n148_;
  assign new_n150_ = ~nn & new_n68_;
  assign new_n151_ = ~no & new_n70_;
  assign new_n152_ = ~nn & new_n73_;
  assign new_n153_ = n71 & new_n152_;
  assign new_n154_ = ~nl & new_n153_;
  assign new_n155_ = new_n52_ & new_n154_;
  assign new_n156_ = ~nm & new_n78_;
  assign new_n157_ = n71 & new_n156_;
  assign new_n158_ = ~nl & new_n157_;
  assign new_n159_ = new_n52_ & new_n158_;
  assign new_n160_ = ~nl & new_n84_;
  assign new_n161_ = new_n52_ & new_n160_;
  assign new_n162_ = ~no & new_n87_;
  assign new_n163_ = n71 & new_n162_;
  assign new_n164_ = ~nl & new_n163_;
  assign new_n165_ = new_n52_ & new_n164_;
  assign new_n166_ = ~nm & new_n92_;
  assign new_n167_ = ~nn & new_n166_;
  assign new_n168_ = ~nl & new_n167_;
  assign new_n169_ = new_n52_ & new_n168_;
  assign new_n170_ = ~nm & new_n97_;
  assign new_n171_ = ~no & new_n170_;
  assign new_n172_ = ~nl & new_n171_;
  assign new_n173_ = new_n52_ & new_n172_;
  assign new_n174_ = ~no & n71;
  assign new_n175_ = ~nm & new_n174_;
  assign new_n176_ = ~nn & new_n175_;
  assign new_n177_ = ~nl & new_n176_;
  assign new_n178_ = new_n52_ & new_n177_;
  assign new_n179_ = ~nn & new_n107_;
  assign new_n180_ = ~no & new_n179_;
  assign new_n181_ = ~nl & new_n180_;
  assign new_n182_ = new_n52_ & new_n181_;
  assign new_n183_ = ~nn & new_n70_;
  assign new_n184_ = n51 & new_n183_;
  assign new_n185_ = ~nm & new_n184_;
  assign new_n186_ = ~nm & new_n116_;
  assign new_n187_ = ~new_n182_ & ~new_n185_;
  assign new_n188_ = ~new_n186_ & new_n187_;
  assign new_n189_ = ~new_n173_ & ~new_n178_;
  assign new_n190_ = ~new_n165_ & ~new_n169_;
  assign new_n191_ = new_n189_ & new_n190_;
  assign new_n192_ = new_n188_ & new_n191_;
  assign new_n193_ = ~new_n159_ & ~new_n161_;
  assign new_n194_ = ~new_n151_ & ~new_n155_;
  assign new_n195_ = new_n193_ & new_n194_;
  assign new_n196_ = ~new_n143_ & ~new_n146_;
  assign new_n197_ = ~new_n149_ & ~new_n150_;
  assign new_n198_ = new_n196_ & new_n197_;
  assign new_n199_ = new_n195_ & new_n198_;
  assign new_n200_ = new_n192_ & new_n199_;
  assign new_n201_ = new_n52_ & ~new_n200_;
  assign new_n202_ = nl & new_n201_;
  assign new_n203_ = ~pc & new_n200_;
  assign new_n204_ = n71 & new_n203_;
  assign new_n205_ = ~new_n202_ & ~new_n204_;
  assign new_n206_ = ~new_n140_ & ~new_n205_;
  assign new_n207_ = ~new_n136_ & new_n206_;
  assign new_n208_ = nm & new_n201_;
  assign new_n209_ = n51 & new_n203_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = new_n206_ & ~new_n210_;
  assign new_n212_ = ~new_n136_ & ~new_n210_;
  assign new_n213_ = ~new_n207_ & ~new_n211_;
  assign new_n214_ = ~new_n212_ & new_n213_;
  assign new_n215_ = new_n53_ & n26;
  assign new_n216_ = new_n214_ & new_n215_;
  assign n46 = new_n52_ & ~new_n140_;
  assign new_n218_ = new_n53_ & ~new_n205_;
  assign new_n219_ = n46 & new_n218_;
  assign new_n220_ = new_n214_ & new_n219_;
  assign new_n221_ = new_n52_ & new_n214_;
  assign new_n222_ = ~new_n210_ & new_n221_;
  assign new_n223_ = new_n53_ & n71;
  assign new_n224_ = pc & new_n223_;
  assign new_n225_ = nh & new_n49_;
  assign new_n226_ = ~new_n140_ & new_n215_;
  assign new_n227_ = ~new_n205_ & new_n226_;
  assign new_n228_ = ~new_n210_ & new_n227_;
  assign new_n229_ = ~new_n216_ & ~new_n220_;
  assign new_n230_ = ~new_n222_ & new_n229_;
  assign new_n231_ = ~new_n224_ & ~new_n225_;
  assign new_n232_ = ~new_n228_ & new_n231_;
  assign pt = ~new_n230_ | ~new_n232_;
  assign new_n234_ = nr & new_n132_;
  assign new_n235_ = n56 & new_n134_;
  assign new_n236_ = ~new_n234_ & ~new_n235_;
  assign n76 = new_n52_ & ~new_n236_;
  assign new_n238_ = nn & new_n201_;
  assign new_n239_ = n56 & new_n203_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = ~new_n214_ & ~new_n240_;
  assign new_n242_ = ~new_n236_ & ~new_n240_;
  assign new_n243_ = ~new_n214_ & ~new_n236_;
  assign new_n244_ = ~new_n241_ & ~new_n242_;
  assign new_n245_ = ~new_n243_ & new_n244_;
  assign new_n246_ = new_n53_ & n76;
  assign new_n247_ = new_n245_ & new_n246_;
  assign new_n248_ = ~pa & ~new_n240_;
  assign n36 = ~new_n52_ | new_n248_;
  assign new_n250_ = new_n53_ & new_n245_;
  assign new_n251_ = ~new_n214_ & new_n250_;
  assign new_n252_ = ~n36 & new_n251_;
  assign new_n253_ = new_n52_ & ~new_n240_;
  assign new_n254_ = new_n245_ & new_n253_;
  assign new_n255_ = new_n53_ & n51;
  assign new_n256_ = pc & new_n255_;
  assign new_n257_ = ni & new_n49_;
  assign new_n258_ = new_n53_ & ~new_n240_;
  assign new_n259_ = n76 & new_n258_;
  assign new_n260_ = ~new_n214_ & new_n259_;
  assign new_n261_ = ~new_n247_ & ~new_n252_;
  assign new_n262_ = ~new_n254_ & new_n261_;
  assign new_n263_ = ~new_n256_ & ~new_n257_;
  assign new_n264_ = ~new_n260_ & new_n263_;
  assign pu = ~new_n262_ | ~new_n264_;
  assign new_n266_ = ns & new_n132_;
  assign new_n267_ = n61 & new_n134_;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign new_n269_ = no & new_n201_;
  assign new_n270_ = n61 & new_n203_;
  assign new_n271_ = ~new_n269_ & ~new_n270_;
  assign new_n272_ = ~pa & ~new_n271_;
  assign n41 = ~new_n52_ | new_n272_;
  assign new_n274_ = ~new_n245_ & new_n268_;
  assign new_n275_ = ~n41 & new_n274_;
  assign n81 = new_n52_ & ~new_n268_;
  assign new_n277_ = ~new_n271_ & n81;
  assign new_n278_ = ~new_n245_ & new_n277_;
  assign new_n279_ = nj & new_n49_;
  assign new_n280_ = new_n245_ & ~new_n268_;
  assign new_n281_ = ~n41 & new_n280_;
  assign new_n282_ = pc & n56;
  assign new_n283_ = new_n52_ & new_n268_;
  assign new_n284_ = ~new_n271_ & new_n283_;
  assign new_n285_ = new_n245_ & new_n284_;
  assign new_n286_ = ~new_n275_ & ~new_n278_;
  assign new_n287_ = ~new_n279_ & new_n286_;
  assign new_n288_ = ~new_n281_ & ~new_n282_;
  assign new_n289_ = ~new_n285_ & new_n288_;
  assign pv = ~new_n287_ | ~new_n289_;
  assign new_n291_ = nk & new_n49_;
  assign new_n292_ = new_n52_ & ~new_n271_;
  assign new_n293_ = ~new_n245_ & new_n292_;
  assign new_n294_ = ~new_n245_ & n81;
  assign new_n295_ = pc & n61;
  assign new_n296_ = ~new_n277_ & ~new_n295_;
  assign new_n297_ = ~new_n291_ & ~new_n293_;
  assign new_n298_ = ~new_n294_ & new_n297_;
  assign pw = ~new_n296_ | ~new_n298_;
  assign new_n300_ = ~pa & ~new_n210_;
  assign n31 = ~new_n52_ | new_n300_;
  assign new_n302_ = ~pa & ~new_n205_;
  assign n66 = ~new_n52_ | new_n302_;
  always @ (posedge clock) begin
    nq <= n26;
    nm <= n31;
    nn <= n36;
    no <= n41;
    np <= n46;
    ni <= n51;
    nj <= n56;
    nk <= n61;
    nl <= n66;
    nh <= n71;
    nr <= n76;
    ns <= n81;
  end
endmodule

