// Benchmark "testing" written by ABC on Thu Oct  8 22:16:46 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A142, A141, A140, A139, A138, A109, A108, A107, A106, A105, A76, A75,
    A74, A73, A72, A43, A42, A41, A40, A39, A6, A7, A8, A9, A10  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A142, A141, A140, A139, A138, A109, A108, A107, A106, A105, A76, A75,
    A74, A73, A72, A43, A42, A41, A40, A39, A6, A7, A8, A9, A10;
  wire \new_[50]_ , \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ ,
    \new_[55]_ , \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ ,
    \new_[60]_ , \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ ,
    \new_[65]_ , \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ ,
    \new_[70]_ , \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ ,
    \new_[75]_ , \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ ,
    \new_[80]_ , \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ ,
    \new_[85]_ , \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ ,
    \new_[90]_ , \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ ,
    \new_[95]_ , \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ ,
    \new_[100]_ , \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ ,
    \new_[105]_ , \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ ,
    \new_[110]_ , \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ ,
    \new_[115]_ , \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ ,
    \new_[120]_ , \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ ,
    \new_[125]_ , \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ ,
    \new_[130]_ , \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ ,
    \new_[135]_ , \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ ,
    \new_[140]_ , \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ ,
    \new_[145]_ , \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ ,
    \new_[150]_ , \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ ,
    \new_[155]_ , \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ , \new_[176]_ ,
    \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ , \new_[181]_ ,
    \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ , \new_[186]_ ,
    \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ , \new_[191]_ ,
    \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ , \new_[196]_ ,
    \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ , \new_[201]_ ,
    \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ , \new_[206]_ ,
    \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ , \new_[211]_ ,
    \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ , \new_[216]_ ,
    \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ , \new_[221]_ ,
    \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ , \new_[226]_ ,
    \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ , \new_[231]_ ,
    \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ , \new_[236]_ ,
    \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ , \new_[241]_ ,
    \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ , \new_[246]_ ,
    \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ , \new_[252]_ ,
    \new_[253]_ , \new_[254]_ , \new_[255]_ , \new_[256]_ , \new_[257]_ ,
    \new_[258]_ , \new_[259]_ , \new_[260]_ , \new_[261]_ , \new_[262]_ ,
    \new_[263]_ , \new_[264]_ , \new_[265]_ , \new_[266]_ , \new_[267]_ ,
    \new_[268]_ , \new_[269]_ , \new_[270]_ , \new_[271]_ , \new_[272]_ ,
    \new_[273]_ , \new_[274]_ , \new_[275]_ , \new_[276]_ , \new_[277]_ ,
    \new_[278]_ , \new_[279]_ , \new_[280]_ , \new_[281]_ , \new_[282]_ ,
    \new_[283]_ , \new_[284]_ , \new_[285]_ , \new_[286]_ , \new_[287]_ ,
    \new_[288]_ , \new_[289]_ , \new_[290]_ , \new_[291]_ , \new_[292]_ ,
    \new_[293]_ , \new_[294]_ , \new_[295]_ , \new_[296]_ , \new_[297]_ ,
    \new_[298]_ , \new_[299]_ , \new_[300]_ , \new_[301]_ , \new_[302]_ ,
    \new_[303]_ , \new_[304]_ , \new_[305]_ , \new_[306]_ , \new_[307]_ ,
    \new_[308]_ , \new_[309]_ , \new_[310]_ , \new_[311]_ , \new_[312]_ ,
    \new_[314]_ , \new_[315]_ , \new_[316]_ , \new_[317]_ , \new_[318]_ ,
    \new_[320]_ , \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ ,
    \new_[325]_ , \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ ,
    \new_[330]_ , \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ ,
    \new_[335]_ , \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ ,
    \new_[340]_ , \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ ,
    \new_[345]_ , \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ ,
    \new_[350]_ , \new_[351]_ , \new_[352]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[406]_ ,
    \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ , \new_[412]_ ,
    \new_[413]_ , \new_[414]_ , \new_[415]_ , \new_[416]_ , \new_[417]_ ,
    \new_[418]_ , \new_[419]_ , \new_[420]_ , \new_[421]_ , \new_[422]_ ,
    \new_[423]_ , \new_[424]_ , \new_[425]_ , \new_[426]_ , \new_[427]_ ,
    \new_[428]_ , \new_[429]_ , \new_[430]_ , \new_[431]_ , \new_[432]_ ,
    \new_[433]_ , \new_[434]_ , \new_[435]_ , \new_[436]_ , \new_[437]_ ,
    \new_[438]_ , \new_[439]_ , \new_[440]_ , \new_[441]_ , \new_[442]_ ,
    \new_[443]_ , \new_[444]_ , \new_[445]_ , \new_[446]_ , \new_[447]_ ,
    \new_[448]_ , \new_[449]_ , \new_[450]_ , \new_[451]_ , \new_[452]_ ,
    \new_[453]_ , \new_[454]_ , \new_[455]_ , \new_[457]_ , \new_[458]_ ,
    \new_[459]_ , \new_[460]_ , \new_[461]_ , \new_[462]_ , \new_[463]_ ,
    \new_[464]_ , \new_[465]_ , \new_[466]_ , \new_[467]_ , \new_[468]_ ,
    \new_[469]_ , \new_[470]_ , \new_[471]_ , \new_[472]_ , \new_[473]_ ,
    \new_[474]_ , \new_[475]_ , \new_[476]_ , \new_[477]_ , \new_[478]_ ,
    \new_[479]_ , \new_[480]_ , \new_[481]_ , \new_[482]_ , \new_[483]_ ,
    \new_[484]_ , \new_[485]_ , \new_[486]_ , \new_[487]_ , \new_[488]_ ,
    \new_[489]_ , \new_[490]_ , \new_[491]_ , \new_[492]_ , \new_[493]_ ,
    \new_[494]_ , \new_[495]_ , \new_[496]_ , \new_[497]_ , \new_[498]_ ,
    \new_[499]_ , \new_[500]_ , \new_[501]_ , \new_[502]_ , \new_[503]_ ,
    \new_[504]_ , \new_[505]_ , \new_[506]_ , \new_[507]_ , \new_[508]_ ,
    \new_[509]_ , \new_[510]_ , \new_[511]_ , \new_[512]_ , \new_[513]_ ,
    \new_[514]_ , \new_[515]_ , \new_[516]_ , \new_[517]_ , \new_[518]_ ,
    \new_[519]_ , \new_[520]_ , \new_[521]_ , \new_[522]_ , \new_[523]_ ,
    \new_[524]_ , \new_[525]_ , \new_[526]_ , \new_[527]_ , \new_[528]_ ,
    \new_[529]_ , \new_[530]_ , \new_[531]_ , \new_[532]_ , \new_[533]_ ,
    \new_[534]_ , \new_[535]_ , \new_[536]_ , \new_[538]_ , \new_[539]_ ,
    \new_[540]_ , \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ ,
    \new_[545]_ , \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ ,
    \new_[550]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[656]_ ,
    \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ , \new_[661]_ ,
    \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ , \new_[666]_ ,
    \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ , \new_[671]_ ,
    \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ , \new_[676]_ ,
    \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ , \new_[681]_ ,
    \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ , \new_[686]_ ,
    \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ , \new_[691]_ ,
    \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ , \new_[696]_ ,
    \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ , \new_[701]_ ,
    \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ , \new_[706]_ ,
    \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ , \new_[711]_ ,
    \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ , \new_[716]_ ,
    \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ , \new_[721]_ ,
    \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ , \new_[726]_ ,
    \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ , \new_[731]_ ,
    \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[736]_ , \new_[737]_ ,
    \new_[738]_ , \new_[739]_ , \new_[740]_ , \new_[741]_ , \new_[742]_ ,
    \new_[743]_ , \new_[744]_ , \new_[745]_ , \new_[746]_ , \new_[747]_ ,
    \new_[748]_ , \new_[749]_ , \new_[750]_ , \new_[751]_ , \new_[752]_ ,
    \new_[753]_ , \new_[754]_ , \new_[755]_ , \new_[756]_ , \new_[757]_ ,
    \new_[758]_ , \new_[759]_ , \new_[760]_ , \new_[761]_ , \new_[762]_ ,
    \new_[763]_ , \new_[764]_ , \new_[765]_ , \new_[766]_ , \new_[767]_ ,
    \new_[768]_ , \new_[769]_ , \new_[770]_ , \new_[771]_ , \new_[772]_ ,
    \new_[773]_ , \new_[774]_ , \new_[775]_ , \new_[776]_ , \new_[777]_ ,
    \new_[778]_ , \new_[779]_ , \new_[780]_ , \new_[781]_ , \new_[782]_ ,
    \new_[783]_ , \new_[784]_ , \new_[785]_ , \new_[786]_ , \new_[787]_ ,
    \new_[788]_ , \new_[789]_ , \new_[790]_ , \new_[791]_ , \new_[792]_ ,
    \new_[793]_ , \new_[794]_ , \new_[795]_ , \new_[796]_ , \new_[797]_ ,
    \new_[798]_ , \new_[799]_ , \new_[800]_ , \new_[801]_ , \new_[802]_ ,
    \new_[803]_ , \new_[804]_ , \new_[805]_ , \new_[806]_ , \new_[808]_ ,
    \new_[809]_ , \new_[810]_ , \new_[811]_ , \new_[812]_ , \new_[813]_ ,
    \new_[814]_ , \new_[815]_ , \new_[816]_ , \new_[817]_ , \new_[818]_ ,
    \new_[819]_ , \new_[820]_ , \new_[821]_ , \new_[822]_ , \new_[823]_ ,
    \new_[824]_ , \new_[825]_ , \new_[826]_ , \new_[827]_ , \new_[828]_ ,
    \new_[829]_ , \new_[830]_ , \new_[831]_ , \new_[832]_ , \new_[833]_ ,
    \new_[834]_ , \new_[835]_ , \new_[836]_ , \new_[837]_ , \new_[839]_ ,
    \new_[840]_ , \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ ,
    \new_[845]_ , \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ ,
    \new_[850]_ , \new_[851]_ , \new_[852]_ , \new_[853]_ ;
  assign \new_[50]_  = ~A169 & A170;
  assign \new_[51]_  = ~A166 & A167;
  assign \new_[52]_  = A166 & ~A167;
  assign \new_[53]_  = ~\new_[51]_  & ~\new_[52]_ ;
  assign \new_[54]_  = ~A200 & A199;
  assign \new_[55]_  = A200 & ~A199;
  assign \new_[56]_  = ~\new_[54]_  & ~\new_[55]_ ;
  assign \new_[57]_  = ~A203 & ~A202;
  assign \new_[58]_  = A201 & ~\new_[57]_ ;
  assign \new_[59]_  = ~A203 & ~A201;
  assign \new_[60]_  = ~A202 & \new_[59]_ ;
  assign \new_[61]_  = ~\new_[58]_  & ~\new_[60]_ ;
  assign \new_[62]_  = ~\new_[56]_  & ~\new_[61]_ ;
  assign \new_[63]_  = A168 & ~\new_[53]_ ;
  assign \new_[64]_  = \new_[62]_  & \new_[63]_ ;
  assign \new_[65]_  = ~A201 & ~\new_[57]_ ;
  assign \new_[66]_  = ~A203 & A201;
  assign \new_[67]_  = ~A202 & \new_[66]_ ;
  assign \new_[68]_  = A200 & A199;
  assign \new_[69]_  = ~A200 & ~A199;
  assign \new_[70]_  = ~\new_[68]_  & ~\new_[69]_ ;
  assign \new_[71]_  = ~\new_[67]_  & \new_[70]_ ;
  assign \new_[72]_  = ~\new_[65]_  & \new_[71]_ ;
  assign \new_[73]_  = ~A168 & ~\new_[72]_ ;
  assign \new_[74]_  = ~\new_[64]_  & ~\new_[73]_ ;
  assign \new_[75]_  = ~\new_[50]_  & ~\new_[74]_ ;
  assign \new_[76]_  = ~\new_[53]_  & ~\new_[56]_ ;
  assign \new_[77]_  = A201 & ~A168;
  assign \new_[78]_  = \new_[76]_  & \new_[77]_ ;
  assign \new_[79]_  = ~A201 & A168;
  assign \new_[80]_  = ~\new_[78]_  & ~\new_[79]_ ;
  assign \new_[81]_  = \new_[50]_  & ~\new_[80]_ ;
  assign \new_[82]_  = A166 & A167;
  assign \new_[83]_  = ~A166 & ~A167;
  assign \new_[84]_  = ~\new_[82]_  & ~\new_[83]_ ;
  assign \new_[85]_  = ~A201 & ~\new_[84]_ ;
  assign \new_[86]_  = ~\new_[81]_  & ~\new_[85]_ ;
  assign \new_[87]_  = ~\new_[57]_  & ~\new_[86]_ ;
  assign \new_[88]_  = A168 & \new_[50]_ ;
  assign \new_[89]_  = \new_[84]_  & ~\new_[88]_ ;
  assign \new_[90]_  = ~\new_[71]_  & ~\new_[89]_ ;
  assign \new_[91]_  = ~A201 & ~A168;
  assign \new_[92]_  = \new_[57]_  & \new_[91]_ ;
  assign \new_[93]_  = \new_[50]_  & \new_[92]_ ;
  assign \new_[94]_  = \new_[76]_  & \new_[93]_ ;
  assign \new_[95]_  = ~A236 & ~A235;
  assign \new_[96]_  = A299 & ~A298;
  assign \new_[97]_  = ~A299 & A298;
  assign \new_[98]_  = ~\new_[96]_  & ~\new_[97]_ ;
  assign \new_[99]_  = ~A302 & ~A301;
  assign \new_[100]_  = A300 & ~\new_[99]_ ;
  assign \new_[101]_  = ~A302 & ~A300;
  assign \new_[102]_  = ~A301 & \new_[101]_ ;
  assign \new_[103]_  = ~\new_[100]_  & ~\new_[102]_ ;
  assign \new_[104]_  = ~\new_[98]_  & ~\new_[103]_ ;
  assign \new_[105]_  = A266 & ~A265;
  assign \new_[106]_  = ~A266 & A265;
  assign \new_[107]_  = ~\new_[105]_  & ~\new_[106]_ ;
  assign \new_[108]_  = ~A269 & ~A268;
  assign \new_[109]_  = A267 & ~\new_[108]_ ;
  assign \new_[110]_  = ~A269 & ~A267;
  assign \new_[111]_  = ~A268 & \new_[110]_ ;
  assign \new_[112]_  = ~\new_[109]_  & ~\new_[111]_ ;
  assign \new_[113]_  = ~\new_[107]_  & ~\new_[112]_ ;
  assign \new_[114]_  = ~\new_[104]_  & ~\new_[113]_ ;
  assign \new_[115]_  = ~A234 & ~\new_[114]_ ;
  assign \new_[116]_  = ~A233 & A232;
  assign \new_[117]_  = A233 & ~A232;
  assign \new_[118]_  = ~\new_[116]_  & ~\new_[117]_ ;
  assign \new_[119]_  = ~A267 & ~\new_[108]_ ;
  assign \new_[120]_  = ~A269 & A267;
  assign \new_[121]_  = ~A268 & \new_[120]_ ;
  assign \new_[122]_  = A266 & A265;
  assign \new_[123]_  = ~A266 & ~A265;
  assign \new_[124]_  = ~\new_[122]_  & ~\new_[123]_ ;
  assign \new_[125]_  = ~\new_[121]_  & \new_[124]_ ;
  assign \new_[126]_  = ~\new_[119]_  & \new_[125]_ ;
  assign \new_[127]_  = ~A300 & ~\new_[99]_ ;
  assign \new_[128]_  = ~A302 & A300;
  assign \new_[129]_  = ~A301 & \new_[128]_ ;
  assign \new_[130]_  = A299 & A298;
  assign \new_[131]_  = ~A299 & ~A298;
  assign \new_[132]_  = ~\new_[130]_  & ~\new_[131]_ ;
  assign \new_[133]_  = ~\new_[129]_  & \new_[132]_ ;
  assign \new_[134]_  = ~\new_[127]_  & \new_[133]_ ;
  assign \new_[135]_  = ~\new_[126]_  & ~\new_[134]_ ;
  assign \new_[136]_  = ~\new_[118]_  & \new_[135]_ ;
  assign \new_[137]_  = A234 & \new_[136]_ ;
  assign \new_[138]_  = ~\new_[115]_  & ~\new_[137]_ ;
  assign \new_[139]_  = ~\new_[95]_  & ~\new_[138]_ ;
  assign \new_[140]_  = ~A236 & A234;
  assign \new_[141]_  = ~A235 & \new_[140]_ ;
  assign \new_[142]_  = A233 & A232;
  assign \new_[143]_  = ~A233 & ~A232;
  assign \new_[144]_  = ~\new_[142]_  & ~\new_[143]_ ;
  assign \new_[145]_  = ~\new_[141]_  & \new_[144]_ ;
  assign \new_[146]_  = ~\new_[98]_  & ~\new_[145]_ ;
  assign \new_[147]_  = ~\new_[103]_  & \new_[146]_ ;
  assign \new_[148]_  = ~\new_[107]_  & ~\new_[145]_ ;
  assign \new_[149]_  = ~\new_[112]_  & \new_[148]_ ;
  assign \new_[150]_  = ~A236 & ~A234;
  assign \new_[151]_  = ~A235 & \new_[150]_ ;
  assign \new_[152]_  = \new_[136]_  & \new_[151]_ ;
  assign \new_[153]_  = ~\new_[90]_  & ~\new_[94]_ ;
  assign \new_[154]_  = ~\new_[149]_  & \new_[153]_ ;
  assign \new_[155]_  = ~\new_[147]_  & \new_[154]_ ;
  assign \new_[156]_  = ~\new_[152]_  & \new_[155]_ ;
  assign \new_[157]_  = ~\new_[75]_  & \new_[156]_ ;
  assign \new_[158]_  = ~\new_[87]_  & \new_[157]_ ;
  assign A142 = ~\new_[139]_  & \new_[158]_ ;
  assign \new_[160]_  = A168 & ~\new_[50]_ ;
  assign \new_[161]_  = ~A168 & \new_[50]_ ;
  assign \new_[162]_  = ~\new_[160]_  & ~\new_[161]_ ;
  assign \new_[163]_  = ~A234 & ~\new_[95]_ ;
  assign \new_[164]_  = \new_[145]_  & ~\new_[163]_ ;
  assign \new_[165]_  = ~\new_[62]_  & \new_[164]_ ;
  assign \new_[166]_  = ~\new_[135]_  & \new_[165]_ ;
  assign \new_[167]_  = ~\new_[53]_  & ~\new_[162]_ ;
  assign \new_[168]_  = ~\new_[166]_  & \new_[167]_ ;
  assign \new_[169]_  = ~A168 & ~\new_[50]_ ;
  assign \new_[170]_  = \new_[89]_  & ~\new_[169]_ ;
  assign \new_[171]_  = ~\new_[72]_  & ~\new_[170]_ ;
  assign A141 = ~\new_[168]_  & ~\new_[171]_ ;
  assign \new_[173]_  = A234 & ~\new_[95]_ ;
  assign \new_[174]_  = ~\new_[151]_  & ~\new_[173]_ ;
  assign \new_[175]_  = ~\new_[118]_  & ~\new_[174]_ ;
  assign \new_[176]_  = ~\new_[61]_  & \new_[175]_ ;
  assign \new_[177]_  = ~\new_[61]_  & \new_[104]_ ;
  assign \new_[178]_  = ~\new_[170]_  & \new_[177]_ ;
  assign \new_[179]_  = ~\new_[176]_  & ~\new_[178]_ ;
  assign \new_[180]_  = ~\new_[56]_  & ~\new_[179]_ ;
  assign \new_[181]_  = ~\new_[162]_  & \new_[175]_ ;
  assign \new_[182]_  = \new_[104]_  & ~\new_[162]_ ;
  assign \new_[183]_  = ~\new_[72]_  & \new_[182]_ ;
  assign \new_[184]_  = ~\new_[181]_  & ~\new_[183]_ ;
  assign \new_[185]_  = ~\new_[53]_  & ~\new_[184]_ ;
  assign \new_[186]_  = ~\new_[113]_  & ~\new_[185]_ ;
  assign \new_[187]_  = ~\new_[180]_  & \new_[186]_ ;
  assign \new_[188]_  = ~A267 & ~A168;
  assign \new_[189]_  = \new_[104]_  & \new_[188]_ ;
  assign \new_[190]_  = A168 & ~\new_[107]_ ;
  assign \new_[191]_  = ~\new_[53]_  & \new_[190]_ ;
  assign \new_[192]_  = ~\new_[134]_  & \new_[191]_ ;
  assign \new_[193]_  = A267 & \new_[192]_ ;
  assign \new_[194]_  = ~\new_[189]_  & ~\new_[193]_ ;
  assign \new_[195]_  = ~\new_[108]_  & ~\new_[194]_ ;
  assign \new_[196]_  = ~A168 & ~\new_[98]_ ;
  assign \new_[197]_  = ~\new_[125]_  & \new_[196]_ ;
  assign \new_[198]_  = ~\new_[103]_  & \new_[197]_ ;
  assign \new_[199]_  = \new_[111]_  & \new_[192]_ ;
  assign \new_[200]_  = ~\new_[198]_  & ~\new_[199]_ ;
  assign \new_[201]_  = ~\new_[195]_  & \new_[200]_ ;
  assign \new_[202]_  = ~\new_[50]_  & ~\new_[201]_ ;
  assign \new_[203]_  = ~\new_[89]_  & \new_[104]_ ;
  assign \new_[204]_  = ~\new_[126]_  & \new_[203]_ ;
  assign \new_[205]_  = ~\new_[107]_  & \new_[161]_ ;
  assign \new_[206]_  = ~\new_[53]_  & \new_[205]_ ;
  assign \new_[207]_  = ~\new_[112]_  & \new_[206]_ ;
  assign \new_[208]_  = ~\new_[134]_  & \new_[207]_ ;
  assign \new_[209]_  = ~\new_[204]_  & ~\new_[208]_ ;
  assign \new_[210]_  = ~\new_[202]_  & \new_[209]_ ;
  assign \new_[211]_  = ~\new_[61]_  & ~\new_[210]_ ;
  assign \new_[212]_  = ~\new_[176]_  & ~\new_[211]_ ;
  assign \new_[213]_  = ~\new_[56]_  & ~\new_[212]_ ;
  assign \new_[214]_  = ~\new_[72]_  & ~\new_[126]_ ;
  assign \new_[215]_  = \new_[182]_  & \new_[214]_ ;
  assign \new_[216]_  = ~\new_[181]_  & ~\new_[215]_ ;
  assign \new_[217]_  = ~\new_[53]_  & ~\new_[216]_ ;
  assign \new_[218]_  = \new_[113]_  & ~\new_[134]_ ;
  assign \new_[219]_  = \new_[171]_  & \new_[218]_ ;
  assign \new_[220]_  = ~\new_[217]_  & ~\new_[219]_ ;
  assign \new_[221]_  = ~\new_[213]_  & \new_[220]_ ;
  assign \new_[222]_  = ~\new_[98]_  & ~\new_[118]_ ;
  assign \new_[223]_  = ~\new_[126]_  & \new_[222]_ ;
  assign \new_[224]_  = A234 & \new_[223]_ ;
  assign \new_[225]_  = A300 & \new_[224]_ ;
  assign \new_[226]_  = ~A300 & ~A234;
  assign \new_[227]_  = ~\new_[225]_  & ~\new_[226]_ ;
  assign \new_[228]_  = ~\new_[99]_  & ~\new_[227]_ ;
  assign \new_[229]_  = ~A300 & \new_[224]_ ;
  assign \new_[230]_  = A300 & ~A234;
  assign \new_[231]_  = ~\new_[229]_  & ~\new_[230]_ ;
  assign \new_[232]_  = \new_[99]_  & ~\new_[231]_ ;
  assign \new_[233]_  = ~\new_[113]_  & \new_[132]_ ;
  assign \new_[234]_  = ~A234 & ~\new_[233]_ ;
  assign \new_[235]_  = ~\new_[232]_  & ~\new_[234]_ ;
  assign \new_[236]_  = ~\new_[228]_  & \new_[235]_ ;
  assign \new_[237]_  = ~\new_[95]_  & ~\new_[236]_ ;
  assign \new_[238]_  = ~A300 & ~\new_[145]_ ;
  assign \new_[239]_  = \new_[151]_  & \new_[223]_ ;
  assign \new_[240]_  = A300 & \new_[239]_ ;
  assign \new_[241]_  = ~\new_[238]_  & ~\new_[240]_ ;
  assign \new_[242]_  = ~\new_[99]_  & ~\new_[241]_ ;
  assign \new_[243]_  = ~\new_[113]_  & \new_[133]_ ;
  assign \new_[244]_  = ~\new_[145]_  & ~\new_[243]_ ;
  assign \new_[245]_  = \new_[102]_  & \new_[239]_ ;
  assign \new_[246]_  = \new_[153]_  & ~\new_[244]_ ;
  assign \new_[247]_  = ~\new_[245]_  & \new_[246]_ ;
  assign \new_[248]_  = ~\new_[75]_  & \new_[247]_ ;
  assign \new_[249]_  = ~\new_[87]_  & \new_[248]_ ;
  assign \new_[250]_  = ~\new_[242]_  & \new_[249]_ ;
  assign A138 = ~\new_[237]_  & \new_[250]_ ;
  assign \new_[252]_  = A234 & ~A233;
  assign \new_[253]_  = ~\new_[95]_  & \new_[252]_ ;
  assign \new_[254]_  = A232 & ~\new_[253]_ ;
  assign \new_[255]_  = ~\new_[143]_  & ~\new_[254]_ ;
  assign \new_[256]_  = A300 & \new_[97]_ ;
  assign \new_[257]_  = ~\new_[99]_  & \new_[256]_ ;
  assign \new_[258]_  = A267 & \new_[106]_ ;
  assign \new_[259]_  = ~\new_[108]_  & \new_[258]_ ;
  assign \new_[260]_  = ~\new_[96]_  & ~\new_[105]_ ;
  assign \new_[261]_  = ~\new_[259]_  & \new_[260]_ ;
  assign \new_[262]_  = ~\new_[257]_  & \new_[261]_ ;
  assign \new_[263]_  = ~\new_[255]_  & ~\new_[262]_ ;
  assign \new_[264]_  = A169 & ~A170;
  assign \new_[265]_  = ~A167 & \new_[264]_ ;
  assign \new_[266]_  = A167 & \new_[50]_ ;
  assign \new_[267]_  = ~\new_[265]_  & ~\new_[266]_ ;
  assign \new_[268]_  = ~A166 & ~\new_[267]_ ;
  assign \new_[269]_  = A166 & \new_[264]_ ;
  assign \new_[270]_  = ~A168 & ~\new_[269]_ ;
  assign \new_[271]_  = A167 & ~\new_[270]_ ;
  assign \new_[272]_  = ~A167 & \new_[50]_ ;
  assign \new_[273]_  = ~A168 & ~\new_[272]_ ;
  assign \new_[274]_  = A166 & ~\new_[273]_ ;
  assign \new_[275]_  = ~\new_[271]_  & ~\new_[274]_ ;
  assign \new_[276]_  = ~\new_[268]_  & \new_[275]_ ;
  assign \new_[277]_  = A201 & \new_[54]_ ;
  assign \new_[278]_  = ~\new_[57]_  & \new_[277]_ ;
  assign \new_[279]_  = ~\new_[55]_  & ~\new_[278]_ ;
  assign \new_[280]_  = ~\new_[276]_  & ~\new_[279]_ ;
  assign \new_[281]_  = A201 & ~A200;
  assign \new_[282]_  = ~\new_[57]_  & \new_[281]_ ;
  assign \new_[283]_  = A199 & ~\new_[282]_ ;
  assign \new_[284]_  = ~\new_[69]_  & ~\new_[283]_ ;
  assign \new_[285]_  = ~A167 & A169;
  assign \new_[286]_  = A167 & ~A169;
  assign \new_[287]_  = ~\new_[285]_  & ~\new_[286]_ ;
  assign \new_[288]_  = A166 & ~\new_[287]_ ;
  assign \new_[289]_  = ~A170 & ~\new_[51]_ ;
  assign \new_[290]_  = A169 & ~\new_[289]_ ;
  assign \new_[291]_  = ~A169 & ~A170;
  assign \new_[292]_  = ~\new_[290]_  & ~\new_[291]_ ;
  assign \new_[293]_  = ~\new_[288]_  & \new_[292]_ ;
  assign \new_[294]_  = ~A168 & ~\new_[293]_ ;
  assign \new_[295]_  = \new_[83]_  & ~\new_[264]_ ;
  assign \new_[296]_  = ~\new_[294]_  & ~\new_[295]_ ;
  assign \new_[297]_  = ~\new_[284]_  & ~\new_[296]_ ;
  assign \new_[298]_  = A234 & \new_[116]_ ;
  assign \new_[299]_  = ~\new_[95]_  & \new_[298]_ ;
  assign \new_[300]_  = ~\new_[117]_  & ~\new_[299]_ ;
  assign \new_[301]_  = A267 & A265;
  assign \new_[302]_  = ~\new_[108]_  & \new_[301]_ ;
  assign \new_[303]_  = ~A266 & ~\new_[302]_ ;
  assign \new_[304]_  = ~\new_[122]_  & ~\new_[303]_ ;
  assign \new_[305]_  = A300 & A298;
  assign \new_[306]_  = ~\new_[99]_  & \new_[305]_ ;
  assign \new_[307]_  = ~A299 & ~\new_[306]_ ;
  assign \new_[308]_  = ~\new_[130]_  & ~\new_[307]_ ;
  assign \new_[309]_  = ~\new_[304]_  & ~\new_[308]_ ;
  assign \new_[310]_  = ~\new_[300]_  & \new_[309]_ ;
  assign \new_[311]_  = ~\new_[263]_  & ~\new_[310]_ ;
  assign \new_[312]_  = ~\new_[280]_  & \new_[311]_ ;
  assign A109 = ~\new_[297]_  & \new_[312]_ ;
  assign \new_[314]_  = ~\new_[55]_  & ~\new_[143]_ ;
  assign \new_[315]_  = ~\new_[254]_  & \new_[314]_ ;
  assign \new_[316]_  = ~\new_[278]_  & \new_[315]_ ;
  assign \new_[317]_  = ~\new_[309]_  & \new_[316]_ ;
  assign \new_[318]_  = ~\new_[276]_  & ~\new_[317]_ ;
  assign A108 = ~\new_[297]_  & ~\new_[318]_ ;
  assign \new_[320]_  = ~\new_[96]_  & ~\new_[257]_ ;
  assign \new_[321]_  = ~\new_[296]_  & ~\new_[320]_ ;
  assign \new_[322]_  = \new_[300]_  & ~\new_[321]_ ;
  assign \new_[323]_  = ~\new_[279]_  & ~\new_[322]_ ;
  assign \new_[324]_  = ~\new_[284]_  & ~\new_[320]_ ;
  assign \new_[325]_  = \new_[300]_  & ~\new_[324]_ ;
  assign \new_[326]_  = ~\new_[276]_  & ~\new_[325]_ ;
  assign \new_[327]_  = ~\new_[105]_  & ~\new_[259]_ ;
  assign \new_[328]_  = ~\new_[326]_  & \new_[327]_ ;
  assign \new_[329]_  = ~\new_[323]_  & \new_[328]_ ;
  assign \new_[330]_  = ~\new_[308]_  & ~\new_[327]_ ;
  assign \new_[331]_  = ~\new_[276]_  & \new_[330]_ ;
  assign \new_[332]_  = ~\new_[304]_  & ~\new_[320]_ ;
  assign \new_[333]_  = ~\new_[296]_  & \new_[332]_ ;
  assign \new_[334]_  = \new_[300]_  & ~\new_[331]_ ;
  assign \new_[335]_  = ~\new_[333]_  & \new_[334]_ ;
  assign \new_[336]_  = ~\new_[279]_  & ~\new_[335]_ ;
  assign \new_[337]_  = ~\new_[284]_  & ~\new_[304]_ ;
  assign \new_[338]_  = ~\new_[320]_  & \new_[337]_ ;
  assign \new_[339]_  = \new_[300]_  & ~\new_[338]_ ;
  assign \new_[340]_  = ~\new_[276]_  & ~\new_[339]_ ;
  assign \new_[341]_  = ~\new_[284]_  & ~\new_[308]_ ;
  assign \new_[342]_  = ~\new_[327]_  & \new_[341]_ ;
  assign \new_[343]_  = ~\new_[296]_  & \new_[342]_ ;
  assign \new_[344]_  = ~\new_[340]_  & ~\new_[343]_ ;
  assign \new_[345]_  = ~\new_[336]_  & \new_[344]_ ;
  assign \new_[346]_  = ~\new_[105]_  & ~\new_[130]_ ;
  assign \new_[347]_  = ~\new_[307]_  & \new_[346]_ ;
  assign \new_[348]_  = ~\new_[259]_  & \new_[347]_ ;
  assign \new_[349]_  = ~\new_[255]_  & ~\new_[348]_ ;
  assign \new_[350]_  = ~\new_[300]_  & \new_[332]_ ;
  assign \new_[351]_  = ~\new_[349]_  & ~\new_[350]_ ;
  assign \new_[352]_  = ~\new_[280]_  & \new_[351]_ ;
  assign A105 = ~\new_[297]_  & \new_[352]_ ;
  assign \new_[354]_  = A236 & ~\new_[142]_ ;
  assign \new_[355]_  = ~A234 & ~\new_[354]_ ;
  assign \new_[356]_  = ~\new_[143]_  & ~\new_[355]_ ;
  assign \new_[357]_  = A302 & ~\new_[98]_ ;
  assign \new_[358]_  = A300 & ~\new_[131]_ ;
  assign \new_[359]_  = A269 & ~\new_[107]_ ;
  assign \new_[360]_  = A267 & ~\new_[123]_ ;
  assign \new_[361]_  = ~A301 & ~A268;
  assign \new_[362]_  = ~\new_[360]_  & \new_[361]_ ;
  assign \new_[363]_  = ~\new_[358]_  & \new_[362]_ ;
  assign \new_[364]_  = ~\new_[357]_  & ~\new_[359]_ ;
  assign \new_[365]_  = \new_[363]_  & \new_[364]_ ;
  assign \new_[366]_  = ~A235 & ~\new_[356]_ ;
  assign \new_[367]_  = ~\new_[365]_  & \new_[366]_ ;
  assign \new_[368]_  = A170 & ~\new_[82]_ ;
  assign \new_[369]_  = ~A168 & ~\new_[368]_ ;
  assign \new_[370]_  = ~\new_[83]_  & ~\new_[369]_ ;
  assign \new_[371]_  = A203 & ~\new_[68]_ ;
  assign \new_[372]_  = ~A201 & ~\new_[371]_ ;
  assign \new_[373]_  = ~\new_[69]_  & ~\new_[372]_ ;
  assign \new_[374]_  = ~A202 & ~A169;
  assign \new_[375]_  = ~\new_[373]_  & \new_[374]_ ;
  assign \new_[376]_  = ~\new_[370]_  & \new_[375]_ ;
  assign \new_[377]_  = ~A167 & A170;
  assign \new_[378]_  = ~A168 & ~\new_[377]_ ;
  assign \new_[379]_  = A166 & ~\new_[378]_ ;
  assign \new_[380]_  = ~A166 & A170;
  assign \new_[381]_  = ~A168 & ~\new_[380]_ ;
  assign \new_[382]_  = A167 & ~\new_[381]_ ;
  assign \new_[383]_  = ~A169 & ~\new_[382]_ ;
  assign \new_[384]_  = ~\new_[379]_  & \new_[383]_ ;
  assign \new_[385]_  = A203 & ~\new_[56]_ ;
  assign \new_[386]_  = A201 & ~\new_[69]_ ;
  assign \new_[387]_  = ~A202 & ~\new_[386]_ ;
  assign \new_[388]_  = ~\new_[385]_  & \new_[387]_ ;
  assign \new_[389]_  = ~\new_[384]_  & ~\new_[388]_ ;
  assign \new_[390]_  = A269 & ~\new_[122]_ ;
  assign \new_[391]_  = ~A267 & ~\new_[390]_ ;
  assign \new_[392]_  = ~\new_[123]_  & ~\new_[391]_ ;
  assign \new_[393]_  = A302 & ~\new_[130]_ ;
  assign \new_[394]_  = ~A300 & ~\new_[393]_ ;
  assign \new_[395]_  = ~\new_[131]_  & ~\new_[394]_ ;
  assign \new_[396]_  = A236 & ~\new_[118]_ ;
  assign \new_[397]_  = A234 & ~\new_[143]_ ;
  assign \new_[398]_  = ~A235 & ~\new_[397]_ ;
  assign \new_[399]_  = ~\new_[396]_  & \new_[398]_ ;
  assign \new_[400]_  = \new_[361]_  & ~\new_[399]_ ;
  assign \new_[401]_  = ~\new_[392]_  & ~\new_[395]_ ;
  assign \new_[402]_  = \new_[400]_  & \new_[401]_ ;
  assign \new_[403]_  = ~\new_[389]_  & ~\new_[402]_ ;
  assign \new_[404]_  = ~\new_[367]_  & ~\new_[376]_ ;
  assign A76 = \new_[403]_  & \new_[404]_ ;
  assign \new_[406]_  = \new_[361]_  & ~\new_[395]_ ;
  assign \new_[407]_  = ~\new_[392]_  & \new_[406]_ ;
  assign \new_[408]_  = ~\new_[366]_  & \new_[388]_ ;
  assign \new_[409]_  = ~\new_[407]_  & \new_[408]_ ;
  assign \new_[410]_  = ~\new_[384]_  & ~\new_[409]_ ;
  assign A75 = ~\new_[376]_  & ~\new_[410]_ ;
  assign \new_[412]_  = ~A301 & ~\new_[358]_ ;
  assign \new_[413]_  = ~\new_[357]_  & \new_[412]_ ;
  assign \new_[414]_  = ~A169 & ~\new_[413]_ ;
  assign \new_[415]_  = ~\new_[370]_  & \new_[414]_ ;
  assign \new_[416]_  = \new_[399]_  & ~\new_[415]_ ;
  assign \new_[417]_  = ~\new_[388]_  & ~\new_[416]_ ;
  assign \new_[418]_  = ~A202 & ~\new_[413]_ ;
  assign \new_[419]_  = ~\new_[373]_  & \new_[418]_ ;
  assign \new_[420]_  = \new_[399]_  & ~\new_[419]_ ;
  assign \new_[421]_  = ~\new_[384]_  & ~\new_[420]_ ;
  assign \new_[422]_  = ~A268 & ~\new_[360]_ ;
  assign \new_[423]_  = ~\new_[359]_  & \new_[422]_ ;
  assign \new_[424]_  = ~\new_[421]_  & \new_[423]_ ;
  assign \new_[425]_  = ~\new_[417]_  & \new_[424]_ ;
  assign \new_[426]_  = ~\new_[392]_  & ~\new_[413]_ ;
  assign \new_[427]_  = ~A268 & ~A169;
  assign \new_[428]_  = ~\new_[370]_  & \new_[427]_ ;
  assign \new_[429]_  = \new_[426]_  & \new_[428]_ ;
  assign \new_[430]_  = ~A301 & ~\new_[423]_ ;
  assign \new_[431]_  = ~\new_[395]_  & \new_[430]_ ;
  assign \new_[432]_  = ~\new_[384]_  & \new_[431]_ ;
  assign \new_[433]_  = \new_[399]_  & ~\new_[429]_ ;
  assign \new_[434]_  = ~\new_[432]_  & \new_[433]_ ;
  assign \new_[435]_  = ~\new_[388]_  & ~\new_[434]_ ;
  assign \new_[436]_  = ~A268 & ~A202;
  assign \new_[437]_  = ~\new_[373]_  & \new_[436]_ ;
  assign \new_[438]_  = \new_[426]_  & \new_[437]_ ;
  assign \new_[439]_  = \new_[399]_  & ~\new_[438]_ ;
  assign \new_[440]_  = ~\new_[384]_  & ~\new_[439]_ ;
  assign \new_[441]_  = ~A301 & \new_[374]_ ;
  assign \new_[442]_  = ~\new_[423]_  & \new_[441]_ ;
  assign \new_[443]_  = ~\new_[373]_  & ~\new_[395]_ ;
  assign \new_[444]_  = ~\new_[370]_  & \new_[443]_ ;
  assign \new_[445]_  = \new_[442]_  & \new_[444]_ ;
  assign \new_[446]_  = ~\new_[440]_  & ~\new_[445]_ ;
  assign \new_[447]_  = ~\new_[435]_  & \new_[446]_ ;
  assign \new_[448]_  = ~A301 & ~\new_[395]_ ;
  assign \new_[449]_  = \new_[423]_  & ~\new_[448]_ ;
  assign \new_[450]_  = \new_[366]_  & ~\new_[449]_ ;
  assign \new_[451]_  = ~A268 & ~\new_[413]_ ;
  assign \new_[452]_  = ~\new_[392]_  & ~\new_[399]_ ;
  assign \new_[453]_  = \new_[451]_  & \new_[452]_ ;
  assign \new_[454]_  = ~\new_[389]_  & ~\new_[453]_ ;
  assign \new_[455]_  = ~\new_[376]_  & \new_[454]_ ;
  assign A72 = ~\new_[450]_  & \new_[455]_ ;
  assign \new_[457]_  = ~A203 & A202;
  assign \new_[458]_  = ~\new_[70]_  & \new_[457]_ ;
  assign \new_[459]_  = ~A202 & \new_[385]_ ;
  assign \new_[460]_  = ~\new_[386]_  & ~\new_[458]_ ;
  assign \new_[461]_  = ~\new_[459]_  & \new_[460]_ ;
  assign \new_[462]_  = A168 & ~\new_[291]_ ;
  assign \new_[463]_  = \new_[52]_  & \new_[462]_ ;
  assign \new_[464]_  = ~\new_[51]_  & ~\new_[463]_ ;
  assign \new_[465]_  = ~\new_[461]_  & ~\new_[464]_ ;
  assign \new_[466]_  = A166 & \new_[462]_ ;
  assign \new_[467]_  = ~A167 & ~\new_[466]_ ;
  assign \new_[468]_  = ~\new_[82]_  & ~\new_[467]_ ;
  assign \new_[469]_  = A203 & ~A202;
  assign \new_[470]_  = ~\new_[56]_  & ~\new_[469]_ ;
  assign \new_[471]_  = \new_[68]_  & ~\new_[457]_ ;
  assign \new_[472]_  = ~\new_[470]_  & ~\new_[471]_ ;
  assign \new_[473]_  = ~\new_[468]_  & ~\new_[472]_ ;
  assign \new_[474]_  = ~A201 & \new_[473]_ ;
  assign \new_[475]_  = \new_[69]_  & ~\new_[457]_ ;
  assign \new_[476]_  = ~\new_[468]_  & \new_[475]_ ;
  assign \new_[477]_  = A236 & ~A235;
  assign \new_[478]_  = ~A302 & A301;
  assign \new_[479]_  = ~\new_[132]_  & \new_[478]_ ;
  assign \new_[480]_  = ~A301 & \new_[357]_ ;
  assign \new_[481]_  = ~A269 & A268;
  assign \new_[482]_  = ~\new_[124]_  & \new_[481]_ ;
  assign \new_[483]_  = ~A268 & \new_[359]_ ;
  assign \new_[484]_  = ~\new_[360]_  & ~\new_[482]_ ;
  assign \new_[485]_  = ~\new_[483]_  & \new_[484]_ ;
  assign \new_[486]_  = ~\new_[358]_  & ~\new_[479]_ ;
  assign \new_[487]_  = ~\new_[480]_  & \new_[486]_ ;
  assign \new_[488]_  = \new_[485]_  & \new_[487]_ ;
  assign \new_[489]_  = ~A234 & ~\new_[477]_ ;
  assign \new_[490]_  = ~\new_[488]_  & \new_[489]_ ;
  assign \new_[491]_  = A269 & ~A268;
  assign \new_[492]_  = A302 & ~A301;
  assign \new_[493]_  = ~\new_[98]_  & ~\new_[492]_ ;
  assign \new_[494]_  = \new_[130]_  & ~\new_[478]_ ;
  assign \new_[495]_  = ~\new_[493]_  & ~\new_[494]_ ;
  assign \new_[496]_  = ~\new_[107]_  & ~\new_[491]_ ;
  assign \new_[497]_  = ~\new_[495]_  & \new_[496]_ ;
  assign \new_[498]_  = \new_[122]_  & ~\new_[481]_ ;
  assign \new_[499]_  = ~\new_[495]_  & \new_[498]_ ;
  assign \new_[500]_  = ~\new_[497]_  & ~\new_[499]_ ;
  assign \new_[501]_  = ~A300 & ~\new_[500]_ ;
  assign \new_[502]_  = ~\new_[496]_  & ~\new_[498]_ ;
  assign \new_[503]_  = \new_[131]_  & ~\new_[478]_ ;
  assign \new_[504]_  = ~\new_[502]_  & \new_[503]_ ;
  assign \new_[505]_  = ~\new_[501]_  & ~\new_[504]_ ;
  assign \new_[506]_  = ~A267 & ~\new_[505]_ ;
  assign \new_[507]_  = ~A300 & ~\new_[495]_ ;
  assign \new_[508]_  = ~\new_[503]_  & ~\new_[507]_ ;
  assign \new_[509]_  = \new_[123]_  & ~\new_[481]_ ;
  assign \new_[510]_  = ~\new_[508]_  & \new_[509]_ ;
  assign \new_[511]_  = ~\new_[506]_  & ~\new_[510]_ ;
  assign \new_[512]_  = \new_[477]_  & ~\new_[511]_ ;
  assign \new_[513]_  = ~\new_[490]_  & ~\new_[512]_ ;
  assign \new_[514]_  = ~\new_[118]_  & ~\new_[513]_ ;
  assign \new_[515]_  = ~A234 & \new_[142]_ ;
  assign \new_[516]_  = ~\new_[143]_  & ~\new_[515]_ ;
  assign \new_[517]_  = ~A236 & A235;
  assign \new_[518]_  = ~\new_[516]_  & ~\new_[517]_ ;
  assign \new_[519]_  = ~\new_[488]_  & \new_[518]_ ;
  assign \new_[520]_  = ~\new_[144]_  & \new_[517]_ ;
  assign \new_[521]_  = ~\new_[397]_  & ~\new_[520]_ ;
  assign \new_[522]_  = ~A300 & ~\new_[521]_ ;
  assign \new_[523]_  = ~\new_[500]_  & \new_[522]_ ;
  assign \new_[524]_  = ~\new_[502]_  & ~\new_[521]_ ;
  assign \new_[525]_  = \new_[503]_  & \new_[524]_ ;
  assign \new_[526]_  = ~\new_[523]_  & ~\new_[525]_ ;
  assign \new_[527]_  = ~A267 & ~\new_[526]_ ;
  assign \new_[528]_  = ~\new_[495]_  & \new_[522]_ ;
  assign \new_[529]_  = \new_[503]_  & ~\new_[521]_ ;
  assign \new_[530]_  = ~\new_[528]_  & ~\new_[529]_ ;
  assign \new_[531]_  = \new_[509]_  & ~\new_[530]_ ;
  assign \new_[532]_  = ~\new_[465]_  & ~\new_[476]_ ;
  assign \new_[533]_  = ~\new_[519]_  & \new_[532]_ ;
  assign \new_[534]_  = ~\new_[474]_  & \new_[533]_ ;
  assign \new_[535]_  = ~\new_[531]_  & \new_[534]_ ;
  assign \new_[536]_  = ~\new_[527]_  & \new_[535]_ ;
  assign A43 = ~\new_[514]_  & \new_[536]_ ;
  assign \new_[538]_  = ~\new_[118]_  & ~\new_[477]_ ;
  assign \new_[539]_  = \new_[142]_  & ~\new_[517]_ ;
  assign \new_[540]_  = ~\new_[538]_  & ~\new_[539]_ ;
  assign \new_[541]_  = ~A234 & ~\new_[540]_ ;
  assign \new_[542]_  = ~\new_[464]_  & \new_[541]_ ;
  assign \new_[543]_  = \new_[143]_  & ~\new_[517]_ ;
  assign \new_[544]_  = ~\new_[386]_  & ~\new_[543]_ ;
  assign \new_[545]_  = ~\new_[458]_  & \new_[544]_ ;
  assign \new_[546]_  = ~\new_[459]_  & \new_[545]_ ;
  assign \new_[547]_  = \new_[511]_  & \new_[546]_ ;
  assign \new_[548]_  = ~\new_[464]_  & ~\new_[547]_ ;
  assign \new_[549]_  = ~\new_[476]_  & ~\new_[542]_ ;
  assign \new_[550]_  = ~\new_[474]_  & \new_[549]_ ;
  assign A42 = ~\new_[548]_  & \new_[550]_ ;
  assign \new_[552]_  = ~A235 & \new_[396]_ ;
  assign \new_[553]_  = \new_[521]_  & ~\new_[552]_ ;
  assign \new_[554]_  = \new_[460]_  & \new_[464]_ ;
  assign \new_[555]_  = ~\new_[459]_  & \new_[554]_ ;
  assign \new_[556]_  = ~\new_[553]_  & ~\new_[555]_ ;
  assign \new_[557]_  = ~\new_[468]_  & ~\new_[487]_ ;
  assign \new_[558]_  = ~\new_[461]_  & \new_[557]_ ;
  assign \new_[559]_  = ~\new_[464]_  & ~\new_[472]_ ;
  assign \new_[560]_  = ~\new_[487]_  & \new_[559]_ ;
  assign \new_[561]_  = ~A201 & \new_[560]_ ;
  assign \new_[562]_  = ~\new_[464]_  & ~\new_[487]_ ;
  assign \new_[563]_  = \new_[475]_  & \new_[562]_ ;
  assign \new_[564]_  = \new_[485]_  & ~\new_[563]_ ;
  assign \new_[565]_  = ~\new_[558]_  & ~\new_[561]_ ;
  assign \new_[566]_  = ~\new_[556]_  & \new_[565]_ ;
  assign \new_[567]_  = \new_[564]_  & \new_[566]_ ;
  assign \new_[568]_  = ~\new_[464]_  & \new_[507]_ ;
  assign \new_[569]_  = ~\new_[464]_  & \new_[503]_ ;
  assign \new_[570]_  = ~\new_[568]_  & ~\new_[569]_ ;
  assign \new_[571]_  = ~\new_[485]_  & ~\new_[570]_ ;
  assign \new_[572]_  = ~A267 & ~\new_[502]_ ;
  assign \new_[573]_  = ~\new_[468]_  & \new_[572]_ ;
  assign \new_[574]_  = ~\new_[487]_  & \new_[573]_ ;
  assign \new_[575]_  = \new_[509]_  & \new_[557]_ ;
  assign \new_[576]_  = ~\new_[574]_  & ~\new_[575]_ ;
  assign \new_[577]_  = ~\new_[571]_  & \new_[576]_ ;
  assign \new_[578]_  = ~\new_[461]_  & ~\new_[577]_ ;
  assign \new_[579]_  = ~A300 & \new_[491]_ ;
  assign \new_[580]_  = ~\new_[492]_  & \new_[579]_ ;
  assign \new_[581]_  = \new_[473]_  & \new_[580]_ ;
  assign \new_[582]_  = A302 & ~A267;
  assign \new_[583]_  = ~A301 & \new_[582]_ ;
  assign \new_[584]_  = ~\new_[491]_  & \new_[583]_ ;
  assign \new_[585]_  = \new_[559]_  & \new_[584]_ ;
  assign \new_[586]_  = ~\new_[581]_  & ~\new_[585]_ ;
  assign \new_[587]_  = ~\new_[98]_  & ~\new_[586]_ ;
  assign \new_[588]_  = ~A300 & \new_[130]_ ;
  assign \new_[589]_  = ~\new_[131]_  & ~\new_[588]_ ;
  assign \new_[590]_  = ~\new_[478]_  & \new_[491]_ ;
  assign \new_[591]_  = ~\new_[589]_  & \new_[590]_ ;
  assign \new_[592]_  = \new_[473]_  & \new_[591]_ ;
  assign \new_[593]_  = ~A267 & ~\new_[491]_ ;
  assign \new_[594]_  = ~\new_[486]_  & \new_[593]_ ;
  assign \new_[595]_  = \new_[559]_  & \new_[594]_ ;
  assign \new_[596]_  = ~\new_[592]_  & ~\new_[595]_ ;
  assign \new_[597]_  = ~\new_[587]_  & \new_[596]_ ;
  assign \new_[598]_  = ~\new_[107]_  & ~\new_[597]_ ;
  assign \new_[599]_  = ~A267 & \new_[122]_ ;
  assign \new_[600]_  = ~\new_[123]_  & ~\new_[599]_ ;
  assign \new_[601]_  = ~\new_[481]_  & ~\new_[600]_ ;
  assign \new_[602]_  = \new_[560]_  & \new_[601]_ ;
  assign \new_[603]_  = \new_[470]_  & ~\new_[495]_ ;
  assign \new_[604]_  = \new_[471]_  & ~\new_[495]_ ;
  assign \new_[605]_  = ~\new_[603]_  & ~\new_[604]_ ;
  assign \new_[606]_  = ~A300 & ~\new_[484]_ ;
  assign \new_[607]_  = ~\new_[468]_  & \new_[606]_ ;
  assign \new_[608]_  = ~\new_[605]_  & \new_[607]_ ;
  assign \new_[609]_  = ~\new_[484]_  & \new_[503]_ ;
  assign \new_[610]_  = ~\new_[472]_  & \new_[609]_ ;
  assign \new_[611]_  = ~\new_[468]_  & \new_[610]_ ;
  assign \new_[612]_  = ~\new_[608]_  & ~\new_[611]_ ;
  assign \new_[613]_  = ~\new_[602]_  & \new_[612]_ ;
  assign \new_[614]_  = ~\new_[598]_  & \new_[613]_ ;
  assign \new_[615]_  = ~A201 & ~\new_[614]_ ;
  assign \new_[616]_  = ~\new_[468]_  & \new_[580]_ ;
  assign \new_[617]_  = ~\new_[464]_  & \new_[584]_ ;
  assign \new_[618]_  = ~\new_[616]_  & ~\new_[617]_ ;
  assign \new_[619]_  = ~\new_[98]_  & ~\new_[618]_ ;
  assign \new_[620]_  = ~\new_[468]_  & \new_[591]_ ;
  assign \new_[621]_  = ~\new_[464]_  & \new_[594]_ ;
  assign \new_[622]_  = ~\new_[620]_  & ~\new_[621]_ ;
  assign \new_[623]_  = ~\new_[619]_  & \new_[622]_ ;
  assign \new_[624]_  = ~\new_[107]_  & ~\new_[623]_ ;
  assign \new_[625]_  = \new_[562]_  & \new_[601]_ ;
  assign \new_[626]_  = ~\new_[495]_  & \new_[606]_ ;
  assign \new_[627]_  = ~\new_[468]_  & \new_[626]_ ;
  assign \new_[628]_  = ~\new_[468]_  & \new_[609]_ ;
  assign \new_[629]_  = ~\new_[627]_  & ~\new_[628]_ ;
  assign \new_[630]_  = ~\new_[625]_  & \new_[629]_ ;
  assign \new_[631]_  = ~\new_[624]_  & \new_[630]_ ;
  assign \new_[632]_  = \new_[475]_  & ~\new_[631]_ ;
  assign \new_[633]_  = ~\new_[556]_  & ~\new_[578]_ ;
  assign \new_[634]_  = ~\new_[632]_  & \new_[633]_ ;
  assign \new_[635]_  = ~\new_[615]_  & \new_[634]_ ;
  assign \new_[636]_  = \new_[485]_  & ~\new_[503]_ ;
  assign \new_[637]_  = ~\new_[507]_  & \new_[636]_ ;
  assign \new_[638]_  = \new_[489]_  & ~\new_[637]_ ;
  assign \new_[639]_  = ~\new_[487]_  & \new_[572]_ ;
  assign \new_[640]_  = ~\new_[487]_  & \new_[509]_ ;
  assign \new_[641]_  = ~\new_[639]_  & ~\new_[640]_ ;
  assign \new_[642]_  = \new_[477]_  & ~\new_[641]_ ;
  assign \new_[643]_  = ~\new_[638]_  & ~\new_[642]_ ;
  assign \new_[644]_  = ~\new_[118]_  & ~\new_[643]_ ;
  assign \new_[645]_  = \new_[518]_  & ~\new_[637]_ ;
  assign \new_[646]_  = ~A267 & ~\new_[487]_ ;
  assign \new_[647]_  = \new_[524]_  & \new_[646]_ ;
  assign \new_[648]_  = \new_[509]_  & ~\new_[521]_ ;
  assign \new_[649]_  = ~\new_[487]_  & \new_[648]_ ;
  assign \new_[650]_  = ~\new_[476]_  & ~\new_[649]_ ;
  assign \new_[651]_  = ~\new_[465]_  & \new_[650]_ ;
  assign \new_[652]_  = ~\new_[474]_  & ~\new_[647]_ ;
  assign \new_[653]_  = \new_[651]_  & \new_[652]_ ;
  assign \new_[654]_  = ~\new_[645]_  & \new_[653]_ ;
  assign A39 = ~\new_[644]_  & \new_[654]_ ;
  assign \new_[656]_  = A300 & ~\new_[492]_ ;
  assign \new_[657]_  = A302 & ~A300;
  assign \new_[658]_  = ~A301 & \new_[657]_ ;
  assign \new_[659]_  = ~\new_[656]_  & ~\new_[658]_ ;
  assign \new_[660]_  = ~\new_[98]_  & ~\new_[107]_ ;
  assign \new_[661]_  = ~\new_[659]_  & \new_[660]_ ;
  assign \new_[662]_  = A267 & \new_[661]_ ;
  assign \new_[663]_  = ~A300 & ~\new_[492]_ ;
  assign \new_[664]_  = A302 & A300;
  assign \new_[665]_  = ~A301 & \new_[664]_ ;
  assign \new_[666]_  = \new_[132]_  & ~\new_[665]_ ;
  assign \new_[667]_  = ~\new_[663]_  & \new_[666]_ ;
  assign \new_[668]_  = ~A267 & ~\new_[667]_ ;
  assign \new_[669]_  = ~\new_[662]_  & ~\new_[668]_ ;
  assign \new_[670]_  = ~\new_[491]_  & ~\new_[669]_ ;
  assign \new_[671]_  = ~A267 & ~\new_[107]_ ;
  assign \new_[672]_  = ~\new_[98]_  & \new_[671]_ ;
  assign \new_[673]_  = A300 & \new_[672]_ ;
  assign \new_[674]_  = ~A300 & A267;
  assign \new_[675]_  = ~\new_[673]_  & ~\new_[674]_ ;
  assign \new_[676]_  = \new_[491]_  & ~\new_[675]_ ;
  assign \new_[677]_  = ~A300 & ~\new_[124]_ ;
  assign \new_[678]_  = ~\new_[676]_  & ~\new_[677]_ ;
  assign \new_[679]_  = ~\new_[492]_  & ~\new_[678]_ ;
  assign \new_[680]_  = A269 & A267;
  assign \new_[681]_  = ~A268 & \new_[680]_ ;
  assign \new_[682]_  = \new_[124]_  & ~\new_[681]_ ;
  assign \new_[683]_  = ~\new_[666]_  & ~\new_[682]_ ;
  assign \new_[684]_  = \new_[491]_  & \new_[658]_ ;
  assign \new_[685]_  = \new_[672]_  & \new_[684]_ ;
  assign \new_[686]_  = A201 & ~\new_[469]_ ;
  assign \new_[687]_  = A203 & ~A201;
  assign \new_[688]_  = ~A202 & \new_[687]_ ;
  assign \new_[689]_  = ~\new_[686]_  & ~\new_[688]_ ;
  assign \new_[690]_  = ~\new_[56]_  & ~\new_[689]_ ;
  assign \new_[691]_  = ~A168 & ~\new_[291]_ ;
  assign \new_[692]_  = A168 & \new_[291]_ ;
  assign \new_[693]_  = \new_[84]_  & ~\new_[692]_ ;
  assign \new_[694]_  = ~\new_[691]_  & \new_[693]_ ;
  assign \new_[695]_  = ~\new_[690]_  & \new_[694]_ ;
  assign \new_[696]_  = ~A234 & ~\new_[695]_ ;
  assign \new_[697]_  = ~A168 & \new_[291]_ ;
  assign \new_[698]_  = ~\new_[462]_  & ~\new_[697]_ ;
  assign \new_[699]_  = ~A201 & ~\new_[469]_ ;
  assign \new_[700]_  = A203 & A201;
  assign \new_[701]_  = ~A202 & \new_[700]_ ;
  assign \new_[702]_  = \new_[70]_  & ~\new_[701]_ ;
  assign \new_[703]_  = ~\new_[699]_  & \new_[702]_ ;
  assign \new_[704]_  = A234 & ~\new_[118]_ ;
  assign \new_[705]_  = ~\new_[53]_  & \new_[704]_ ;
  assign \new_[706]_  = ~\new_[698]_  & \new_[705]_ ;
  assign \new_[707]_  = ~\new_[703]_  & \new_[706]_ ;
  assign \new_[708]_  = ~\new_[696]_  & ~\new_[707]_ ;
  assign \new_[709]_  = ~\new_[477]_  & ~\new_[708]_ ;
  assign \new_[710]_  = A236 & A234;
  assign \new_[711]_  = ~A235 & \new_[710]_ ;
  assign \new_[712]_  = \new_[144]_  & ~\new_[711]_ ;
  assign \new_[713]_  = ~\new_[56]_  & ~\new_[712]_ ;
  assign \new_[714]_  = ~\new_[689]_  & \new_[713]_ ;
  assign \new_[715]_  = ~A168 & ~\new_[712]_ ;
  assign \new_[716]_  = ~\new_[53]_  & ~\new_[118]_ ;
  assign \new_[717]_  = ~\new_[703]_  & \new_[716]_ ;
  assign \new_[718]_  = ~A234 & A168;
  assign \new_[719]_  = \new_[477]_  & \new_[718]_ ;
  assign \new_[720]_  = \new_[717]_  & \new_[719]_ ;
  assign \new_[721]_  = ~\new_[715]_  & ~\new_[720]_ ;
  assign \new_[722]_  = ~\new_[291]_  & ~\new_[721]_ ;
  assign \new_[723]_  = ~\new_[693]_  & ~\new_[712]_ ;
  assign \new_[724]_  = ~A234 & ~A168;
  assign \new_[725]_  = \new_[477]_  & \new_[724]_ ;
  assign \new_[726]_  = \new_[291]_  & \new_[725]_ ;
  assign \new_[727]_  = \new_[717]_  & \new_[726]_ ;
  assign \new_[728]_  = ~\new_[683]_  & ~\new_[723]_ ;
  assign \new_[729]_  = ~\new_[714]_  & \new_[728]_ ;
  assign \new_[730]_  = ~\new_[685]_  & \new_[729]_ ;
  assign \new_[731]_  = ~\new_[727]_  & \new_[730]_ ;
  assign \new_[732]_  = ~\new_[670]_  & \new_[731]_ ;
  assign \new_[733]_  = ~\new_[709]_  & ~\new_[722]_ ;
  assign \new_[734]_  = \new_[732]_  & \new_[733]_ ;
  assign A6 = ~\new_[679]_  & \new_[734]_ ;
  assign \new_[736]_  = ~\new_[53]_  & ~\new_[698]_ ;
  assign \new_[737]_  = \new_[703]_  & ~\new_[736]_ ;
  assign \new_[738]_  = ~A267 & ~\new_[737]_ ;
  assign \new_[739]_  = ~\new_[489]_  & \new_[712]_ ;
  assign \new_[740]_  = ~\new_[694]_  & ~\new_[739]_ ;
  assign \new_[741]_  = A267 & ~\new_[107]_ ;
  assign \new_[742]_  = \new_[740]_  & \new_[741]_ ;
  assign \new_[743]_  = ~\new_[738]_  & ~\new_[742]_ ;
  assign \new_[744]_  = ~A300 & ~\new_[743]_ ;
  assign \new_[745]_  = ~\new_[53]_  & ~\new_[107]_ ;
  assign \new_[746]_  = A267 & A168;
  assign \new_[747]_  = \new_[745]_  & \new_[746]_ ;
  assign \new_[748]_  = ~\new_[188]_  & ~\new_[747]_ ;
  assign \new_[749]_  = ~\new_[291]_  & ~\new_[739]_ ;
  assign \new_[750]_  = ~\new_[748]_  & \new_[749]_ ;
  assign \new_[751]_  = A267 & ~A168;
  assign \new_[752]_  = \new_[745]_  & \new_[751]_ ;
  assign \new_[753]_  = ~A267 & A168;
  assign \new_[754]_  = ~\new_[752]_  & ~\new_[753]_ ;
  assign \new_[755]_  = \new_[291]_  & ~\new_[754]_ ;
  assign \new_[756]_  = ~A267 & ~\new_[84]_ ;
  assign \new_[757]_  = ~\new_[755]_  & ~\new_[756]_ ;
  assign \new_[758]_  = ~\new_[739]_  & ~\new_[757]_ ;
  assign \new_[759]_  = ~\new_[750]_  & ~\new_[758]_ ;
  assign \new_[760]_  = ~\new_[98]_  & ~\new_[759]_ ;
  assign \new_[761]_  = A300 & \new_[760]_ ;
  assign \new_[762]_  = ~\new_[744]_  & ~\new_[761]_ ;
  assign \new_[763]_  = ~\new_[492]_  & ~\new_[762]_ ;
  assign \new_[764]_  = ~\new_[666]_  & ~\new_[743]_ ;
  assign \new_[765]_  = \new_[658]_  & \new_[760]_ ;
  assign \new_[766]_  = ~\new_[764]_  & ~\new_[765]_ ;
  assign \new_[767]_  = ~\new_[763]_  & \new_[766]_ ;
  assign \new_[768]_  = ~\new_[491]_  & ~\new_[767]_ ;
  assign \new_[769]_  = ~A300 & ~\new_[737]_ ;
  assign \new_[770]_  = ~\new_[98]_  & \new_[740]_ ;
  assign \new_[771]_  = A300 & \new_[770]_ ;
  assign \new_[772]_  = ~\new_[769]_  & ~\new_[771]_ ;
  assign \new_[773]_  = ~\new_[492]_  & ~\new_[772]_ ;
  assign \new_[774]_  = ~\new_[666]_  & ~\new_[737]_ ;
  assign \new_[775]_  = \new_[658]_  & \new_[770]_ ;
  assign \new_[776]_  = ~\new_[774]_  & ~\new_[775]_ ;
  assign \new_[777]_  = ~\new_[773]_  & \new_[776]_ ;
  assign \new_[778]_  = ~\new_[682]_  & ~\new_[777]_ ;
  assign \new_[779]_  = \new_[690]_  & ~\new_[739]_ ;
  assign \new_[780]_  = A269 & ~A267;
  assign \new_[781]_  = ~A268 & \new_[780]_ ;
  assign \new_[782]_  = ~\new_[98]_  & \new_[781]_ ;
  assign \new_[783]_  = ~\new_[107]_  & \new_[782]_ ;
  assign \new_[784]_  = ~\new_[659]_  & \new_[783]_ ;
  assign \new_[785]_  = ~\new_[739]_  & \new_[784]_ ;
  assign \new_[786]_  = ~\new_[779]_  & ~\new_[785]_ ;
  assign \new_[787]_  = \new_[63]_  & ~\new_[786]_ ;
  assign \new_[788]_  = ~\new_[107]_  & \new_[781]_ ;
  assign \new_[789]_  = ~\new_[667]_  & \new_[788]_ ;
  assign \new_[790]_  = \new_[703]_  & ~\new_[789]_ ;
  assign \new_[791]_  = ~A168 & ~\new_[739]_ ;
  assign \new_[792]_  = ~\new_[790]_  & \new_[791]_ ;
  assign \new_[793]_  = ~\new_[787]_  & ~\new_[792]_ ;
  assign \new_[794]_  = ~\new_[291]_  & ~\new_[793]_ ;
  assign \new_[795]_  = \new_[661]_  & \new_[781]_ ;
  assign \new_[796]_  = ~\new_[690]_  & ~\new_[795]_ ;
  assign \new_[797]_  = ~A168 & ~\new_[53]_ ;
  assign \new_[798]_  = ~\new_[796]_  & \new_[797]_ ;
  assign \new_[799]_  = A168 & ~\new_[790]_ ;
  assign \new_[800]_  = ~\new_[798]_  & ~\new_[799]_ ;
  assign \new_[801]_  = \new_[291]_  & ~\new_[800]_ ;
  assign \new_[802]_  = ~\new_[84]_  & ~\new_[790]_ ;
  assign \new_[803]_  = ~\new_[801]_  & ~\new_[802]_ ;
  assign \new_[804]_  = ~\new_[739]_  & ~\new_[803]_ ;
  assign \new_[805]_  = ~\new_[794]_  & ~\new_[804]_ ;
  assign \new_[806]_  = ~\new_[778]_  & \new_[805]_ ;
  assign A7 = ~\new_[768]_  & \new_[806]_ ;
  assign \new_[808]_  = A234 & ~\new_[477]_ ;
  assign \new_[809]_  = A236 & ~A234;
  assign \new_[810]_  = ~A235 & \new_[809]_ ;
  assign \new_[811]_  = ~\new_[808]_  & ~\new_[810]_ ;
  assign \new_[812]_  = ~\new_[98]_  & ~\new_[811]_ ;
  assign \new_[813]_  = ~\new_[659]_  & \new_[812]_ ;
  assign \new_[814]_  = A267 & ~\new_[491]_ ;
  assign \new_[815]_  = ~\new_[781]_  & ~\new_[814]_ ;
  assign \new_[816]_  = ~\new_[107]_  & ~\new_[815]_ ;
  assign \new_[817]_  = ~\new_[811]_  & \new_[816]_ ;
  assign \new_[818]_  = ~\new_[813]_  & ~\new_[817]_ ;
  assign \new_[819]_  = ~\new_[118]_  & ~\new_[818]_ ;
  assign \new_[820]_  = ~\new_[593]_  & \new_[682]_ ;
  assign \new_[821]_  = ~\new_[98]_  & ~\new_[659]_ ;
  assign \new_[822]_  = ~\new_[820]_  & \new_[821]_ ;
  assign \new_[823]_  = ~\new_[667]_  & \new_[816]_ ;
  assign \new_[824]_  = ~\new_[822]_  & ~\new_[823]_ ;
  assign \new_[825]_  = \new_[736]_  & ~\new_[824]_ ;
  assign \new_[826]_  = ~\new_[690]_  & ~\new_[825]_ ;
  assign \new_[827]_  = ~\new_[819]_  & \new_[826]_ ;
  assign \new_[828]_  = ~\new_[694]_  & ~\new_[703]_ ;
  assign \new_[829]_  = ~\new_[489]_  & ~\new_[663]_ ;
  assign \new_[830]_  = \new_[712]_  & \new_[829]_ ;
  assign \new_[831]_  = \new_[666]_  & \new_[830]_ ;
  assign \new_[832]_  = ~\new_[828]_  & \new_[831]_ ;
  assign \new_[833]_  = ~A267 & ~\new_[832]_ ;
  assign \new_[834]_  = ~\new_[662]_  & ~\new_[833]_ ;
  assign \new_[835]_  = ~\new_[491]_  & ~\new_[834]_ ;
  assign \new_[836]_  = ~\new_[682]_  & ~\new_[832]_ ;
  assign \new_[837]_  = ~\new_[795]_  & ~\new_[836]_ ;
  assign A9 = ~\new_[835]_  & \new_[837]_ ;
  assign \new_[839]_  = ~\new_[690]_  & ~\new_[736]_ ;
  assign \new_[840]_  = ~A234 & ~\new_[839]_ ;
  assign \new_[841]_  = ~\new_[118]_  & \new_[828]_ ;
  assign \new_[842]_  = A234 & \new_[841]_ ;
  assign \new_[843]_  = ~\new_[840]_  & ~\new_[842]_ ;
  assign \new_[844]_  = ~\new_[477]_  & ~\new_[843]_ ;
  assign \new_[845]_  = ~\new_[53]_  & ~\new_[712]_ ;
  assign \new_[846]_  = ~\new_[698]_  & \new_[845]_ ;
  assign \new_[847]_  = \new_[810]_  & \new_[841]_ ;
  assign \new_[848]_  = ~\new_[683]_  & ~\new_[846]_ ;
  assign \new_[849]_  = ~\new_[685]_  & ~\new_[714]_ ;
  assign \new_[850]_  = \new_[848]_  & \new_[849]_ ;
  assign \new_[851]_  = ~\new_[847]_  & \new_[850]_ ;
  assign \new_[852]_  = ~\new_[670]_  & \new_[851]_ ;
  assign \new_[853]_  = ~\new_[844]_  & \new_[852]_ ;
  assign A10 = ~\new_[679]_  & \new_[853]_ ;
  assign A140 = ~\new_[187]_ ;
  assign A139 = ~\new_[221]_ ;
  assign A107 = ~\new_[329]_ ;
  assign A106 = ~\new_[345]_ ;
  assign A74 = ~\new_[425]_ ;
  assign A73 = ~\new_[447]_ ;
  assign A41 = ~\new_[567]_ ;
  assign A40 = ~\new_[635]_ ;
  assign A8 = ~\new_[827]_ ;
endmodule


