module top ( clock, 
    p_30, p_20, p_10, p_12, p_23, p_34, p_11, p_24, p_33, pclk, p_14, p_21,
    p_32, p_13, p_22, p_31, p_16, p_27, p_15, p_28, p_9, p_18, p_25, p_8,
    p_17, p_26, p_7, p_6, p_19, p_5, p_29, p_4, p_3, p_1,
    p_68  );
  input  clock;
  input  p_30, p_20, p_10, p_12, p_23, p_34, p_11, p_24, p_33, pclk,
    p_14, p_21, p_32, p_13, p_22, p_31, p_16, p_27, p_15, p_28, p_9, p_18,
    p_25, p_8, p_17, p_26, p_7, p_6, p_19, p_5, p_29, p_4, p_3, p_1;
  output p_68;
  reg n_44, n_40, n_41, n_42, n_43, n_36, n_37, n_38, n_39, n_2, n_45, n_56,
    n_46, n_55, n_47, n_58, n_65, n_48, n_57, n_66, n_49, n_60, n_50, n_59,
    n_51, n_62, n_52, n_61, n_53, n_64, n_54, n_63;
  wire new_n132_1_, new_n133_, new_n134_, new_n136_, new_n137_1_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_1_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_1_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_1_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_1_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_1_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_1_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_1_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_1_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_1_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_1_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_1_,
    new_n193_, new_n194_, new_n195_, new_n197_1_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_1_, new_n203_, new_n204_, new_n205_,
    new_n207_1_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_1_,
    new_n213_, new_n214_, new_n215_, new_n217_1_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_1_, new_n223_, new_n224_, new_n225_,
    new_n227_1_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, n72, n77, n82, n87, n92, n97, n102, n107, n112, n117, n122,
    n127, n132, n137, n142, n147, n152, n157, n162, n167, n172, n177, n182,
    n187, n192, n197, n202, n207, n212, n217, n222, n227;
  assign new_n132_1_ = p_3 & p_1;
  assign new_n133_ = ~n_36 & new_n132_1_;
  assign new_n134_ = n_36 & ~new_n132_1_;
  assign p_68 = new_n133_ | new_n134_;
  assign new_n136_ = p_11 & p_1;
  assign new_n137_1_ = n_44 & new_n136_;
  assign new_n138_ = p_10 & p_1;
  assign new_n139_ = n_43 & new_n138_;
  assign new_n140_ = p_9 & p_1;
  assign new_n141_ = n_42 & new_n140_;
  assign new_n142_1_ = p_8 & p_1;
  assign new_n143_ = n_41 & new_n142_1_;
  assign new_n144_ = p_7 & p_1;
  assign new_n145_ = n_40 & new_n144_;
  assign new_n146_ = p_6 & p_1;
  assign new_n147_1_ = n_39 & new_n146_;
  assign new_n148_ = p_5 & p_1;
  assign new_n149_ = n_38 & new_n148_;
  assign new_n150_ = p_4 & p_1;
  assign new_n151_ = n_37 & new_n150_;
  assign new_n152_1_ = n_36 & new_n132_1_;
  assign new_n153_ = n_37 & new_n152_1_;
  assign new_n154_ = new_n150_ & new_n152_1_;
  assign new_n155_ = ~new_n151_ & ~new_n153_;
  assign new_n156_ = ~new_n154_ & new_n155_;
  assign new_n157_1_ = n_38 & ~new_n156_;
  assign new_n158_ = new_n148_ & ~new_n156_;
  assign new_n159_ = ~new_n149_ & ~new_n157_1_;
  assign new_n160_ = ~new_n158_ & new_n159_;
  assign new_n161_ = n_39 & ~new_n160_;
  assign new_n162_1_ = new_n146_ & ~new_n160_;
  assign new_n163_ = ~new_n147_1_ & ~new_n161_;
  assign new_n164_ = ~new_n162_1_ & new_n163_;
  assign new_n165_ = n_40 & ~new_n164_;
  assign new_n166_ = new_n144_ & ~new_n164_;
  assign new_n167_1_ = ~new_n145_ & ~new_n165_;
  assign new_n168_ = ~new_n166_ & new_n167_1_;
  assign new_n169_ = n_41 & ~new_n168_;
  assign new_n170_ = new_n142_1_ & ~new_n168_;
  assign new_n171_ = ~new_n143_ & ~new_n169_;
  assign new_n172_1_ = ~new_n170_ & new_n171_;
  assign new_n173_ = n_42 & ~new_n172_1_;
  assign new_n174_ = new_n140_ & ~new_n172_1_;
  assign new_n175_ = ~new_n141_ & ~new_n173_;
  assign new_n176_ = ~new_n174_ & new_n175_;
  assign new_n177_1_ = n_43 & ~new_n176_;
  assign new_n178_ = new_n138_ & ~new_n176_;
  assign new_n179_ = ~new_n139_ & ~new_n177_1_;
  assign new_n180_ = ~new_n178_ & new_n179_;
  assign new_n181_ = n_44 & ~new_n180_;
  assign new_n182_1_ = new_n136_ & ~new_n180_;
  assign new_n183_ = ~new_n137_1_ & ~new_n181_;
  assign new_n184_ = ~new_n182_1_ & new_n183_;
  assign new_n185_ = p_12 & p_1;
  assign new_n186_ = ~new_n184_ & new_n185_;
  assign new_n187_1_ = n_45 & new_n186_;
  assign new_n188_ = new_n184_ & new_n185_;
  assign new_n189_ = ~n_45 & new_n188_;
  assign new_n190_ = new_n184_ & ~new_n185_;
  assign new_n191_ = n_45 & new_n190_;
  assign new_n192_1_ = ~new_n184_ & ~new_n185_;
  assign new_n193_ = ~n_45 & new_n192_1_;
  assign new_n194_ = ~new_n191_ & ~new_n193_;
  assign new_n195_ = ~new_n187_1_ & ~new_n189_;
  assign n72 = ~new_n194_ | ~new_n195_;
  assign new_n197_1_ = n_41 & new_n170_;
  assign new_n198_ = new_n142_1_ & new_n168_;
  assign new_n199_ = ~n_41 & new_n198_;
  assign new_n200_ = ~new_n142_1_ & new_n168_;
  assign new_n201_ = n_41 & new_n200_;
  assign new_n202_1_ = ~new_n142_1_ & ~new_n168_;
  assign new_n203_ = ~n_41 & new_n202_1_;
  assign new_n204_ = ~new_n201_ & ~new_n203_;
  assign new_n205_ = ~new_n197_1_ & ~new_n199_;
  assign n77 = ~new_n204_ | ~new_n205_;
  assign new_n207_1_ = n_42 & new_n174_;
  assign new_n208_ = new_n140_ & new_n172_1_;
  assign new_n209_ = ~n_42 & new_n208_;
  assign new_n210_ = ~new_n140_ & new_n172_1_;
  assign new_n211_ = n_42 & new_n210_;
  assign new_n212_1_ = ~new_n140_ & ~new_n172_1_;
  assign new_n213_ = ~n_42 & new_n212_1_;
  assign new_n214_ = ~new_n211_ & ~new_n213_;
  assign new_n215_ = ~new_n207_1_ & ~new_n209_;
  assign n82 = ~new_n214_ | ~new_n215_;
  assign new_n217_1_ = n_43 & new_n178_;
  assign new_n218_ = new_n138_ & new_n176_;
  assign new_n219_ = ~n_43 & new_n218_;
  assign new_n220_ = ~new_n138_ & new_n176_;
  assign new_n221_ = n_43 & new_n220_;
  assign new_n222_1_ = ~new_n138_ & ~new_n176_;
  assign new_n223_ = ~n_43 & new_n222_1_;
  assign new_n224_ = ~new_n221_ & ~new_n223_;
  assign new_n225_ = ~new_n217_1_ & ~new_n219_;
  assign n87 = ~new_n224_ | ~new_n225_;
  assign new_n227_1_ = n_44 & new_n182_1_;
  assign new_n228_ = new_n136_ & new_n180_;
  assign new_n229_ = ~n_44 & new_n228_;
  assign new_n230_ = ~new_n136_ & new_n180_;
  assign new_n231_ = n_44 & new_n230_;
  assign new_n232_ = ~new_n136_ & ~new_n180_;
  assign new_n233_ = ~n_44 & new_n232_;
  assign new_n234_ = ~new_n231_ & ~new_n233_;
  assign new_n235_ = ~new_n227_1_ & ~new_n229_;
  assign n92 = ~new_n234_ | ~new_n235_;
  assign new_n237_ = n_37 & new_n154_;
  assign new_n238_ = new_n150_ & ~new_n152_1_;
  assign new_n239_ = ~n_37 & new_n238_;
  assign new_n240_ = ~new_n150_ & ~new_n152_1_;
  assign new_n241_ = n_37 & new_n240_;
  assign new_n242_ = ~new_n150_ & new_n152_1_;
  assign new_n243_ = ~n_37 & new_n242_;
  assign new_n244_ = ~new_n241_ & ~new_n243_;
  assign new_n245_ = ~new_n237_ & ~new_n239_;
  assign n97 = ~new_n244_ | ~new_n245_;
  assign new_n247_ = n_38 & new_n158_;
  assign new_n248_ = new_n148_ & new_n156_;
  assign new_n249_ = ~n_38 & new_n248_;
  assign new_n250_ = ~new_n148_ & new_n156_;
  assign new_n251_ = n_38 & new_n250_;
  assign new_n252_ = ~new_n148_ & ~new_n156_;
  assign new_n253_ = ~n_38 & new_n252_;
  assign new_n254_ = ~new_n251_ & ~new_n253_;
  assign new_n255_ = ~new_n247_ & ~new_n249_;
  assign n102 = ~new_n254_ | ~new_n255_;
  assign new_n257_ = n_39 & new_n162_1_;
  assign new_n258_ = new_n146_ & new_n160_;
  assign new_n259_ = ~n_39 & new_n258_;
  assign new_n260_ = ~new_n146_ & new_n160_;
  assign new_n261_ = n_39 & new_n260_;
  assign new_n262_ = ~new_n146_ & ~new_n160_;
  assign new_n263_ = ~n_39 & new_n262_;
  assign new_n264_ = ~new_n261_ & ~new_n263_;
  assign new_n265_ = ~new_n257_ & ~new_n259_;
  assign n107 = ~new_n264_ | ~new_n265_;
  assign new_n267_ = n_40 & new_n166_;
  assign new_n268_ = new_n144_ & new_n164_;
  assign new_n269_ = ~n_40 & new_n268_;
  assign new_n270_ = ~new_n144_ & new_n164_;
  assign new_n271_ = n_40 & new_n270_;
  assign new_n272_ = ~new_n144_ & ~new_n164_;
  assign new_n273_ = ~n_40 & new_n272_;
  assign new_n274_ = ~new_n271_ & ~new_n273_;
  assign new_n275_ = ~new_n267_ & ~new_n269_;
  assign n112 = ~new_n274_ | ~new_n275_;
  assign new_n277_ = p_33 & p_1;
  assign new_n278_ = n_66 & new_n277_;
  assign new_n279_ = p_32 & p_1;
  assign new_n280_ = n_65 & new_n279_;
  assign new_n281_ = p_31 & p_1;
  assign new_n282_ = n_64 & new_n281_;
  assign new_n283_ = p_30 & p_1;
  assign new_n284_ = n_63 & new_n283_;
  assign new_n285_ = p_29 & p_1;
  assign new_n286_ = n_62 & new_n285_;
  assign new_n287_ = p_28 & p_1;
  assign new_n288_ = n_61 & new_n287_;
  assign new_n289_ = p_27 & p_1;
  assign new_n290_ = n_60 & new_n289_;
  assign new_n291_ = p_26 & p_1;
  assign new_n292_ = n_59 & new_n291_;
  assign new_n293_ = p_25 & p_1;
  assign new_n294_ = n_58 & new_n293_;
  assign new_n295_ = p_24 & p_1;
  assign new_n296_ = n_57 & new_n295_;
  assign new_n297_ = p_23 & p_1;
  assign new_n298_ = n_56 & new_n297_;
  assign new_n299_ = p_22 & p_1;
  assign new_n300_ = n_55 & new_n299_;
  assign new_n301_ = p_21 & p_1;
  assign new_n302_ = n_54 & new_n301_;
  assign new_n303_ = p_20 & p_1;
  assign new_n304_ = n_53 & new_n303_;
  assign new_n305_ = p_19 & p_1;
  assign new_n306_ = n_52 & new_n305_;
  assign new_n307_ = p_18 & p_1;
  assign new_n308_ = n_51 & new_n307_;
  assign new_n309_ = p_17 & p_1;
  assign new_n310_ = n_50 & new_n309_;
  assign new_n311_ = p_16 & p_1;
  assign new_n312_ = n_49 & new_n311_;
  assign new_n313_ = p_15 & p_1;
  assign new_n314_ = n_48 & new_n313_;
  assign new_n315_ = p_14 & p_1;
  assign new_n316_ = n_47 & new_n315_;
  assign new_n317_ = p_13 & p_1;
  assign new_n318_ = n_46 & new_n317_;
  assign new_n319_ = n_45 & new_n185_;
  assign new_n320_ = n_45 & ~new_n184_;
  assign new_n321_ = ~new_n319_ & ~new_n320_;
  assign new_n322_ = ~new_n186_ & new_n321_;
  assign new_n323_ = n_46 & ~new_n322_;
  assign new_n324_ = new_n317_ & ~new_n322_;
  assign new_n325_ = ~new_n318_ & ~new_n323_;
  assign new_n326_ = ~new_n324_ & new_n325_;
  assign new_n327_ = n_47 & ~new_n326_;
  assign new_n328_ = new_n315_ & ~new_n326_;
  assign new_n329_ = ~new_n316_ & ~new_n327_;
  assign new_n330_ = ~new_n328_ & new_n329_;
  assign new_n331_ = n_48 & ~new_n330_;
  assign new_n332_ = new_n313_ & ~new_n330_;
  assign new_n333_ = ~new_n314_ & ~new_n331_;
  assign new_n334_ = ~new_n332_ & new_n333_;
  assign new_n335_ = n_49 & ~new_n334_;
  assign new_n336_ = new_n311_ & ~new_n334_;
  assign new_n337_ = ~new_n312_ & ~new_n335_;
  assign new_n338_ = ~new_n336_ & new_n337_;
  assign new_n339_ = n_50 & ~new_n338_;
  assign new_n340_ = new_n309_ & ~new_n338_;
  assign new_n341_ = ~new_n310_ & ~new_n339_;
  assign new_n342_ = ~new_n340_ & new_n341_;
  assign new_n343_ = n_51 & ~new_n342_;
  assign new_n344_ = new_n307_ & ~new_n342_;
  assign new_n345_ = ~new_n308_ & ~new_n343_;
  assign new_n346_ = ~new_n344_ & new_n345_;
  assign new_n347_ = n_52 & ~new_n346_;
  assign new_n348_ = new_n305_ & ~new_n346_;
  assign new_n349_ = ~new_n306_ & ~new_n347_;
  assign new_n350_ = ~new_n348_ & new_n349_;
  assign new_n351_ = n_53 & ~new_n350_;
  assign new_n352_ = new_n303_ & ~new_n350_;
  assign new_n353_ = ~new_n304_ & ~new_n351_;
  assign new_n354_ = ~new_n352_ & new_n353_;
  assign new_n355_ = n_54 & ~new_n354_;
  assign new_n356_ = new_n301_ & ~new_n354_;
  assign new_n357_ = ~new_n302_ & ~new_n355_;
  assign new_n358_ = ~new_n356_ & new_n357_;
  assign new_n359_ = n_55 & ~new_n358_;
  assign new_n360_ = new_n299_ & ~new_n358_;
  assign new_n361_ = ~new_n300_ & ~new_n359_;
  assign new_n362_ = ~new_n360_ & new_n361_;
  assign new_n363_ = n_56 & ~new_n362_;
  assign new_n364_ = new_n297_ & ~new_n362_;
  assign new_n365_ = ~new_n298_ & ~new_n363_;
  assign new_n366_ = ~new_n364_ & new_n365_;
  assign new_n367_ = n_57 & ~new_n366_;
  assign new_n368_ = new_n295_ & ~new_n366_;
  assign new_n369_ = ~new_n296_ & ~new_n367_;
  assign new_n370_ = ~new_n368_ & new_n369_;
  assign new_n371_ = n_58 & ~new_n370_;
  assign new_n372_ = new_n293_ & ~new_n370_;
  assign new_n373_ = ~new_n294_ & ~new_n371_;
  assign new_n374_ = ~new_n372_ & new_n373_;
  assign new_n375_ = n_59 & ~new_n374_;
  assign new_n376_ = new_n291_ & ~new_n374_;
  assign new_n377_ = ~new_n292_ & ~new_n375_;
  assign new_n378_ = ~new_n376_ & new_n377_;
  assign new_n379_ = n_60 & ~new_n378_;
  assign new_n380_ = new_n289_ & ~new_n378_;
  assign new_n381_ = ~new_n290_ & ~new_n379_;
  assign new_n382_ = ~new_n380_ & new_n381_;
  assign new_n383_ = n_61 & ~new_n382_;
  assign new_n384_ = new_n287_ & ~new_n382_;
  assign new_n385_ = ~new_n288_ & ~new_n383_;
  assign new_n386_ = ~new_n384_ & new_n385_;
  assign new_n387_ = n_62 & ~new_n386_;
  assign new_n388_ = new_n285_ & ~new_n386_;
  assign new_n389_ = ~new_n286_ & ~new_n387_;
  assign new_n390_ = ~new_n388_ & new_n389_;
  assign new_n391_ = n_63 & ~new_n390_;
  assign new_n392_ = new_n283_ & ~new_n390_;
  assign new_n393_ = ~new_n284_ & ~new_n391_;
  assign new_n394_ = ~new_n392_ & new_n393_;
  assign new_n395_ = n_64 & ~new_n394_;
  assign new_n396_ = new_n281_ & ~new_n394_;
  assign new_n397_ = ~new_n282_ & ~new_n395_;
  assign new_n398_ = ~new_n396_ & new_n397_;
  assign new_n399_ = n_65 & ~new_n398_;
  assign new_n400_ = new_n279_ & ~new_n398_;
  assign new_n401_ = ~new_n280_ & ~new_n399_;
  assign new_n402_ = ~new_n400_ & new_n401_;
  assign new_n403_ = n_66 & ~new_n402_;
  assign new_n404_ = new_n277_ & ~new_n402_;
  assign new_n405_ = ~new_n278_ & ~new_n403_;
  assign new_n406_ = ~new_n404_ & new_n405_;
  assign new_n407_ = p_34 & p_1;
  assign new_n408_ = n_2 & new_n407_;
  assign new_n409_ = new_n406_ & new_n408_;
  assign new_n410_ = n_2 & ~new_n407_;
  assign new_n411_ = ~new_n406_ & new_n410_;
  assign new_n412_ = ~new_n409_ & ~new_n411_;
  assign new_n413_ = ~n_2 & new_n407_;
  assign new_n414_ = ~new_n406_ & new_n413_;
  assign new_n415_ = ~new_n406_ & new_n408_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign n117 = ~new_n412_ | ~new_n416_;
  assign new_n418_ = n_46 & new_n324_;
  assign new_n419_ = new_n317_ & new_n322_;
  assign new_n420_ = ~n_46 & new_n419_;
  assign new_n421_ = ~new_n317_ & new_n322_;
  assign new_n422_ = n_46 & new_n421_;
  assign new_n423_ = ~new_n317_ & ~new_n322_;
  assign new_n424_ = ~n_46 & new_n423_;
  assign new_n425_ = ~new_n422_ & ~new_n424_;
  assign new_n426_ = ~new_n418_ & ~new_n420_;
  assign n122 = ~new_n425_ | ~new_n426_;
  assign new_n428_ = n_57 & new_n368_;
  assign new_n429_ = new_n295_ & new_n366_;
  assign new_n430_ = ~n_57 & new_n429_;
  assign new_n431_ = ~new_n295_ & new_n366_;
  assign new_n432_ = n_57 & new_n431_;
  assign new_n433_ = ~new_n295_ & ~new_n366_;
  assign new_n434_ = ~n_57 & new_n433_;
  assign new_n435_ = ~new_n432_ & ~new_n434_;
  assign new_n436_ = ~new_n428_ & ~new_n430_;
  assign n127 = ~new_n435_ | ~new_n436_;
  assign new_n438_ = n_47 & new_n328_;
  assign new_n439_ = new_n315_ & new_n326_;
  assign new_n440_ = ~n_47 & new_n439_;
  assign new_n441_ = ~new_n315_ & new_n326_;
  assign new_n442_ = n_47 & new_n441_;
  assign new_n443_ = ~new_n315_ & ~new_n326_;
  assign new_n444_ = ~n_47 & new_n443_;
  assign new_n445_ = ~new_n442_ & ~new_n444_;
  assign new_n446_ = ~new_n438_ & ~new_n440_;
  assign n132 = ~new_n445_ | ~new_n446_;
  assign new_n448_ = n_56 & new_n364_;
  assign new_n449_ = new_n297_ & new_n362_;
  assign new_n450_ = ~n_56 & new_n449_;
  assign new_n451_ = ~new_n297_ & new_n362_;
  assign new_n452_ = n_56 & new_n451_;
  assign new_n453_ = ~new_n297_ & ~new_n362_;
  assign new_n454_ = ~n_56 & new_n453_;
  assign new_n455_ = ~new_n452_ & ~new_n454_;
  assign new_n456_ = ~new_n448_ & ~new_n450_;
  assign n137 = ~new_n455_ | ~new_n456_;
  assign new_n458_ = n_48 & new_n332_;
  assign new_n459_ = new_n313_ & new_n330_;
  assign new_n460_ = ~n_48 & new_n459_;
  assign new_n461_ = ~new_n313_ & new_n330_;
  assign new_n462_ = n_48 & new_n461_;
  assign new_n463_ = ~new_n313_ & ~new_n330_;
  assign new_n464_ = ~n_48 & new_n463_;
  assign new_n465_ = ~new_n462_ & ~new_n464_;
  assign new_n466_ = ~new_n458_ & ~new_n460_;
  assign n142 = ~new_n465_ | ~new_n466_;
  assign new_n468_ = n_59 & new_n376_;
  assign new_n469_ = new_n291_ & new_n374_;
  assign new_n470_ = ~n_59 & new_n469_;
  assign new_n471_ = ~new_n291_ & new_n374_;
  assign new_n472_ = n_59 & new_n471_;
  assign new_n473_ = ~new_n291_ & ~new_n374_;
  assign new_n474_ = ~n_59 & new_n473_;
  assign new_n475_ = ~new_n472_ & ~new_n474_;
  assign new_n476_ = ~new_n468_ & ~new_n470_;
  assign n147 = ~new_n475_ | ~new_n476_;
  assign new_n478_ = n_66 & new_n404_;
  assign new_n479_ = new_n277_ & new_n402_;
  assign new_n480_ = ~n_66 & new_n479_;
  assign new_n481_ = ~new_n277_ & new_n402_;
  assign new_n482_ = n_66 & new_n481_;
  assign new_n483_ = ~new_n277_ & ~new_n402_;
  assign new_n484_ = ~n_66 & new_n483_;
  assign new_n485_ = ~new_n482_ & ~new_n484_;
  assign new_n486_ = ~new_n478_ & ~new_n480_;
  assign n152 = ~new_n485_ | ~new_n486_;
  assign new_n488_ = n_49 & new_n336_;
  assign new_n489_ = new_n311_ & new_n334_;
  assign new_n490_ = ~n_49 & new_n489_;
  assign new_n491_ = ~new_n311_ & new_n334_;
  assign new_n492_ = n_49 & new_n491_;
  assign new_n493_ = ~new_n311_ & ~new_n334_;
  assign new_n494_ = ~n_49 & new_n493_;
  assign new_n495_ = ~new_n492_ & ~new_n494_;
  assign new_n496_ = ~new_n488_ & ~new_n490_;
  assign n157 = ~new_n495_ | ~new_n496_;
  assign new_n498_ = n_58 & new_n372_;
  assign new_n499_ = new_n293_ & new_n370_;
  assign new_n500_ = ~n_58 & new_n499_;
  assign new_n501_ = ~new_n293_ & new_n370_;
  assign new_n502_ = n_58 & new_n501_;
  assign new_n503_ = ~new_n293_ & ~new_n370_;
  assign new_n504_ = ~n_58 & new_n503_;
  assign new_n505_ = ~new_n502_ & ~new_n504_;
  assign new_n506_ = ~new_n498_ & ~new_n500_;
  assign n162 = ~new_n505_ | ~new_n506_;
  assign new_n508_ = ~new_n406_ & ~new_n407_;
  assign new_n509_ = new_n406_ & new_n407_;
  assign new_n510_ = ~new_n508_ & ~new_n509_;
  assign new_n511_ = ~n_2 & ~new_n510_;
  assign new_n512_ = n_2 & new_n510_;
  assign n167 = new_n511_ | new_n512_;
  assign new_n514_ = n_50 & new_n340_;
  assign new_n515_ = new_n309_ & new_n338_;
  assign new_n516_ = ~n_50 & new_n515_;
  assign new_n517_ = ~new_n309_ & new_n338_;
  assign new_n518_ = n_50 & new_n517_;
  assign new_n519_ = ~new_n309_ & ~new_n338_;
  assign new_n520_ = ~n_50 & new_n519_;
  assign new_n521_ = ~new_n518_ & ~new_n520_;
  assign new_n522_ = ~new_n514_ & ~new_n516_;
  assign n172 = ~new_n521_ | ~new_n522_;
  assign new_n524_ = n_61 & new_n384_;
  assign new_n525_ = new_n287_ & new_n382_;
  assign new_n526_ = ~n_61 & new_n525_;
  assign new_n527_ = ~new_n287_ & new_n382_;
  assign new_n528_ = n_61 & new_n527_;
  assign new_n529_ = ~new_n287_ & ~new_n382_;
  assign new_n530_ = ~n_61 & new_n529_;
  assign new_n531_ = ~new_n528_ & ~new_n530_;
  assign new_n532_ = ~new_n524_ & ~new_n526_;
  assign n177 = ~new_n531_ | ~new_n532_;
  assign new_n534_ = n_51 & new_n344_;
  assign new_n535_ = new_n307_ & new_n342_;
  assign new_n536_ = ~n_51 & new_n535_;
  assign new_n537_ = ~new_n307_ & new_n342_;
  assign new_n538_ = n_51 & new_n537_;
  assign new_n539_ = ~new_n307_ & ~new_n342_;
  assign new_n540_ = ~n_51 & new_n539_;
  assign new_n541_ = ~new_n538_ & ~new_n540_;
  assign new_n542_ = ~new_n534_ & ~new_n536_;
  assign n182 = ~new_n541_ | ~new_n542_;
  assign new_n544_ = n_60 & new_n380_;
  assign new_n545_ = new_n289_ & new_n378_;
  assign new_n546_ = ~n_60 & new_n545_;
  assign new_n547_ = ~new_n289_ & new_n378_;
  assign new_n548_ = n_60 & new_n547_;
  assign new_n549_ = ~new_n289_ & ~new_n378_;
  assign new_n550_ = ~n_60 & new_n549_;
  assign new_n551_ = ~new_n548_ & ~new_n550_;
  assign new_n552_ = ~new_n544_ & ~new_n546_;
  assign n187 = ~new_n551_ | ~new_n552_;
  assign new_n554_ = n_52 & new_n348_;
  assign new_n555_ = new_n305_ & new_n346_;
  assign new_n556_ = ~n_52 & new_n555_;
  assign new_n557_ = ~new_n305_ & new_n346_;
  assign new_n558_ = n_52 & new_n557_;
  assign new_n559_ = ~new_n305_ & ~new_n346_;
  assign new_n560_ = ~n_52 & new_n559_;
  assign new_n561_ = ~new_n558_ & ~new_n560_;
  assign new_n562_ = ~new_n554_ & ~new_n556_;
  assign n192 = ~new_n561_ | ~new_n562_;
  assign new_n564_ = n_63 & new_n392_;
  assign new_n565_ = new_n283_ & new_n390_;
  assign new_n566_ = ~n_63 & new_n565_;
  assign new_n567_ = ~new_n283_ & new_n390_;
  assign new_n568_ = n_63 & new_n567_;
  assign new_n569_ = ~new_n283_ & ~new_n390_;
  assign new_n570_ = ~n_63 & new_n569_;
  assign new_n571_ = ~new_n568_ & ~new_n570_;
  assign new_n572_ = ~new_n564_ & ~new_n566_;
  assign n197 = ~new_n571_ | ~new_n572_;
  assign new_n574_ = n_53 & new_n352_;
  assign new_n575_ = new_n303_ & new_n350_;
  assign new_n576_ = ~n_53 & new_n575_;
  assign new_n577_ = ~new_n303_ & new_n350_;
  assign new_n578_ = n_53 & new_n577_;
  assign new_n579_ = ~new_n303_ & ~new_n350_;
  assign new_n580_ = ~n_53 & new_n579_;
  assign new_n581_ = ~new_n578_ & ~new_n580_;
  assign new_n582_ = ~new_n574_ & ~new_n576_;
  assign n202 = ~new_n581_ | ~new_n582_;
  assign new_n584_ = n_62 & new_n388_;
  assign new_n585_ = new_n285_ & new_n386_;
  assign new_n586_ = ~n_62 & new_n585_;
  assign new_n587_ = ~new_n285_ & new_n386_;
  assign new_n588_ = n_62 & new_n587_;
  assign new_n589_ = ~new_n285_ & ~new_n386_;
  assign new_n590_ = ~n_62 & new_n589_;
  assign new_n591_ = ~new_n588_ & ~new_n590_;
  assign new_n592_ = ~new_n584_ & ~new_n586_;
  assign n207 = ~new_n591_ | ~new_n592_;
  assign new_n594_ = n_54 & new_n356_;
  assign new_n595_ = new_n301_ & new_n354_;
  assign new_n596_ = ~n_54 & new_n595_;
  assign new_n597_ = ~new_n301_ & new_n354_;
  assign new_n598_ = n_54 & new_n597_;
  assign new_n599_ = ~new_n301_ & ~new_n354_;
  assign new_n600_ = ~n_54 & new_n599_;
  assign new_n601_ = ~new_n598_ & ~new_n600_;
  assign new_n602_ = ~new_n594_ & ~new_n596_;
  assign n212 = ~new_n601_ | ~new_n602_;
  assign new_n604_ = n_65 & new_n400_;
  assign new_n605_ = new_n279_ & new_n398_;
  assign new_n606_ = ~n_65 & new_n605_;
  assign new_n607_ = ~new_n279_ & new_n398_;
  assign new_n608_ = n_65 & new_n607_;
  assign new_n609_ = ~new_n279_ & ~new_n398_;
  assign new_n610_ = ~n_65 & new_n609_;
  assign new_n611_ = ~new_n608_ & ~new_n610_;
  assign new_n612_ = ~new_n604_ & ~new_n606_;
  assign n217 = ~new_n611_ | ~new_n612_;
  assign new_n614_ = n_55 & new_n360_;
  assign new_n615_ = new_n299_ & new_n358_;
  assign new_n616_ = ~n_55 & new_n615_;
  assign new_n617_ = ~new_n299_ & new_n358_;
  assign new_n618_ = n_55 & new_n617_;
  assign new_n619_ = ~new_n299_ & ~new_n358_;
  assign new_n620_ = ~n_55 & new_n619_;
  assign new_n621_ = ~new_n618_ & ~new_n620_;
  assign new_n622_ = ~new_n614_ & ~new_n616_;
  assign n222 = ~new_n621_ | ~new_n622_;
  assign new_n624_ = n_64 & new_n396_;
  assign new_n625_ = new_n281_ & new_n394_;
  assign new_n626_ = ~n_64 & new_n625_;
  assign new_n627_ = ~new_n281_ & new_n394_;
  assign new_n628_ = n_64 & new_n627_;
  assign new_n629_ = ~new_n281_ & ~new_n394_;
  assign new_n630_ = ~n_64 & new_n629_;
  assign new_n631_ = ~new_n628_ & ~new_n630_;
  assign new_n632_ = ~new_n624_ & ~new_n626_;
  assign n227 = ~new_n631_ | ~new_n632_;
  always @ (posedge clock) begin
    n_44 <= n72;
    n_40 <= n77;
    n_41 <= n82;
    n_42 <= n87;
    n_43 <= n92;
    n_36 <= n97;
    n_37 <= n102;
    n_38 <= n107;
    n_39 <= n112;
    n_2 <= n117;
    n_45 <= n122;
    n_56 <= n127;
    n_46 <= n132;
    n_55 <= n137;
    n_47 <= n142;
    n_58 <= n147;
    n_65 <= n152;
    n_48 <= n157;
    n_57 <= n162;
    n_66 <= n167;
    n_49 <= n172;
    n_60 <= n177;
    n_50 <= n182;
    n_59 <= n187;
    n_51 <= n192;
    n_62 <= n197;
    n_52 <= n202;
    n_61 <= n207;
    n_53 <= n212;
    n_64 <= n217;
    n_54 <= n222;
    n_63 <= n227;
  end
endmodule

