module top ( clock, 
    pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_,
    pkey_243_, pcount_2_, pkey_4_, pkey_132_, pkey_143_, pkey_158_,
    pkey_169_, pkey_231_, pkey_242_, pcount_1_, pkey_7_, pkey_146_,
    pkey_159_, pkey_168_, pkey_245_, pcount_0_, pkey_6_, pkey_130_,
    pkey_145_, pkey_167_, pkey_244_, pkey_9_, pkey_16_, pkey_27_, pkey_38_,
    pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_, pkey_221_,
    pkey_247_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_39_, pkey_48_,
    pkey_110_, pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_,
    pkey_246_, pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_47_,
    pkey_111_, pkey_120_, pkey_155_, pkey_164_, pkey_210_, pkey_249_,
    pkey_254_, pkey_19_, pkey_28_, pkey_37_, pkey_46_, pkey_112_,
    pkey_149_, pkey_156_, pkey_163_, pkey_211_, pkey_248_, pkey_255_,
    pkey_56_, pkey_67_, pkey_78_, pkey_89_, pkey_113_, pkey_126_,
    pkey_139_, pkey_162_, pkey_212_, pkey_225_, pkey_238_, pkey_57_,
    pkey_66_, pkey_79_, pkey_88_, pkey_114_, pkey_125_, pkey_150_,
    pkey_161_, pkey_213_, pkey_224_, pkey_239_, pkey_58_, pkey_69_,
    pkey_76_, pkey_87_, pkey_115_, pkey_124_, pkey_137_, pkey_151_,
    pkey_160_, pkey_214_, pkey_223_, pkey_236_, pkey_250_, pkey_59_,
    pkey_68_, pkey_77_, pkey_86_, pkey_116_, pkey_123_, pkey_138_,
    pkey_152_, pkey_215_, pkey_222_, pkey_237_, pkey_251_, pkey_1_,
    pkey_96_, pkey_117_, pkey_135_, pkey_140_, pkey_216_, pkey_229_,
    pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_,
    pkey_217_, pkey_228_, pkey_235_, pkey_3_, pkey_98_, pkey_119_,
    pkey_128_, pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_,
    pkey_241_, pkey_2_, pkey_99_, pkey_127_, pkey_134_, pkey_141_,
    pkey_219_, pkey_226_, pkey_233_, pkey_240_, pkey_70_, pkey_81_,
    pkey_92_, pkey_108_, pkey_180_, pkey_193_, pkey_207_, pkey_71_,
    pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, pclk, pkey_50_,
    pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_, pstart_0_,
    pkey_51_, pkey_60_, pkey_95_, pkey_109_, pkey_181_, pkey_196_,
    pkey_208_, pkey_52_, pkey_63_, pkey_74_, pkey_85_, pkey_104_,
    pkey_171_, pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_,
    pkey_75_, pkey_84_, pkey_103_, pkey_172_, pkey_198_, pkey_202_,
    pkey_54_, pkey_65_, pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_199_,
    pkey_205_, pkey_55_, pkey_64_, pkey_73_, pkey_82_, pkey_91_, pkey_105_,
    pkey_170_, pkey_204_, pkey_12_, pkey_23_, pkey_34_, pkey_45_,
    pkey_100_, pkey_175_, pkey_188_, pkey_13_, pkey_22_, pkey_35_,
    pkey_44_, pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_,
    pkey_102_, pkey_173_, pkey_201_, pkey_15_, pkey_24_, pkey_33_,
    pkey_42_, pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_,
    pkey_41_, pkey_179_, pkey_184_, pkey_31_, pkey_40_, pkey_183_,
    pkey_190_, pkey_10_, pkey_21_, pkey_177_, pkey_186_, pkey_191_,
    pkey_11_, pkey_20_, pkey_178_, pkey_185_, pkey_192_,
    pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_, pksi_115_,
    pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_, pksi_82_,
    pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_, pksi_63_,
    pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_, pksi_62_,
    pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_, pksi_65_,
    pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_, pksi_191_,
    pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_, pksi_56_,
    pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_, pksi_57_,
    pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_,
    pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_,
    pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_,
    pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_,
    pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_,
    pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_,
    pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_,
    pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_,
    pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_,
    pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_,
    pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_,
    pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_,
    pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_,
    pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_,
    pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_,
    pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_,
    pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_,
    pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_,
    pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_,
    pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_,
    pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_,
    pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_,
    pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_,
    pksi_161_  );
  input  clock;
  input  pcount_3_, pkey_5_, pkey_131_, pkey_144_, pkey_157_, pkey_230_,
    pkey_243_, pcount_2_, pkey_4_, pkey_132_, pkey_143_, pkey_158_,
    pkey_169_, pkey_231_, pkey_242_, pcount_1_, pkey_7_, pkey_146_,
    pkey_159_, pkey_168_, pkey_245_, pcount_0_, pkey_6_, pkey_130_,
    pkey_145_, pkey_167_, pkey_244_, pkey_9_, pkey_16_, pkey_27_, pkey_38_,
    pkey_49_, pkey_122_, pkey_148_, pkey_153_, pkey_166_, pkey_221_,
    pkey_247_, pkey_252_, pkey_8_, pkey_17_, pkey_26_, pkey_39_, pkey_48_,
    pkey_110_, pkey_121_, pkey_147_, pkey_154_, pkey_165_, pkey_220_,
    pkey_246_, pkey_253_, pkey_18_, pkey_29_, pkey_36_, pkey_47_,
    pkey_111_, pkey_120_, pkey_155_, pkey_164_, pkey_210_, pkey_249_,
    pkey_254_, pkey_19_, pkey_28_, pkey_37_, pkey_46_, pkey_112_,
    pkey_149_, pkey_156_, pkey_163_, pkey_211_, pkey_248_, pkey_255_,
    pkey_56_, pkey_67_, pkey_78_, pkey_89_, pkey_113_, pkey_126_,
    pkey_139_, pkey_162_, pkey_212_, pkey_225_, pkey_238_, pkey_57_,
    pkey_66_, pkey_79_, pkey_88_, pkey_114_, pkey_125_, pkey_150_,
    pkey_161_, pkey_213_, pkey_224_, pkey_239_, pkey_58_, pkey_69_,
    pkey_76_, pkey_87_, pkey_115_, pkey_124_, pkey_137_, pkey_151_,
    pkey_160_, pkey_214_, pkey_223_, pkey_236_, pkey_250_, pkey_59_,
    pkey_68_, pkey_77_, pkey_86_, pkey_116_, pkey_123_, pkey_138_,
    pkey_152_, pkey_215_, pkey_222_, pkey_237_, pkey_251_, pkey_1_,
    pkey_96_, pkey_117_, pkey_135_, pkey_140_, pkey_216_, pkey_229_,
    pkey_234_, pkey_0_, pkey_97_, pkey_118_, pkey_129_, pkey_136_,
    pkey_217_, pkey_228_, pkey_235_, pkey_3_, pkey_98_, pkey_119_,
    pkey_128_, pkey_133_, pkey_142_, pkey_218_, pkey_227_, pkey_232_,
    pkey_241_, pkey_2_, pkey_99_, pkey_127_, pkey_134_, pkey_141_,
    pkey_219_, pkey_226_, pkey_233_, pkey_240_, pkey_70_, pkey_81_,
    pkey_92_, pkey_108_, pkey_180_, pkey_193_, pkey_207_, pkey_71_,
    pkey_80_, pkey_93_, pkey_107_, pkey_194_, pkey_206_, pclk, pkey_50_,
    pkey_61_, pkey_94_, pkey_182_, pkey_195_, pkey_209_, pstart_0_,
    pkey_51_, pkey_60_, pkey_95_, pkey_109_, pkey_181_, pkey_196_,
    pkey_208_, pkey_52_, pkey_63_, pkey_74_, pkey_85_, pkey_104_,
    pkey_171_, pkey_197_, pkey_203_, pencrypt_0_, pkey_53_, pkey_62_,
    pkey_75_, pkey_84_, pkey_103_, pkey_172_, pkey_198_, pkey_202_,
    pkey_54_, pkey_65_, pkey_72_, pkey_83_, pkey_90_, pkey_106_, pkey_199_,
    pkey_205_, pkey_55_, pkey_64_, pkey_73_, pkey_82_, pkey_91_, pkey_105_,
    pkey_170_, pkey_204_, pkey_12_, pkey_23_, pkey_34_, pkey_45_,
    pkey_100_, pkey_175_, pkey_188_, pkey_13_, pkey_22_, pkey_35_,
    pkey_44_, pkey_176_, pkey_187_, pkey_14_, pkey_25_, pkey_32_, pkey_43_,
    pkey_102_, pkey_173_, pkey_201_, pkey_15_, pkey_24_, pkey_33_,
    pkey_42_, pkey_101_, pkey_174_, pkey_189_, pkey_200_, pkey_30_,
    pkey_41_, pkey_179_, pkey_184_, pkey_31_, pkey_40_, pkey_183_,
    pkey_190_, pkey_10_, pkey_21_, pkey_177_, pkey_186_, pkey_191_,
    pkey_11_, pkey_20_, pkey_178_, pkey_185_, pkey_192_;
  output pksi_50_, pksi_61_, pksi_72_, pksi_83_, pksi_94_, pksi_102_,
    pksi_115_, pksi_128_, pdata_ready_0_, pksi_51_, pksi_60_, pksi_73_,
    pksi_82_, pksi_95_, pksi_101_, pksi_116_, pksi_127_, pksi_52_,
    pksi_63_, pksi_70_, pksi_81_, pksi_96_, pksi_100_, pksi_113_, pksi_53_,
    pksi_62_, pksi_71_, pksi_80_, pksi_97_, pksi_114_, pksi_129_, pksi_54_,
    pksi_65_, pksi_76_, pksi_87_, pksi_90_, pksi_119_, pksi_124_,
    pksi_191_, pksi_55_, pksi_64_, pksi_77_, pksi_86_, pksi_91_, pksi_123_,
    pksi_56_, pksi_67_, pksi_74_, pksi_85_, pksi_92_, pksi_117_, pksi_126_,
    pksi_57_, pksi_66_, pksi_75_, pksi_84_, pksi_93_, pksi_118_, pksi_125_,
    pksi_190_, pksi_14_, pksi_25_, pksi_36_, pksi_47_, pksi_120_, pksi_15_,
    pksi_24_, pksi_37_, pksi_46_, pksi_109_, pnew_count_3_, pksi_16_,
    pksi_27_, pksi_34_, pksi_45_, pksi_108_, pksi_122_, pksi_17_, pksi_26_,
    pksi_35_, pksi_44_, pksi_107_, pksi_121_, pksi_10_, pksi_21_, pksi_32_,
    pksi_43_, pksi_106_, pksi_111_, pnew_count_0_, pksi_11_, pksi_20_,
    pksi_33_, pksi_42_, pksi_105_, pksi_112_, pksi_12_, pksi_23_, pksi_30_,
    pksi_41_, pksi_104_, pnew_count_2_, pksi_13_, pksi_22_, pksi_31_,
    pksi_40_, pksi_103_, pksi_110_, pnew_count_1_, pksi_3_, pksi_151_,
    pksi_164_, pksi_177_, pksi_2_, pksi_152_, pksi_163_, pksi_178_,
    pksi_189_, pksi_1_, pksi_166_, pksi_179_, pksi_188_, pksi_0_,
    pksi_150_, pksi_165_, pksi_187_, pksi_18_, pksi_29_, pksi_142_,
    pksi_168_, pksi_173_, pksi_186_, pksi_19_, pksi_28_, pksi_130_,
    pksi_141_, pksi_167_, pksi_174_, pksi_185_, pksi_38_, pksi_49_,
    pksi_131_, pksi_140_, pksi_175_, pksi_184_, pksi_39_, pksi_48_,
    pksi_132_, pksi_169_, pksi_176_, pksi_183_, pksi_58_, pksi_69_,
    pksi_133_, pksi_146_, pksi_159_, pksi_182_, pksi_59_, pksi_68_,
    pksi_134_, pksi_145_, pksi_170_, pksi_181_, pksi_9_, pksi_78_,
    pksi_89_, pksi_135_, pksi_144_, pksi_157_, pksi_171_, pksi_180_,
    pksi_8_, pksi_79_, pksi_88_, pksi_136_, pksi_143_, pksi_158_,
    pksi_172_, pksi_7_, pksi_98_, pksi_137_, pksi_155_, pksi_160_, pksi_6_,
    pksi_99_, pksi_138_, pksi_149_, pksi_156_, pksi_5_, pksi_139_,
    pksi_148_, pksi_153_, pksi_162_, pksi_4_, pksi_147_, pksi_154_,
    pksi_161_;
  reg n_n2365, n_n2375, n_n2879, n_n2392, n_n2402, n_n2411, n_n2448,
    n_n2982, n_n2366, n_n2865, n_n2881, n_n2391, n_n2403, n_n2917, n_n2449,
    n_n2457, n_n2367, n_n2377, n_n2384, n_n2390, n_n2419, n_n2429, n_n2450,
    n_n2459, n_n2465, n_n2368, n_n2376, n_n2877, n_n2389, n_n2420, n_n2428,
    n_n2451, n_n2458, n_n2285, n_n2362, n_n2372, n_n2382, n_n2889, n_n2435,
    n_n2444, n_n2454, n_n2463, n_n2363, n_n2371, n_n2383, n_n2388, n_n2954,
    n_n2964, n_n2445, n_n2464, n_n2364, n_n2374, n_n2380, n_n2387, n_n2446,
    n_n2456, n_n2853, n_n2373, n_n2381, n_n2885, n_n2447, n_n2455, n_n2462,
    n_n2282, n_n2395, n_n2909, n_n2413, n_n2423, n_n2432, n_n2441, n_n2741,
    n_n2396, n_n2404, n_n2414, n_n2422, n_n2433, n_n2440, n_n2283, n_n2899,
    n_n2406, n_n2412, n_n2421, n_n2950, n_n2443, n_n2284, n_n2397, n_n2405,
    n_n2921, n_n2931, n_n2434, n_n2442, n_n2279, n_n2369, n_n2379, n_n2398,
    n_n2408, n_n2417, n_n2427, n_n2430, n_n2437, n_n2452, n_n2460, n_n2280,
    n_n2370, n_n2378, n_n2399, n_n2407, n_n2418, n_n2426, n_n2943, n_n2436,
    n_n2453, n_n2986, n_n2737, n_n2385, n_n2394, n_n2400, n_n2410, n_n2415,
    n_n2425, n_n2945, n_n2439, n_n2976, n_n2281, n_n2386, n_n2393, n_n2401,
    n_n2409, n_n2416, n_n2424, n_n2431, n_n2438, n_n2461, n_n2319, n_n2329,
    n_n2338, n_n2348, n_n2843, n_n2320, n_n2328, n_n2339, n_n2347, n_n2357,
    n_n2321, n_n2330, n_n2336, n_n2346, n_n2358, n_n2278, n_n2322, n_n2806,
    n_n2337, n_n2345, n_n2359, n_n2746, n_n2294, n_n2304, n_n2313, n_n2360,
    n_n2286, n_n2293, n_n2305, n_n2312, n_n2361, n_n2749, n_n2296, n_n2303,
    n_n2311, n_n2287, n_n2295, n_n2770, n_n2310, n_n2288, n_n2298, n_n2307,
    n_n2789, n_n2327, n_n2335, n_n2289, n_n2297, n_n2308, n_n2316, n_n2802,
    n_n2334, n_n2290, n_n2300, n_n2774, n_n2315, n_n2343, n_n2353, n_n2291,
    n_n2299, n_n2306, n_n2314, n_n2344, n_n2352, n_n2292, n_n2302, n_n2323,
    n_n2332, n_n2341, n_n2834, n_n2838, n_n2757, n_n2301, n_n2324, n_n2331,
    n_n2342, n_n2351, n_n2354, n_n2779, n_n2318, n_n2325, n_n2333, n_n2340,
    n_n2350, n_n2355, n_n2309, n_n2317, n_n2326, n_n2811, n_n2821, n_n2349,
    n_n2356;
  wire new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_1_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_1_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_1_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_1_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_1_, new_n1158_,
    new_n1159_, new_n1161_, new_n1162_1_, new_n1163_, new_n1164_,
    new_n1165_, new_n1167_1_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_1_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_1_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_1_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_1_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_1_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_1_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_1_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_1_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_1_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_1_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_1_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_1_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_1_,
    new_n1243_, new_n1245_, new_n1246_, new_n1247_1_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_1_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_1_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_1_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_1_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_1_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_1_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_1_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_1_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_1_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_1_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_1_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_1_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_1_, new_n1318_, new_n1319_, new_n1321_,
    new_n1322_1_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_1_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_1_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_1_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_1_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_1_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_1_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_1_, new_n1359_, new_n1360_, new_n1361_, new_n1362_1_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_1_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_1_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_1_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_1_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_1_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_1_,
    new_n1393_, new_n1394_, new_n1395_, new_n1397_1_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_1_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_1_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_1_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_1_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_1_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_1_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_1_, new_n1433_,
    new_n1435_, new_n1436_, new_n1437_1_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_1_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_1_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_1_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_1_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_1_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_1_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_1_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_1_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_1_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_1_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_1_, new_n1498_, new_n1499_, new_n1500_, new_n1501_,
    new_n1502_1_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_1_, new_n1508_, new_n1509_, new_n1511_, new_n1512_1_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_1_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_1_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_1_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_1_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_1_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_1_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_1_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_1_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_1_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_1_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_1_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_1_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_1_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_1_, new_n1583_,
    new_n1584_, new_n1585_, new_n1587_1_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_1_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_1_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_1_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_1_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_1_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_1_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_1_, new_n1623_, new_n1625_,
    new_n1626_, new_n1627_1_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_1_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_1_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_1_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_1_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_1_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_1_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_1_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_1_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_1_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_1_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_1_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_1_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_1_, new_n1698_, new_n1699_, new_n1701_, new_n1702_1_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_1_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_1_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_1_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_1_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_1_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_1_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_1_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_1_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_1_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_1_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_1_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_1_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_1_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_1_, new_n1773_,
    new_n1774_, new_n1775_, new_n1777_1_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_1_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_1_, new_n1788_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_1_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_1_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_1_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_1_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_1_, new_n1813_, new_n1815_,
    new_n1816_, new_n1817_1_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_1_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_1_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_1_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_1_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_1_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_1_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_1_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_1_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_1_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_1_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_1_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_1_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_1_, new_n1888_, new_n1889_, new_n1891_, new_n1892_1_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_1_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_1_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_1_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_1_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_1_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_1_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_1_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_1_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_1_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_1_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_1_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_1_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_1_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_1_, new_n1963_,
    new_n1964_, new_n1965_, new_n1967_1_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_1_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_1_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_1_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_1_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_1_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_1_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_1_, new_n2003_, new_n2005_,
    new_n2006_, new_n2007_1_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_1_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_1_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_1_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_1_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_1_, new_n2033_, new_n2034_, new_n2035_,
    new_n2036_, new_n2037_1_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_,
    new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_,
    new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_,
    new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_,
    new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_,
    new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_,
    new_n2078_, new_n2079_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3113_, new_n3114_,
    new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_,
    new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_,
    new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_,
    new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_,
    new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_,
    new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_,
    new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3265_, new_n3266_, new_n3267_, new_n3268_,
    new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_,
    new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3549_, new_n3550_, new_n3551_, new_n3552_,
    new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_,
    new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_,
    new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_,
    new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_,
    new_n3577_, new_n3578_, new_n3579_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_,
    new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_,
    new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_,
    new_n3731_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3921_, new_n3922_,
    new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_,
    new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_,
    new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_,
    new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_,
    new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_,
    new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4073_, new_n4074_, new_n4075_, new_n4076_,
    new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_,
    new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_,
    new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_,
    new_n4107_, new_n4108_, new_n4109_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4149_, new_n4150_,
    new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4301_, new_n4302_, new_n4303_, new_n4304_,
    new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_,
    new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_,
    new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_,
    new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_,
    new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_,
    new_n4335_, new_n4336_, new_n4337_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_,
    new_n4483_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4599_, new_n4600_,
    new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_,
    new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_,
    new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_,
    new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_,
    new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_,
    new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4733_, new_n4734_, new_n4735_, new_n4736_,
    new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_,
    new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_,
    new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_,
    new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_,
    new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_,
    new_n4767_, new_n4768_, new_n4769_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_,
    new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_,
    new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_,
    new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_,
    new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_,
    new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_,
    new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_,
    new_n4989_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_,
    new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_,
    new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_,
    new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_,
    new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_,
    new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_,
    new_n5199_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_,
    new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_,
    new_n5415_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_,
    new_n5489_, new_n5490_, new_n5491_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_,
    new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_,
    new_n5643_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5683_, new_n5684_, new_n5685_, new_n5686_,
    new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_,
    new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_,
    new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_,
    new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_,
    new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_,
    new_n5717_, new_n5718_, new_n5719_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_,
    new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_,
    new_n5939_, new_n5940_, new_n5941_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5981_, new_n5982_,
    new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_,
    new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_,
    new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_,
    new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_,
    new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_,
    new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_,
    new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6127_, new_n6128_, new_n6129_, new_n6130_,
    new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_,
    new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_,
    new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_,
    new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_,
    new_n6155_, new_n6156_, new_n6157_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_,
    new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_,
    new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_,
    new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_,
    new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_,
    new_n6285_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_,
    new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_,
    new_n6316_, new_n6317_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_,
    new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_,
    new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_,
    new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_,
    new_n6347_, new_n6348_, new_n6349_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6383_, new_n6384_,
    new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_,
    new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_,
    new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_,
    new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_,
    new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_,
    new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_,
    new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_,
    new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_,
    new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_,
    new_n6477_, new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_,
    new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6511_, new_n6512_, new_n6513_, new_n6514_,
    new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_,
    new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_,
    new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_,
    new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_,
    new_n6539_, new_n6540_, new_n6541_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6575_, new_n6576_,
    new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_,
    new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_,
    new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_,
    new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_,
    new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_,
    new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6703_, new_n6704_, new_n6705_, new_n6706_,
    new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_,
    new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_,
    new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_,
    new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_,
    new_n6731_, new_n6732_, new_n6733_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6767_, new_n6768_,
    new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_,
    new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_,
    new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_,
    new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_,
    new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_,
    new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_,
    new_n6892_, new_n6893_, new_n6895_, new_n6896_, new_n6897_, new_n6898_,
    new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_,
    new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_,
    new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_,
    new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_,
    new_n6923_, new_n6924_, new_n6925_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_,
    new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_,
    new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7151_, new_n7152_,
    new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_,
    new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_,
    new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_,
    new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_,
    new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7279_, new_n7280_, new_n7281_, new_n7282_,
    new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_,
    new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_,
    new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_,
    new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_,
    new_n7307_, new_n7308_, new_n7309_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7343_, new_n7344_,
    new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_,
    new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7471_, new_n7472_, new_n7473_, new_n7474_,
    new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_,
    new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_,
    new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_,
    new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_,
    new_n7499_, new_n7500_, new_n7501_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_,
    new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_,
    new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7535_, new_n7536_,
    new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_,
    new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_,
    new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_,
    new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7727_, new_n7728_,
    new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_,
    new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_,
    new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_,
    new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_,
    new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7919_, new_n7920_,
    new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_,
    new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_,
    new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_,
    new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_,
    new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_,
    new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_,
    new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_,
    new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_,
    new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_,
    new_n8013_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8111_, new_n8112_,
    new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_,
    new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_,
    new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_,
    new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_,
    new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_,
    new_n8205_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_,
    new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_,
    new_n8236_, new_n8237_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8303_, new_n8304_,
    new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_,
    new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_,
    new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_,
    new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_,
    new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_,
    new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_,
    new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_,
    new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_,
    new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_,
    new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_,
    new_n8397_, new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_,
    new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_,
    new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_,
    new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_,
    new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_,
    new_n8428_, new_n8429_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_,
    new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_,
    new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_,
    new_n8459_, new_n8460_, new_n8461_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_,
    new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_,
    new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_,
    new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_,
    new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_,
    new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_,
    new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_,
    new_n8589_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_,
    new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_,
    new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_,
    new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_,
    new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_,
    new_n8781_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8815_, new_n8816_, new_n8817_, new_n8818_,
    new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_,
    new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_,
    new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_,
    new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_,
    new_n8843_, new_n8844_, new_n8845_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_,
    new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_,
    new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_,
    new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_,
    new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_,
    new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_,
    new_n8973_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9007_, new_n9008_, new_n9009_, new_n9010_,
    new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_,
    new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_,
    new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_,
    new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_,
    new_n9035_, new_n9036_, new_n9037_, n922, n927, n932, n937, n942, n947,
    n952, n957, n962, n967, n972, n977, n982, n987, n992, n997, n1002,
    n1007, n1012, n1017, n1022, n1027, n1032, n1037, n1042, n1047, n1052,
    n1057, n1062, n1067, n1072, n1077, n1082, n1087, n1092, n1097, n1102,
    n1107, n1112, n1117, n1122, n1127, n1132, n1137, n1142, n1147, n1152,
    n1157, n1162, n1167, n1172, n1177, n1182, n1187, n1192, n1197, n1202,
    n1207, n1212, n1217, n1222, n1227, n1232, n1237, n1242, n1247, n1252,
    n1257, n1262, n1267, n1272, n1277, n1282, n1287, n1292, n1297, n1302,
    n1307, n1312, n1317, n1322, n1327, n1332, n1337, n1342, n1347, n1352,
    n1357, n1362, n1367, n1372, n1377, n1382, n1387, n1392, n1397, n1402,
    n1407, n1412, n1417, n1422, n1427, n1432, n1437, n1442, n1447, n1452,
    n1457, n1462, n1467, n1472, n1477, n1482, n1487, n1492, n1497, n1502,
    n1507, n1512, n1517, n1522, n1527, n1532, n1537, n1542, n1547, n1552,
    n1557, n1562, n1567, n1572, n1577, n1582, n1587, n1592, n1597, n1602,
    n1607, n1612, n1617, n1622, n1627, n1632, n1637, n1642, n1647, n1652,
    n1657, n1662, n1667, n1672, n1677, n1682, n1687, n1692, n1697, n1702,
    n1707, n1712, n1717, n1722, n1727, n1732, n1737, n1742, n1747, n1752,
    n1757, n1762, n1767, n1772, n1777, n1782, n1787, n1792, n1797, n1802,
    n1807, n1812, n1817, n1822, n1827, n1832, n1837, n1842, n1847, n1852,
    n1857, n1862, n1867, n1872, n1877, n1882, n1887, n1892, n1897, n1902,
    n1907, n1912, n1917, n1922, n1927, n1932, n1937, n1942, n1947, n1952,
    n1957, n1962, n1967, n1972, n1977, n1982, n1987, n1992, n1997, n2002,
    n2007, n2012, n2017, n2022, n2027, n2032, n2037;
  assign new_n1133_ = ~pcount_2_ & ~pcount_1_;
  assign new_n1134_ = ~pencrypt_0_ & new_n1133_;
  assign new_n1135_ = ~pcount_0_ & new_n1134_;
  assign new_n1136_ = ~pstart_0_ & new_n1135_;
  assign new_n1137_1_ = ~pcount_3_ & new_n1136_;
  assign new_n1138_ = pcount_2_ & pcount_1_;
  assign new_n1139_ = pencrypt_0_ & new_n1138_;
  assign new_n1140_ = pcount_0_ & new_n1139_;
  assign new_n1141_ = ~pstart_0_ & new_n1140_;
  assign new_n1142_1_ = pcount_3_ & new_n1141_;
  assign pdata_ready_0_ = new_n1137_1_ | new_n1142_1_;
  assign new_n1144_ = ~pcount_1_ & ~pcount_0_;
  assign new_n1145_ = ~pcount_2_ & new_n1144_;
  assign new_n1146_ = ~pcount_3_ & new_n1145_;
  assign new_n1147_1_ = pcount_3_ & ~new_n1145_;
  assign new_n1148_ = ~new_n1146_ & ~new_n1147_1_;
  assign new_n1149_ = ~pencrypt_0_ & ~new_n1148_;
  assign new_n1150_ = ~pstart_0_ & new_n1149_;
  assign new_n1151_ = pcount_1_ & pcount_0_;
  assign new_n1152_1_ = pcount_2_ & new_n1151_;
  assign new_n1153_ = pcount_3_ & ~new_n1152_1_;
  assign new_n1154_ = ~pcount_3_ & new_n1152_1_;
  assign new_n1155_ = ~new_n1153_ & ~new_n1154_;
  assign new_n1156_ = pencrypt_0_ & ~new_n1155_;
  assign new_n1157_1_ = ~pstart_0_ & new_n1156_;
  assign new_n1158_ = pstart_0_ & ~pencrypt_0_;
  assign new_n1159_ = ~new_n1150_ & ~new_n1157_1_;
  assign pnew_count_3_ = new_n1158_ | ~new_n1159_;
  assign new_n1161_ = ~pcount_0_ & ~pencrypt_0_;
  assign new_n1162_1_ = ~pstart_0_ & new_n1161_;
  assign new_n1163_ = ~pcount_0_ & pencrypt_0_;
  assign new_n1164_ = ~pstart_0_ & new_n1163_;
  assign new_n1165_ = ~new_n1162_1_ & ~new_n1164_;
  assign pnew_count_0_ = new_n1158_ | ~new_n1165_;
  assign new_n1167_1_ = pcount_2_ & ~new_n1144_;
  assign new_n1168_ = ~new_n1145_ & ~new_n1167_1_;
  assign new_n1169_ = ~pencrypt_0_ & ~new_n1168_;
  assign new_n1170_ = ~pstart_0_ & new_n1169_;
  assign new_n1171_ = pcount_2_ & ~new_n1151_;
  assign new_n1172_1_ = ~pcount_2_ & new_n1151_;
  assign new_n1173_ = ~new_n1171_ & ~new_n1172_1_;
  assign new_n1174_ = pencrypt_0_ & ~new_n1173_;
  assign new_n1175_ = ~pstart_0_ & new_n1174_;
  assign new_n1176_ = ~new_n1170_ & ~new_n1175_;
  assign pnew_count_2_ = new_n1158_ | ~new_n1176_;
  assign new_n1178_ = ~new_n1144_ & ~new_n1151_;
  assign new_n1179_ = ~pencrypt_0_ & ~new_n1178_;
  assign new_n1180_ = ~pstart_0_ & new_n1179_;
  assign new_n1181_ = pcount_1_ & ~pcount_0_;
  assign new_n1182_1_ = ~pcount_1_ & pcount_0_;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_1_;
  assign new_n1184_ = pencrypt_0_ & ~new_n1183_;
  assign new_n1185_ = ~pstart_0_ & new_n1184_;
  assign new_n1186_ = ~new_n1180_ & ~new_n1185_;
  assign pnew_count_1_ = new_n1158_ | ~new_n1186_;
  assign new_n1188_ = ~pcount_3_ & ~pcount_1_;
  assign new_n1189_ = ~pcount_2_ & new_n1188_;
  assign new_n1190_ = ~pcount_0_ & new_n1189_;
  assign new_n1191_ = pcount_3_ & ~pcount_1_;
  assign new_n1192_1_ = ~pcount_2_ & new_n1191_;
  assign new_n1193_ = ~pcount_0_ & new_n1192_1_;
  assign new_n1194_ = pcount_0_ & new_n1189_;
  assign new_n1195_ = pcount_3_ & pcount_1_;
  assign new_n1196_ = pcount_2_ & new_n1195_;
  assign new_n1197_1_ = pcount_0_ & new_n1196_;
  assign new_n1198_ = ~new_n1190_ & ~new_n1193_;
  assign new_n1199_ = ~new_n1194_ & ~new_n1197_1_;
  assign new_n1200_ = new_n1198_ & new_n1199_;
  assign new_n1201_ = ~pencrypt_0_ & n_n2459;
  assign new_n1202_1_ = new_n1200_ & new_n1201_;
  assign new_n1203_ = ~pstart_0_ & new_n1202_1_;
  assign new_n1204_ = n_n2365 & n_n2459;
  assign new_n1205_ = ~pencrypt_0_ & new_n1204_;
  assign new_n1206_ = ~new_n1200_ & new_n1205_;
  assign new_n1207_1_ = ~pstart_0_ & new_n1206_;
  assign new_n1208_ = pkey_57_ & pencrypt_0_;
  assign new_n1209_ = pstart_0_ & new_n1208_;
  assign new_n1210_ = ~pencrypt_0_ & n_n2365;
  assign new_n1211_ = new_n1200_ & new_n1210_;
  assign new_n1212_1_ = ~pstart_0_ & new_n1211_;
  assign new_n1213_ = pkey_0_ & ~pencrypt_0_;
  assign new_n1214_ = pstart_0_ & new_n1213_;
  assign new_n1215_ = ~pcount_3_ & pcount_1_;
  assign new_n1216_ = pcount_2_ & new_n1215_;
  assign new_n1217_1_ = pcount_0_ & new_n1216_;
  assign new_n1218_ = ~pcount_0_ & new_n1196_;
  assign new_n1219_ = ~new_n1190_ & ~new_n1217_1_;
  assign new_n1220_ = ~new_n1218_ & new_n1219_;
  assign new_n1221_ = n_n2459 & new_n1220_;
  assign new_n1222_1_ = pencrypt_0_ & new_n1221_;
  assign new_n1223_ = ~n_n2365 & new_n1222_1_;
  assign new_n1224_ = ~pstart_0_ & new_n1223_;
  assign new_n1225_ = ~n_n2459 & new_n1220_;
  assign new_n1226_ = pencrypt_0_ & new_n1225_;
  assign new_n1227_1_ = n_n2365 & new_n1226_;
  assign new_n1228_ = ~pstart_0_ & new_n1227_1_;
  assign new_n1229_ = ~n_n2365 & ~n_n2459;
  assign new_n1230_ = ~pencrypt_0_ & new_n1229_;
  assign new_n1231_ = ~new_n1200_ & new_n1230_;
  assign new_n1232_1_ = ~pstart_0_ & new_n1231_;
  assign new_n1233_ = n_n2459 & ~new_n1220_;
  assign new_n1234_ = pencrypt_0_ & new_n1233_;
  assign new_n1235_ = n_n2365 & new_n1234_;
  assign new_n1236_ = ~pstart_0_ & new_n1235_;
  assign new_n1237_1_ = ~new_n1232_1_ & ~new_n1236_;
  assign new_n1238_ = ~new_n1224_ & ~new_n1228_;
  assign new_n1239_ = new_n1237_1_ & new_n1238_;
  assign new_n1240_ = ~new_n1212_1_ & ~new_n1214_;
  assign new_n1241_ = ~new_n1203_ & ~new_n1207_1_;
  assign new_n1242_1_ = ~new_n1209_ & new_n1241_;
  assign new_n1243_ = new_n1240_ & new_n1242_1_;
  assign n922 = ~new_n1239_ | ~new_n1243_;
  assign new_n1245_ = ~pencrypt_0_ & n_n2737;
  assign new_n1246_ = ~new_n1200_ & new_n1245_;
  assign new_n1247_1_ = ~pstart_0_ & new_n1246_;
  assign new_n1248_ = n_n2375 & n_n2737;
  assign new_n1249_ = ~pencrypt_0_ & new_n1248_;
  assign new_n1250_ = new_n1200_ & new_n1249_;
  assign new_n1251_ = ~pstart_0_ & new_n1250_;
  assign new_n1252_1_ = pkey_211_ & pencrypt_0_;
  assign new_n1253_ = pstart_0_ & new_n1252_1_;
  assign new_n1254_ = ~pencrypt_0_ & n_n2375;
  assign new_n1255_ = ~new_n1200_ & new_n1254_;
  assign new_n1256_ = ~pstart_0_ & new_n1255_;
  assign new_n1257_1_ = pkey_219_ & ~pencrypt_0_;
  assign new_n1258_ = pstart_0_ & new_n1257_1_;
  assign new_n1259_ = ~n_n2737 & ~new_n1220_;
  assign new_n1260_ = pencrypt_0_ & new_n1259_;
  assign new_n1261_ = n_n2375 & new_n1260_;
  assign new_n1262_1_ = ~pstart_0_ & new_n1261_;
  assign new_n1263_ = n_n2737 & new_n1220_;
  assign new_n1264_ = pencrypt_0_ & new_n1263_;
  assign new_n1265_ = n_n2375 & new_n1264_;
  assign new_n1266_ = ~pstart_0_ & new_n1265_;
  assign new_n1267_1_ = ~n_n2375 & ~n_n2737;
  assign new_n1268_ = ~pencrypt_0_ & new_n1267_1_;
  assign new_n1269_ = new_n1200_ & new_n1268_;
  assign new_n1270_ = ~pstart_0_ & new_n1269_;
  assign new_n1271_ = n_n2737 & ~new_n1220_;
  assign new_n1272_1_ = pencrypt_0_ & new_n1271_;
  assign new_n1273_ = ~n_n2375 & new_n1272_1_;
  assign new_n1274_ = ~pstart_0_ & new_n1273_;
  assign new_n1275_ = ~new_n1270_ & ~new_n1274_;
  assign new_n1276_ = ~new_n1262_1_ & ~new_n1266_;
  assign new_n1277_1_ = new_n1275_ & new_n1276_;
  assign new_n1278_ = ~new_n1256_ & ~new_n1258_;
  assign new_n1279_ = ~new_n1247_1_ & ~new_n1251_;
  assign new_n1280_ = ~new_n1253_ & new_n1279_;
  assign new_n1281_ = new_n1278_ & new_n1280_;
  assign n927 = ~new_n1277_1_ | ~new_n1281_;
  assign new_n1283_ = ~pencrypt_0_ & n_n2288;
  assign new_n1284_ = ~new_n1200_ & new_n1283_;
  assign new_n1285_ = ~pstart_0_ & new_n1284_;
  assign new_n1286_ = n_n2879 & n_n2288;
  assign new_n1287_1_ = ~pencrypt_0_ & new_n1286_;
  assign new_n1288_ = new_n1200_ & new_n1287_1_;
  assign new_n1289_ = ~pstart_0_ & new_n1288_;
  assign new_n1290_ = pencrypt_0_ & pkey_205_;
  assign new_n1291_ = pstart_0_ & new_n1290_;
  assign new_n1292_1_ = ~pencrypt_0_ & n_n2879;
  assign new_n1293_ = ~new_n1200_ & new_n1292_1_;
  assign new_n1294_ = ~pstart_0_ & new_n1293_;
  assign new_n1295_ = pkey_213_ & ~pencrypt_0_;
  assign new_n1296_ = pstart_0_ & new_n1295_;
  assign new_n1297_1_ = ~n_n2288 & ~new_n1220_;
  assign new_n1298_ = pencrypt_0_ & new_n1297_1_;
  assign new_n1299_ = n_n2879 & new_n1298_;
  assign new_n1300_ = ~pstart_0_ & new_n1299_;
  assign new_n1301_ = n_n2288 & new_n1220_;
  assign new_n1302_1_ = pencrypt_0_ & new_n1301_;
  assign new_n1303_ = n_n2879 & new_n1302_1_;
  assign new_n1304_ = ~pstart_0_ & new_n1303_;
  assign new_n1305_ = ~n_n2879 & ~n_n2288;
  assign new_n1306_ = ~pencrypt_0_ & new_n1305_;
  assign new_n1307_1_ = new_n1200_ & new_n1306_;
  assign new_n1308_ = ~pstart_0_ & new_n1307_1_;
  assign new_n1309_ = n_n2288 & ~new_n1220_;
  assign new_n1310_ = pencrypt_0_ & new_n1309_;
  assign new_n1311_ = ~n_n2879 & new_n1310_;
  assign new_n1312_1_ = ~pstart_0_ & new_n1311_;
  assign new_n1313_ = ~new_n1308_ & ~new_n1312_1_;
  assign new_n1314_ = ~new_n1300_ & ~new_n1304_;
  assign new_n1315_ = new_n1313_ & new_n1314_;
  assign new_n1316_ = ~new_n1294_ & ~new_n1296_;
  assign new_n1317_1_ = ~new_n1285_ & ~new_n1289_;
  assign new_n1318_ = ~new_n1291_ & new_n1317_1_;
  assign new_n1319_ = new_n1316_ & new_n1318_;
  assign n932 = ~new_n1315_ | ~new_n1319_;
  assign new_n1321_ = ~pencrypt_0_ & n_n2298;
  assign new_n1322_1_ = ~new_n1200_ & new_n1321_;
  assign new_n1323_ = ~pstart_0_ & new_n1322_1_;
  assign new_n1324_ = n_n2392 & n_n2298;
  assign new_n1325_ = ~pencrypt_0_ & new_n1324_;
  assign new_n1326_ = new_n1200_ & new_n1325_;
  assign new_n1327_1_ = ~pstart_0_ & new_n1326_;
  assign new_n1328_ = pkey_230_ & pencrypt_0_;
  assign new_n1329_ = pstart_0_ & new_n1328_;
  assign new_n1330_ = ~pencrypt_0_ & n_n2392;
  assign new_n1331_ = ~new_n1200_ & new_n1330_;
  assign new_n1332_1_ = ~pstart_0_ & new_n1331_;
  assign new_n1333_ = pkey_238_ & ~pencrypt_0_;
  assign new_n1334_ = pstart_0_ & new_n1333_;
  assign new_n1335_ = ~n_n2298 & ~new_n1220_;
  assign new_n1336_ = pencrypt_0_ & new_n1335_;
  assign new_n1337_1_ = n_n2392 & new_n1336_;
  assign new_n1338_ = ~pstart_0_ & new_n1337_1_;
  assign new_n1339_ = n_n2298 & new_n1220_;
  assign new_n1340_ = pencrypt_0_ & new_n1339_;
  assign new_n1341_ = n_n2392 & new_n1340_;
  assign new_n1342_1_ = ~pstart_0_ & new_n1341_;
  assign new_n1343_ = ~n_n2392 & ~n_n2298;
  assign new_n1344_ = ~pencrypt_0_ & new_n1343_;
  assign new_n1345_ = new_n1200_ & new_n1344_;
  assign new_n1346_ = ~pstart_0_ & new_n1345_;
  assign new_n1347_1_ = n_n2298 & ~new_n1220_;
  assign new_n1348_ = pencrypt_0_ & new_n1347_1_;
  assign new_n1349_ = ~n_n2392 & new_n1348_;
  assign new_n1350_ = ~pstart_0_ & new_n1349_;
  assign new_n1351_ = ~new_n1346_ & ~new_n1350_;
  assign new_n1352_1_ = ~new_n1338_ & ~new_n1342_1_;
  assign new_n1353_ = new_n1351_ & new_n1352_1_;
  assign new_n1354_ = ~new_n1332_1_ & ~new_n1334_;
  assign new_n1355_ = ~new_n1323_ & ~new_n1327_1_;
  assign new_n1356_ = ~new_n1329_ & new_n1355_;
  assign new_n1357_1_ = new_n1354_ & new_n1356_;
  assign n937 = ~new_n1353_ | ~new_n1357_1_;
  assign new_n1359_ = ~pencrypt_0_ & n_n2307;
  assign new_n1360_ = ~new_n1200_ & new_n1359_;
  assign new_n1361_ = ~pstart_0_ & new_n1360_;
  assign new_n1362_1_ = n_n2402 & n_n2307;
  assign new_n1363_ = ~pencrypt_0_ & new_n1362_1_;
  assign new_n1364_ = new_n1200_ & new_n1363_;
  assign new_n1365_ = ~pstart_0_ & new_n1364_;
  assign new_n1366_ = pkey_156_ & pencrypt_0_;
  assign new_n1367_1_ = pstart_0_ & new_n1366_;
  assign new_n1368_ = ~pencrypt_0_ & n_n2402;
  assign new_n1369_ = ~new_n1200_ & new_n1368_;
  assign new_n1370_ = ~pstart_0_ & new_n1369_;
  assign new_n1371_ = pkey_164_ & ~pencrypt_0_;
  assign new_n1372_1_ = pstart_0_ & new_n1371_;
  assign new_n1373_ = ~n_n2307 & ~new_n1220_;
  assign new_n1374_ = pencrypt_0_ & new_n1373_;
  assign new_n1375_ = n_n2402 & new_n1374_;
  assign new_n1376_ = ~pstart_0_ & new_n1375_;
  assign new_n1377_1_ = n_n2307 & new_n1220_;
  assign new_n1378_ = pencrypt_0_ & new_n1377_1_;
  assign new_n1379_ = n_n2402 & new_n1378_;
  assign new_n1380_ = ~pstart_0_ & new_n1379_;
  assign new_n1381_ = ~n_n2402 & ~n_n2307;
  assign new_n1382_1_ = ~pencrypt_0_ & new_n1381_;
  assign new_n1383_ = new_n1200_ & new_n1382_1_;
  assign new_n1384_ = ~pstart_0_ & new_n1383_;
  assign new_n1385_ = n_n2307 & ~new_n1220_;
  assign new_n1386_ = pencrypt_0_ & new_n1385_;
  assign new_n1387_1_ = ~n_n2402 & new_n1386_;
  assign new_n1388_ = ~pstart_0_ & new_n1387_1_;
  assign new_n1389_ = ~new_n1384_ & ~new_n1388_;
  assign new_n1390_ = ~new_n1376_ & ~new_n1380_;
  assign new_n1391_ = new_n1389_ & new_n1390_;
  assign new_n1392_1_ = ~new_n1370_ & ~new_n1372_1_;
  assign new_n1393_ = ~new_n1361_ & ~new_n1365_;
  assign new_n1394_ = ~new_n1367_1_ & new_n1393_;
  assign new_n1395_ = new_n1392_1_ & new_n1394_;
  assign n942 = ~new_n1391_ | ~new_n1395_;
  assign new_n1397_1_ = ~pencrypt_0_ & n_n2789;
  assign new_n1398_ = ~new_n1200_ & new_n1397_1_;
  assign new_n1399_ = ~pstart_0_ & new_n1398_;
  assign new_n1400_ = n_n2411 & n_n2789;
  assign new_n1401_ = ~pencrypt_0_ & new_n1400_;
  assign new_n1402_1_ = new_n1200_ & new_n1401_;
  assign new_n1403_ = ~pstart_0_ & new_n1402_1_;
  assign new_n1404_ = pkey_181_ & pencrypt_0_;
  assign new_n1405_ = pstart_0_ & new_n1404_;
  assign new_n1406_ = ~pencrypt_0_ & n_n2411;
  assign new_n1407_1_ = ~new_n1200_ & new_n1406_;
  assign new_n1408_ = ~pstart_0_ & new_n1407_1_;
  assign new_n1409_ = ~pencrypt_0_ & pkey_189_;
  assign new_n1410_ = pstart_0_ & new_n1409_;
  assign new_n1411_ = ~n_n2789 & ~new_n1220_;
  assign new_n1412_1_ = pencrypt_0_ & new_n1411_;
  assign new_n1413_ = n_n2411 & new_n1412_1_;
  assign new_n1414_ = ~pstart_0_ & new_n1413_;
  assign new_n1415_ = n_n2789 & new_n1220_;
  assign new_n1416_ = pencrypt_0_ & new_n1415_;
  assign new_n1417_1_ = n_n2411 & new_n1416_;
  assign new_n1418_ = ~pstart_0_ & new_n1417_1_;
  assign new_n1419_ = ~n_n2411 & ~n_n2789;
  assign new_n1420_ = ~pencrypt_0_ & new_n1419_;
  assign new_n1421_ = new_n1200_ & new_n1420_;
  assign new_n1422_1_ = ~pstart_0_ & new_n1421_;
  assign new_n1423_ = n_n2789 & ~new_n1220_;
  assign new_n1424_ = pencrypt_0_ & new_n1423_;
  assign new_n1425_ = ~n_n2411 & new_n1424_;
  assign new_n1426_ = ~pstart_0_ & new_n1425_;
  assign new_n1427_1_ = ~new_n1422_1_ & ~new_n1426_;
  assign new_n1428_ = ~new_n1414_ & ~new_n1418_;
  assign new_n1429_ = new_n1427_1_ & new_n1428_;
  assign new_n1430_ = ~new_n1408_ & ~new_n1410_;
  assign new_n1431_ = ~new_n1399_ & ~new_n1403_;
  assign new_n1432_1_ = ~new_n1405_ & new_n1431_;
  assign new_n1433_ = new_n1430_ & new_n1432_1_;
  assign n947 = ~new_n1429_ | ~new_n1433_;
  assign new_n1435_ = ~pencrypt_0_ & n_n2354;
  assign new_n1436_ = ~new_n1200_ & new_n1435_;
  assign new_n1437_1_ = ~pstart_0_ & new_n1436_;
  assign new_n1438_ = n_n2448 & n_n2354;
  assign new_n1439_ = ~pencrypt_0_ & new_n1438_;
  assign new_n1440_ = new_n1200_ & new_n1439_;
  assign new_n1441_ = ~pstart_0_ & new_n1440_;
  assign new_n1442_1_ = pencrypt_0_ & pkey_20_;
  assign new_n1443_ = pstart_0_ & new_n1442_1_;
  assign new_n1444_ = ~pencrypt_0_ & n_n2448;
  assign new_n1445_ = ~new_n1200_ & new_n1444_;
  assign new_n1446_ = ~pstart_0_ & new_n1445_;
  assign new_n1447_1_ = pkey_28_ & ~pencrypt_0_;
  assign new_n1448_ = pstart_0_ & new_n1447_1_;
  assign new_n1449_ = ~n_n2354 & ~new_n1220_;
  assign new_n1450_ = pencrypt_0_ & new_n1449_;
  assign new_n1451_ = n_n2448 & new_n1450_;
  assign new_n1452_1_ = ~pstart_0_ & new_n1451_;
  assign new_n1453_ = n_n2354 & new_n1220_;
  assign new_n1454_ = pencrypt_0_ & new_n1453_;
  assign new_n1455_ = n_n2448 & new_n1454_;
  assign new_n1456_ = ~pstart_0_ & new_n1455_;
  assign new_n1457_1_ = ~n_n2448 & ~n_n2354;
  assign new_n1458_ = ~pencrypt_0_ & new_n1457_1_;
  assign new_n1459_ = new_n1200_ & new_n1458_;
  assign new_n1460_ = ~pstart_0_ & new_n1459_;
  assign new_n1461_ = n_n2354 & ~new_n1220_;
  assign new_n1462_1_ = pencrypt_0_ & new_n1461_;
  assign new_n1463_ = ~n_n2448 & new_n1462_1_;
  assign new_n1464_ = ~pstart_0_ & new_n1463_;
  assign new_n1465_ = ~new_n1460_ & ~new_n1464_;
  assign new_n1466_ = ~new_n1452_1_ & ~new_n1456_;
  assign new_n1467_1_ = new_n1465_ & new_n1466_;
  assign new_n1468_ = ~new_n1446_ & ~new_n1448_;
  assign new_n1469_ = ~new_n1437_1_ & ~new_n1441_;
  assign new_n1470_ = ~new_n1443_ & new_n1469_;
  assign new_n1471_ = new_n1468_ & new_n1470_;
  assign n952 = ~new_n1467_1_ | ~new_n1471_;
  assign new_n1473_ = ~pencrypt_0_ & n_n2364;
  assign new_n1474_ = ~new_n1200_ & new_n1473_;
  assign new_n1475_ = ~pstart_0_ & new_n1474_;
  assign new_n1476_ = n_n2982 & n_n2364;
  assign new_n1477_1_ = ~pencrypt_0_ & new_n1476_;
  assign new_n1478_ = new_n1200_ & new_n1477_1_;
  assign new_n1479_ = ~pstart_0_ & new_n1478_;
  assign new_n1480_ = pencrypt_0_ & pkey_45_;
  assign new_n1481_ = pstart_0_ & new_n1480_;
  assign new_n1482_1_ = ~pencrypt_0_ & n_n2982;
  assign new_n1483_ = ~new_n1200_ & new_n1482_1_;
  assign new_n1484_ = ~pstart_0_ & new_n1483_;
  assign new_n1485_ = ~pencrypt_0_ & pkey_53_;
  assign new_n1486_ = pstart_0_ & new_n1485_;
  assign new_n1487_1_ = ~n_n2364 & ~new_n1220_;
  assign new_n1488_ = pencrypt_0_ & new_n1487_1_;
  assign new_n1489_ = n_n2982 & new_n1488_;
  assign new_n1490_ = ~pstart_0_ & new_n1489_;
  assign new_n1491_ = n_n2364 & new_n1220_;
  assign new_n1492_1_ = pencrypt_0_ & new_n1491_;
  assign new_n1493_ = n_n2982 & new_n1492_1_;
  assign new_n1494_ = ~pstart_0_ & new_n1493_;
  assign new_n1495_ = ~n_n2982 & ~n_n2364;
  assign new_n1496_ = ~pencrypt_0_ & new_n1495_;
  assign new_n1497_1_ = new_n1200_ & new_n1496_;
  assign new_n1498_ = ~pstart_0_ & new_n1497_1_;
  assign new_n1499_ = n_n2364 & ~new_n1220_;
  assign new_n1500_ = pencrypt_0_ & new_n1499_;
  assign new_n1501_ = ~n_n2982 & new_n1500_;
  assign new_n1502_1_ = ~pstart_0_ & new_n1501_;
  assign new_n1503_ = ~new_n1498_ & ~new_n1502_1_;
  assign new_n1504_ = ~new_n1490_ & ~new_n1494_;
  assign new_n1505_ = new_n1503_ & new_n1504_;
  assign new_n1506_ = ~new_n1484_ & ~new_n1486_;
  assign new_n1507_1_ = ~new_n1475_ & ~new_n1479_;
  assign new_n1508_ = ~new_n1481_ & new_n1507_1_;
  assign new_n1509_ = new_n1506_ & new_n1508_;
  assign n957 = ~new_n1505_ | ~new_n1509_;
  assign new_n1511_ = ~pencrypt_0_ & n_n2986;
  assign new_n1512_1_ = new_n1200_ & new_n1511_;
  assign new_n1513_ = ~pstart_0_ & new_n1512_1_;
  assign new_n1514_ = n_n2366 & n_n2986;
  assign new_n1515_ = ~pencrypt_0_ & new_n1514_;
  assign new_n1516_ = ~new_n1200_ & new_n1515_;
  assign new_n1517_1_ = ~pstart_0_ & new_n1516_;
  assign new_n1518_ = pkey_0_ & pencrypt_0_;
  assign new_n1519_ = pstart_0_ & new_n1518_;
  assign new_n1520_ = ~pencrypt_0_ & n_n2366;
  assign new_n1521_ = new_n1200_ & new_n1520_;
  assign new_n1522_1_ = ~pstart_0_ & new_n1521_;
  assign new_n1523_ = pkey_8_ & ~pencrypt_0_;
  assign new_n1524_ = pstart_0_ & new_n1523_;
  assign new_n1525_ = n_n2986 & new_n1220_;
  assign new_n1526_ = pencrypt_0_ & new_n1525_;
  assign new_n1527_1_ = ~n_n2366 & new_n1526_;
  assign new_n1528_ = ~pstart_0_ & new_n1527_1_;
  assign new_n1529_ = ~n_n2986 & new_n1220_;
  assign new_n1530_ = pencrypt_0_ & new_n1529_;
  assign new_n1531_ = n_n2366 & new_n1530_;
  assign new_n1532_1_ = ~pstart_0_ & new_n1531_;
  assign new_n1533_ = ~n_n2366 & ~n_n2986;
  assign new_n1534_ = ~pencrypt_0_ & new_n1533_;
  assign new_n1535_ = ~new_n1200_ & new_n1534_;
  assign new_n1536_ = ~pstart_0_ & new_n1535_;
  assign new_n1537_1_ = n_n2986 & ~new_n1220_;
  assign new_n1538_ = pencrypt_0_ & new_n1537_1_;
  assign new_n1539_ = n_n2366 & new_n1538_;
  assign new_n1540_ = ~pstart_0_ & new_n1539_;
  assign new_n1541_ = ~new_n1536_ & ~new_n1540_;
  assign new_n1542_1_ = ~new_n1528_ & ~new_n1532_1_;
  assign new_n1543_ = new_n1541_ & new_n1542_1_;
  assign new_n1544_ = ~new_n1522_1_ & ~new_n1524_;
  assign new_n1545_ = ~new_n1513_ & ~new_n1517_1_;
  assign new_n1546_ = ~new_n1519_ & new_n1545_;
  assign new_n1547_1_ = new_n1544_ & new_n1546_;
  assign n962 = ~new_n1543_ | ~new_n1547_1_;
  assign new_n1549_ = ~pencrypt_0_ & n_n2280;
  assign new_n1550_ = ~new_n1200_ & new_n1549_;
  assign new_n1551_ = ~pstart_0_ & new_n1550_;
  assign new_n1552_1_ = n_n2865 & n_n2280;
  assign new_n1553_ = ~pencrypt_0_ & new_n1552_1_;
  assign new_n1554_ = new_n1200_ & new_n1553_;
  assign new_n1555_ = ~pstart_0_ & new_n1554_;
  assign new_n1556_ = pkey_203_ & pencrypt_0_;
  assign new_n1557_1_ = pstart_0_ & new_n1556_;
  assign new_n1558_ = ~pencrypt_0_ & n_n2865;
  assign new_n1559_ = ~new_n1200_ & new_n1558_;
  assign new_n1560_ = ~pstart_0_ & new_n1559_;
  assign new_n1561_ = pkey_211_ & ~pencrypt_0_;
  assign new_n1562_1_ = pstart_0_ & new_n1561_;
  assign new_n1563_ = ~n_n2280 & ~new_n1220_;
  assign new_n1564_ = pencrypt_0_ & new_n1563_;
  assign new_n1565_ = n_n2865 & new_n1564_;
  assign new_n1566_ = ~pstart_0_ & new_n1565_;
  assign new_n1567_1_ = n_n2280 & new_n1220_;
  assign new_n1568_ = pencrypt_0_ & new_n1567_1_;
  assign new_n1569_ = n_n2865 & new_n1568_;
  assign new_n1570_ = ~pstart_0_ & new_n1569_;
  assign new_n1571_ = ~n_n2865 & ~n_n2280;
  assign new_n1572_1_ = ~pencrypt_0_ & new_n1571_;
  assign new_n1573_ = new_n1200_ & new_n1572_1_;
  assign new_n1574_ = ~pstart_0_ & new_n1573_;
  assign new_n1575_ = n_n2280 & ~new_n1220_;
  assign new_n1576_ = pencrypt_0_ & new_n1575_;
  assign new_n1577_1_ = ~n_n2865 & new_n1576_;
  assign new_n1578_ = ~pstart_0_ & new_n1577_1_;
  assign new_n1579_ = ~new_n1574_ & ~new_n1578_;
  assign new_n1580_ = ~new_n1566_ & ~new_n1570_;
  assign new_n1581_ = new_n1579_ & new_n1580_;
  assign new_n1582_1_ = ~new_n1560_ & ~new_n1562_1_;
  assign new_n1583_ = ~new_n1551_ & ~new_n1555_;
  assign new_n1584_ = ~new_n1557_1_ & new_n1583_;
  assign new_n1585_ = new_n1582_1_ & new_n1584_;
  assign n967 = ~new_n1581_ | ~new_n1585_;
  assign new_n1587_1_ = ~pencrypt_0_ & n_n2289;
  assign new_n1588_ = ~new_n1200_ & new_n1587_1_;
  assign new_n1589_ = ~pstart_0_ & new_n1588_;
  assign new_n1590_ = n_n2881 & n_n2289;
  assign new_n1591_ = ~pencrypt_0_ & new_n1590_;
  assign new_n1592_1_ = new_n1200_ & new_n1591_;
  assign new_n1593_ = ~pstart_0_ & new_n1592_1_;
  assign new_n1594_ = pkey_213_ & pencrypt_0_;
  assign new_n1595_ = pstart_0_ & new_n1594_;
  assign new_n1596_ = ~pencrypt_0_ & n_n2881;
  assign new_n1597_1_ = ~new_n1200_ & new_n1596_;
  assign new_n1598_ = ~pstart_0_ & new_n1597_1_;
  assign new_n1599_ = pkey_221_ & ~pencrypt_0_;
  assign new_n1600_ = pstart_0_ & new_n1599_;
  assign new_n1601_ = ~n_n2289 & ~new_n1220_;
  assign new_n1602_1_ = pencrypt_0_ & new_n1601_;
  assign new_n1603_ = n_n2881 & new_n1602_1_;
  assign new_n1604_ = ~pstart_0_ & new_n1603_;
  assign new_n1605_ = n_n2289 & new_n1220_;
  assign new_n1606_ = pencrypt_0_ & new_n1605_;
  assign new_n1607_1_ = n_n2881 & new_n1606_;
  assign new_n1608_ = ~pstart_0_ & new_n1607_1_;
  assign new_n1609_ = ~n_n2881 & ~n_n2289;
  assign new_n1610_ = ~pencrypt_0_ & new_n1609_;
  assign new_n1611_ = new_n1200_ & new_n1610_;
  assign new_n1612_1_ = ~pstart_0_ & new_n1611_;
  assign new_n1613_ = n_n2289 & ~new_n1220_;
  assign new_n1614_ = pencrypt_0_ & new_n1613_;
  assign new_n1615_ = ~n_n2881 & new_n1614_;
  assign new_n1616_ = ~pstart_0_ & new_n1615_;
  assign new_n1617_1_ = ~new_n1612_1_ & ~new_n1616_;
  assign new_n1618_ = ~new_n1604_ & ~new_n1608_;
  assign new_n1619_ = new_n1617_1_ & new_n1618_;
  assign new_n1620_ = ~new_n1598_ & ~new_n1600_;
  assign new_n1621_ = ~new_n1589_ & ~new_n1593_;
  assign new_n1622_1_ = ~new_n1595_ & new_n1621_;
  assign new_n1623_ = new_n1620_ & new_n1622_1_;
  assign n972 = ~new_n1619_ | ~new_n1623_;
  assign new_n1625_ = ~pencrypt_0_ & n_n2297;
  assign new_n1626_ = ~new_n1200_ & new_n1625_;
  assign new_n1627_1_ = ~pstart_0_ & new_n1626_;
  assign new_n1628_ = n_n2391 & n_n2297;
  assign new_n1629_ = ~pencrypt_0_ & new_n1628_;
  assign new_n1630_ = new_n1200_ & new_n1629_;
  assign new_n1631_ = ~pstart_0_ & new_n1630_;
  assign new_n1632_1_ = pkey_222_ & pencrypt_0_;
  assign new_n1633_ = pstart_0_ & new_n1632_1_;
  assign new_n1634_ = ~pencrypt_0_ & n_n2391;
  assign new_n1635_ = ~new_n1200_ & new_n1634_;
  assign new_n1636_ = ~pstart_0_ & new_n1635_;
  assign new_n1637_1_ = pkey_230_ & ~pencrypt_0_;
  assign new_n1638_ = pstart_0_ & new_n1637_1_;
  assign new_n1639_ = ~n_n2297 & ~new_n1220_;
  assign new_n1640_ = pencrypt_0_ & new_n1639_;
  assign new_n1641_ = n_n2391 & new_n1640_;
  assign new_n1642_1_ = ~pstart_0_ & new_n1641_;
  assign new_n1643_ = n_n2297 & new_n1220_;
  assign new_n1644_ = pencrypt_0_ & new_n1643_;
  assign new_n1645_ = n_n2391 & new_n1644_;
  assign new_n1646_ = ~pstart_0_ & new_n1645_;
  assign new_n1647_1_ = ~n_n2391 & ~n_n2297;
  assign new_n1648_ = ~pencrypt_0_ & new_n1647_1_;
  assign new_n1649_ = new_n1200_ & new_n1648_;
  assign new_n1650_ = ~pstart_0_ & new_n1649_;
  assign new_n1651_ = n_n2297 & ~new_n1220_;
  assign new_n1652_1_ = pencrypt_0_ & new_n1651_;
  assign new_n1653_ = ~n_n2391 & new_n1652_1_;
  assign new_n1654_ = ~pstart_0_ & new_n1653_;
  assign new_n1655_ = ~new_n1650_ & ~new_n1654_;
  assign new_n1656_ = ~new_n1642_1_ & ~new_n1646_;
  assign new_n1657_1_ = new_n1655_ & new_n1656_;
  assign new_n1658_ = ~new_n1636_ & ~new_n1638_;
  assign new_n1659_ = ~new_n1627_1_ & ~new_n1631_;
  assign new_n1660_ = ~new_n1633_ & new_n1659_;
  assign new_n1661_ = new_n1658_ & new_n1660_;
  assign n977 = ~new_n1657_1_ | ~new_n1661_;
  assign new_n1663_ = ~pencrypt_0_ & n_n2308;
  assign new_n1664_ = ~new_n1200_ & new_n1663_;
  assign new_n1665_ = ~pstart_0_ & new_n1664_;
  assign new_n1666_ = n_n2403 & n_n2308;
  assign new_n1667_1_ = ~pencrypt_0_ & new_n1666_;
  assign new_n1668_ = new_n1200_ & new_n1667_1_;
  assign new_n1669_ = ~pstart_0_ & new_n1668_;
  assign new_n1670_ = pkey_164_ & pencrypt_0_;
  assign new_n1671_ = pstart_0_ & new_n1670_;
  assign new_n1672_1_ = ~pencrypt_0_ & n_n2403;
  assign new_n1673_ = ~new_n1200_ & new_n1672_1_;
  assign new_n1674_ = ~pstart_0_ & new_n1673_;
  assign new_n1675_ = ~pencrypt_0_ & pkey_172_;
  assign new_n1676_ = pstart_0_ & new_n1675_;
  assign new_n1677_1_ = ~n_n2308 & ~new_n1220_;
  assign new_n1678_ = pencrypt_0_ & new_n1677_1_;
  assign new_n1679_ = n_n2403 & new_n1678_;
  assign new_n1680_ = ~pstart_0_ & new_n1679_;
  assign new_n1681_ = n_n2308 & new_n1220_;
  assign new_n1682_1_ = pencrypt_0_ & new_n1681_;
  assign new_n1683_ = n_n2403 & new_n1682_1_;
  assign new_n1684_ = ~pstart_0_ & new_n1683_;
  assign new_n1685_ = ~n_n2403 & ~n_n2308;
  assign new_n1686_ = ~pencrypt_0_ & new_n1685_;
  assign new_n1687_1_ = new_n1200_ & new_n1686_;
  assign new_n1688_ = ~pstart_0_ & new_n1687_1_;
  assign new_n1689_ = n_n2308 & ~new_n1220_;
  assign new_n1690_ = pencrypt_0_ & new_n1689_;
  assign new_n1691_ = ~n_n2403 & new_n1690_;
  assign new_n1692_1_ = ~pstart_0_ & new_n1691_;
  assign new_n1693_ = ~new_n1688_ & ~new_n1692_1_;
  assign new_n1694_ = ~new_n1680_ & ~new_n1684_;
  assign new_n1695_ = new_n1693_ & new_n1694_;
  assign new_n1696_ = ~new_n1674_ & ~new_n1676_;
  assign new_n1697_1_ = ~new_n1665_ & ~new_n1669_;
  assign new_n1698_ = ~new_n1671_ & new_n1697_1_;
  assign new_n1699_ = new_n1696_ & new_n1698_;
  assign n982 = ~new_n1695_ | ~new_n1699_;
  assign new_n1701_ = ~pencrypt_0_ & n_n2316;
  assign new_n1702_1_ = ~new_n1200_ & new_n1701_;
  assign new_n1703_ = ~pstart_0_ & new_n1702_1_;
  assign new_n1704_ = n_n2917 & n_n2316;
  assign new_n1705_ = ~pencrypt_0_ & new_n1704_;
  assign new_n1706_ = new_n1200_ & new_n1705_;
  assign new_n1707_1_ = ~pstart_0_ & new_n1706_;
  assign new_n1708_ = pencrypt_0_ & pkey_173_;
  assign new_n1709_ = pstart_0_ & new_n1708_;
  assign new_n1710_ = ~pencrypt_0_ & n_n2917;
  assign new_n1711_ = ~new_n1200_ & new_n1710_;
  assign new_n1712_1_ = ~pstart_0_ & new_n1711_;
  assign new_n1713_ = pkey_181_ & ~pencrypt_0_;
  assign new_n1714_ = pstart_0_ & new_n1713_;
  assign new_n1715_ = ~n_n2316 & ~new_n1220_;
  assign new_n1716_ = pencrypt_0_ & new_n1715_;
  assign new_n1717_1_ = n_n2917 & new_n1716_;
  assign new_n1718_ = ~pstart_0_ & new_n1717_1_;
  assign new_n1719_ = n_n2316 & new_n1220_;
  assign new_n1720_ = pencrypt_0_ & new_n1719_;
  assign new_n1721_ = n_n2917 & new_n1720_;
  assign new_n1722_1_ = ~pstart_0_ & new_n1721_;
  assign new_n1723_ = ~n_n2917 & ~n_n2316;
  assign new_n1724_ = ~pencrypt_0_ & new_n1723_;
  assign new_n1725_ = new_n1200_ & new_n1724_;
  assign new_n1726_ = ~pstart_0_ & new_n1725_;
  assign new_n1727_1_ = n_n2316 & ~new_n1220_;
  assign new_n1728_ = pencrypt_0_ & new_n1727_1_;
  assign new_n1729_ = ~n_n2917 & new_n1728_;
  assign new_n1730_ = ~pstart_0_ & new_n1729_;
  assign new_n1731_ = ~new_n1726_ & ~new_n1730_;
  assign new_n1732_1_ = ~new_n1718_ & ~new_n1722_1_;
  assign new_n1733_ = new_n1731_ & new_n1732_1_;
  assign new_n1734_ = ~new_n1712_1_ & ~new_n1714_;
  assign new_n1735_ = ~new_n1703_ & ~new_n1707_1_;
  assign new_n1736_ = ~new_n1709_ & new_n1735_;
  assign new_n1737_1_ = new_n1734_ & new_n1736_;
  assign n987 = ~new_n1733_ | ~new_n1737_1_;
  assign new_n1739_ = ~pencrypt_0_ & n_n2355;
  assign new_n1740_ = ~new_n1200_ & new_n1739_;
  assign new_n1741_ = ~pstart_0_ & new_n1740_;
  assign new_n1742_1_ = n_n2449 & n_n2355;
  assign new_n1743_ = ~pencrypt_0_ & new_n1742_1_;
  assign new_n1744_ = new_n1200_ & new_n1743_;
  assign new_n1745_ = ~pstart_0_ & new_n1744_;
  assign new_n1746_ = pkey_28_ & pencrypt_0_;
  assign new_n1747_1_ = pstart_0_ & new_n1746_;
  assign new_n1748_ = ~pencrypt_0_ & n_n2449;
  assign new_n1749_ = ~new_n1200_ & new_n1748_;
  assign new_n1750_ = ~pstart_0_ & new_n1749_;
  assign new_n1751_ = pkey_36_ & ~pencrypt_0_;
  assign new_n1752_1_ = pstart_0_ & new_n1751_;
  assign new_n1753_ = ~n_n2355 & ~new_n1220_;
  assign new_n1754_ = pencrypt_0_ & new_n1753_;
  assign new_n1755_ = n_n2449 & new_n1754_;
  assign new_n1756_ = ~pstart_0_ & new_n1755_;
  assign new_n1757_1_ = n_n2355 & new_n1220_;
  assign new_n1758_ = pencrypt_0_ & new_n1757_1_;
  assign new_n1759_ = n_n2449 & new_n1758_;
  assign new_n1760_ = ~pstart_0_ & new_n1759_;
  assign new_n1761_ = ~n_n2449 & ~n_n2355;
  assign new_n1762_1_ = ~pencrypt_0_ & new_n1761_;
  assign new_n1763_ = new_n1200_ & new_n1762_1_;
  assign new_n1764_ = ~pstart_0_ & new_n1763_;
  assign new_n1765_ = n_n2355 & ~new_n1220_;
  assign new_n1766_ = pencrypt_0_ & new_n1765_;
  assign new_n1767_1_ = ~n_n2449 & new_n1766_;
  assign new_n1768_ = ~pstart_0_ & new_n1767_1_;
  assign new_n1769_ = ~new_n1764_ & ~new_n1768_;
  assign new_n1770_ = ~new_n1756_ & ~new_n1760_;
  assign new_n1771_ = new_n1769_ & new_n1770_;
  assign new_n1772_1_ = ~new_n1750_ & ~new_n1752_1_;
  assign new_n1773_ = ~new_n1741_ & ~new_n1745_;
  assign new_n1774_ = ~new_n1747_1_ & new_n1773_;
  assign new_n1775_ = new_n1772_1_ & new_n1774_;
  assign n992 = ~new_n1771_ | ~new_n1775_;
  assign new_n1777_1_ = ~pencrypt_0_ & n_n2363;
  assign new_n1778_ = ~new_n1200_ & new_n1777_1_;
  assign new_n1779_ = ~pstart_0_ & new_n1778_;
  assign new_n1780_ = n_n2457 & n_n2363;
  assign new_n1781_ = ~pencrypt_0_ & new_n1780_;
  assign new_n1782_1_ = new_n1200_ & new_n1781_;
  assign new_n1783_ = ~pstart_0_ & new_n1782_1_;
  assign new_n1784_ = pkey_37_ & pencrypt_0_;
  assign new_n1785_ = pstart_0_ & new_n1784_;
  assign new_n1786_ = ~pencrypt_0_ & n_n2457;
  assign new_n1787_1_ = ~new_n1200_ & new_n1786_;
  assign new_n1788_ = ~pstart_0_ & new_n1787_1_;
  assign new_n1789_ = ~pencrypt_0_ & pkey_45_;
  assign new_n1790_ = pstart_0_ & new_n1789_;
  assign new_n1791_ = ~n_n2363 & ~new_n1220_;
  assign new_n1792_1_ = pencrypt_0_ & new_n1791_;
  assign new_n1793_ = n_n2457 & new_n1792_1_;
  assign new_n1794_ = ~pstart_0_ & new_n1793_;
  assign new_n1795_ = n_n2363 & new_n1220_;
  assign new_n1796_ = pencrypt_0_ & new_n1795_;
  assign new_n1797_1_ = n_n2457 & new_n1796_;
  assign new_n1798_ = ~pstart_0_ & new_n1797_1_;
  assign new_n1799_ = ~n_n2457 & ~n_n2363;
  assign new_n1800_ = ~pencrypt_0_ & new_n1799_;
  assign new_n1801_ = new_n1200_ & new_n1800_;
  assign new_n1802_1_ = ~pstart_0_ & new_n1801_;
  assign new_n1803_ = n_n2363 & ~new_n1220_;
  assign new_n1804_ = pencrypt_0_ & new_n1803_;
  assign new_n1805_ = ~n_n2457 & new_n1804_;
  assign new_n1806_ = ~pstart_0_ & new_n1805_;
  assign new_n1807_1_ = ~new_n1802_1_ & ~new_n1806_;
  assign new_n1808_ = ~new_n1794_ & ~new_n1798_;
  assign new_n1809_ = new_n1807_1_ & new_n1808_;
  assign new_n1810_ = ~new_n1788_ & ~new_n1790_;
  assign new_n1811_ = ~new_n1779_ & ~new_n1783_;
  assign new_n1812_1_ = ~new_n1785_ & new_n1811_;
  assign new_n1813_ = new_n1810_ & new_n1812_1_;
  assign n997 = ~new_n1809_ | ~new_n1813_;
  assign new_n1815_ = ~pencrypt_0_ & n_n2460;
  assign new_n1816_ = new_n1200_ & new_n1815_;
  assign new_n1817_1_ = ~pstart_0_ & new_n1816_;
  assign new_n1818_ = n_n2367 & n_n2460;
  assign new_n1819_ = ~pencrypt_0_ & new_n1818_;
  assign new_n1820_ = ~new_n1200_ & new_n1819_;
  assign new_n1821_ = ~pstart_0_ & new_n1820_;
  assign new_n1822_1_ = pkey_8_ & pencrypt_0_;
  assign new_n1823_ = pstart_0_ & new_n1822_1_;
  assign new_n1824_ = ~pencrypt_0_ & n_n2367;
  assign new_n1825_ = new_n1200_ & new_n1824_;
  assign new_n1826_ = ~pstart_0_ & new_n1825_;
  assign new_n1827_1_ = pkey_16_ & ~pencrypt_0_;
  assign new_n1828_ = pstart_0_ & new_n1827_1_;
  assign new_n1829_ = n_n2460 & new_n1220_;
  assign new_n1830_ = pencrypt_0_ & new_n1829_;
  assign new_n1831_ = ~n_n2367 & new_n1830_;
  assign new_n1832_1_ = ~pstart_0_ & new_n1831_;
  assign new_n1833_ = ~n_n2460 & new_n1220_;
  assign new_n1834_ = pencrypt_0_ & new_n1833_;
  assign new_n1835_ = n_n2367 & new_n1834_;
  assign new_n1836_ = ~pstart_0_ & new_n1835_;
  assign new_n1837_1_ = ~n_n2367 & ~n_n2460;
  assign new_n1838_ = ~pencrypt_0_ & new_n1837_1_;
  assign new_n1839_ = ~new_n1200_ & new_n1838_;
  assign new_n1840_ = ~pstart_0_ & new_n1839_;
  assign new_n1841_ = n_n2460 & ~new_n1220_;
  assign new_n1842_1_ = pencrypt_0_ & new_n1841_;
  assign new_n1843_ = n_n2367 & new_n1842_1_;
  assign new_n1844_ = ~pstart_0_ & new_n1843_;
  assign new_n1845_ = ~new_n1840_ & ~new_n1844_;
  assign new_n1846_ = ~new_n1832_1_ & ~new_n1836_;
  assign new_n1847_1_ = new_n1845_ & new_n1846_;
  assign new_n1848_ = ~new_n1826_ & ~new_n1828_;
  assign new_n1849_ = ~new_n1817_1_ & ~new_n1821_;
  assign new_n1850_ = ~new_n1823_ & new_n1849_;
  assign new_n1851_ = new_n1848_ & new_n1850_;
  assign n1002 = ~new_n1847_1_ | ~new_n1851_;
  assign new_n1853_ = ~pencrypt_0_ & n_n2282;
  assign new_n1854_ = ~new_n1200_ & new_n1853_;
  assign new_n1855_ = ~pstart_0_ & new_n1854_;
  assign new_n1856_ = n_n2377 & n_n2282;
  assign new_n1857_1_ = ~pencrypt_0_ & new_n1856_;
  assign new_n1858_ = new_n1200_ & new_n1857_1_;
  assign new_n1859_ = ~pstart_0_ & new_n1858_;
  assign new_n1860_ = pkey_196_ & pencrypt_0_;
  assign new_n1861_ = pstart_0_ & new_n1860_;
  assign new_n1862_1_ = ~pencrypt_0_ & n_n2377;
  assign new_n1863_ = ~new_n1200_ & new_n1862_1_;
  assign new_n1864_ = ~pstart_0_ & new_n1863_;
  assign new_n1865_ = ~pencrypt_0_ & pkey_204_;
  assign new_n1866_ = pstart_0_ & new_n1865_;
  assign new_n1867_1_ = ~n_n2282 & ~new_n1220_;
  assign new_n1868_ = pencrypt_0_ & new_n1867_1_;
  assign new_n1869_ = n_n2377 & new_n1868_;
  assign new_n1870_ = ~pstart_0_ & new_n1869_;
  assign new_n1871_ = n_n2282 & new_n1220_;
  assign new_n1872_1_ = pencrypt_0_ & new_n1871_;
  assign new_n1873_ = n_n2377 & new_n1872_1_;
  assign new_n1874_ = ~pstart_0_ & new_n1873_;
  assign new_n1875_ = ~n_n2377 & ~n_n2282;
  assign new_n1876_ = ~pencrypt_0_ & new_n1875_;
  assign new_n1877_1_ = new_n1200_ & new_n1876_;
  assign new_n1878_ = ~pstart_0_ & new_n1877_1_;
  assign new_n1879_ = n_n2282 & ~new_n1220_;
  assign new_n1880_ = pencrypt_0_ & new_n1879_;
  assign new_n1881_ = ~n_n2377 & new_n1880_;
  assign new_n1882_1_ = ~pstart_0_ & new_n1881_;
  assign new_n1883_ = ~new_n1878_ & ~new_n1882_1_;
  assign new_n1884_ = ~new_n1870_ & ~new_n1874_;
  assign new_n1885_ = new_n1883_ & new_n1884_;
  assign new_n1886_ = ~new_n1864_ & ~new_n1866_;
  assign new_n1887_1_ = ~new_n1855_ & ~new_n1859_;
  assign new_n1888_ = ~new_n1861_ & new_n1887_1_;
  assign new_n1889_ = new_n1886_ & new_n1888_;
  assign n1007 = ~new_n1885_ | ~new_n1889_;
  assign new_n1891_ = ~pencrypt_0_ & n_n2749;
  assign new_n1892_1_ = ~new_n1200_ & new_n1891_;
  assign new_n1893_ = ~pstart_0_ & new_n1892_1_;
  assign new_n1894_ = n_n2384 & n_n2749;
  assign new_n1895_ = ~pencrypt_0_ & new_n1894_;
  assign new_n1896_ = new_n1200_ & new_n1895_;
  assign new_n1897_1_ = ~pstart_0_ & new_n1896_;
  assign new_n1898_ = pkey_252_ & pencrypt_0_;
  assign new_n1899_ = pstart_0_ & new_n1898_;
  assign new_n1900_ = ~pencrypt_0_ & n_n2384;
  assign new_n1901_ = ~new_n1200_ & new_n1900_;
  assign new_n1902_1_ = ~pstart_0_ & new_n1901_;
  assign new_n1903_ = pkey_197_ & ~pencrypt_0_;
  assign new_n1904_ = pstart_0_ & new_n1903_;
  assign new_n1905_ = ~n_n2749 & ~new_n1220_;
  assign new_n1906_ = pencrypt_0_ & new_n1905_;
  assign new_n1907_1_ = n_n2384 & new_n1906_;
  assign new_n1908_ = ~pstart_0_ & new_n1907_1_;
  assign new_n1909_ = n_n2749 & new_n1220_;
  assign new_n1910_ = pencrypt_0_ & new_n1909_;
  assign new_n1911_ = n_n2384 & new_n1910_;
  assign new_n1912_1_ = ~pstart_0_ & new_n1911_;
  assign new_n1913_ = ~n_n2384 & ~n_n2749;
  assign new_n1914_ = ~pencrypt_0_ & new_n1913_;
  assign new_n1915_ = new_n1200_ & new_n1914_;
  assign new_n1916_ = ~pstart_0_ & new_n1915_;
  assign new_n1917_1_ = n_n2749 & ~new_n1220_;
  assign new_n1918_ = pencrypt_0_ & new_n1917_1_;
  assign new_n1919_ = ~n_n2384 & new_n1918_;
  assign new_n1920_ = ~pstart_0_ & new_n1919_;
  assign new_n1921_ = ~new_n1916_ & ~new_n1920_;
  assign new_n1922_1_ = ~new_n1908_ & ~new_n1912_1_;
  assign new_n1923_ = new_n1921_ & new_n1922_1_;
  assign new_n1924_ = ~new_n1902_1_ & ~new_n1904_;
  assign new_n1925_ = ~new_n1893_ & ~new_n1897_1_;
  assign new_n1926_ = ~new_n1899_ & new_n1925_;
  assign new_n1927_1_ = new_n1924_ & new_n1926_;
  assign n1012 = ~new_n1923_ | ~new_n1927_1_;
  assign new_n1929_ = ~pencrypt_0_ & n_n2296;
  assign new_n1930_ = ~new_n1200_ & new_n1929_;
  assign new_n1931_ = ~pstart_0_ & new_n1930_;
  assign new_n1932_1_ = n_n2390 & n_n2296;
  assign new_n1933_ = ~pencrypt_0_ & new_n1932_1_;
  assign new_n1934_ = new_n1200_ & new_n1933_;
  assign new_n1935_ = ~pstart_0_ & new_n1934_;
  assign new_n1936_ = pkey_214_ & pencrypt_0_;
  assign new_n1937_1_ = pstart_0_ & new_n1936_;
  assign new_n1938_ = ~pencrypt_0_ & n_n2390;
  assign new_n1939_ = ~new_n1200_ & new_n1938_;
  assign new_n1940_ = ~pstart_0_ & new_n1939_;
  assign new_n1941_ = pkey_222_ & ~pencrypt_0_;
  assign new_n1942_1_ = pstart_0_ & new_n1941_;
  assign new_n1943_ = ~n_n2296 & ~new_n1220_;
  assign new_n1944_ = pencrypt_0_ & new_n1943_;
  assign new_n1945_ = n_n2390 & new_n1944_;
  assign new_n1946_ = ~pstart_0_ & new_n1945_;
  assign new_n1947_1_ = n_n2296 & new_n1220_;
  assign new_n1948_ = pencrypt_0_ & new_n1947_1_;
  assign new_n1949_ = n_n2390 & new_n1948_;
  assign new_n1950_ = ~pstart_0_ & new_n1949_;
  assign new_n1951_ = ~n_n2390 & ~n_n2296;
  assign new_n1952_1_ = ~pencrypt_0_ & new_n1951_;
  assign new_n1953_ = new_n1200_ & new_n1952_1_;
  assign new_n1954_ = ~pstart_0_ & new_n1953_;
  assign new_n1955_ = n_n2296 & ~new_n1220_;
  assign new_n1956_ = pencrypt_0_ & new_n1955_;
  assign new_n1957_1_ = ~n_n2390 & new_n1956_;
  assign new_n1958_ = ~pstart_0_ & new_n1957_1_;
  assign new_n1959_ = ~new_n1954_ & ~new_n1958_;
  assign new_n1960_ = ~new_n1946_ & ~new_n1950_;
  assign new_n1961_ = new_n1959_ & new_n1960_;
  assign new_n1962_1_ = ~new_n1940_ & ~new_n1942_1_;
  assign new_n1963_ = ~new_n1931_ & ~new_n1935_;
  assign new_n1964_ = ~new_n1937_1_ & new_n1963_;
  assign new_n1965_ = new_n1962_1_ & new_n1964_;
  assign n1017 = ~new_n1961_ | ~new_n1965_;
  assign new_n1967_1_ = ~pencrypt_0_ & n_n2325;
  assign new_n1968_ = ~new_n1200_ & new_n1967_1_;
  assign new_n1969_ = ~pstart_0_ & new_n1968_;
  assign new_n1970_ = n_n2419 & n_n2325;
  assign new_n1971_ = ~pencrypt_0_ & new_n1970_;
  assign new_n1972_1_ = new_n1200_ & new_n1971_;
  assign new_n1973_ = ~pstart_0_ & new_n1972_1_;
  assign new_n1974_ = pencrypt_0_ & pkey_190_;
  assign new_n1975_ = pstart_0_ & new_n1974_;
  assign new_n1976_ = ~pencrypt_0_ & n_n2419;
  assign new_n1977_1_ = ~new_n1200_ & new_n1976_;
  assign new_n1978_ = ~pstart_0_ & new_n1977_1_;
  assign new_n1979_ = pkey_67_ & ~pencrypt_0_;
  assign new_n1980_ = pstart_0_ & new_n1979_;
  assign new_n1981_ = ~n_n2325 & ~new_n1220_;
  assign new_n1982_1_ = pencrypt_0_ & new_n1981_;
  assign new_n1983_ = n_n2419 & new_n1982_1_;
  assign new_n1984_ = ~pstart_0_ & new_n1983_;
  assign new_n1985_ = n_n2325 & new_n1220_;
  assign new_n1986_ = pencrypt_0_ & new_n1985_;
  assign new_n1987_1_ = n_n2419 & new_n1986_;
  assign new_n1988_ = ~pstart_0_ & new_n1987_1_;
  assign new_n1989_ = ~n_n2419 & ~n_n2325;
  assign new_n1990_ = ~pencrypt_0_ & new_n1989_;
  assign new_n1991_ = new_n1200_ & new_n1990_;
  assign new_n1992_1_ = ~pstart_0_ & new_n1991_;
  assign new_n1993_ = n_n2325 & ~new_n1220_;
  assign new_n1994_ = pencrypt_0_ & new_n1993_;
  assign new_n1995_ = ~n_n2419 & new_n1994_;
  assign new_n1996_ = ~pstart_0_ & new_n1995_;
  assign new_n1997_1_ = ~new_n1992_1_ & ~new_n1996_;
  assign new_n1998_ = ~new_n1984_ & ~new_n1988_;
  assign new_n1999_ = new_n1997_1_ & new_n1998_;
  assign new_n2000_ = ~new_n1978_ & ~new_n1980_;
  assign new_n2001_ = ~new_n1969_ & ~new_n1973_;
  assign new_n2002_1_ = ~new_n1975_ & new_n2001_;
  assign new_n2003_ = new_n2000_ & new_n2002_1_;
  assign n1022 = ~new_n1999_ | ~new_n2003_;
  assign new_n2005_ = ~pencrypt_0_ & n_n2333;
  assign new_n2006_ = ~new_n1200_ & new_n2005_;
  assign new_n2007_1_ = ~pstart_0_ & new_n2006_;
  assign new_n2008_ = n_n2429 & n_n2333;
  assign new_n2009_ = ~pencrypt_0_ & new_n2008_;
  assign new_n2010_ = new_n1200_ & new_n2009_;
  assign new_n2011_ = ~pstart_0_ & new_n2010_;
  assign new_n2012_1_ = pkey_116_ & pencrypt_0_;
  assign new_n2013_ = pstart_0_ & new_n2012_1_;
  assign new_n2014_ = ~pencrypt_0_ & n_n2429;
  assign new_n2015_ = ~new_n1200_ & new_n2014_;
  assign new_n2016_ = ~pstart_0_ & new_n2015_;
  assign new_n2017_1_ = pkey_124_ & ~pencrypt_0_;
  assign new_n2018_ = pstart_0_ & new_n2017_1_;
  assign new_n2019_ = ~n_n2333 & ~new_n1220_;
  assign new_n2020_ = pencrypt_0_ & new_n2019_;
  assign new_n2021_ = n_n2429 & new_n2020_;
  assign new_n2022_1_ = ~pstart_0_ & new_n2021_;
  assign new_n2023_ = n_n2333 & new_n1220_;
  assign new_n2024_ = pencrypt_0_ & new_n2023_;
  assign new_n2025_ = n_n2429 & new_n2024_;
  assign new_n2026_ = ~pstart_0_ & new_n2025_;
  assign new_n2027_1_ = ~n_n2429 & ~n_n2333;
  assign new_n2028_ = ~pencrypt_0_ & new_n2027_1_;
  assign new_n2029_ = new_n1200_ & new_n2028_;
  assign new_n2030_ = ~pstart_0_ & new_n2029_;
  assign new_n2031_ = n_n2333 & ~new_n1220_;
  assign new_n2032_1_ = pencrypt_0_ & new_n2031_;
  assign new_n2033_ = ~n_n2429 & new_n2032_1_;
  assign new_n2034_ = ~pstart_0_ & new_n2033_;
  assign new_n2035_ = ~new_n2030_ & ~new_n2034_;
  assign new_n2036_ = ~new_n2022_1_ & ~new_n2026_;
  assign new_n2037_1_ = new_n2035_ & new_n2036_;
  assign new_n2038_ = ~new_n2016_ & ~new_n2018_;
  assign new_n2039_ = ~new_n2007_1_ & ~new_n2011_;
  assign new_n2040_ = ~new_n2013_ & new_n2039_;
  assign new_n2041_ = new_n2038_ & new_n2040_;
  assign n1027 = ~new_n2037_1_ | ~new_n2041_;
  assign new_n2043_ = ~pencrypt_0_ & n_n2356;
  assign new_n2044_ = ~new_n1200_ & new_n2043_;
  assign new_n2045_ = ~pstart_0_ & new_n2044_;
  assign new_n2046_ = n_n2450 & n_n2356;
  assign new_n2047_ = ~pencrypt_0_ & new_n2046_;
  assign new_n2048_ = new_n1200_ & new_n2047_;
  assign new_n2049_ = ~pstart_0_ & new_n2048_;
  assign new_n2050_ = pkey_36_ & pencrypt_0_;
  assign new_n2051_ = pstart_0_ & new_n2050_;
  assign new_n2052_ = ~pencrypt_0_ & n_n2450;
  assign new_n2053_ = ~new_n1200_ & new_n2052_;
  assign new_n2054_ = ~pstart_0_ & new_n2053_;
  assign new_n2055_ = ~pencrypt_0_ & pkey_44_;
  assign new_n2056_ = pstart_0_ & new_n2055_;
  assign new_n2057_ = ~n_n2356 & ~new_n1220_;
  assign new_n2058_ = pencrypt_0_ & new_n2057_;
  assign new_n2059_ = n_n2450 & new_n2058_;
  assign new_n2060_ = ~pstart_0_ & new_n2059_;
  assign new_n2061_ = n_n2356 & new_n1220_;
  assign new_n2062_ = pencrypt_0_ & new_n2061_;
  assign new_n2063_ = n_n2450 & new_n2062_;
  assign new_n2064_ = ~pstart_0_ & new_n2063_;
  assign new_n2065_ = ~n_n2450 & ~n_n2356;
  assign new_n2066_ = ~pencrypt_0_ & new_n2065_;
  assign new_n2067_ = new_n1200_ & new_n2066_;
  assign new_n2068_ = ~pstart_0_ & new_n2067_;
  assign new_n2069_ = n_n2356 & ~new_n1220_;
  assign new_n2070_ = pencrypt_0_ & new_n2069_;
  assign new_n2071_ = ~n_n2450 & new_n2070_;
  assign new_n2072_ = ~pstart_0_ & new_n2071_;
  assign new_n2073_ = ~new_n2068_ & ~new_n2072_;
  assign new_n2074_ = ~new_n2060_ & ~new_n2064_;
  assign new_n2075_ = new_n2073_ & new_n2074_;
  assign new_n2076_ = ~new_n2054_ & ~new_n2056_;
  assign new_n2077_ = ~new_n2045_ & ~new_n2049_;
  assign new_n2078_ = ~new_n2051_ & new_n2077_;
  assign new_n2079_ = new_n2076_ & new_n2078_;
  assign n1032 = ~new_n2075_ | ~new_n2079_;
  assign new_n2081_ = ~new_n1200_ & new_n1210_;
  assign new_n2082_ = ~pstart_0_ & new_n2081_;
  assign new_n2083_ = new_n1200_ & new_n1205_;
  assign new_n2084_ = ~pstart_0_ & new_n2083_;
  assign new_n2085_ = pkey_61_ & pencrypt_0_;
  assign new_n2086_ = pstart_0_ & new_n2085_;
  assign new_n2087_ = ~new_n1200_ & new_n1201_;
  assign new_n2088_ = ~pstart_0_ & new_n2087_;
  assign new_n2089_ = pkey_6_ & ~pencrypt_0_;
  assign new_n2090_ = pstart_0_ & new_n2089_;
  assign new_n2091_ = ~n_n2365 & ~new_n1220_;
  assign new_n2092_ = pencrypt_0_ & new_n2091_;
  assign new_n2093_ = n_n2459 & new_n2092_;
  assign new_n2094_ = ~pstart_0_ & new_n2093_;
  assign new_n2095_ = n_n2365 & new_n1220_;
  assign new_n2096_ = pencrypt_0_ & new_n2095_;
  assign new_n2097_ = n_n2459 & new_n2096_;
  assign new_n2098_ = ~pstart_0_ & new_n2097_;
  assign new_n2099_ = new_n1200_ & new_n1230_;
  assign new_n2100_ = ~pstart_0_ & new_n2099_;
  assign new_n2101_ = n_n2365 & ~new_n1220_;
  assign new_n2102_ = pencrypt_0_ & new_n2101_;
  assign new_n2103_ = ~n_n2459 & new_n2102_;
  assign new_n2104_ = ~pstart_0_ & new_n2103_;
  assign new_n2105_ = ~new_n2100_ & ~new_n2104_;
  assign new_n2106_ = ~new_n2094_ & ~new_n2098_;
  assign new_n2107_ = new_n2105_ & new_n2106_;
  assign new_n2108_ = ~new_n2088_ & ~new_n2090_;
  assign new_n2109_ = ~new_n2082_ & ~new_n2084_;
  assign new_n2110_ = ~new_n2086_ & new_n2109_;
  assign new_n2111_ = new_n2108_ & new_n2110_;
  assign n1037 = ~new_n2107_ | ~new_n2111_;
  assign new_n2113_ = ~pencrypt_0_ & n_n2372;
  assign new_n2114_ = ~new_n1200_ & new_n2113_;
  assign new_n2115_ = ~pstart_0_ & new_n2114_;
  assign new_n2116_ = n_n2465 & n_n2372;
  assign new_n2117_ = ~pencrypt_0_ & new_n2116_;
  assign new_n2118_ = new_n1200_ & new_n2117_;
  assign new_n2119_ = ~pstart_0_ & new_n2118_;
  assign new_n2120_ = pencrypt_0_ & pkey_54_;
  assign new_n2121_ = pstart_0_ & new_n2120_;
  assign new_n2122_ = ~pencrypt_0_ & n_n2465;
  assign new_n2123_ = ~new_n1200_ & new_n2122_;
  assign new_n2124_ = ~pstart_0_ & new_n2123_;
  assign new_n2125_ = ~pencrypt_0_ & pkey_62_;
  assign new_n2126_ = pstart_0_ & new_n2125_;
  assign new_n2127_ = ~n_n2372 & ~new_n1220_;
  assign new_n2128_ = pencrypt_0_ & new_n2127_;
  assign new_n2129_ = n_n2465 & new_n2128_;
  assign new_n2130_ = ~pstart_0_ & new_n2129_;
  assign new_n2131_ = n_n2372 & new_n1220_;
  assign new_n2132_ = pencrypt_0_ & new_n2131_;
  assign new_n2133_ = n_n2465 & new_n2132_;
  assign new_n2134_ = ~pstart_0_ & new_n2133_;
  assign new_n2135_ = ~n_n2465 & ~n_n2372;
  assign new_n2136_ = ~pencrypt_0_ & new_n2135_;
  assign new_n2137_ = new_n1200_ & new_n2136_;
  assign new_n2138_ = ~pstart_0_ & new_n2137_;
  assign new_n2139_ = n_n2372 & ~new_n1220_;
  assign new_n2140_ = pencrypt_0_ & new_n2139_;
  assign new_n2141_ = ~n_n2465 & new_n2140_;
  assign new_n2142_ = ~pstart_0_ & new_n2141_;
  assign new_n2143_ = ~new_n2138_ & ~new_n2142_;
  assign new_n2144_ = ~new_n2130_ & ~new_n2134_;
  assign new_n2145_ = new_n2143_ & new_n2144_;
  assign new_n2146_ = ~new_n2124_ & ~new_n2126_;
  assign new_n2147_ = ~new_n2115_ & ~new_n2119_;
  assign new_n2148_ = ~new_n2121_ & new_n2147_;
  assign new_n2149_ = new_n2146_ & new_n2148_;
  assign n1042 = ~new_n2145_ | ~new_n2149_;
  assign new_n2151_ = ~pencrypt_0_ & n_n2461;
  assign new_n2152_ = new_n1200_ & new_n2151_;
  assign new_n2153_ = ~pstart_0_ & new_n2152_;
  assign new_n2154_ = n_n2368 & n_n2461;
  assign new_n2155_ = ~pencrypt_0_ & new_n2154_;
  assign new_n2156_ = ~new_n1200_ & new_n2155_;
  assign new_n2157_ = ~pstart_0_ & new_n2156_;
  assign new_n2158_ = pkey_16_ & pencrypt_0_;
  assign new_n2159_ = pstart_0_ & new_n2158_;
  assign new_n2160_ = ~pencrypt_0_ & n_n2368;
  assign new_n2161_ = new_n1200_ & new_n2160_;
  assign new_n2162_ = ~pstart_0_ & new_n2161_;
  assign new_n2163_ = ~pencrypt_0_ & pkey_24_;
  assign new_n2164_ = pstart_0_ & new_n2163_;
  assign new_n2165_ = n_n2461 & new_n1220_;
  assign new_n2166_ = pencrypt_0_ & new_n2165_;
  assign new_n2167_ = ~n_n2368 & new_n2166_;
  assign new_n2168_ = ~pstart_0_ & new_n2167_;
  assign new_n2169_ = ~n_n2461 & new_n1220_;
  assign new_n2170_ = pencrypt_0_ & new_n2169_;
  assign new_n2171_ = n_n2368 & new_n2170_;
  assign new_n2172_ = ~pstart_0_ & new_n2171_;
  assign new_n2173_ = ~n_n2368 & ~n_n2461;
  assign new_n2174_ = ~pencrypt_0_ & new_n2173_;
  assign new_n2175_ = ~new_n1200_ & new_n2174_;
  assign new_n2176_ = ~pstart_0_ & new_n2175_;
  assign new_n2177_ = n_n2461 & ~new_n1220_;
  assign new_n2178_ = pencrypt_0_ & new_n2177_;
  assign new_n2179_ = n_n2368 & new_n2178_;
  assign new_n2180_ = ~pstart_0_ & new_n2179_;
  assign new_n2181_ = ~new_n2176_ & ~new_n2180_;
  assign new_n2182_ = ~new_n2168_ & ~new_n2172_;
  assign new_n2183_ = new_n2181_ & new_n2182_;
  assign new_n2184_ = ~new_n2162_ & ~new_n2164_;
  assign new_n2185_ = ~new_n2153_ & ~new_n2157_;
  assign new_n2186_ = ~new_n2159_ & new_n2185_;
  assign new_n2187_ = new_n2184_ & new_n2186_;
  assign n1047 = ~new_n2183_ | ~new_n2187_;
  assign new_n2189_ = ~pencrypt_0_ & n_n2281;
  assign new_n2190_ = ~new_n1200_ & new_n2189_;
  assign new_n2191_ = ~pstart_0_ & new_n2190_;
  assign new_n2192_ = n_n2376 & n_n2281;
  assign new_n2193_ = ~pencrypt_0_ & new_n2192_;
  assign new_n2194_ = new_n1200_ & new_n2193_;
  assign new_n2195_ = ~pstart_0_ & new_n2194_;
  assign new_n2196_ = pkey_219_ & pencrypt_0_;
  assign new_n2197_ = pstart_0_ & new_n2196_;
  assign new_n2198_ = ~pencrypt_0_ & n_n2376;
  assign new_n2199_ = ~new_n1200_ & new_n2198_;
  assign new_n2200_ = ~pstart_0_ & new_n2199_;
  assign new_n2201_ = pkey_196_ & ~pencrypt_0_;
  assign new_n2202_ = pstart_0_ & new_n2201_;
  assign new_n2203_ = ~n_n2281 & ~new_n1220_;
  assign new_n2204_ = pencrypt_0_ & new_n2203_;
  assign new_n2205_ = n_n2376 & new_n2204_;
  assign new_n2206_ = ~pstart_0_ & new_n2205_;
  assign new_n2207_ = n_n2281 & new_n1220_;
  assign new_n2208_ = pencrypt_0_ & new_n2207_;
  assign new_n2209_ = n_n2376 & new_n2208_;
  assign new_n2210_ = ~pstart_0_ & new_n2209_;
  assign new_n2211_ = ~n_n2376 & ~n_n2281;
  assign new_n2212_ = ~pencrypt_0_ & new_n2211_;
  assign new_n2213_ = new_n1200_ & new_n2212_;
  assign new_n2214_ = ~pstart_0_ & new_n2213_;
  assign new_n2215_ = n_n2281 & ~new_n1220_;
  assign new_n2216_ = pencrypt_0_ & new_n2215_;
  assign new_n2217_ = ~n_n2376 & new_n2216_;
  assign new_n2218_ = ~pstart_0_ & new_n2217_;
  assign new_n2219_ = ~new_n2214_ & ~new_n2218_;
  assign new_n2220_ = ~new_n2206_ & ~new_n2210_;
  assign new_n2221_ = new_n2219_ & new_n2220_;
  assign new_n2222_ = ~new_n2200_ & ~new_n2202_;
  assign new_n2223_ = ~new_n2191_ & ~new_n2195_;
  assign new_n2224_ = ~new_n2197_ & new_n2223_;
  assign new_n2225_ = new_n2222_ & new_n2224_;
  assign n1052 = ~new_n2221_ | ~new_n2225_;
  assign new_n2227_ = ~pencrypt_0_ & n_n2287;
  assign new_n2228_ = ~new_n1200_ & new_n2227_;
  assign new_n2229_ = ~pstart_0_ & new_n2228_;
  assign new_n2230_ = n_n2877 & n_n2287;
  assign new_n2231_ = ~pencrypt_0_ & new_n2230_;
  assign new_n2232_ = new_n1200_ & new_n2231_;
  assign new_n2233_ = ~pstart_0_ & new_n2232_;
  assign new_n2234_ = pkey_197_ & pencrypt_0_;
  assign new_n2235_ = pstart_0_ & new_n2234_;
  assign new_n2236_ = ~pencrypt_0_ & n_n2877;
  assign new_n2237_ = ~new_n1200_ & new_n2236_;
  assign new_n2238_ = ~pstart_0_ & new_n2237_;
  assign new_n2239_ = ~pencrypt_0_ & pkey_205_;
  assign new_n2240_ = pstart_0_ & new_n2239_;
  assign new_n2241_ = ~n_n2287 & ~new_n1220_;
  assign new_n2242_ = pencrypt_0_ & new_n2241_;
  assign new_n2243_ = n_n2877 & new_n2242_;
  assign new_n2244_ = ~pstart_0_ & new_n2243_;
  assign new_n2245_ = n_n2287 & new_n1220_;
  assign new_n2246_ = pencrypt_0_ & new_n2245_;
  assign new_n2247_ = n_n2877 & new_n2246_;
  assign new_n2248_ = ~pstart_0_ & new_n2247_;
  assign new_n2249_ = ~n_n2877 & ~n_n2287;
  assign new_n2250_ = ~pencrypt_0_ & new_n2249_;
  assign new_n2251_ = new_n1200_ & new_n2250_;
  assign new_n2252_ = ~pstart_0_ & new_n2251_;
  assign new_n2253_ = n_n2287 & ~new_n1220_;
  assign new_n2254_ = pencrypt_0_ & new_n2253_;
  assign new_n2255_ = ~n_n2877 & new_n2254_;
  assign new_n2256_ = ~pstart_0_ & new_n2255_;
  assign new_n2257_ = ~new_n2252_ & ~new_n2256_;
  assign new_n2258_ = ~new_n2244_ & ~new_n2248_;
  assign new_n2259_ = new_n2257_ & new_n2258_;
  assign new_n2260_ = ~new_n2238_ & ~new_n2240_;
  assign new_n2261_ = ~new_n2229_ & ~new_n2233_;
  assign new_n2262_ = ~new_n2235_ & new_n2261_;
  assign new_n2263_ = new_n2260_ & new_n2262_;
  assign n1057 = ~new_n2259_ | ~new_n2263_;
  assign new_n2265_ = ~pencrypt_0_ & n_n2295;
  assign new_n2266_ = ~new_n1200_ & new_n2265_;
  assign new_n2267_ = ~pstart_0_ & new_n2266_;
  assign new_n2268_ = n_n2389 & n_n2295;
  assign new_n2269_ = ~pencrypt_0_ & new_n2268_;
  assign new_n2270_ = new_n1200_ & new_n2269_;
  assign new_n2271_ = ~pstart_0_ & new_n2270_;
  assign new_n2272_ = pkey_206_ & pencrypt_0_;
  assign new_n2273_ = pstart_0_ & new_n2272_;
  assign new_n2274_ = ~pencrypt_0_ & n_n2389;
  assign new_n2275_ = ~new_n1200_ & new_n2274_;
  assign new_n2276_ = ~pstart_0_ & new_n2275_;
  assign new_n2277_ = pkey_214_ & ~pencrypt_0_;
  assign new_n2278_ = pstart_0_ & new_n2277_;
  assign new_n2279_ = ~n_n2295 & ~new_n1220_;
  assign new_n2280_ = pencrypt_0_ & new_n2279_;
  assign new_n2281_ = n_n2389 & new_n2280_;
  assign new_n2282_ = ~pstart_0_ & new_n2281_;
  assign new_n2283_ = n_n2295 & new_n1220_;
  assign new_n2284_ = pencrypt_0_ & new_n2283_;
  assign new_n2285_ = n_n2389 & new_n2284_;
  assign new_n2286_ = ~pstart_0_ & new_n2285_;
  assign new_n2287_ = ~n_n2389 & ~n_n2295;
  assign new_n2288_ = ~pencrypt_0_ & new_n2287_;
  assign new_n2289_ = new_n1200_ & new_n2288_;
  assign new_n2290_ = ~pstart_0_ & new_n2289_;
  assign new_n2291_ = n_n2295 & ~new_n1220_;
  assign new_n2292_ = pencrypt_0_ & new_n2291_;
  assign new_n2293_ = ~n_n2389 & new_n2292_;
  assign new_n2294_ = ~pstart_0_ & new_n2293_;
  assign new_n2295_ = ~new_n2290_ & ~new_n2294_;
  assign new_n2296_ = ~new_n2282_ & ~new_n2286_;
  assign new_n2297_ = new_n2295_ & new_n2296_;
  assign new_n2298_ = ~new_n2276_ & ~new_n2278_;
  assign new_n2299_ = ~new_n2267_ & ~new_n2271_;
  assign new_n2300_ = ~new_n2273_ & new_n2299_;
  assign new_n2301_ = new_n2298_ & new_n2300_;
  assign n1062 = ~new_n2297_ | ~new_n2301_;
  assign new_n2303_ = ~pencrypt_0_ & n_n2326;
  assign new_n2304_ = ~new_n1200_ & new_n2303_;
  assign new_n2305_ = ~pstart_0_ & new_n2304_;
  assign new_n2306_ = n_n2420 & n_n2326;
  assign new_n2307_ = ~pencrypt_0_ & new_n2306_;
  assign new_n2308_ = new_n1200_ & new_n2307_;
  assign new_n2309_ = ~pstart_0_ & new_n2308_;
  assign new_n2310_ = pkey_67_ & pencrypt_0_;
  assign new_n2311_ = pstart_0_ & new_n2310_;
  assign new_n2312_ = ~pencrypt_0_ & n_n2420;
  assign new_n2313_ = ~new_n1200_ & new_n2312_;
  assign new_n2314_ = ~pstart_0_ & new_n2313_;
  assign new_n2315_ = ~pencrypt_0_ & pkey_75_;
  assign new_n2316_ = pstart_0_ & new_n2315_;
  assign new_n2317_ = ~n_n2326 & ~new_n1220_;
  assign new_n2318_ = pencrypt_0_ & new_n2317_;
  assign new_n2319_ = n_n2420 & new_n2318_;
  assign new_n2320_ = ~pstart_0_ & new_n2319_;
  assign new_n2321_ = n_n2326 & new_n1220_;
  assign new_n2322_ = pencrypt_0_ & new_n2321_;
  assign new_n2323_ = n_n2420 & new_n2322_;
  assign new_n2324_ = ~pstart_0_ & new_n2323_;
  assign new_n2325_ = ~n_n2420 & ~n_n2326;
  assign new_n2326_ = ~pencrypt_0_ & new_n2325_;
  assign new_n2327_ = new_n1200_ & new_n2326_;
  assign new_n2328_ = ~pstart_0_ & new_n2327_;
  assign new_n2329_ = n_n2326 & ~new_n1220_;
  assign new_n2330_ = pencrypt_0_ & new_n2329_;
  assign new_n2331_ = ~n_n2420 & new_n2330_;
  assign new_n2332_ = ~pstart_0_ & new_n2331_;
  assign new_n2333_ = ~new_n2328_ & ~new_n2332_;
  assign new_n2334_ = ~new_n2320_ & ~new_n2324_;
  assign new_n2335_ = new_n2333_ & new_n2334_;
  assign new_n2336_ = ~new_n2314_ & ~new_n2316_;
  assign new_n2337_ = ~new_n2305_ & ~new_n2309_;
  assign new_n2338_ = ~new_n2311_ & new_n2337_;
  assign new_n2339_ = new_n2336_ & new_n2338_;
  assign n1067 = ~new_n2335_ | ~new_n2339_;
  assign new_n2341_ = ~pencrypt_0_ & n_n2811;
  assign new_n2342_ = ~new_n1200_ & new_n2341_;
  assign new_n2343_ = ~pstart_0_ & new_n2342_;
  assign new_n2344_ = n_n2428 & n_n2811;
  assign new_n2345_ = ~pencrypt_0_ & new_n2344_;
  assign new_n2346_ = new_n1200_ & new_n2345_;
  assign new_n2347_ = ~pstart_0_ & new_n2346_;
  assign new_n2348_ = pencrypt_0_ & pkey_44_;
  assign new_n2349_ = pstart_0_ & new_n2348_;
  assign new_n2350_ = ~pencrypt_0_ & n_n2428;
  assign new_n2351_ = ~new_n1200_ & new_n2350_;
  assign new_n2352_ = ~pstart_0_ & new_n2351_;
  assign new_n2353_ = pkey_116_ & ~pencrypt_0_;
  assign new_n2354_ = pstart_0_ & new_n2353_;
  assign new_n2355_ = ~n_n2811 & ~new_n1220_;
  assign new_n2356_ = pencrypt_0_ & new_n2355_;
  assign new_n2357_ = n_n2428 & new_n2356_;
  assign new_n2358_ = ~pstart_0_ & new_n2357_;
  assign new_n2359_ = n_n2811 & new_n1220_;
  assign new_n2360_ = pencrypt_0_ & new_n2359_;
  assign new_n2361_ = n_n2428 & new_n2360_;
  assign new_n2362_ = ~pstart_0_ & new_n2361_;
  assign new_n2363_ = ~n_n2428 & ~n_n2811;
  assign new_n2364_ = ~pencrypt_0_ & new_n2363_;
  assign new_n2365_ = new_n1200_ & new_n2364_;
  assign new_n2366_ = ~pstart_0_ & new_n2365_;
  assign new_n2367_ = n_n2811 & ~new_n1220_;
  assign new_n2368_ = pencrypt_0_ & new_n2367_;
  assign new_n2369_ = ~n_n2428 & new_n2368_;
  assign new_n2370_ = ~pstart_0_ & new_n2369_;
  assign new_n2371_ = ~new_n2366_ & ~new_n2370_;
  assign new_n2372_ = ~new_n2358_ & ~new_n2362_;
  assign new_n2373_ = new_n2371_ & new_n2372_;
  assign new_n2374_ = ~new_n2352_ & ~new_n2354_;
  assign new_n2375_ = ~new_n2343_ & ~new_n2347_;
  assign new_n2376_ = ~new_n2349_ & new_n2375_;
  assign new_n2377_ = new_n2374_ & new_n2376_;
  assign n1072 = ~new_n2373_ | ~new_n2377_;
  assign new_n2379_ = ~pencrypt_0_ & n_n2843;
  assign new_n2380_ = ~new_n1200_ & new_n2379_;
  assign new_n2381_ = ~pstart_0_ & new_n2380_;
  assign new_n2382_ = n_n2451 & n_n2843;
  assign new_n2383_ = ~pencrypt_0_ & new_n2382_;
  assign new_n2384_ = new_n1200_ & new_n2383_;
  assign new_n2385_ = ~pstart_0_ & new_n2384_;
  assign new_n2386_ = ~pencrypt_0_ & n_n2451;
  assign new_n2387_ = ~new_n1200_ & new_n2386_;
  assign new_n2388_ = ~pstart_0_ & new_n2387_;
  assign new_n2389_ = pkey_52_ & ~pencrypt_0_;
  assign new_n2390_ = pstart_0_ & new_n2389_;
  assign new_n2391_ = ~n_n2843 & ~new_n1220_;
  assign new_n2392_ = pencrypt_0_ & new_n2391_;
  assign new_n2393_ = n_n2451 & new_n2392_;
  assign new_n2394_ = ~pstart_0_ & new_n2393_;
  assign new_n2395_ = n_n2843 & new_n1220_;
  assign new_n2396_ = pencrypt_0_ & new_n2395_;
  assign new_n2397_ = n_n2451 & new_n2396_;
  assign new_n2398_ = ~pstart_0_ & new_n2397_;
  assign new_n2399_ = ~n_n2451 & ~n_n2843;
  assign new_n2400_ = ~pencrypt_0_ & new_n2399_;
  assign new_n2401_ = new_n1200_ & new_n2400_;
  assign new_n2402_ = ~pstart_0_ & new_n2401_;
  assign new_n2403_ = n_n2843 & ~new_n1220_;
  assign new_n2404_ = pencrypt_0_ & new_n2403_;
  assign new_n2405_ = ~n_n2451 & new_n2404_;
  assign new_n2406_ = ~pstart_0_ & new_n2405_;
  assign new_n2407_ = ~new_n2402_ & ~new_n2406_;
  assign new_n2408_ = ~new_n2394_ & ~new_n2398_;
  assign new_n2409_ = new_n2407_ & new_n2408_;
  assign new_n2410_ = ~new_n2388_ & ~new_n2390_;
  assign new_n2411_ = ~new_n2381_ & ~new_n2385_;
  assign new_n2412_ = ~new_n2349_ & new_n2411_;
  assign new_n2413_ = new_n2410_ & new_n2412_;
  assign n1077 = ~new_n2409_ | ~new_n2413_;
  assign new_n2415_ = ~pencrypt_0_ & n_n2853;
  assign new_n2416_ = ~new_n1200_ & new_n2415_;
  assign new_n2417_ = ~pstart_0_ & new_n2416_;
  assign new_n2418_ = n_n2458 & n_n2853;
  assign new_n2419_ = ~pencrypt_0_ & new_n2418_;
  assign new_n2420_ = new_n1200_ & new_n2419_;
  assign new_n2421_ = ~pstart_0_ & new_n2420_;
  assign new_n2422_ = pencrypt_0_ & pkey_53_;
  assign new_n2423_ = pstart_0_ & new_n2422_;
  assign new_n2424_ = ~pencrypt_0_ & n_n2458;
  assign new_n2425_ = ~new_n1200_ & new_n2424_;
  assign new_n2426_ = ~pstart_0_ & new_n2425_;
  assign new_n2427_ = pkey_61_ & ~pencrypt_0_;
  assign new_n2428_ = pstart_0_ & new_n2427_;
  assign new_n2429_ = ~n_n2853 & ~new_n1220_;
  assign new_n2430_ = pencrypt_0_ & new_n2429_;
  assign new_n2431_ = n_n2458 & new_n2430_;
  assign new_n2432_ = ~pstart_0_ & new_n2431_;
  assign new_n2433_ = n_n2853 & new_n1220_;
  assign new_n2434_ = pencrypt_0_ & new_n2433_;
  assign new_n2435_ = n_n2458 & new_n2434_;
  assign new_n2436_ = ~pstart_0_ & new_n2435_;
  assign new_n2437_ = ~n_n2458 & ~n_n2853;
  assign new_n2438_ = ~pencrypt_0_ & new_n2437_;
  assign new_n2439_ = new_n1200_ & new_n2438_;
  assign new_n2440_ = ~pstart_0_ & new_n2439_;
  assign new_n2441_ = n_n2853 & ~new_n1220_;
  assign new_n2442_ = pencrypt_0_ & new_n2441_;
  assign new_n2443_ = ~n_n2458 & new_n2442_;
  assign new_n2444_ = ~pstart_0_ & new_n2443_;
  assign new_n2445_ = ~new_n2440_ & ~new_n2444_;
  assign new_n2446_ = ~new_n2432_ & ~new_n2436_;
  assign new_n2447_ = new_n2445_ & new_n2446_;
  assign new_n2448_ = ~new_n2426_ & ~new_n2428_;
  assign new_n2449_ = ~new_n2417_ & ~new_n2421_;
  assign new_n2450_ = ~new_n2423_ & new_n2449_;
  assign new_n2451_ = new_n2448_ & new_n2450_;
  assign n1082 = ~new_n2447_ | ~new_n2451_;
  assign new_n2453_ = ~pencrypt_0_ & n_n2381;
  assign new_n2454_ = new_n1200_ & new_n2453_;
  assign new_n2455_ = ~pstart_0_ & new_n2454_;
  assign new_n2456_ = n_n2285 & n_n2381;
  assign new_n2457_ = ~pencrypt_0_ & new_n2456_;
  assign new_n2458_ = ~new_n1200_ & new_n2457_;
  assign new_n2459_ = ~pstart_0_ & new_n2458_;
  assign new_n2460_ = pkey_226_ & pencrypt_0_;
  assign new_n2461_ = pstart_0_ & new_n2460_;
  assign new_n2462_ = ~pencrypt_0_ & n_n2285;
  assign new_n2463_ = new_n1200_ & new_n2462_;
  assign new_n2464_ = ~pstart_0_ & new_n2463_;
  assign new_n2465_ = pkey_234_ & ~pencrypt_0_;
  assign new_n2466_ = pstart_0_ & new_n2465_;
  assign new_n2467_ = n_n2381 & new_n1220_;
  assign new_n2468_ = pencrypt_0_ & new_n2467_;
  assign new_n2469_ = ~n_n2285 & new_n2468_;
  assign new_n2470_ = ~pstart_0_ & new_n2469_;
  assign new_n2471_ = ~n_n2381 & new_n1220_;
  assign new_n2472_ = pencrypt_0_ & new_n2471_;
  assign new_n2473_ = n_n2285 & new_n2472_;
  assign new_n2474_ = ~pstart_0_ & new_n2473_;
  assign new_n2475_ = ~n_n2285 & ~n_n2381;
  assign new_n2476_ = ~pencrypt_0_ & new_n2475_;
  assign new_n2477_ = ~new_n1200_ & new_n2476_;
  assign new_n2478_ = ~pstart_0_ & new_n2477_;
  assign new_n2479_ = n_n2381 & ~new_n1220_;
  assign new_n2480_ = pencrypt_0_ & new_n2479_;
  assign new_n2481_ = n_n2285 & new_n2480_;
  assign new_n2482_ = ~pstart_0_ & new_n2481_;
  assign new_n2483_ = ~new_n2478_ & ~new_n2482_;
  assign new_n2484_ = ~new_n2470_ & ~new_n2474_;
  assign new_n2485_ = new_n2483_ & new_n2484_;
  assign new_n2486_ = ~new_n2464_ & ~new_n2466_;
  assign new_n2487_ = ~new_n2455_ & ~new_n2459_;
  assign new_n2488_ = ~new_n2461_ & new_n2487_;
  assign new_n2489_ = new_n2486_ & new_n2488_;
  assign n1087 = ~new_n2485_ | ~new_n2489_;
  assign new_n2491_ = ~pencrypt_0_ & n_n2456;
  assign new_n2492_ = new_n1200_ & new_n2491_;
  assign new_n2493_ = ~pstart_0_ & new_n2492_;
  assign new_n2494_ = n_n2362 & n_n2456;
  assign new_n2495_ = ~pencrypt_0_ & new_n2494_;
  assign new_n2496_ = ~new_n1200_ & new_n2495_;
  assign new_n2497_ = ~pstart_0_ & new_n2496_;
  assign new_n2498_ = pencrypt_0_ & pkey_25_;
  assign new_n2499_ = pstart_0_ & new_n2498_;
  assign new_n2500_ = ~pencrypt_0_ & n_n2362;
  assign new_n2501_ = new_n1200_ & new_n2500_;
  assign new_n2502_ = ~pstart_0_ & new_n2501_;
  assign new_n2503_ = ~pencrypt_0_ & pkey_33_;
  assign new_n2504_ = pstart_0_ & new_n2503_;
  assign new_n2505_ = n_n2456 & new_n1220_;
  assign new_n2506_ = pencrypt_0_ & new_n2505_;
  assign new_n2507_ = ~n_n2362 & new_n2506_;
  assign new_n2508_ = ~pstart_0_ & new_n2507_;
  assign new_n2509_ = ~n_n2456 & new_n1220_;
  assign new_n2510_ = pencrypt_0_ & new_n2509_;
  assign new_n2511_ = n_n2362 & new_n2510_;
  assign new_n2512_ = ~pstart_0_ & new_n2511_;
  assign new_n2513_ = ~n_n2362 & ~n_n2456;
  assign new_n2514_ = ~pencrypt_0_ & new_n2513_;
  assign new_n2515_ = ~new_n1200_ & new_n2514_;
  assign new_n2516_ = ~pstart_0_ & new_n2515_;
  assign new_n2517_ = n_n2456 & ~new_n1220_;
  assign new_n2518_ = pencrypt_0_ & new_n2517_;
  assign new_n2519_ = n_n2362 & new_n2518_;
  assign new_n2520_ = ~pstart_0_ & new_n2519_;
  assign new_n2521_ = ~new_n2516_ & ~new_n2520_;
  assign new_n2522_ = ~new_n2508_ & ~new_n2512_;
  assign new_n2523_ = new_n2521_ & new_n2522_;
  assign new_n2524_ = ~new_n2502_ & ~new_n2504_;
  assign new_n2525_ = ~new_n2493_ & ~new_n2497_;
  assign new_n2526_ = ~new_n2499_ & new_n2525_;
  assign new_n2527_ = new_n2524_ & new_n2526_;
  assign n1092 = ~new_n2523_ | ~new_n2527_;
  assign new_n2529_ = new_n1200_ & new_n2122_;
  assign new_n2530_ = ~pstart_0_ & new_n2529_;
  assign new_n2531_ = ~new_n1200_ & new_n2117_;
  assign new_n2532_ = ~pstart_0_ & new_n2531_;
  assign new_n2533_ = pkey_48_ & pencrypt_0_;
  assign new_n2534_ = pstart_0_ & new_n2533_;
  assign new_n2535_ = new_n1200_ & new_n2113_;
  assign new_n2536_ = ~pstart_0_ & new_n2535_;
  assign new_n2537_ = pkey_56_ & ~pencrypt_0_;
  assign new_n2538_ = pstart_0_ & new_n2537_;
  assign new_n2539_ = n_n2465 & new_n1220_;
  assign new_n2540_ = pencrypt_0_ & new_n2539_;
  assign new_n2541_ = ~n_n2372 & new_n2540_;
  assign new_n2542_ = ~pstart_0_ & new_n2541_;
  assign new_n2543_ = ~n_n2465 & new_n1220_;
  assign new_n2544_ = pencrypt_0_ & new_n2543_;
  assign new_n2545_ = n_n2372 & new_n2544_;
  assign new_n2546_ = ~pstart_0_ & new_n2545_;
  assign new_n2547_ = ~new_n1200_ & new_n2136_;
  assign new_n2548_ = ~pstart_0_ & new_n2547_;
  assign new_n2549_ = n_n2465 & ~new_n1220_;
  assign new_n2550_ = pencrypt_0_ & new_n2549_;
  assign new_n2551_ = n_n2372 & new_n2550_;
  assign new_n2552_ = ~pstart_0_ & new_n2551_;
  assign new_n2553_ = ~new_n2548_ & ~new_n2552_;
  assign new_n2554_ = ~new_n2542_ & ~new_n2546_;
  assign new_n2555_ = new_n2553_ & new_n2554_;
  assign new_n2556_ = ~new_n2536_ & ~new_n2538_;
  assign new_n2557_ = ~new_n2530_ & ~new_n2532_;
  assign new_n2558_ = ~new_n2534_ & new_n2557_;
  assign new_n2559_ = new_n2556_ & new_n2558_;
  assign n1097 = ~new_n2555_ | ~new_n2559_;
  assign new_n2561_ = ~pencrypt_0_ & n_n2746;
  assign new_n2562_ = ~new_n1200_ & new_n2561_;
  assign new_n2563_ = ~pstart_0_ & new_n2562_;
  assign new_n2564_ = n_n2382 & n_n2746;
  assign new_n2565_ = ~pencrypt_0_ & new_n2564_;
  assign new_n2566_ = new_n1200_ & new_n2565_;
  assign new_n2567_ = ~pstart_0_ & new_n2566_;
  assign new_n2568_ = pencrypt_0_ & pkey_172_;
  assign new_n2569_ = pstart_0_ & new_n2568_;
  assign new_n2570_ = ~pencrypt_0_ & n_n2382;
  assign new_n2571_ = ~new_n1200_ & new_n2570_;
  assign new_n2572_ = ~pstart_0_ & new_n2571_;
  assign new_n2573_ = pkey_244_ & ~pencrypt_0_;
  assign new_n2574_ = pstart_0_ & new_n2573_;
  assign new_n2575_ = ~n_n2746 & ~new_n1220_;
  assign new_n2576_ = pencrypt_0_ & new_n2575_;
  assign new_n2577_ = n_n2382 & new_n2576_;
  assign new_n2578_ = ~pstart_0_ & new_n2577_;
  assign new_n2579_ = n_n2746 & new_n1220_;
  assign new_n2580_ = pencrypt_0_ & new_n2579_;
  assign new_n2581_ = n_n2382 & new_n2580_;
  assign new_n2582_ = ~pstart_0_ & new_n2581_;
  assign new_n2583_ = ~n_n2382 & ~n_n2746;
  assign new_n2584_ = ~pencrypt_0_ & new_n2583_;
  assign new_n2585_ = new_n1200_ & new_n2584_;
  assign new_n2586_ = ~pstart_0_ & new_n2585_;
  assign new_n2587_ = n_n2746 & ~new_n1220_;
  assign new_n2588_ = pencrypt_0_ & new_n2587_;
  assign new_n2589_ = ~n_n2382 & new_n2588_;
  assign new_n2590_ = ~pstart_0_ & new_n2589_;
  assign new_n2591_ = ~new_n2586_ & ~new_n2590_;
  assign new_n2592_ = ~new_n2578_ & ~new_n2582_;
  assign new_n2593_ = new_n2591_ & new_n2592_;
  assign new_n2594_ = ~new_n2572_ & ~new_n2574_;
  assign new_n2595_ = ~new_n2563_ & ~new_n2567_;
  assign new_n2596_ = ~new_n2569_ & new_n2595_;
  assign new_n2597_ = new_n2594_ & new_n2596_;
  assign n1102 = ~new_n2593_ | ~new_n2597_;
  assign new_n2599_ = ~pencrypt_0_ & n_n2294;
  assign new_n2600_ = ~new_n1200_ & new_n2599_;
  assign new_n2601_ = ~pstart_0_ & new_n2600_;
  assign new_n2602_ = n_n2889 & n_n2294;
  assign new_n2603_ = ~pencrypt_0_ & new_n2602_;
  assign new_n2604_ = new_n1200_ & new_n2603_;
  assign new_n2605_ = ~pstart_0_ & new_n2604_;
  assign new_n2606_ = pencrypt_0_ & pkey_198_;
  assign new_n2607_ = pstart_0_ & new_n2606_;
  assign new_n2608_ = ~pencrypt_0_ & n_n2889;
  assign new_n2609_ = ~new_n1200_ & new_n2608_;
  assign new_n2610_ = ~pstart_0_ & new_n2609_;
  assign new_n2611_ = pkey_206_ & ~pencrypt_0_;
  assign new_n2612_ = pstart_0_ & new_n2611_;
  assign new_n2613_ = ~n_n2294 & ~new_n1220_;
  assign new_n2614_ = pencrypt_0_ & new_n2613_;
  assign new_n2615_ = n_n2889 & new_n2614_;
  assign new_n2616_ = ~pstart_0_ & new_n2615_;
  assign new_n2617_ = n_n2294 & new_n1220_;
  assign new_n2618_ = pencrypt_0_ & new_n2617_;
  assign new_n2619_ = n_n2889 & new_n2618_;
  assign new_n2620_ = ~pstart_0_ & new_n2619_;
  assign new_n2621_ = ~n_n2889 & ~n_n2294;
  assign new_n2622_ = ~pencrypt_0_ & new_n2621_;
  assign new_n2623_ = new_n1200_ & new_n2622_;
  assign new_n2624_ = ~pstart_0_ & new_n2623_;
  assign new_n2625_ = n_n2294 & ~new_n1220_;
  assign new_n2626_ = pencrypt_0_ & new_n2625_;
  assign new_n2627_ = ~n_n2889 & new_n2626_;
  assign new_n2628_ = ~pstart_0_ & new_n2627_;
  assign new_n2629_ = ~new_n2624_ & ~new_n2628_;
  assign new_n2630_ = ~new_n2616_ & ~new_n2620_;
  assign new_n2631_ = new_n2629_ & new_n2630_;
  assign new_n2632_ = ~new_n2610_ & ~new_n2612_;
  assign new_n2633_ = ~new_n2601_ & ~new_n2605_;
  assign new_n2634_ = ~new_n2607_ & new_n2633_;
  assign new_n2635_ = new_n2632_ & new_n2634_;
  assign n1107 = ~new_n2631_ | ~new_n2635_;
  assign new_n2637_ = ~pencrypt_0_ & n_n2341;
  assign new_n2638_ = ~new_n1200_ & new_n2637_;
  assign new_n2639_ = ~pstart_0_ & new_n2638_;
  assign new_n2640_ = n_n2435 & n_n2341;
  assign new_n2641_ = ~pencrypt_0_ & new_n2640_;
  assign new_n2642_ = new_n1200_ & new_n2641_;
  assign new_n2643_ = ~pstart_0_ & new_n2642_;
  assign new_n2644_ = pkey_125_ & pencrypt_0_;
  assign new_n2645_ = pstart_0_ & new_n2644_;
  assign new_n2646_ = ~pencrypt_0_ & n_n2435;
  assign new_n2647_ = ~new_n1200_ & new_n2646_;
  assign new_n2648_ = ~pstart_0_ & new_n2647_;
  assign new_n2649_ = pkey_70_ & ~pencrypt_0_;
  assign new_n2650_ = pstart_0_ & new_n2649_;
  assign new_n2651_ = ~n_n2341 & ~new_n1220_;
  assign new_n2652_ = pencrypt_0_ & new_n2651_;
  assign new_n2653_ = n_n2435 & new_n2652_;
  assign new_n2654_ = ~pstart_0_ & new_n2653_;
  assign new_n2655_ = n_n2341 & new_n1220_;
  assign new_n2656_ = pencrypt_0_ & new_n2655_;
  assign new_n2657_ = n_n2435 & new_n2656_;
  assign new_n2658_ = ~pstart_0_ & new_n2657_;
  assign new_n2659_ = ~n_n2435 & ~n_n2341;
  assign new_n2660_ = ~pencrypt_0_ & new_n2659_;
  assign new_n2661_ = new_n1200_ & new_n2660_;
  assign new_n2662_ = ~pstart_0_ & new_n2661_;
  assign new_n2663_ = n_n2341 & ~new_n1220_;
  assign new_n2664_ = pencrypt_0_ & new_n2663_;
  assign new_n2665_ = ~n_n2435 & new_n2664_;
  assign new_n2666_ = ~pstart_0_ & new_n2665_;
  assign new_n2667_ = ~new_n2662_ & ~new_n2666_;
  assign new_n2668_ = ~new_n2654_ & ~new_n2658_;
  assign new_n2669_ = new_n2667_ & new_n2668_;
  assign new_n2670_ = ~new_n2648_ & ~new_n2650_;
  assign new_n2671_ = ~new_n2639_ & ~new_n2643_;
  assign new_n2672_ = ~new_n2645_ & new_n2671_;
  assign new_n2673_ = new_n2670_ & new_n2672_;
  assign n1112 = ~new_n2669_ | ~new_n2673_;
  assign new_n2675_ = ~pencrypt_0_ & n_n2834;
  assign new_n2676_ = ~new_n1200_ & new_n2675_;
  assign new_n2677_ = ~pstart_0_ & new_n2676_;
  assign new_n2678_ = n_n2444 & n_n2834;
  assign new_n2679_ = ~pencrypt_0_ & new_n2678_;
  assign new_n2680_ = new_n1200_ & new_n2679_;
  assign new_n2681_ = ~pstart_0_ & new_n2680_;
  assign new_n2682_ = pkey_19_ & pencrypt_0_;
  assign new_n2683_ = pstart_0_ & new_n2682_;
  assign new_n2684_ = ~pencrypt_0_ & n_n2444;
  assign new_n2685_ = ~new_n1200_ & new_n2684_;
  assign new_n2686_ = ~pstart_0_ & new_n2685_;
  assign new_n2687_ = pkey_27_ & ~pencrypt_0_;
  assign new_n2688_ = pstart_0_ & new_n2687_;
  assign new_n2689_ = ~n_n2834 & ~new_n1220_;
  assign new_n2690_ = pencrypt_0_ & new_n2689_;
  assign new_n2691_ = n_n2444 & new_n2690_;
  assign new_n2692_ = ~pstart_0_ & new_n2691_;
  assign new_n2693_ = n_n2834 & new_n1220_;
  assign new_n2694_ = pencrypt_0_ & new_n2693_;
  assign new_n2695_ = n_n2444 & new_n2694_;
  assign new_n2696_ = ~pstart_0_ & new_n2695_;
  assign new_n2697_ = ~n_n2444 & ~n_n2834;
  assign new_n2698_ = ~pencrypt_0_ & new_n2697_;
  assign new_n2699_ = new_n1200_ & new_n2698_;
  assign new_n2700_ = ~pstart_0_ & new_n2699_;
  assign new_n2701_ = n_n2834 & ~new_n1220_;
  assign new_n2702_ = pencrypt_0_ & new_n2701_;
  assign new_n2703_ = ~n_n2444 & new_n2702_;
  assign new_n2704_ = ~pstart_0_ & new_n2703_;
  assign new_n2705_ = ~new_n2700_ & ~new_n2704_;
  assign new_n2706_ = ~new_n2692_ & ~new_n2696_;
  assign new_n2707_ = new_n2705_ & new_n2706_;
  assign new_n2708_ = ~new_n2686_ & ~new_n2688_;
  assign new_n2709_ = ~new_n2677_ & ~new_n2681_;
  assign new_n2710_ = ~new_n2683_ & new_n2709_;
  assign new_n2711_ = new_n2708_ & new_n2710_;
  assign n1117 = ~new_n2707_ | ~new_n2711_;
  assign new_n2713_ = ~pencrypt_0_ & n_n2360;
  assign new_n2714_ = ~new_n1200_ & new_n2713_;
  assign new_n2715_ = ~pstart_0_ & new_n2714_;
  assign new_n2716_ = n_n2454 & n_n2360;
  assign new_n2717_ = ~pencrypt_0_ & new_n2716_;
  assign new_n2718_ = new_n1200_ & new_n2717_;
  assign new_n2719_ = ~pstart_0_ & new_n2718_;
  assign new_n2720_ = pencrypt_0_ & pkey_13_;
  assign new_n2721_ = pstart_0_ & new_n2720_;
  assign new_n2722_ = ~pencrypt_0_ & n_n2454;
  assign new_n2723_ = ~new_n1200_ & new_n2722_;
  assign new_n2724_ = ~pstart_0_ & new_n2723_;
  assign new_n2725_ = ~pencrypt_0_ & pkey_21_;
  assign new_n2726_ = pstart_0_ & new_n2725_;
  assign new_n2727_ = ~n_n2360 & ~new_n1220_;
  assign new_n2728_ = pencrypt_0_ & new_n2727_;
  assign new_n2729_ = n_n2454 & new_n2728_;
  assign new_n2730_ = ~pstart_0_ & new_n2729_;
  assign new_n2731_ = n_n2360 & new_n1220_;
  assign new_n2732_ = pencrypt_0_ & new_n2731_;
  assign new_n2733_ = n_n2454 & new_n2732_;
  assign new_n2734_ = ~pstart_0_ & new_n2733_;
  assign new_n2735_ = ~n_n2454 & ~n_n2360;
  assign new_n2736_ = ~pencrypt_0_ & new_n2735_;
  assign new_n2737_ = new_n1200_ & new_n2736_;
  assign new_n2738_ = ~pstart_0_ & new_n2737_;
  assign new_n2739_ = n_n2360 & ~new_n1220_;
  assign new_n2740_ = pencrypt_0_ & new_n2739_;
  assign new_n2741_ = ~n_n2454 & new_n2740_;
  assign new_n2742_ = ~pstart_0_ & new_n2741_;
  assign new_n2743_ = ~new_n2738_ & ~new_n2742_;
  assign new_n2744_ = ~new_n2730_ & ~new_n2734_;
  assign new_n2745_ = new_n2743_ & new_n2744_;
  assign new_n2746_ = ~new_n2724_ & ~new_n2726_;
  assign new_n2747_ = ~new_n2715_ & ~new_n2719_;
  assign new_n2748_ = ~new_n2721_ & new_n2747_;
  assign new_n2749_ = new_n2746_ & new_n2748_;
  assign n1122 = ~new_n2745_ | ~new_n2749_;
  assign new_n2751_ = ~pencrypt_0_ & n_n2370;
  assign new_n2752_ = ~new_n1200_ & new_n2751_;
  assign new_n2753_ = ~pstart_0_ & new_n2752_;
  assign new_n2754_ = n_n2463 & n_n2370;
  assign new_n2755_ = ~pencrypt_0_ & new_n2754_;
  assign new_n2756_ = new_n1200_ & new_n2755_;
  assign new_n2757_ = ~pstart_0_ & new_n2756_;
  assign new_n2758_ = pkey_38_ & pencrypt_0_;
  assign new_n2759_ = pstart_0_ & new_n2758_;
  assign new_n2760_ = ~pencrypt_0_ & n_n2463;
  assign new_n2761_ = ~new_n1200_ & new_n2760_;
  assign new_n2762_ = ~pstart_0_ & new_n2761_;
  assign new_n2763_ = pkey_46_ & ~pencrypt_0_;
  assign new_n2764_ = pstart_0_ & new_n2763_;
  assign new_n2765_ = ~n_n2370 & ~new_n1220_;
  assign new_n2766_ = pencrypt_0_ & new_n2765_;
  assign new_n2767_ = n_n2463 & new_n2766_;
  assign new_n2768_ = ~pstart_0_ & new_n2767_;
  assign new_n2769_ = n_n2370 & new_n1220_;
  assign new_n2770_ = pencrypt_0_ & new_n2769_;
  assign new_n2771_ = n_n2463 & new_n2770_;
  assign new_n2772_ = ~pstart_0_ & new_n2771_;
  assign new_n2773_ = ~n_n2463 & ~n_n2370;
  assign new_n2774_ = ~pencrypt_0_ & new_n2773_;
  assign new_n2775_ = new_n1200_ & new_n2774_;
  assign new_n2776_ = ~pstart_0_ & new_n2775_;
  assign new_n2777_ = n_n2370 & ~new_n1220_;
  assign new_n2778_ = pencrypt_0_ & new_n2777_;
  assign new_n2779_ = ~n_n2463 & new_n2778_;
  assign new_n2780_ = ~pstart_0_ & new_n2779_;
  assign new_n2781_ = ~new_n2776_ & ~new_n2780_;
  assign new_n2782_ = ~new_n2768_ & ~new_n2772_;
  assign new_n2783_ = new_n2781_ & new_n2782_;
  assign new_n2784_ = ~new_n2762_ & ~new_n2764_;
  assign new_n2785_ = ~new_n2753_ & ~new_n2757_;
  assign new_n2786_ = ~new_n2759_ & new_n2785_;
  assign new_n2787_ = new_n2784_ & new_n2786_;
  assign n1127 = ~new_n2783_ | ~new_n2787_;
  assign new_n2789_ = new_n1200_ & new_n1786_;
  assign new_n2790_ = ~pstart_0_ & new_n2789_;
  assign new_n2791_ = ~new_n1200_ & new_n1781_;
  assign new_n2792_ = ~pstart_0_ & new_n2791_;
  assign new_n2793_ = pencrypt_0_ & pkey_33_;
  assign new_n2794_ = pstart_0_ & new_n2793_;
  assign new_n2795_ = new_n1200_ & new_n1777_1_;
  assign new_n2796_ = ~pstart_0_ & new_n2795_;
  assign new_n2797_ = ~pencrypt_0_ & pkey_41_;
  assign new_n2798_ = pstart_0_ & new_n2797_;
  assign new_n2799_ = n_n2457 & new_n1220_;
  assign new_n2800_ = pencrypt_0_ & new_n2799_;
  assign new_n2801_ = ~n_n2363 & new_n2800_;
  assign new_n2802_ = ~pstart_0_ & new_n2801_;
  assign new_n2803_ = ~n_n2457 & new_n1220_;
  assign new_n2804_ = pencrypt_0_ & new_n2803_;
  assign new_n2805_ = n_n2363 & new_n2804_;
  assign new_n2806_ = ~pstart_0_ & new_n2805_;
  assign new_n2807_ = ~new_n1200_ & new_n1800_;
  assign new_n2808_ = ~pstart_0_ & new_n2807_;
  assign new_n2809_ = n_n2457 & ~new_n1220_;
  assign new_n2810_ = pencrypt_0_ & new_n2809_;
  assign new_n2811_ = n_n2363 & new_n2810_;
  assign new_n2812_ = ~pstart_0_ & new_n2811_;
  assign new_n2813_ = ~new_n2808_ & ~new_n2812_;
  assign new_n2814_ = ~new_n2802_ & ~new_n2806_;
  assign new_n2815_ = new_n2813_ & new_n2814_;
  assign new_n2816_ = ~new_n2796_ & ~new_n2798_;
  assign new_n2817_ = ~new_n2790_ & ~new_n2792_;
  assign new_n2818_ = ~new_n2794_ & new_n2817_;
  assign new_n2819_ = new_n2816_ & new_n2818_;
  assign n1132 = ~new_n2815_ | ~new_n2819_;
  assign new_n2821_ = ~pencrypt_0_ & n_n2464;
  assign new_n2822_ = new_n1200_ & new_n2821_;
  assign new_n2823_ = ~pstart_0_ & new_n2822_;
  assign new_n2824_ = n_n2371 & n_n2464;
  assign new_n2825_ = ~pencrypt_0_ & new_n2824_;
  assign new_n2826_ = ~new_n1200_ & new_n2825_;
  assign new_n2827_ = ~pstart_0_ & new_n2826_;
  assign new_n2828_ = pencrypt_0_ & pkey_40_;
  assign new_n2829_ = pstart_0_ & new_n2828_;
  assign new_n2830_ = ~pencrypt_0_ & n_n2371;
  assign new_n2831_ = new_n1200_ & new_n2830_;
  assign new_n2832_ = ~pstart_0_ & new_n2831_;
  assign new_n2833_ = pkey_48_ & ~pencrypt_0_;
  assign new_n2834_ = pstart_0_ & new_n2833_;
  assign new_n2835_ = n_n2464 & new_n1220_;
  assign new_n2836_ = pencrypt_0_ & new_n2835_;
  assign new_n2837_ = ~n_n2371 & new_n2836_;
  assign new_n2838_ = ~pstart_0_ & new_n2837_;
  assign new_n2839_ = ~n_n2464 & new_n1220_;
  assign new_n2840_ = pencrypt_0_ & new_n2839_;
  assign new_n2841_ = n_n2371 & new_n2840_;
  assign new_n2842_ = ~pstart_0_ & new_n2841_;
  assign new_n2843_ = ~n_n2371 & ~n_n2464;
  assign new_n2844_ = ~pencrypt_0_ & new_n2843_;
  assign new_n2845_ = ~new_n1200_ & new_n2844_;
  assign new_n2846_ = ~pstart_0_ & new_n2845_;
  assign new_n2847_ = n_n2464 & ~new_n1220_;
  assign new_n2848_ = pencrypt_0_ & new_n2847_;
  assign new_n2849_ = n_n2371 & new_n2848_;
  assign new_n2850_ = ~pstart_0_ & new_n2849_;
  assign new_n2851_ = ~new_n2846_ & ~new_n2850_;
  assign new_n2852_ = ~new_n2838_ & ~new_n2842_;
  assign new_n2853_ = new_n2851_ & new_n2852_;
  assign new_n2854_ = ~new_n2832_ & ~new_n2834_;
  assign new_n2855_ = ~new_n2823_ & ~new_n2827_;
  assign new_n2856_ = ~new_n2829_ & new_n2855_;
  assign new_n2857_ = new_n2854_ & new_n2856_;
  assign n1137 = ~new_n2853_ | ~new_n2857_;
  assign new_n2859_ = ~pencrypt_0_ & n_n2286;
  assign new_n2860_ = ~new_n1200_ & new_n2859_;
  assign new_n2861_ = ~pstart_0_ & new_n2860_;
  assign new_n2862_ = n_n2383 & n_n2286;
  assign new_n2863_ = ~pencrypt_0_ & new_n2862_;
  assign new_n2864_ = new_n1200_ & new_n2863_;
  assign new_n2865_ = ~pstart_0_ & new_n2864_;
  assign new_n2866_ = pkey_244_ & pencrypt_0_;
  assign new_n2867_ = pstart_0_ & new_n2866_;
  assign new_n2868_ = ~pencrypt_0_ & n_n2383;
  assign new_n2869_ = ~new_n1200_ & new_n2868_;
  assign new_n2870_ = ~pstart_0_ & new_n2869_;
  assign new_n2871_ = pkey_252_ & ~pencrypt_0_;
  assign new_n2872_ = pstart_0_ & new_n2871_;
  assign new_n2873_ = ~n_n2286 & ~new_n1220_;
  assign new_n2874_ = pencrypt_0_ & new_n2873_;
  assign new_n2875_ = n_n2383 & new_n2874_;
  assign new_n2876_ = ~pstart_0_ & new_n2875_;
  assign new_n2877_ = n_n2286 & new_n1220_;
  assign new_n2878_ = pencrypt_0_ & new_n2877_;
  assign new_n2879_ = n_n2383 & new_n2878_;
  assign new_n2880_ = ~pstart_0_ & new_n2879_;
  assign new_n2881_ = ~n_n2383 & ~n_n2286;
  assign new_n2882_ = ~pencrypt_0_ & new_n2881_;
  assign new_n2883_ = new_n1200_ & new_n2882_;
  assign new_n2884_ = ~pstart_0_ & new_n2883_;
  assign new_n2885_ = n_n2286 & ~new_n1220_;
  assign new_n2886_ = pencrypt_0_ & new_n2885_;
  assign new_n2887_ = ~n_n2383 & new_n2886_;
  assign new_n2888_ = ~pstart_0_ & new_n2887_;
  assign new_n2889_ = ~new_n2884_ & ~new_n2888_;
  assign new_n2890_ = ~new_n2876_ & ~new_n2880_;
  assign new_n2891_ = new_n2889_ & new_n2890_;
  assign new_n2892_ = ~new_n2870_ & ~new_n2872_;
  assign new_n2893_ = ~new_n2861_ & ~new_n2865_;
  assign new_n2894_ = ~new_n2867_ & new_n2893_;
  assign new_n2895_ = new_n2892_ & new_n2894_;
  assign n1142 = ~new_n2891_ | ~new_n2895_;
  assign new_n2897_ = ~pencrypt_0_ & n_n2293;
  assign new_n2898_ = ~new_n1200_ & new_n2897_;
  assign new_n2899_ = ~pstart_0_ & new_n2898_;
  assign new_n2900_ = n_n2388 & n_n2293;
  assign new_n2901_ = ~pencrypt_0_ & new_n2900_;
  assign new_n2902_ = new_n1200_ & new_n2901_;
  assign new_n2903_ = ~pstart_0_ & new_n2902_;
  assign new_n2904_ = pkey_253_ & pencrypt_0_;
  assign new_n2905_ = pstart_0_ & new_n2904_;
  assign new_n2906_ = ~pencrypt_0_ & n_n2388;
  assign new_n2907_ = ~new_n1200_ & new_n2906_;
  assign new_n2908_ = ~pstart_0_ & new_n2907_;
  assign new_n2909_ = ~pencrypt_0_ & pkey_198_;
  assign new_n2910_ = pstart_0_ & new_n2909_;
  assign new_n2911_ = ~n_n2293 & ~new_n1220_;
  assign new_n2912_ = pencrypt_0_ & new_n2911_;
  assign new_n2913_ = n_n2388 & new_n2912_;
  assign new_n2914_ = ~pstart_0_ & new_n2913_;
  assign new_n2915_ = n_n2293 & new_n1220_;
  assign new_n2916_ = pencrypt_0_ & new_n2915_;
  assign new_n2917_ = n_n2388 & new_n2916_;
  assign new_n2918_ = ~pstart_0_ & new_n2917_;
  assign new_n2919_ = ~n_n2388 & ~n_n2293;
  assign new_n2920_ = ~pencrypt_0_ & new_n2919_;
  assign new_n2921_ = new_n1200_ & new_n2920_;
  assign new_n2922_ = ~pstart_0_ & new_n2921_;
  assign new_n2923_ = n_n2293 & ~new_n1220_;
  assign new_n2924_ = pencrypt_0_ & new_n2923_;
  assign new_n2925_ = ~n_n2388 & new_n2924_;
  assign new_n2926_ = ~pstart_0_ & new_n2925_;
  assign new_n2927_ = ~new_n2922_ & ~new_n2926_;
  assign new_n2928_ = ~new_n2914_ & ~new_n2918_;
  assign new_n2929_ = new_n2927_ & new_n2928_;
  assign new_n2930_ = ~new_n2908_ & ~new_n2910_;
  assign new_n2931_ = ~new_n2899_ & ~new_n2903_;
  assign new_n2932_ = ~new_n2905_ & new_n2931_;
  assign new_n2933_ = new_n2930_ & new_n2932_;
  assign n1147 = ~new_n2929_ | ~new_n2933_;
  assign new_n2935_ = ~pencrypt_0_ & n_n2342;
  assign new_n2936_ = ~new_n1200_ & new_n2935_;
  assign new_n2937_ = ~pstart_0_ & new_n2936_;
  assign new_n2938_ = n_n2954 & n_n2342;
  assign new_n2939_ = ~pencrypt_0_ & new_n2938_;
  assign new_n2940_ = new_n1200_ & new_n2939_;
  assign new_n2941_ = ~pstart_0_ & new_n2940_;
  assign new_n2942_ = pkey_70_ & pencrypt_0_;
  assign new_n2943_ = pstart_0_ & new_n2942_;
  assign new_n2944_ = ~pencrypt_0_ & n_n2954;
  assign new_n2945_ = ~new_n1200_ & new_n2944_;
  assign new_n2946_ = ~pstart_0_ & new_n2945_;
  assign new_n2947_ = pkey_78_ & ~pencrypt_0_;
  assign new_n2948_ = pstart_0_ & new_n2947_;
  assign new_n2949_ = ~n_n2342 & ~new_n1220_;
  assign new_n2950_ = pencrypt_0_ & new_n2949_;
  assign new_n2951_ = n_n2954 & new_n2950_;
  assign new_n2952_ = ~pstart_0_ & new_n2951_;
  assign new_n2953_ = n_n2342 & new_n1220_;
  assign new_n2954_ = pencrypt_0_ & new_n2953_;
  assign new_n2955_ = n_n2954 & new_n2954_;
  assign new_n2956_ = ~pstart_0_ & new_n2955_;
  assign new_n2957_ = ~n_n2954 & ~n_n2342;
  assign new_n2958_ = ~pencrypt_0_ & new_n2957_;
  assign new_n2959_ = new_n1200_ & new_n2958_;
  assign new_n2960_ = ~pstart_0_ & new_n2959_;
  assign new_n2961_ = n_n2342 & ~new_n1220_;
  assign new_n2962_ = pencrypt_0_ & new_n2961_;
  assign new_n2963_ = ~n_n2954 & new_n2962_;
  assign new_n2964_ = ~pstart_0_ & new_n2963_;
  assign new_n2965_ = ~new_n2960_ & ~new_n2964_;
  assign new_n2966_ = ~new_n2952_ & ~new_n2956_;
  assign new_n2967_ = new_n2965_ & new_n2966_;
  assign new_n2968_ = ~new_n2946_ & ~new_n2948_;
  assign new_n2969_ = ~new_n2937_ & ~new_n2941_;
  assign new_n2970_ = ~new_n2943_ & new_n2969_;
  assign new_n2971_ = new_n2968_ & new_n2970_;
  assign n1152 = ~new_n2967_ | ~new_n2971_;
  assign new_n2973_ = ~pencrypt_0_ & n_n2351;
  assign new_n2974_ = ~new_n1200_ & new_n2973_;
  assign new_n2975_ = ~pstart_0_ & new_n2974_;
  assign new_n2976_ = n_n2964 & n_n2351;
  assign new_n2977_ = ~pencrypt_0_ & new_n2976_;
  assign new_n2978_ = new_n1200_ & new_n2977_;
  assign new_n2979_ = ~pstart_0_ & new_n2978_;
  assign new_n2980_ = pencrypt_0_ & pkey_11_;
  assign new_n2981_ = pstart_0_ & new_n2980_;
  assign new_n2982_ = ~pencrypt_0_ & n_n2964;
  assign new_n2983_ = ~new_n1200_ & new_n2982_;
  assign new_n2984_ = ~pstart_0_ & new_n2983_;
  assign new_n2985_ = pkey_19_ & ~pencrypt_0_;
  assign new_n2986_ = pstart_0_ & new_n2985_;
  assign new_n2987_ = ~n_n2351 & ~new_n1220_;
  assign new_n2988_ = pencrypt_0_ & new_n2987_;
  assign new_n2989_ = n_n2964 & new_n2988_;
  assign new_n2990_ = ~pstart_0_ & new_n2989_;
  assign new_n2991_ = n_n2351 & new_n1220_;
  assign new_n2992_ = pencrypt_0_ & new_n2991_;
  assign new_n2993_ = n_n2964 & new_n2992_;
  assign new_n2994_ = ~pstart_0_ & new_n2993_;
  assign new_n2995_ = ~n_n2964 & ~n_n2351;
  assign new_n2996_ = ~pencrypt_0_ & new_n2995_;
  assign new_n2997_ = new_n1200_ & new_n2996_;
  assign new_n2998_ = ~pstart_0_ & new_n2997_;
  assign new_n2999_ = n_n2351 & ~new_n1220_;
  assign new_n3000_ = pencrypt_0_ & new_n2999_;
  assign new_n3001_ = ~n_n2964 & new_n3000_;
  assign new_n3002_ = ~pstart_0_ & new_n3001_;
  assign new_n3003_ = ~new_n2998_ & ~new_n3002_;
  assign new_n3004_ = ~new_n2990_ & ~new_n2994_;
  assign new_n3005_ = new_n3003_ & new_n3004_;
  assign new_n3006_ = ~new_n2984_ & ~new_n2986_;
  assign new_n3007_ = ~new_n2975_ & ~new_n2979_;
  assign new_n3008_ = ~new_n2981_ & new_n3007_;
  assign new_n3009_ = new_n3006_ & new_n3008_;
  assign n1157 = ~new_n3005_ | ~new_n3009_;
  assign new_n3011_ = ~pencrypt_0_ & n_n2352;
  assign new_n3012_ = ~new_n1200_ & new_n3011_;
  assign new_n3013_ = ~pstart_0_ & new_n3012_;
  assign new_n3014_ = n_n2445 & n_n2352;
  assign new_n3015_ = ~pencrypt_0_ & new_n3014_;
  assign new_n3016_ = new_n1200_ & new_n3015_;
  assign new_n3017_ = ~pstart_0_ & new_n3016_;
  assign new_n3018_ = pkey_27_ & pencrypt_0_;
  assign new_n3019_ = pstart_0_ & new_n3018_;
  assign new_n3020_ = ~pencrypt_0_ & n_n2445;
  assign new_n3021_ = ~new_n1200_ & new_n3020_;
  assign new_n3022_ = ~pstart_0_ & new_n3021_;
  assign new_n3023_ = pkey_4_ & ~pencrypt_0_;
  assign new_n3024_ = pstart_0_ & new_n3023_;
  assign new_n3025_ = ~n_n2352 & ~new_n1220_;
  assign new_n3026_ = pencrypt_0_ & new_n3025_;
  assign new_n3027_ = n_n2445 & new_n3026_;
  assign new_n3028_ = ~pstart_0_ & new_n3027_;
  assign new_n3029_ = n_n2352 & new_n1220_;
  assign new_n3030_ = pencrypt_0_ & new_n3029_;
  assign new_n3031_ = n_n2445 & new_n3030_;
  assign new_n3032_ = ~pstart_0_ & new_n3031_;
  assign new_n3033_ = ~n_n2445 & ~n_n2352;
  assign new_n3034_ = ~pencrypt_0_ & new_n3033_;
  assign new_n3035_ = new_n1200_ & new_n3034_;
  assign new_n3036_ = ~pstart_0_ & new_n3035_;
  assign new_n3037_ = n_n2352 & ~new_n1220_;
  assign new_n3038_ = pencrypt_0_ & new_n3037_;
  assign new_n3039_ = ~n_n2445 & new_n3038_;
  assign new_n3040_ = ~pstart_0_ & new_n3039_;
  assign new_n3041_ = ~new_n3036_ & ~new_n3040_;
  assign new_n3042_ = ~new_n3028_ & ~new_n3032_;
  assign new_n3043_ = new_n3041_ & new_n3042_;
  assign new_n3044_ = ~new_n3022_ & ~new_n3024_;
  assign new_n3045_ = ~new_n3013_ & ~new_n3017_;
  assign new_n3046_ = ~new_n3019_ & new_n3045_;
  assign new_n3047_ = new_n3044_ & new_n3046_;
  assign n1162 = ~new_n3043_ | ~new_n3047_;
  assign new_n3049_ = ~new_n1200_ & new_n2830_;
  assign new_n3050_ = ~pstart_0_ & new_n3049_;
  assign new_n3051_ = new_n1200_ & new_n2825_;
  assign new_n3052_ = ~pstart_0_ & new_n3051_;
  assign new_n3053_ = pkey_46_ & pencrypt_0_;
  assign new_n3054_ = pstart_0_ & new_n3053_;
  assign new_n3055_ = ~new_n1200_ & new_n2821_;
  assign new_n3056_ = ~pstart_0_ & new_n3055_;
  assign new_n3057_ = ~pencrypt_0_ & pkey_54_;
  assign new_n3058_ = pstart_0_ & new_n3057_;
  assign new_n3059_ = ~n_n2371 & ~new_n1220_;
  assign new_n3060_ = pencrypt_0_ & new_n3059_;
  assign new_n3061_ = n_n2464 & new_n3060_;
  assign new_n3062_ = ~pstart_0_ & new_n3061_;
  assign new_n3063_ = n_n2371 & new_n1220_;
  assign new_n3064_ = pencrypt_0_ & new_n3063_;
  assign new_n3065_ = n_n2464 & new_n3064_;
  assign new_n3066_ = ~pstart_0_ & new_n3065_;
  assign new_n3067_ = new_n1200_ & new_n2844_;
  assign new_n3068_ = ~pstart_0_ & new_n3067_;
  assign new_n3069_ = n_n2371 & ~new_n1220_;
  assign new_n3070_ = pencrypt_0_ & new_n3069_;
  assign new_n3071_ = ~n_n2464 & new_n3070_;
  assign new_n3072_ = ~pstart_0_ & new_n3071_;
  assign new_n3073_ = ~new_n3068_ & ~new_n3072_;
  assign new_n3074_ = ~new_n3062_ & ~new_n3066_;
  assign new_n3075_ = new_n3073_ & new_n3074_;
  assign new_n3076_ = ~new_n3056_ & ~new_n3058_;
  assign new_n3077_ = ~new_n3050_ & ~new_n3052_;
  assign new_n3078_ = ~new_n3054_ & new_n3077_;
  assign new_n3079_ = new_n3076_ & new_n3078_;
  assign n1167 = ~new_n3075_ | ~new_n3079_;
  assign new_n3081_ = new_n1200_ & new_n1482_1_;
  assign new_n3082_ = ~pstart_0_ & new_n3081_;
  assign new_n3083_ = ~new_n1200_ & new_n1477_1_;
  assign new_n3084_ = ~pstart_0_ & new_n3083_;
  assign new_n3085_ = pencrypt_0_ & pkey_41_;
  assign new_n3086_ = pstart_0_ & new_n3085_;
  assign new_n3087_ = new_n1200_ & new_n1473_;
  assign new_n3088_ = ~pstart_0_ & new_n3087_;
  assign new_n3089_ = pkey_49_ & ~pencrypt_0_;
  assign new_n3090_ = pstart_0_ & new_n3089_;
  assign new_n3091_ = n_n2982 & new_n1220_;
  assign new_n3092_ = pencrypt_0_ & new_n3091_;
  assign new_n3093_ = ~n_n2364 & new_n3092_;
  assign new_n3094_ = ~pstart_0_ & new_n3093_;
  assign new_n3095_ = ~n_n2982 & new_n1220_;
  assign new_n3096_ = pencrypt_0_ & new_n3095_;
  assign new_n3097_ = n_n2364 & new_n3096_;
  assign new_n3098_ = ~pstart_0_ & new_n3097_;
  assign new_n3099_ = ~new_n1200_ & new_n1496_;
  assign new_n3100_ = ~pstart_0_ & new_n3099_;
  assign new_n3101_ = n_n2982 & ~new_n1220_;
  assign new_n3102_ = pencrypt_0_ & new_n3101_;
  assign new_n3103_ = n_n2364 & new_n3102_;
  assign new_n3104_ = ~pstart_0_ & new_n3103_;
  assign new_n3105_ = ~new_n3100_ & ~new_n3104_;
  assign new_n3106_ = ~new_n3094_ & ~new_n3098_;
  assign new_n3107_ = new_n3105_ & new_n3106_;
  assign new_n3108_ = ~new_n3088_ & ~new_n3090_;
  assign new_n3109_ = ~new_n3082_ & ~new_n3084_;
  assign new_n3110_ = ~new_n3086_ & new_n3109_;
  assign new_n3111_ = new_n3108_ & new_n3110_;
  assign n1172 = ~new_n3107_ | ~new_n3111_;
  assign new_n3113_ = ~pencrypt_0_ & n_n2279;
  assign new_n3114_ = ~new_n1200_ & new_n3113_;
  assign new_n3115_ = ~pstart_0_ & new_n3114_;
  assign new_n3116_ = n_n2374 & n_n2279;
  assign new_n3117_ = ~pencrypt_0_ & new_n3116_;
  assign new_n3118_ = new_n1200_ & new_n3117_;
  assign new_n3119_ = ~pstart_0_ & new_n3118_;
  assign new_n3120_ = pkey_195_ & pencrypt_0_;
  assign new_n3121_ = pstart_0_ & new_n3120_;
  assign new_n3122_ = ~pencrypt_0_ & n_n2374;
  assign new_n3123_ = ~new_n1200_ & new_n3122_;
  assign new_n3124_ = ~pstart_0_ & new_n3123_;
  assign new_n3125_ = pkey_203_ & ~pencrypt_0_;
  assign new_n3126_ = pstart_0_ & new_n3125_;
  assign new_n3127_ = ~n_n2279 & ~new_n1220_;
  assign new_n3128_ = pencrypt_0_ & new_n3127_;
  assign new_n3129_ = n_n2374 & new_n3128_;
  assign new_n3130_ = ~pstart_0_ & new_n3129_;
  assign new_n3131_ = n_n2279 & new_n1220_;
  assign new_n3132_ = pencrypt_0_ & new_n3131_;
  assign new_n3133_ = n_n2374 & new_n3132_;
  assign new_n3134_ = ~pstart_0_ & new_n3133_;
  assign new_n3135_ = ~n_n2374 & ~n_n2279;
  assign new_n3136_ = ~pencrypt_0_ & new_n3135_;
  assign new_n3137_ = new_n1200_ & new_n3136_;
  assign new_n3138_ = ~pstart_0_ & new_n3137_;
  assign new_n3139_ = n_n2279 & ~new_n1220_;
  assign new_n3140_ = pencrypt_0_ & new_n3139_;
  assign new_n3141_ = ~n_n2374 & new_n3140_;
  assign new_n3142_ = ~pstart_0_ & new_n3141_;
  assign new_n3143_ = ~new_n3138_ & ~new_n3142_;
  assign new_n3144_ = ~new_n3130_ & ~new_n3134_;
  assign new_n3145_ = new_n3143_ & new_n3144_;
  assign new_n3146_ = ~new_n3124_ & ~new_n3126_;
  assign new_n3147_ = ~new_n3115_ & ~new_n3119_;
  assign new_n3148_ = ~new_n3121_ & new_n3147_;
  assign new_n3149_ = new_n3146_ & new_n3148_;
  assign n1177 = ~new_n3145_ | ~new_n3149_;
  assign new_n3151_ = ~pencrypt_0_ & n_n2284;
  assign new_n3152_ = ~new_n1200_ & new_n3151_;
  assign new_n3153_ = ~pstart_0_ & new_n3152_;
  assign new_n3154_ = n_n2380 & n_n2284;
  assign new_n3155_ = ~pencrypt_0_ & new_n3154_;
  assign new_n3156_ = new_n1200_ & new_n3155_;
  assign new_n3157_ = ~pstart_0_ & new_n3156_;
  assign new_n3158_ = pkey_220_ & pencrypt_0_;
  assign new_n3159_ = pstart_0_ & new_n3158_;
  assign new_n3160_ = ~pencrypt_0_ & n_n2380;
  assign new_n3161_ = ~new_n1200_ & new_n3160_;
  assign new_n3162_ = ~pstart_0_ & new_n3161_;
  assign new_n3163_ = pkey_228_ & ~pencrypt_0_;
  assign new_n3164_ = pstart_0_ & new_n3163_;
  assign new_n3165_ = ~n_n2284 & ~new_n1220_;
  assign new_n3166_ = pencrypt_0_ & new_n3165_;
  assign new_n3167_ = n_n2380 & new_n3166_;
  assign new_n3168_ = ~pstart_0_ & new_n3167_;
  assign new_n3169_ = n_n2284 & new_n1220_;
  assign new_n3170_ = pencrypt_0_ & new_n3169_;
  assign new_n3171_ = n_n2380 & new_n3170_;
  assign new_n3172_ = ~pstart_0_ & new_n3171_;
  assign new_n3173_ = ~n_n2380 & ~n_n2284;
  assign new_n3174_ = ~pencrypt_0_ & new_n3173_;
  assign new_n3175_ = new_n1200_ & new_n3174_;
  assign new_n3176_ = ~pstart_0_ & new_n3175_;
  assign new_n3177_ = n_n2284 & ~new_n1220_;
  assign new_n3178_ = pencrypt_0_ & new_n3177_;
  assign new_n3179_ = ~n_n2380 & new_n3178_;
  assign new_n3180_ = ~pstart_0_ & new_n3179_;
  assign new_n3181_ = ~new_n3176_ & ~new_n3180_;
  assign new_n3182_ = ~new_n3168_ & ~new_n3172_;
  assign new_n3183_ = new_n3181_ & new_n3182_;
  assign new_n3184_ = ~new_n3162_ & ~new_n3164_;
  assign new_n3185_ = ~new_n3153_ & ~new_n3157_;
  assign new_n3186_ = ~new_n3159_ & new_n3185_;
  assign new_n3187_ = new_n3184_ & new_n3186_;
  assign n1182 = ~new_n3183_ | ~new_n3187_;
  assign new_n3189_ = ~pencrypt_0_ & n_n2757;
  assign new_n3190_ = ~new_n1200_ & new_n3189_;
  assign new_n3191_ = ~pstart_0_ & new_n3190_;
  assign new_n3192_ = n_n2387 & n_n2757;
  assign new_n3193_ = ~pencrypt_0_ & new_n3192_;
  assign new_n3194_ = new_n1200_ & new_n3193_;
  assign new_n3195_ = ~pstart_0_ & new_n3194_;
  assign new_n3196_ = pkey_245_ & pencrypt_0_;
  assign new_n3197_ = pstart_0_ & new_n3196_;
  assign new_n3198_ = ~pencrypt_0_ & n_n2387;
  assign new_n3199_ = ~new_n1200_ & new_n3198_;
  assign new_n3200_ = ~pstart_0_ & new_n3199_;
  assign new_n3201_ = pkey_253_ & ~pencrypt_0_;
  assign new_n3202_ = pstart_0_ & new_n3201_;
  assign new_n3203_ = ~n_n2757 & ~new_n1220_;
  assign new_n3204_ = pencrypt_0_ & new_n3203_;
  assign new_n3205_ = n_n2387 & new_n3204_;
  assign new_n3206_ = ~pstart_0_ & new_n3205_;
  assign new_n3207_ = n_n2757 & new_n1220_;
  assign new_n3208_ = pencrypt_0_ & new_n3207_;
  assign new_n3209_ = n_n2387 & new_n3208_;
  assign new_n3210_ = ~pstart_0_ & new_n3209_;
  assign new_n3211_ = ~n_n2387 & ~n_n2757;
  assign new_n3212_ = ~pencrypt_0_ & new_n3211_;
  assign new_n3213_ = new_n1200_ & new_n3212_;
  assign new_n3214_ = ~pstart_0_ & new_n3213_;
  assign new_n3215_ = n_n2757 & ~new_n1220_;
  assign new_n3216_ = pencrypt_0_ & new_n3215_;
  assign new_n3217_ = ~n_n2387 & new_n3216_;
  assign new_n3218_ = ~pstart_0_ & new_n3217_;
  assign new_n3219_ = ~new_n3214_ & ~new_n3218_;
  assign new_n3220_ = ~new_n3206_ & ~new_n3210_;
  assign new_n3221_ = new_n3219_ & new_n3220_;
  assign new_n3222_ = ~new_n3200_ & ~new_n3202_;
  assign new_n3223_ = ~new_n3191_ & ~new_n3195_;
  assign new_n3224_ = ~new_n3197_ & new_n3223_;
  assign new_n3225_ = new_n3222_ & new_n3224_;
  assign n1187 = ~new_n3221_ | ~new_n3225_;
  assign new_n3227_ = ~pencrypt_0_ & n_n2353;
  assign new_n3228_ = ~new_n1200_ & new_n3227_;
  assign new_n3229_ = ~pstart_0_ & new_n3228_;
  assign new_n3230_ = n_n2446 & n_n2353;
  assign new_n3231_ = ~pencrypt_0_ & new_n3230_;
  assign new_n3232_ = new_n1200_ & new_n3231_;
  assign new_n3233_ = ~pstart_0_ & new_n3232_;
  assign new_n3234_ = pkey_4_ & pencrypt_0_;
  assign new_n3235_ = pstart_0_ & new_n3234_;
  assign new_n3236_ = ~pencrypt_0_ & n_n2446;
  assign new_n3237_ = ~new_n1200_ & new_n3236_;
  assign new_n3238_ = ~pstart_0_ & new_n3237_;
  assign new_n3239_ = ~pencrypt_0_ & pkey_12_;
  assign new_n3240_ = pstart_0_ & new_n3239_;
  assign new_n3241_ = ~n_n2353 & ~new_n1220_;
  assign new_n3242_ = pencrypt_0_ & new_n3241_;
  assign new_n3243_ = n_n2446 & new_n3242_;
  assign new_n3244_ = ~pstart_0_ & new_n3243_;
  assign new_n3245_ = n_n2353 & new_n1220_;
  assign new_n3246_ = pencrypt_0_ & new_n3245_;
  assign new_n3247_ = n_n2446 & new_n3246_;
  assign new_n3248_ = ~pstart_0_ & new_n3247_;
  assign new_n3249_ = ~n_n2446 & ~n_n2353;
  assign new_n3250_ = ~pencrypt_0_ & new_n3249_;
  assign new_n3251_ = new_n1200_ & new_n3250_;
  assign new_n3252_ = ~pstart_0_ & new_n3251_;
  assign new_n3253_ = n_n2353 & ~new_n1220_;
  assign new_n3254_ = pencrypt_0_ & new_n3253_;
  assign new_n3255_ = ~n_n2446 & new_n3254_;
  assign new_n3256_ = ~pstart_0_ & new_n3255_;
  assign new_n3257_ = ~new_n3252_ & ~new_n3256_;
  assign new_n3258_ = ~new_n3244_ & ~new_n3248_;
  assign new_n3259_ = new_n3257_ & new_n3258_;
  assign new_n3260_ = ~new_n3238_ & ~new_n3240_;
  assign new_n3261_ = ~new_n3229_ & ~new_n3233_;
  assign new_n3262_ = ~new_n3235_ & new_n3261_;
  assign new_n3263_ = new_n3260_ & new_n3262_;
  assign n1192 = ~new_n3259_ | ~new_n3263_;
  assign new_n3265_ = ~new_n1200_ & new_n2500_;
  assign new_n3266_ = ~pstart_0_ & new_n3265_;
  assign new_n3267_ = new_n1200_ & new_n2495_;
  assign new_n3268_ = ~pstart_0_ & new_n3267_;
  assign new_n3269_ = pkey_29_ & pencrypt_0_;
  assign new_n3270_ = pstart_0_ & new_n3269_;
  assign new_n3271_ = ~new_n1200_ & new_n2491_;
  assign new_n3272_ = ~pstart_0_ & new_n3271_;
  assign new_n3273_ = pkey_37_ & ~pencrypt_0_;
  assign new_n3274_ = pstart_0_ & new_n3273_;
  assign new_n3275_ = ~n_n2362 & ~new_n1220_;
  assign new_n3276_ = pencrypt_0_ & new_n3275_;
  assign new_n3277_ = n_n2456 & new_n3276_;
  assign new_n3278_ = ~pstart_0_ & new_n3277_;
  assign new_n3279_ = n_n2362 & new_n1220_;
  assign new_n3280_ = pencrypt_0_ & new_n3279_;
  assign new_n3281_ = n_n2456 & new_n3280_;
  assign new_n3282_ = ~pstart_0_ & new_n3281_;
  assign new_n3283_ = new_n1200_ & new_n2514_;
  assign new_n3284_ = ~pstart_0_ & new_n3283_;
  assign new_n3285_ = n_n2362 & ~new_n1220_;
  assign new_n3286_ = pencrypt_0_ & new_n3285_;
  assign new_n3287_ = ~n_n2456 & new_n3286_;
  assign new_n3288_ = ~pstart_0_ & new_n3287_;
  assign new_n3289_ = ~new_n3284_ & ~new_n3288_;
  assign new_n3290_ = ~new_n3278_ & ~new_n3282_;
  assign new_n3291_ = new_n3289_ & new_n3290_;
  assign new_n3292_ = ~new_n3272_ & ~new_n3274_;
  assign new_n3293_ = ~new_n3266_ & ~new_n3268_;
  assign new_n3294_ = ~new_n3270_ & new_n3293_;
  assign new_n3295_ = new_n3292_ & new_n3294_;
  assign n1197 = ~new_n3291_ | ~new_n3295_;
  assign new_n3297_ = new_n1200_ & new_n2424_;
  assign new_n3298_ = ~pstart_0_ & new_n3297_;
  assign new_n3299_ = ~new_n1200_ & new_n2419_;
  assign new_n3300_ = ~pstart_0_ & new_n3299_;
  assign new_n3301_ = pkey_49_ & pencrypt_0_;
  assign new_n3302_ = pstart_0_ & new_n3301_;
  assign new_n3303_ = new_n1200_ & new_n2415_;
  assign new_n3304_ = ~pstart_0_ & new_n3303_;
  assign new_n3305_ = pkey_57_ & ~pencrypt_0_;
  assign new_n3306_ = pstart_0_ & new_n3305_;
  assign new_n3307_ = n_n2458 & new_n1220_;
  assign new_n3308_ = pencrypt_0_ & new_n3307_;
  assign new_n3309_ = ~n_n2853 & new_n3308_;
  assign new_n3310_ = ~pstart_0_ & new_n3309_;
  assign new_n3311_ = ~n_n2458 & new_n1220_;
  assign new_n3312_ = pencrypt_0_ & new_n3311_;
  assign new_n3313_ = n_n2853 & new_n3312_;
  assign new_n3314_ = ~pstart_0_ & new_n3313_;
  assign new_n3315_ = ~new_n1200_ & new_n2438_;
  assign new_n3316_ = ~pstart_0_ & new_n3315_;
  assign new_n3317_ = n_n2458 & ~new_n1220_;
  assign new_n3318_ = pencrypt_0_ & new_n3317_;
  assign new_n3319_ = n_n2853 & new_n3318_;
  assign new_n3320_ = ~pstart_0_ & new_n3319_;
  assign new_n3321_ = ~new_n3316_ & ~new_n3320_;
  assign new_n3322_ = ~new_n3310_ & ~new_n3314_;
  assign new_n3323_ = new_n3321_ & new_n3322_;
  assign new_n3324_ = ~new_n3304_ & ~new_n3306_;
  assign new_n3325_ = ~new_n3298_ & ~new_n3300_;
  assign new_n3326_ = ~new_n3302_ & new_n3325_;
  assign new_n3327_ = new_n3324_ & new_n3326_;
  assign n1202 = ~new_n3323_ | ~new_n3327_;
  assign new_n3329_ = ~pencrypt_0_ & n_n2278;
  assign new_n3330_ = ~new_n1200_ & new_n3329_;
  assign new_n3331_ = ~pstart_0_ & new_n3330_;
  assign new_n3332_ = n_n2373 & n_n2278;
  assign new_n3333_ = ~pencrypt_0_ & new_n3332_;
  assign new_n3334_ = new_n1200_ & new_n3333_;
  assign new_n3335_ = ~pstart_0_ & new_n3334_;
  assign new_n3336_ = pencrypt_0_ & pkey_62_;
  assign new_n3337_ = pstart_0_ & new_n3336_;
  assign new_n3338_ = ~pencrypt_0_ & n_n2373;
  assign new_n3339_ = ~new_n1200_ & new_n3338_;
  assign new_n3340_ = ~pstart_0_ & new_n3339_;
  assign new_n3341_ = pkey_195_ & ~pencrypt_0_;
  assign new_n3342_ = pstart_0_ & new_n3341_;
  assign new_n3343_ = ~n_n2278 & ~new_n1220_;
  assign new_n3344_ = pencrypt_0_ & new_n3343_;
  assign new_n3345_ = n_n2373 & new_n3344_;
  assign new_n3346_ = ~pstart_0_ & new_n3345_;
  assign new_n3347_ = n_n2278 & new_n1220_;
  assign new_n3348_ = pencrypt_0_ & new_n3347_;
  assign new_n3349_ = n_n2373 & new_n3348_;
  assign new_n3350_ = ~pstart_0_ & new_n3349_;
  assign new_n3351_ = ~n_n2373 & ~n_n2278;
  assign new_n3352_ = ~pencrypt_0_ & new_n3351_;
  assign new_n3353_ = new_n1200_ & new_n3352_;
  assign new_n3354_ = ~pstart_0_ & new_n3353_;
  assign new_n3355_ = n_n2278 & ~new_n1220_;
  assign new_n3356_ = pencrypt_0_ & new_n3355_;
  assign new_n3357_ = ~n_n2373 & new_n3356_;
  assign new_n3358_ = ~pstart_0_ & new_n3357_;
  assign new_n3359_ = ~new_n3354_ & ~new_n3358_;
  assign new_n3360_ = ~new_n3346_ & ~new_n3350_;
  assign new_n3361_ = new_n3359_ & new_n3360_;
  assign new_n3362_ = ~new_n3340_ & ~new_n3342_;
  assign new_n3363_ = ~new_n3331_ & ~new_n3335_;
  assign new_n3364_ = ~new_n3337_ & new_n3363_;
  assign new_n3365_ = new_n3362_ & new_n3364_;
  assign n1207 = ~new_n3361_ | ~new_n3365_;
  assign new_n3367_ = ~new_n1200_ & new_n2462_;
  assign new_n3368_ = ~pstart_0_ & new_n3367_;
  assign new_n3369_ = new_n1200_ & new_n2457_;
  assign new_n3370_ = ~pstart_0_ & new_n3369_;
  assign new_n3371_ = pkey_228_ & pencrypt_0_;
  assign new_n3372_ = pstart_0_ & new_n3371_;
  assign new_n3373_ = ~new_n1200_ & new_n2453_;
  assign new_n3374_ = ~pstart_0_ & new_n3373_;
  assign new_n3375_ = ~n_n2285 & ~new_n1220_;
  assign new_n3376_ = pencrypt_0_ & new_n3375_;
  assign new_n3377_ = n_n2381 & new_n3376_;
  assign new_n3378_ = ~pstart_0_ & new_n3377_;
  assign new_n3379_ = n_n2285 & new_n1220_;
  assign new_n3380_ = pencrypt_0_ & new_n3379_;
  assign new_n3381_ = n_n2381 & new_n3380_;
  assign new_n3382_ = ~pstart_0_ & new_n3381_;
  assign new_n3383_ = new_n1200_ & new_n2476_;
  assign new_n3384_ = ~pstart_0_ & new_n3383_;
  assign new_n3385_ = n_n2285 & ~new_n1220_;
  assign new_n3386_ = pencrypt_0_ & new_n3385_;
  assign new_n3387_ = ~n_n2381 & new_n3386_;
  assign new_n3388_ = ~pstart_0_ & new_n3387_;
  assign new_n3389_ = ~new_n3384_ & ~new_n3388_;
  assign new_n3390_ = ~new_n3378_ & ~new_n3382_;
  assign new_n3391_ = new_n3389_ & new_n3390_;
  assign new_n3392_ = ~new_n1676_ & ~new_n3374_;
  assign new_n3393_ = ~new_n3368_ & ~new_n3370_;
  assign new_n3394_ = ~new_n3372_ & new_n3393_;
  assign new_n3395_ = new_n3392_ & new_n3394_;
  assign n1212 = ~new_n3391_ | ~new_n3395_;
  assign new_n3397_ = ~pencrypt_0_ & n_n2292;
  assign new_n3398_ = ~new_n1200_ & new_n3397_;
  assign new_n3399_ = ~pstart_0_ & new_n3398_;
  assign new_n3400_ = n_n2885 & n_n2292;
  assign new_n3401_ = ~pencrypt_0_ & new_n3400_;
  assign new_n3402_ = new_n1200_ & new_n3401_;
  assign new_n3403_ = ~pstart_0_ & new_n3402_;
  assign new_n3404_ = pkey_237_ & pencrypt_0_;
  assign new_n3405_ = pstart_0_ & new_n3404_;
  assign new_n3406_ = ~pencrypt_0_ & n_n2885;
  assign new_n3407_ = ~new_n1200_ & new_n3406_;
  assign new_n3408_ = ~pstart_0_ & new_n3407_;
  assign new_n3409_ = pkey_245_ & ~pencrypt_0_;
  assign new_n3410_ = pstart_0_ & new_n3409_;
  assign new_n3411_ = ~n_n2292 & ~new_n1220_;
  assign new_n3412_ = pencrypt_0_ & new_n3411_;
  assign new_n3413_ = n_n2885 & new_n3412_;
  assign new_n3414_ = ~pstart_0_ & new_n3413_;
  assign new_n3415_ = n_n2292 & new_n1220_;
  assign new_n3416_ = pencrypt_0_ & new_n3415_;
  assign new_n3417_ = n_n2885 & new_n3416_;
  assign new_n3418_ = ~pstart_0_ & new_n3417_;
  assign new_n3419_ = ~n_n2885 & ~n_n2292;
  assign new_n3420_ = ~pencrypt_0_ & new_n3419_;
  assign new_n3421_ = new_n1200_ & new_n3420_;
  assign new_n3422_ = ~pstart_0_ & new_n3421_;
  assign new_n3423_ = n_n2292 & ~new_n1220_;
  assign new_n3424_ = pencrypt_0_ & new_n3423_;
  assign new_n3425_ = ~n_n2885 & new_n3424_;
  assign new_n3426_ = ~pstart_0_ & new_n3425_;
  assign new_n3427_ = ~new_n3422_ & ~new_n3426_;
  assign new_n3428_ = ~new_n3414_ & ~new_n3418_;
  assign new_n3429_ = new_n3427_ & new_n3428_;
  assign new_n3430_ = ~new_n3408_ & ~new_n3410_;
  assign new_n3431_ = ~new_n3399_ & ~new_n3403_;
  assign new_n3432_ = ~new_n3405_ & new_n3431_;
  assign new_n3433_ = new_n3430_ & new_n3432_;
  assign n1217 = ~new_n3429_ | ~new_n3433_;
  assign new_n3435_ = ~pencrypt_0_ & n_n2838;
  assign new_n3436_ = ~new_n1200_ & new_n3435_;
  assign new_n3437_ = ~pstart_0_ & new_n3436_;
  assign new_n3438_ = n_n2447 & n_n2838;
  assign new_n3439_ = ~pencrypt_0_ & new_n3438_;
  assign new_n3440_ = new_n1200_ & new_n3439_;
  assign new_n3441_ = ~pstart_0_ & new_n3440_;
  assign new_n3442_ = pencrypt_0_ & pkey_12_;
  assign new_n3443_ = pstart_0_ & new_n3442_;
  assign new_n3444_ = ~pencrypt_0_ & n_n2447;
  assign new_n3445_ = ~new_n1200_ & new_n3444_;
  assign new_n3446_ = ~pstart_0_ & new_n3445_;
  assign new_n3447_ = ~pencrypt_0_ & pkey_20_;
  assign new_n3448_ = pstart_0_ & new_n3447_;
  assign new_n3449_ = ~n_n2838 & ~new_n1220_;
  assign new_n3450_ = pencrypt_0_ & new_n3449_;
  assign new_n3451_ = n_n2447 & new_n3450_;
  assign new_n3452_ = ~pstart_0_ & new_n3451_;
  assign new_n3453_ = n_n2838 & new_n1220_;
  assign new_n3454_ = pencrypt_0_ & new_n3453_;
  assign new_n3455_ = n_n2447 & new_n3454_;
  assign new_n3456_ = ~pstart_0_ & new_n3455_;
  assign new_n3457_ = ~n_n2447 & ~n_n2838;
  assign new_n3458_ = ~pencrypt_0_ & new_n3457_;
  assign new_n3459_ = new_n1200_ & new_n3458_;
  assign new_n3460_ = ~pstart_0_ & new_n3459_;
  assign new_n3461_ = n_n2838 & ~new_n1220_;
  assign new_n3462_ = pencrypt_0_ & new_n3461_;
  assign new_n3463_ = ~n_n2447 & new_n3462_;
  assign new_n3464_ = ~pstart_0_ & new_n3463_;
  assign new_n3465_ = ~new_n3460_ & ~new_n3464_;
  assign new_n3466_ = ~new_n3452_ & ~new_n3456_;
  assign new_n3467_ = new_n3465_ & new_n3466_;
  assign new_n3468_ = ~new_n3446_ & ~new_n3448_;
  assign new_n3469_ = ~new_n3437_ & ~new_n3441_;
  assign new_n3470_ = ~new_n3443_ & new_n3469_;
  assign new_n3471_ = new_n3468_ & new_n3470_;
  assign n1222 = ~new_n3467_ | ~new_n3471_;
  assign new_n3473_ = ~pencrypt_0_ & n_n2361;
  assign new_n3474_ = ~new_n1200_ & new_n3473_;
  assign new_n3475_ = ~pstart_0_ & new_n3474_;
  assign new_n3476_ = n_n2455 & n_n2361;
  assign new_n3477_ = ~pencrypt_0_ & new_n3476_;
  assign new_n3478_ = new_n1200_ & new_n3477_;
  assign new_n3479_ = ~pstart_0_ & new_n3478_;
  assign new_n3480_ = pencrypt_0_ & pkey_21_;
  assign new_n3481_ = pstart_0_ & new_n3480_;
  assign new_n3482_ = ~pencrypt_0_ & n_n2455;
  assign new_n3483_ = ~new_n1200_ & new_n3482_;
  assign new_n3484_ = ~pstart_0_ & new_n3483_;
  assign new_n3485_ = pkey_29_ & ~pencrypt_0_;
  assign new_n3486_ = pstart_0_ & new_n3485_;
  assign new_n3487_ = ~n_n2361 & ~new_n1220_;
  assign new_n3488_ = pencrypt_0_ & new_n3487_;
  assign new_n3489_ = n_n2455 & new_n3488_;
  assign new_n3490_ = ~pstart_0_ & new_n3489_;
  assign new_n3491_ = n_n2361 & new_n1220_;
  assign new_n3492_ = pencrypt_0_ & new_n3491_;
  assign new_n3493_ = n_n2455 & new_n3492_;
  assign new_n3494_ = ~pstart_0_ & new_n3493_;
  assign new_n3495_ = ~n_n2455 & ~n_n2361;
  assign new_n3496_ = ~pencrypt_0_ & new_n3495_;
  assign new_n3497_ = new_n1200_ & new_n3496_;
  assign new_n3498_ = ~pstart_0_ & new_n3497_;
  assign new_n3499_ = n_n2361 & ~new_n1220_;
  assign new_n3500_ = pencrypt_0_ & new_n3499_;
  assign new_n3501_ = ~n_n2455 & new_n3500_;
  assign new_n3502_ = ~pstart_0_ & new_n3501_;
  assign new_n3503_ = ~new_n3498_ & ~new_n3502_;
  assign new_n3504_ = ~new_n3490_ & ~new_n3494_;
  assign new_n3505_ = new_n3503_ & new_n3504_;
  assign new_n3506_ = ~new_n3484_ & ~new_n3486_;
  assign new_n3507_ = ~new_n3475_ & ~new_n3479_;
  assign new_n3508_ = ~new_n3481_ & new_n3507_;
  assign new_n3509_ = new_n3506_ & new_n3508_;
  assign n1227 = ~new_n3505_ | ~new_n3509_;
  assign new_n3511_ = ~pencrypt_0_ & n_n2369;
  assign new_n3512_ = ~new_n1200_ & new_n3511_;
  assign new_n3513_ = ~pstart_0_ & new_n3512_;
  assign new_n3514_ = n_n2462 & n_n2369;
  assign new_n3515_ = ~pencrypt_0_ & new_n3514_;
  assign new_n3516_ = new_n1200_ & new_n3515_;
  assign new_n3517_ = ~pstart_0_ & new_n3516_;
  assign new_n3518_ = pencrypt_0_ & pkey_30_;
  assign new_n3519_ = pstart_0_ & new_n3518_;
  assign new_n3520_ = ~pencrypt_0_ & n_n2462;
  assign new_n3521_ = ~new_n1200_ & new_n3520_;
  assign new_n3522_ = ~pstart_0_ & new_n3521_;
  assign new_n3523_ = pkey_38_ & ~pencrypt_0_;
  assign new_n3524_ = pstart_0_ & new_n3523_;
  assign new_n3525_ = ~n_n2369 & ~new_n1220_;
  assign new_n3526_ = pencrypt_0_ & new_n3525_;
  assign new_n3527_ = n_n2462 & new_n3526_;
  assign new_n3528_ = ~pstart_0_ & new_n3527_;
  assign new_n3529_ = n_n2369 & new_n1220_;
  assign new_n3530_ = pencrypt_0_ & new_n3529_;
  assign new_n3531_ = n_n2462 & new_n3530_;
  assign new_n3532_ = ~pstart_0_ & new_n3531_;
  assign new_n3533_ = ~n_n2462 & ~n_n2369;
  assign new_n3534_ = ~pencrypt_0_ & new_n3533_;
  assign new_n3535_ = new_n1200_ & new_n3534_;
  assign new_n3536_ = ~pstart_0_ & new_n3535_;
  assign new_n3537_ = n_n2369 & ~new_n1220_;
  assign new_n3538_ = pencrypt_0_ & new_n3537_;
  assign new_n3539_ = ~n_n2462 & new_n3538_;
  assign new_n3540_ = ~pstart_0_ & new_n3539_;
  assign new_n3541_ = ~new_n3536_ & ~new_n3540_;
  assign new_n3542_ = ~new_n3528_ & ~new_n3532_;
  assign new_n3543_ = new_n3541_ & new_n3542_;
  assign new_n3544_ = ~new_n3522_ & ~new_n3524_;
  assign new_n3545_ = ~new_n3513_ & ~new_n3517_;
  assign new_n3546_ = ~new_n3519_ & new_n3545_;
  assign new_n3547_ = new_n3544_ & new_n3546_;
  assign n1232 = ~new_n3543_ | ~new_n3547_;
  assign new_n3549_ = new_n1200_ & new_n1862_1_;
  assign new_n3550_ = ~pstart_0_ & new_n3549_;
  assign new_n3551_ = ~new_n1200_ & new_n1857_1_;
  assign new_n3552_ = ~pstart_0_ & new_n3551_;
  assign new_n3553_ = pkey_194_ & pencrypt_0_;
  assign new_n3554_ = pstart_0_ & new_n3553_;
  assign new_n3555_ = new_n1200_ & new_n1853_;
  assign new_n3556_ = ~pstart_0_ & new_n3555_;
  assign new_n3557_ = ~pencrypt_0_ & pkey_202_;
  assign new_n3558_ = pstart_0_ & new_n3557_;
  assign new_n3559_ = n_n2377 & new_n1220_;
  assign new_n3560_ = pencrypt_0_ & new_n3559_;
  assign new_n3561_ = ~n_n2282 & new_n3560_;
  assign new_n3562_ = ~pstart_0_ & new_n3561_;
  assign new_n3563_ = ~n_n2377 & new_n1220_;
  assign new_n3564_ = pencrypt_0_ & new_n3563_;
  assign new_n3565_ = n_n2282 & new_n3564_;
  assign new_n3566_ = ~pstart_0_ & new_n3565_;
  assign new_n3567_ = ~new_n1200_ & new_n1876_;
  assign new_n3568_ = ~pstart_0_ & new_n3567_;
  assign new_n3569_ = n_n2377 & ~new_n1220_;
  assign new_n3570_ = pencrypt_0_ & new_n3569_;
  assign new_n3571_ = n_n2282 & new_n3570_;
  assign new_n3572_ = ~pstart_0_ & new_n3571_;
  assign new_n3573_ = ~new_n3568_ & ~new_n3572_;
  assign new_n3574_ = ~new_n3562_ & ~new_n3566_;
  assign new_n3575_ = new_n3573_ & new_n3574_;
  assign new_n3576_ = ~new_n3556_ & ~new_n3558_;
  assign new_n3577_ = ~new_n3550_ & ~new_n3552_;
  assign new_n3578_ = ~new_n3554_ & new_n3577_;
  assign new_n3579_ = new_n3576_ & new_n3578_;
  assign n1237 = ~new_n3575_ | ~new_n3579_;
  assign new_n3581_ = ~pencrypt_0_ & n_n2301;
  assign new_n3582_ = ~new_n1200_ & new_n3581_;
  assign new_n3583_ = ~pstart_0_ & new_n3582_;
  assign new_n3584_ = n_n2395 & n_n2301;
  assign new_n3585_ = ~pencrypt_0_ & new_n3584_;
  assign new_n3586_ = new_n1200_ & new_n3585_;
  assign new_n3587_ = ~pstart_0_ & new_n3586_;
  assign new_n3588_ = pkey_254_ & pencrypt_0_;
  assign new_n3589_ = pstart_0_ & new_n3588_;
  assign new_n3590_ = ~pencrypt_0_ & n_n2395;
  assign new_n3591_ = ~new_n1200_ & new_n3590_;
  assign new_n3592_ = ~pstart_0_ & new_n3591_;
  assign new_n3593_ = pkey_131_ & ~pencrypt_0_;
  assign new_n3594_ = pstart_0_ & new_n3593_;
  assign new_n3595_ = ~n_n2301 & ~new_n1220_;
  assign new_n3596_ = pencrypt_0_ & new_n3595_;
  assign new_n3597_ = n_n2395 & new_n3596_;
  assign new_n3598_ = ~pstart_0_ & new_n3597_;
  assign new_n3599_ = n_n2301 & new_n1220_;
  assign new_n3600_ = pencrypt_0_ & new_n3599_;
  assign new_n3601_ = n_n2395 & new_n3600_;
  assign new_n3602_ = ~pstart_0_ & new_n3601_;
  assign new_n3603_ = ~n_n2395 & ~n_n2301;
  assign new_n3604_ = ~pencrypt_0_ & new_n3603_;
  assign new_n3605_ = new_n1200_ & new_n3604_;
  assign new_n3606_ = ~pstart_0_ & new_n3605_;
  assign new_n3607_ = n_n2301 & ~new_n1220_;
  assign new_n3608_ = pencrypt_0_ & new_n3607_;
  assign new_n3609_ = ~n_n2395 & new_n3608_;
  assign new_n3610_ = ~pstart_0_ & new_n3609_;
  assign new_n3611_ = ~new_n3606_ & ~new_n3610_;
  assign new_n3612_ = ~new_n3598_ & ~new_n3602_;
  assign new_n3613_ = new_n3611_ & new_n3612_;
  assign new_n3614_ = ~new_n3592_ & ~new_n3594_;
  assign new_n3615_ = ~new_n3583_ & ~new_n3587_;
  assign new_n3616_ = ~new_n3589_ & new_n3615_;
  assign new_n3617_ = new_n3614_ & new_n3616_;
  assign n1242 = ~new_n3613_ | ~new_n3617_;
  assign new_n3619_ = ~pencrypt_0_ & n_n2309;
  assign new_n3620_ = ~new_n1200_ & new_n3619_;
  assign new_n3621_ = ~pstart_0_ & new_n3620_;
  assign new_n3622_ = n_n2909 & n_n2309;
  assign new_n3623_ = ~pencrypt_0_ & new_n3622_;
  assign new_n3624_ = new_n1200_ & new_n3623_;
  assign new_n3625_ = ~pstart_0_ & new_n3624_;
  assign new_n3626_ = pkey_180_ & pencrypt_0_;
  assign new_n3627_ = pstart_0_ & new_n3626_;
  assign new_n3628_ = ~pencrypt_0_ & n_n2909;
  assign new_n3629_ = ~new_n1200_ & new_n3628_;
  assign new_n3630_ = ~pstart_0_ & new_n3629_;
  assign new_n3631_ = ~pencrypt_0_ & pkey_188_;
  assign new_n3632_ = pstart_0_ & new_n3631_;
  assign new_n3633_ = ~n_n2309 & ~new_n1220_;
  assign new_n3634_ = pencrypt_0_ & new_n3633_;
  assign new_n3635_ = n_n2909 & new_n3634_;
  assign new_n3636_ = ~pstart_0_ & new_n3635_;
  assign new_n3637_ = n_n2309 & new_n1220_;
  assign new_n3638_ = pencrypt_0_ & new_n3637_;
  assign new_n3639_ = n_n2909 & new_n3638_;
  assign new_n3640_ = ~pstart_0_ & new_n3639_;
  assign new_n3641_ = ~n_n2909 & ~n_n2309;
  assign new_n3642_ = ~pencrypt_0_ & new_n3641_;
  assign new_n3643_ = new_n1200_ & new_n3642_;
  assign new_n3644_ = ~pstart_0_ & new_n3643_;
  assign new_n3645_ = n_n2309 & ~new_n1220_;
  assign new_n3646_ = pencrypt_0_ & new_n3645_;
  assign new_n3647_ = ~n_n2909 & new_n3646_;
  assign new_n3648_ = ~pstart_0_ & new_n3647_;
  assign new_n3649_ = ~new_n3644_ & ~new_n3648_;
  assign new_n3650_ = ~new_n3636_ & ~new_n3640_;
  assign new_n3651_ = new_n3649_ & new_n3650_;
  assign new_n3652_ = ~new_n3630_ & ~new_n3632_;
  assign new_n3653_ = ~new_n3621_ & ~new_n3625_;
  assign new_n3654_ = ~new_n3627_ & new_n3653_;
  assign new_n3655_ = new_n3652_ & new_n3654_;
  assign n1247 = ~new_n3651_ | ~new_n3655_;
  assign new_n3657_ = ~pencrypt_0_ & n_n2319;
  assign new_n3658_ = ~new_n1200_ & new_n3657_;
  assign new_n3659_ = ~pstart_0_ & new_n3658_;
  assign new_n3660_ = n_n2413 & n_n2319;
  assign new_n3661_ = ~pencrypt_0_ & new_n3660_;
  assign new_n3662_ = new_n1200_ & new_n3661_;
  assign new_n3663_ = ~pstart_0_ & new_n3662_;
  assign new_n3664_ = pkey_142_ & pencrypt_0_;
  assign new_n3665_ = pstart_0_ & new_n3664_;
  assign new_n3666_ = ~pencrypt_0_ & n_n2413;
  assign new_n3667_ = ~new_n1200_ & new_n3666_;
  assign new_n3668_ = ~pstart_0_ & new_n3667_;
  assign new_n3669_ = pkey_150_ & ~pencrypt_0_;
  assign new_n3670_ = pstart_0_ & new_n3669_;
  assign new_n3671_ = ~n_n2319 & ~new_n1220_;
  assign new_n3672_ = pencrypt_0_ & new_n3671_;
  assign new_n3673_ = n_n2413 & new_n3672_;
  assign new_n3674_ = ~pstart_0_ & new_n3673_;
  assign new_n3675_ = n_n2319 & new_n1220_;
  assign new_n3676_ = pencrypt_0_ & new_n3675_;
  assign new_n3677_ = n_n2413 & new_n3676_;
  assign new_n3678_ = ~pstart_0_ & new_n3677_;
  assign new_n3679_ = ~n_n2413 & ~n_n2319;
  assign new_n3680_ = ~pencrypt_0_ & new_n3679_;
  assign new_n3681_ = new_n1200_ & new_n3680_;
  assign new_n3682_ = ~pstart_0_ & new_n3681_;
  assign new_n3683_ = n_n2319 & ~new_n1220_;
  assign new_n3684_ = pencrypt_0_ & new_n3683_;
  assign new_n3685_ = ~n_n2413 & new_n3684_;
  assign new_n3686_ = ~pstart_0_ & new_n3685_;
  assign new_n3687_ = ~new_n3682_ & ~new_n3686_;
  assign new_n3688_ = ~new_n3674_ & ~new_n3678_;
  assign new_n3689_ = new_n3687_ & new_n3688_;
  assign new_n3690_ = ~new_n3668_ & ~new_n3670_;
  assign new_n3691_ = ~new_n3659_ & ~new_n3663_;
  assign new_n3692_ = ~new_n3665_ & new_n3691_;
  assign new_n3693_ = new_n3690_ & new_n3692_;
  assign n1252 = ~new_n3689_ | ~new_n3693_;
  assign new_n3695_ = ~pencrypt_0_ & n_n2329;
  assign new_n3696_ = ~new_n1200_ & new_n3695_;
  assign new_n3697_ = ~pstart_0_ & new_n3696_;
  assign new_n3698_ = n_n2423 & n_n2329;
  assign new_n3699_ = ~pencrypt_0_ & new_n3698_;
  assign new_n3700_ = new_n1200_ & new_n3699_;
  assign new_n3701_ = ~pstart_0_ & new_n3700_;
  assign new_n3702_ = pkey_68_ & pencrypt_0_;
  assign new_n3703_ = pstart_0_ & new_n3702_;
  assign new_n3704_ = ~pencrypt_0_ & n_n2423;
  assign new_n3705_ = ~new_n1200_ & new_n3704_;
  assign new_n3706_ = ~pstart_0_ & new_n3705_;
  assign new_n3707_ = pkey_76_ & ~pencrypt_0_;
  assign new_n3708_ = pstart_0_ & new_n3707_;
  assign new_n3709_ = ~n_n2329 & ~new_n1220_;
  assign new_n3710_ = pencrypt_0_ & new_n3709_;
  assign new_n3711_ = n_n2423 & new_n3710_;
  assign new_n3712_ = ~pstart_0_ & new_n3711_;
  assign new_n3713_ = n_n2329 & new_n1220_;
  assign new_n3714_ = pencrypt_0_ & new_n3713_;
  assign new_n3715_ = n_n2423 & new_n3714_;
  assign new_n3716_ = ~pstart_0_ & new_n3715_;
  assign new_n3717_ = ~n_n2423 & ~n_n2329;
  assign new_n3718_ = ~pencrypt_0_ & new_n3717_;
  assign new_n3719_ = new_n1200_ & new_n3718_;
  assign new_n3720_ = ~pstart_0_ & new_n3719_;
  assign new_n3721_ = n_n2329 & ~new_n1220_;
  assign new_n3722_ = pencrypt_0_ & new_n3721_;
  assign new_n3723_ = ~n_n2423 & new_n3722_;
  assign new_n3724_ = ~pstart_0_ & new_n3723_;
  assign new_n3725_ = ~new_n3720_ & ~new_n3724_;
  assign new_n3726_ = ~new_n3712_ & ~new_n3716_;
  assign new_n3727_ = new_n3725_ & new_n3726_;
  assign new_n3728_ = ~new_n3706_ & ~new_n3708_;
  assign new_n3729_ = ~new_n3697_ & ~new_n3701_;
  assign new_n3730_ = ~new_n3703_ & new_n3729_;
  assign new_n3731_ = new_n3728_ & new_n3730_;
  assign n1257 = ~new_n3727_ | ~new_n3731_;
  assign new_n3733_ = ~pencrypt_0_ & n_n2338;
  assign new_n3734_ = ~new_n1200_ & new_n3733_;
  assign new_n3735_ = ~pstart_0_ & new_n3734_;
  assign new_n3736_ = n_n2432 & n_n2338;
  assign new_n3737_ = ~pencrypt_0_ & new_n3736_;
  assign new_n3738_ = new_n1200_ & new_n3737_;
  assign new_n3739_ = ~pstart_0_ & new_n3738_;
  assign new_n3740_ = pkey_93_ & pencrypt_0_;
  assign new_n3741_ = pstart_0_ & new_n3740_;
  assign new_n3742_ = ~pencrypt_0_ & n_n2432;
  assign new_n3743_ = ~new_n1200_ & new_n3742_;
  assign new_n3744_ = ~pstart_0_ & new_n3743_;
  assign new_n3745_ = ~pencrypt_0_ & pkey_101_;
  assign new_n3746_ = pstart_0_ & new_n3745_;
  assign new_n3747_ = ~n_n2338 & ~new_n1220_;
  assign new_n3748_ = pencrypt_0_ & new_n3747_;
  assign new_n3749_ = n_n2432 & new_n3748_;
  assign new_n3750_ = ~pstart_0_ & new_n3749_;
  assign new_n3751_ = n_n2338 & new_n1220_;
  assign new_n3752_ = pencrypt_0_ & new_n3751_;
  assign new_n3753_ = n_n2432 & new_n3752_;
  assign new_n3754_ = ~pstart_0_ & new_n3753_;
  assign new_n3755_ = ~n_n2432 & ~n_n2338;
  assign new_n3756_ = ~pencrypt_0_ & new_n3755_;
  assign new_n3757_ = new_n1200_ & new_n3756_;
  assign new_n3758_ = ~pstart_0_ & new_n3757_;
  assign new_n3759_ = n_n2338 & ~new_n1220_;
  assign new_n3760_ = pencrypt_0_ & new_n3759_;
  assign new_n3761_ = ~n_n2432 & new_n3760_;
  assign new_n3762_ = ~pstart_0_ & new_n3761_;
  assign new_n3763_ = ~new_n3758_ & ~new_n3762_;
  assign new_n3764_ = ~new_n3750_ & ~new_n3754_;
  assign new_n3765_ = new_n3763_ & new_n3764_;
  assign new_n3766_ = ~new_n3744_ & ~new_n3746_;
  assign new_n3767_ = ~new_n3735_ & ~new_n3739_;
  assign new_n3768_ = ~new_n3741_ & new_n3767_;
  assign new_n3769_ = new_n3766_ & new_n3768_;
  assign n1262 = ~new_n3765_ | ~new_n3769_;
  assign new_n3771_ = ~pencrypt_0_ & n_n2348;
  assign new_n3772_ = ~new_n1200_ & new_n3771_;
  assign new_n3773_ = ~pstart_0_ & new_n3772_;
  assign new_n3774_ = n_n2441 & n_n2348;
  assign new_n3775_ = ~pencrypt_0_ & new_n3774_;
  assign new_n3776_ = new_n1200_ & new_n3775_;
  assign new_n3777_ = ~pstart_0_ & new_n3776_;
  assign new_n3778_ = pkey_118_ & pencrypt_0_;
  assign new_n3779_ = pstart_0_ & new_n3778_;
  assign new_n3780_ = ~pencrypt_0_ & n_n2441;
  assign new_n3781_ = ~new_n1200_ & new_n3780_;
  assign new_n3782_ = ~pstart_0_ & new_n3781_;
  assign new_n3783_ = pkey_126_ & ~pencrypt_0_;
  assign new_n3784_ = pstart_0_ & new_n3783_;
  assign new_n3785_ = ~n_n2348 & ~new_n1220_;
  assign new_n3786_ = pencrypt_0_ & new_n3785_;
  assign new_n3787_ = n_n2441 & new_n3786_;
  assign new_n3788_ = ~pstart_0_ & new_n3787_;
  assign new_n3789_ = n_n2348 & new_n1220_;
  assign new_n3790_ = pencrypt_0_ & new_n3789_;
  assign new_n3791_ = n_n2441 & new_n3790_;
  assign new_n3792_ = ~pstart_0_ & new_n3791_;
  assign new_n3793_ = ~n_n2441 & ~n_n2348;
  assign new_n3794_ = ~pencrypt_0_ & new_n3793_;
  assign new_n3795_ = new_n1200_ & new_n3794_;
  assign new_n3796_ = ~pstart_0_ & new_n3795_;
  assign new_n3797_ = n_n2348 & ~new_n1220_;
  assign new_n3798_ = pencrypt_0_ & new_n3797_;
  assign new_n3799_ = ~n_n2441 & new_n3798_;
  assign new_n3800_ = ~pstart_0_ & new_n3799_;
  assign new_n3801_ = ~new_n3796_ & ~new_n3800_;
  assign new_n3802_ = ~new_n3788_ & ~new_n3792_;
  assign new_n3803_ = new_n3801_ & new_n3802_;
  assign new_n3804_ = ~new_n3782_ & ~new_n3784_;
  assign new_n3805_ = ~new_n3773_ & ~new_n3777_;
  assign new_n3806_ = ~new_n3779_ & new_n3805_;
  assign new_n3807_ = new_n3804_ & new_n3806_;
  assign n1267 = ~new_n3803_ | ~new_n3807_;
  assign new_n3809_ = ~pencrypt_0_ & n_n2378;
  assign new_n3810_ = new_n1200_ & new_n3809_;
  assign new_n3811_ = ~pstart_0_ & new_n3810_;
  assign new_n3812_ = n_n2741 & n_n2378;
  assign new_n3813_ = ~pencrypt_0_ & new_n3812_;
  assign new_n3814_ = ~new_n1200_ & new_n3813_;
  assign new_n3815_ = ~pstart_0_ & new_n3814_;
  assign new_n3816_ = pencrypt_0_ & pkey_202_;
  assign new_n3817_ = pstart_0_ & new_n3816_;
  assign new_n3818_ = ~pencrypt_0_ & n_n2741;
  assign new_n3819_ = new_n1200_ & new_n3818_;
  assign new_n3820_ = ~pstart_0_ & new_n3819_;
  assign new_n3821_ = pkey_210_ & ~pencrypt_0_;
  assign new_n3822_ = pstart_0_ & new_n3821_;
  assign new_n3823_ = n_n2378 & new_n1220_;
  assign new_n3824_ = pencrypt_0_ & new_n3823_;
  assign new_n3825_ = ~n_n2741 & new_n3824_;
  assign new_n3826_ = ~pstart_0_ & new_n3825_;
  assign new_n3827_ = ~n_n2378 & new_n1220_;
  assign new_n3828_ = pencrypt_0_ & new_n3827_;
  assign new_n3829_ = n_n2741 & new_n3828_;
  assign new_n3830_ = ~pstart_0_ & new_n3829_;
  assign new_n3831_ = ~n_n2741 & ~n_n2378;
  assign new_n3832_ = ~pencrypt_0_ & new_n3831_;
  assign new_n3833_ = ~new_n1200_ & new_n3832_;
  assign new_n3834_ = ~pstart_0_ & new_n3833_;
  assign new_n3835_ = n_n2378 & ~new_n1220_;
  assign new_n3836_ = pencrypt_0_ & new_n3835_;
  assign new_n3837_ = n_n2741 & new_n3836_;
  assign new_n3838_ = ~pstart_0_ & new_n3837_;
  assign new_n3839_ = ~new_n3834_ & ~new_n3838_;
  assign new_n3840_ = ~new_n3826_ & ~new_n3830_;
  assign new_n3841_ = new_n3839_ & new_n3840_;
  assign new_n3842_ = ~new_n3820_ & ~new_n3822_;
  assign new_n3843_ = ~new_n3811_ & ~new_n3815_;
  assign new_n3844_ = ~new_n3817_ & new_n3843_;
  assign new_n3845_ = new_n3842_ & new_n3844_;
  assign n1272 = ~new_n3841_ | ~new_n3845_;
  assign new_n3847_ = ~pencrypt_0_ & n_n2302;
  assign new_n3848_ = ~new_n1200_ & new_n3847_;
  assign new_n3849_ = ~pstart_0_ & new_n3848_;
  assign new_n3850_ = n_n2396 & n_n2302;
  assign new_n3851_ = ~pencrypt_0_ & new_n3850_;
  assign new_n3852_ = new_n1200_ & new_n3851_;
  assign new_n3853_ = ~pstart_0_ & new_n3852_;
  assign new_n3854_ = pkey_131_ & pencrypt_0_;
  assign new_n3855_ = pstart_0_ & new_n3854_;
  assign new_n3856_ = ~pencrypt_0_ & n_n2396;
  assign new_n3857_ = ~new_n1200_ & new_n3856_;
  assign new_n3858_ = ~pstart_0_ & new_n3857_;
  assign new_n3859_ = pkey_139_ & ~pencrypt_0_;
  assign new_n3860_ = pstart_0_ & new_n3859_;
  assign new_n3861_ = ~n_n2302 & ~new_n1220_;
  assign new_n3862_ = pencrypt_0_ & new_n3861_;
  assign new_n3863_ = n_n2396 & new_n3862_;
  assign new_n3864_ = ~pstart_0_ & new_n3863_;
  assign new_n3865_ = n_n2302 & new_n1220_;
  assign new_n3866_ = pencrypt_0_ & new_n3865_;
  assign new_n3867_ = n_n2396 & new_n3866_;
  assign new_n3868_ = ~pstart_0_ & new_n3867_;
  assign new_n3869_ = ~n_n2396 & ~n_n2302;
  assign new_n3870_ = ~pencrypt_0_ & new_n3869_;
  assign new_n3871_ = new_n1200_ & new_n3870_;
  assign new_n3872_ = ~pstart_0_ & new_n3871_;
  assign new_n3873_ = n_n2302 & ~new_n1220_;
  assign new_n3874_ = pencrypt_0_ & new_n3873_;
  assign new_n3875_ = ~n_n2396 & new_n3874_;
  assign new_n3876_ = ~pstart_0_ & new_n3875_;
  assign new_n3877_ = ~new_n3872_ & ~new_n3876_;
  assign new_n3878_ = ~new_n3864_ & ~new_n3868_;
  assign new_n3879_ = new_n3877_ & new_n3878_;
  assign new_n3880_ = ~new_n3858_ & ~new_n3860_;
  assign new_n3881_ = ~new_n3849_ & ~new_n3853_;
  assign new_n3882_ = ~new_n3855_ & new_n3881_;
  assign new_n3883_ = new_n3880_ & new_n3882_;
  assign n1277 = ~new_n3879_ | ~new_n3883_;
  assign new_n3885_ = ~pencrypt_0_ & n_n2779;
  assign new_n3886_ = ~new_n1200_ & new_n3885_;
  assign new_n3887_ = ~pstart_0_ & new_n3886_;
  assign new_n3888_ = n_n2404 & n_n2779;
  assign new_n3889_ = ~pencrypt_0_ & new_n3888_;
  assign new_n3890_ = new_n1200_ & new_n3889_;
  assign new_n3891_ = ~pstart_0_ & new_n3890_;
  assign new_n3892_ = ~pencrypt_0_ & n_n2404;
  assign new_n3893_ = ~new_n1200_ & new_n3892_;
  assign new_n3894_ = ~pstart_0_ & new_n3893_;
  assign new_n3895_ = pkey_180_ & ~pencrypt_0_;
  assign new_n3896_ = pstart_0_ & new_n3895_;
  assign new_n3897_ = ~n_n2779 & ~new_n1220_;
  assign new_n3898_ = pencrypt_0_ & new_n3897_;
  assign new_n3899_ = n_n2404 & new_n3898_;
  assign new_n3900_ = ~pstart_0_ & new_n3899_;
  assign new_n3901_ = n_n2779 & new_n1220_;
  assign new_n3902_ = pencrypt_0_ & new_n3901_;
  assign new_n3903_ = n_n2404 & new_n3902_;
  assign new_n3904_ = ~pstart_0_ & new_n3903_;
  assign new_n3905_ = ~n_n2404 & ~n_n2779;
  assign new_n3906_ = ~pencrypt_0_ & new_n3905_;
  assign new_n3907_ = new_n1200_ & new_n3906_;
  assign new_n3908_ = ~pstart_0_ & new_n3907_;
  assign new_n3909_ = n_n2779 & ~new_n1220_;
  assign new_n3910_ = pencrypt_0_ & new_n3909_;
  assign new_n3911_ = ~n_n2404 & new_n3910_;
  assign new_n3912_ = ~pstart_0_ & new_n3911_;
  assign new_n3913_ = ~new_n3908_ & ~new_n3912_;
  assign new_n3914_ = ~new_n3900_ & ~new_n3904_;
  assign new_n3915_ = new_n3913_ & new_n3914_;
  assign new_n3916_ = ~new_n3894_ & ~new_n3896_;
  assign new_n3917_ = ~new_n3887_ & ~new_n3891_;
  assign new_n3918_ = ~new_n2569_ & new_n3917_;
  assign new_n3919_ = new_n3916_ & new_n3918_;
  assign n1282 = ~new_n3915_ | ~new_n3919_;
  assign new_n3921_ = ~pencrypt_0_ & n_n2320;
  assign new_n3922_ = ~new_n1200_ & new_n3921_;
  assign new_n3923_ = ~pstart_0_ & new_n3922_;
  assign new_n3924_ = n_n2414 & n_n2320;
  assign new_n3925_ = ~pencrypt_0_ & new_n3924_;
  assign new_n3926_ = new_n1200_ & new_n3925_;
  assign new_n3927_ = ~pstart_0_ & new_n3926_;
  assign new_n3928_ = pkey_150_ & pencrypt_0_;
  assign new_n3929_ = pstart_0_ & new_n3928_;
  assign new_n3930_ = ~pencrypt_0_ & n_n2414;
  assign new_n3931_ = ~new_n1200_ & new_n3930_;
  assign new_n3932_ = ~pstart_0_ & new_n3931_;
  assign new_n3933_ = pkey_158_ & ~pencrypt_0_;
  assign new_n3934_ = pstart_0_ & new_n3933_;
  assign new_n3935_ = ~n_n2320 & ~new_n1220_;
  assign new_n3936_ = pencrypt_0_ & new_n3935_;
  assign new_n3937_ = n_n2414 & new_n3936_;
  assign new_n3938_ = ~pstart_0_ & new_n3937_;
  assign new_n3939_ = n_n2320 & new_n1220_;
  assign new_n3940_ = pencrypt_0_ & new_n3939_;
  assign new_n3941_ = n_n2414 & new_n3940_;
  assign new_n3942_ = ~pstart_0_ & new_n3941_;
  assign new_n3943_ = ~n_n2414 & ~n_n2320;
  assign new_n3944_ = ~pencrypt_0_ & new_n3943_;
  assign new_n3945_ = new_n1200_ & new_n3944_;
  assign new_n3946_ = ~pstart_0_ & new_n3945_;
  assign new_n3947_ = n_n2320 & ~new_n1220_;
  assign new_n3948_ = pencrypt_0_ & new_n3947_;
  assign new_n3949_ = ~n_n2414 & new_n3948_;
  assign new_n3950_ = ~pstart_0_ & new_n3949_;
  assign new_n3951_ = ~new_n3946_ & ~new_n3950_;
  assign new_n3952_ = ~new_n3938_ & ~new_n3942_;
  assign new_n3953_ = new_n3951_ & new_n3952_;
  assign new_n3954_ = ~new_n3932_ & ~new_n3934_;
  assign new_n3955_ = ~new_n3923_ & ~new_n3927_;
  assign new_n3956_ = ~new_n3929_ & new_n3955_;
  assign new_n3957_ = new_n3954_ & new_n3956_;
  assign n1287 = ~new_n3953_ | ~new_n3957_;
  assign new_n3959_ = ~pencrypt_0_ & n_n2328;
  assign new_n3960_ = ~new_n1200_ & new_n3959_;
  assign new_n3961_ = ~pstart_0_ & new_n3960_;
  assign new_n3962_ = n_n2422 & n_n2328;
  assign new_n3963_ = ~pencrypt_0_ & new_n3962_;
  assign new_n3964_ = new_n1200_ & new_n3963_;
  assign new_n3965_ = ~pstart_0_ & new_n3964_;
  assign new_n3966_ = pencrypt_0_ & pkey_91_;
  assign new_n3967_ = pstart_0_ & new_n3966_;
  assign new_n3968_ = ~pencrypt_0_ & n_n2422;
  assign new_n3969_ = ~new_n1200_ & new_n3968_;
  assign new_n3970_ = ~pstart_0_ & new_n3969_;
  assign new_n3971_ = pkey_68_ & ~pencrypt_0_;
  assign new_n3972_ = pstart_0_ & new_n3971_;
  assign new_n3973_ = ~n_n2328 & ~new_n1220_;
  assign new_n3974_ = pencrypt_0_ & new_n3973_;
  assign new_n3975_ = n_n2422 & new_n3974_;
  assign new_n3976_ = ~pstart_0_ & new_n3975_;
  assign new_n3977_ = n_n2328 & new_n1220_;
  assign new_n3978_ = pencrypt_0_ & new_n3977_;
  assign new_n3979_ = n_n2422 & new_n3978_;
  assign new_n3980_ = ~pstart_0_ & new_n3979_;
  assign new_n3981_ = ~n_n2422 & ~n_n2328;
  assign new_n3982_ = ~pencrypt_0_ & new_n3981_;
  assign new_n3983_ = new_n1200_ & new_n3982_;
  assign new_n3984_ = ~pstart_0_ & new_n3983_;
  assign new_n3985_ = n_n2328 & ~new_n1220_;
  assign new_n3986_ = pencrypt_0_ & new_n3985_;
  assign new_n3987_ = ~n_n2422 & new_n3986_;
  assign new_n3988_ = ~pstart_0_ & new_n3987_;
  assign new_n3989_ = ~new_n3984_ & ~new_n3988_;
  assign new_n3990_ = ~new_n3976_ & ~new_n3980_;
  assign new_n3991_ = new_n3989_ & new_n3990_;
  assign new_n3992_ = ~new_n3970_ & ~new_n3972_;
  assign new_n3993_ = ~new_n3961_ & ~new_n3965_;
  assign new_n3994_ = ~new_n3967_ & new_n3993_;
  assign new_n3995_ = new_n3992_ & new_n3994_;
  assign n1292 = ~new_n3991_ | ~new_n3995_;
  assign new_n3997_ = ~pencrypt_0_ & n_n2339;
  assign new_n3998_ = ~new_n1200_ & new_n3997_;
  assign new_n3999_ = ~pstart_0_ & new_n3998_;
  assign new_n4000_ = n_n2433 & n_n2339;
  assign new_n4001_ = ~pencrypt_0_ & new_n4000_;
  assign new_n4002_ = new_n1200_ & new_n4001_;
  assign new_n4003_ = ~pstart_0_ & new_n4002_;
  assign new_n4004_ = pencrypt_0_ & pkey_101_;
  assign new_n4005_ = pstart_0_ & new_n4004_;
  assign new_n4006_ = ~pencrypt_0_ & n_n2433;
  assign new_n4007_ = ~new_n1200_ & new_n4006_;
  assign new_n4008_ = ~pstart_0_ & new_n4007_;
  assign new_n4009_ = pkey_109_ & ~pencrypt_0_;
  assign new_n4010_ = pstart_0_ & new_n4009_;
  assign new_n4011_ = ~n_n2339 & ~new_n1220_;
  assign new_n4012_ = pencrypt_0_ & new_n4011_;
  assign new_n4013_ = n_n2433 & new_n4012_;
  assign new_n4014_ = ~pstart_0_ & new_n4013_;
  assign new_n4015_ = n_n2339 & new_n1220_;
  assign new_n4016_ = pencrypt_0_ & new_n4015_;
  assign new_n4017_ = n_n2433 & new_n4016_;
  assign new_n4018_ = ~pstart_0_ & new_n4017_;
  assign new_n4019_ = ~n_n2433 & ~n_n2339;
  assign new_n4020_ = ~pencrypt_0_ & new_n4019_;
  assign new_n4021_ = new_n1200_ & new_n4020_;
  assign new_n4022_ = ~pstart_0_ & new_n4021_;
  assign new_n4023_ = n_n2339 & ~new_n1220_;
  assign new_n4024_ = pencrypt_0_ & new_n4023_;
  assign new_n4025_ = ~n_n2433 & new_n4024_;
  assign new_n4026_ = ~pstart_0_ & new_n4025_;
  assign new_n4027_ = ~new_n4022_ & ~new_n4026_;
  assign new_n4028_ = ~new_n4014_ & ~new_n4018_;
  assign new_n4029_ = new_n4027_ & new_n4028_;
  assign new_n4030_ = ~new_n4008_ & ~new_n4010_;
  assign new_n4031_ = ~new_n3999_ & ~new_n4003_;
  assign new_n4032_ = ~new_n4005_ & new_n4031_;
  assign new_n4033_ = new_n4030_ & new_n4032_;
  assign n1297 = ~new_n4029_ | ~new_n4033_;
  assign new_n4035_ = ~pencrypt_0_ & n_n2347;
  assign new_n4036_ = ~new_n1200_ & new_n4035_;
  assign new_n4037_ = ~pstart_0_ & new_n4036_;
  assign new_n4038_ = n_n2440 & n_n2347;
  assign new_n4039_ = ~pencrypt_0_ & new_n4038_;
  assign new_n4040_ = new_n1200_ & new_n4039_;
  assign new_n4041_ = ~pstart_0_ & new_n4040_;
  assign new_n4042_ = pkey_110_ & pencrypt_0_;
  assign new_n4043_ = pstart_0_ & new_n4042_;
  assign new_n4044_ = ~pencrypt_0_ & n_n2440;
  assign new_n4045_ = ~new_n1200_ & new_n4044_;
  assign new_n4046_ = ~pstart_0_ & new_n4045_;
  assign new_n4047_ = pkey_118_ & ~pencrypt_0_;
  assign new_n4048_ = pstart_0_ & new_n4047_;
  assign new_n4049_ = ~n_n2347 & ~new_n1220_;
  assign new_n4050_ = pencrypt_0_ & new_n4049_;
  assign new_n4051_ = n_n2440 & new_n4050_;
  assign new_n4052_ = ~pstart_0_ & new_n4051_;
  assign new_n4053_ = n_n2347 & new_n1220_;
  assign new_n4054_ = pencrypt_0_ & new_n4053_;
  assign new_n4055_ = n_n2440 & new_n4054_;
  assign new_n4056_ = ~pstart_0_ & new_n4055_;
  assign new_n4057_ = ~n_n2440 & ~n_n2347;
  assign new_n4058_ = ~pencrypt_0_ & new_n4057_;
  assign new_n4059_ = new_n1200_ & new_n4058_;
  assign new_n4060_ = ~pstart_0_ & new_n4059_;
  assign new_n4061_ = n_n2347 & ~new_n1220_;
  assign new_n4062_ = pencrypt_0_ & new_n4061_;
  assign new_n4063_ = ~n_n2440 & new_n4062_;
  assign new_n4064_ = ~pstart_0_ & new_n4063_;
  assign new_n4065_ = ~new_n4060_ & ~new_n4064_;
  assign new_n4066_ = ~new_n4052_ & ~new_n4056_;
  assign new_n4067_ = new_n4065_ & new_n4066_;
  assign new_n4068_ = ~new_n4046_ & ~new_n4048_;
  assign new_n4069_ = ~new_n4037_ & ~new_n4041_;
  assign new_n4070_ = ~new_n4043_ & new_n4069_;
  assign new_n4071_ = new_n4068_ & new_n4070_;
  assign n1302 = ~new_n4067_ | ~new_n4071_;
  assign new_n4073_ = ~pencrypt_0_ & n_n2379;
  assign new_n4074_ = new_n1200_ & new_n4073_;
  assign new_n4075_ = ~pstart_0_ & new_n4074_;
  assign new_n4076_ = n_n2283 & n_n2379;
  assign new_n4077_ = ~pencrypt_0_ & new_n4076_;
  assign new_n4078_ = ~new_n1200_ & new_n4077_;
  assign new_n4079_ = ~pstart_0_ & new_n4078_;
  assign new_n4080_ = pkey_210_ & pencrypt_0_;
  assign new_n4081_ = pstart_0_ & new_n4080_;
  assign new_n4082_ = ~pencrypt_0_ & n_n2283;
  assign new_n4083_ = new_n1200_ & new_n4082_;
  assign new_n4084_ = ~pstart_0_ & new_n4083_;
  assign new_n4085_ = pkey_218_ & ~pencrypt_0_;
  assign new_n4086_ = pstart_0_ & new_n4085_;
  assign new_n4087_ = n_n2379 & new_n1220_;
  assign new_n4088_ = pencrypt_0_ & new_n4087_;
  assign new_n4089_ = ~n_n2283 & new_n4088_;
  assign new_n4090_ = ~pstart_0_ & new_n4089_;
  assign new_n4091_ = ~n_n2379 & new_n1220_;
  assign new_n4092_ = pencrypt_0_ & new_n4091_;
  assign new_n4093_ = n_n2283 & new_n4092_;
  assign new_n4094_ = ~pstart_0_ & new_n4093_;
  assign new_n4095_ = ~n_n2283 & ~n_n2379;
  assign new_n4096_ = ~pencrypt_0_ & new_n4095_;
  assign new_n4097_ = ~new_n1200_ & new_n4096_;
  assign new_n4098_ = ~pstart_0_ & new_n4097_;
  assign new_n4099_ = n_n2379 & ~new_n1220_;
  assign new_n4100_ = pencrypt_0_ & new_n4099_;
  assign new_n4101_ = n_n2283 & new_n4100_;
  assign new_n4102_ = ~pstart_0_ & new_n4101_;
  assign new_n4103_ = ~new_n4098_ & ~new_n4102_;
  assign new_n4104_ = ~new_n4090_ & ~new_n4094_;
  assign new_n4105_ = new_n4103_ & new_n4104_;
  assign new_n4106_ = ~new_n4084_ & ~new_n4086_;
  assign new_n4107_ = ~new_n4075_ & ~new_n4079_;
  assign new_n4108_ = ~new_n4081_ & new_n4107_;
  assign new_n4109_ = new_n4106_ & new_n4108_;
  assign n1307 = ~new_n4105_ | ~new_n4109_;
  assign new_n4111_ = ~pencrypt_0_ & n_n2303;
  assign new_n4112_ = ~new_n1200_ & new_n4111_;
  assign new_n4113_ = ~pstart_0_ & new_n4112_;
  assign new_n4114_ = n_n2899 & n_n2303;
  assign new_n4115_ = ~pencrypt_0_ & new_n4114_;
  assign new_n4116_ = new_n1200_ & new_n4115_;
  assign new_n4117_ = ~pstart_0_ & new_n4116_;
  assign new_n4118_ = pkey_139_ & pencrypt_0_;
  assign new_n4119_ = pstart_0_ & new_n4118_;
  assign new_n4120_ = ~pencrypt_0_ & n_n2899;
  assign new_n4121_ = ~new_n1200_ & new_n4120_;
  assign new_n4122_ = ~pstart_0_ & new_n4121_;
  assign new_n4123_ = pkey_147_ & ~pencrypt_0_;
  assign new_n4124_ = pstart_0_ & new_n4123_;
  assign new_n4125_ = ~n_n2303 & ~new_n1220_;
  assign new_n4126_ = pencrypt_0_ & new_n4125_;
  assign new_n4127_ = n_n2899 & new_n4126_;
  assign new_n4128_ = ~pstart_0_ & new_n4127_;
  assign new_n4129_ = n_n2303 & new_n1220_;
  assign new_n4130_ = pencrypt_0_ & new_n4129_;
  assign new_n4131_ = n_n2899 & new_n4130_;
  assign new_n4132_ = ~pstart_0_ & new_n4131_;
  assign new_n4133_ = ~n_n2899 & ~n_n2303;
  assign new_n4134_ = ~pencrypt_0_ & new_n4133_;
  assign new_n4135_ = new_n1200_ & new_n4134_;
  assign new_n4136_ = ~pstart_0_ & new_n4135_;
  assign new_n4137_ = n_n2303 & ~new_n1220_;
  assign new_n4138_ = pencrypt_0_ & new_n4137_;
  assign new_n4139_ = ~n_n2899 & new_n4138_;
  assign new_n4140_ = ~pstart_0_ & new_n4139_;
  assign new_n4141_ = ~new_n4136_ & ~new_n4140_;
  assign new_n4142_ = ~new_n4128_ & ~new_n4132_;
  assign new_n4143_ = new_n4141_ & new_n4142_;
  assign new_n4144_ = ~new_n4122_ & ~new_n4124_;
  assign new_n4145_ = ~new_n4113_ & ~new_n4117_;
  assign new_n4146_ = ~new_n4119_ & new_n4145_;
  assign new_n4147_ = new_n4144_ & new_n4146_;
  assign n1312 = ~new_n4143_ | ~new_n4147_;
  assign new_n4149_ = ~pencrypt_0_ & n_n2311;
  assign new_n4150_ = ~new_n1200_ & new_n4149_;
  assign new_n4151_ = ~pstart_0_ & new_n4150_;
  assign new_n4152_ = n_n2406 & n_n2311;
  assign new_n4153_ = ~pencrypt_0_ & new_n4152_;
  assign new_n4154_ = new_n1200_ & new_n4153_;
  assign new_n4155_ = ~pstart_0_ & new_n4154_;
  assign new_n4156_ = pkey_133_ & pencrypt_0_;
  assign new_n4157_ = pstart_0_ & new_n4156_;
  assign new_n4158_ = ~pencrypt_0_ & n_n2406;
  assign new_n4159_ = ~new_n1200_ & new_n4158_;
  assign new_n4160_ = ~pstart_0_ & new_n4159_;
  assign new_n4161_ = pkey_141_ & ~pencrypt_0_;
  assign new_n4162_ = pstart_0_ & new_n4161_;
  assign new_n4163_ = ~n_n2311 & ~new_n1220_;
  assign new_n4164_ = pencrypt_0_ & new_n4163_;
  assign new_n4165_ = n_n2406 & new_n4164_;
  assign new_n4166_ = ~pstart_0_ & new_n4165_;
  assign new_n4167_ = n_n2311 & new_n1220_;
  assign new_n4168_ = pencrypt_0_ & new_n4167_;
  assign new_n4169_ = n_n2406 & new_n4168_;
  assign new_n4170_ = ~pstart_0_ & new_n4169_;
  assign new_n4171_ = ~n_n2406 & ~n_n2311;
  assign new_n4172_ = ~pencrypt_0_ & new_n4171_;
  assign new_n4173_ = new_n1200_ & new_n4172_;
  assign new_n4174_ = ~pstart_0_ & new_n4173_;
  assign new_n4175_ = n_n2311 & ~new_n1220_;
  assign new_n4176_ = pencrypt_0_ & new_n4175_;
  assign new_n4177_ = ~n_n2406 & new_n4176_;
  assign new_n4178_ = ~pstart_0_ & new_n4177_;
  assign new_n4179_ = ~new_n4174_ & ~new_n4178_;
  assign new_n4180_ = ~new_n4166_ & ~new_n4170_;
  assign new_n4181_ = new_n4179_ & new_n4180_;
  assign new_n4182_ = ~new_n4160_ & ~new_n4162_;
  assign new_n4183_ = ~new_n4151_ & ~new_n4155_;
  assign new_n4184_ = ~new_n4157_ & new_n4183_;
  assign new_n4185_ = new_n4182_ & new_n4184_;
  assign n1317 = ~new_n4181_ | ~new_n4185_;
  assign new_n4187_ = ~pencrypt_0_ & n_n2317;
  assign new_n4188_ = ~new_n1200_ & new_n4187_;
  assign new_n4189_ = ~pstart_0_ & new_n4188_;
  assign new_n4190_ = n_n2412 & n_n2317;
  assign new_n4191_ = ~pencrypt_0_ & new_n4190_;
  assign new_n4192_ = new_n1200_ & new_n4191_;
  assign new_n4193_ = ~pstart_0_ & new_n4192_;
  assign new_n4194_ = pencrypt_0_ & pkey_189_;
  assign new_n4195_ = pstart_0_ & new_n4194_;
  assign new_n4196_ = ~pencrypt_0_ & n_n2412;
  assign new_n4197_ = ~new_n1200_ & new_n4196_;
  assign new_n4198_ = ~pstart_0_ & new_n4197_;
  assign new_n4199_ = pkey_134_ & ~pencrypt_0_;
  assign new_n4200_ = pstart_0_ & new_n4199_;
  assign new_n4201_ = ~n_n2317 & ~new_n1220_;
  assign new_n4202_ = pencrypt_0_ & new_n4201_;
  assign new_n4203_ = n_n2412 & new_n4202_;
  assign new_n4204_ = ~pstart_0_ & new_n4203_;
  assign new_n4205_ = n_n2317 & new_n1220_;
  assign new_n4206_ = pencrypt_0_ & new_n4205_;
  assign new_n4207_ = n_n2412 & new_n4206_;
  assign new_n4208_ = ~pstart_0_ & new_n4207_;
  assign new_n4209_ = ~n_n2412 & ~n_n2317;
  assign new_n4210_ = ~pencrypt_0_ & new_n4209_;
  assign new_n4211_ = new_n1200_ & new_n4210_;
  assign new_n4212_ = ~pstart_0_ & new_n4211_;
  assign new_n4213_ = n_n2317 & ~new_n1220_;
  assign new_n4214_ = pencrypt_0_ & new_n4213_;
  assign new_n4215_ = ~n_n2412 & new_n4214_;
  assign new_n4216_ = ~pstart_0_ & new_n4215_;
  assign new_n4217_ = ~new_n4212_ & ~new_n4216_;
  assign new_n4218_ = ~new_n4204_ & ~new_n4208_;
  assign new_n4219_ = new_n4217_ & new_n4218_;
  assign new_n4220_ = ~new_n4198_ & ~new_n4200_;
  assign new_n4221_ = ~new_n4189_ & ~new_n4193_;
  assign new_n4222_ = ~new_n4195_ & new_n4221_;
  assign new_n4223_ = new_n4220_ & new_n4222_;
  assign n1322 = ~new_n4219_ | ~new_n4223_;
  assign new_n4225_ = ~pencrypt_0_ & n_n2802;
  assign new_n4226_ = ~new_n1200_ & new_n4225_;
  assign new_n4227_ = ~pstart_0_ & new_n4226_;
  assign new_n4228_ = n_n2421 & n_n2802;
  assign new_n4229_ = ~pencrypt_0_ & new_n4228_;
  assign new_n4230_ = new_n1200_ & new_n4229_;
  assign new_n4231_ = ~pstart_0_ & new_n4230_;
  assign new_n4232_ = pencrypt_0_ & pkey_83_;
  assign new_n4233_ = pstart_0_ & new_n4232_;
  assign new_n4234_ = ~pencrypt_0_ & n_n2421;
  assign new_n4235_ = ~new_n1200_ & new_n4234_;
  assign new_n4236_ = ~pstart_0_ & new_n4235_;
  assign new_n4237_ = ~pencrypt_0_ & pkey_91_;
  assign new_n4238_ = pstart_0_ & new_n4237_;
  assign new_n4239_ = ~n_n2802 & ~new_n1220_;
  assign new_n4240_ = pencrypt_0_ & new_n4239_;
  assign new_n4241_ = n_n2421 & new_n4240_;
  assign new_n4242_ = ~pstart_0_ & new_n4241_;
  assign new_n4243_ = n_n2802 & new_n1220_;
  assign new_n4244_ = pencrypt_0_ & new_n4243_;
  assign new_n4245_ = n_n2421 & new_n4244_;
  assign new_n4246_ = ~pstart_0_ & new_n4245_;
  assign new_n4247_ = ~n_n2421 & ~n_n2802;
  assign new_n4248_ = ~pencrypt_0_ & new_n4247_;
  assign new_n4249_ = new_n1200_ & new_n4248_;
  assign new_n4250_ = ~pstart_0_ & new_n4249_;
  assign new_n4251_ = n_n2802 & ~new_n1220_;
  assign new_n4252_ = pencrypt_0_ & new_n4251_;
  assign new_n4253_ = ~n_n2421 & new_n4252_;
  assign new_n4254_ = ~pstart_0_ & new_n4253_;
  assign new_n4255_ = ~new_n4250_ & ~new_n4254_;
  assign new_n4256_ = ~new_n4242_ & ~new_n4246_;
  assign new_n4257_ = new_n4255_ & new_n4256_;
  assign new_n4258_ = ~new_n4236_ & ~new_n4238_;
  assign new_n4259_ = ~new_n4227_ & ~new_n4231_;
  assign new_n4260_ = ~new_n4233_ & new_n4259_;
  assign new_n4261_ = new_n4258_ & new_n4260_;
  assign n1327 = ~new_n4257_ | ~new_n4261_;
  assign new_n4263_ = ~pencrypt_0_ & n_n2340;
  assign new_n4264_ = ~new_n1200_ & new_n4263_;
  assign new_n4265_ = ~pstart_0_ & new_n4264_;
  assign new_n4266_ = n_n2950 & n_n2340;
  assign new_n4267_ = ~pencrypt_0_ & new_n4266_;
  assign new_n4268_ = new_n1200_ & new_n4267_;
  assign new_n4269_ = ~pstart_0_ & new_n4268_;
  assign new_n4270_ = pkey_109_ & pencrypt_0_;
  assign new_n4271_ = pstart_0_ & new_n4270_;
  assign new_n4272_ = ~pencrypt_0_ & n_n2950;
  assign new_n4273_ = ~new_n1200_ & new_n4272_;
  assign new_n4274_ = ~pstart_0_ & new_n4273_;
  assign new_n4275_ = pkey_117_ & ~pencrypt_0_;
  assign new_n4276_ = pstart_0_ & new_n4275_;
  assign new_n4277_ = ~n_n2340 & ~new_n1220_;
  assign new_n4278_ = pencrypt_0_ & new_n4277_;
  assign new_n4279_ = n_n2950 & new_n4278_;
  assign new_n4280_ = ~pstart_0_ & new_n4279_;
  assign new_n4281_ = n_n2340 & new_n1220_;
  assign new_n4282_ = pencrypt_0_ & new_n4281_;
  assign new_n4283_ = n_n2950 & new_n4282_;
  assign new_n4284_ = ~pstart_0_ & new_n4283_;
  assign new_n4285_ = ~n_n2950 & ~n_n2340;
  assign new_n4286_ = ~pencrypt_0_ & new_n4285_;
  assign new_n4287_ = new_n1200_ & new_n4286_;
  assign new_n4288_ = ~pstart_0_ & new_n4287_;
  assign new_n4289_ = n_n2340 & ~new_n1220_;
  assign new_n4290_ = pencrypt_0_ & new_n4289_;
  assign new_n4291_ = ~n_n2950 & new_n4290_;
  assign new_n4292_ = ~pstart_0_ & new_n4291_;
  assign new_n4293_ = ~new_n4288_ & ~new_n4292_;
  assign new_n4294_ = ~new_n4280_ & ~new_n4284_;
  assign new_n4295_ = new_n4293_ & new_n4294_;
  assign new_n4296_ = ~new_n4274_ & ~new_n4276_;
  assign new_n4297_ = ~new_n4265_ & ~new_n4269_;
  assign new_n4298_ = ~new_n4271_ & new_n4297_;
  assign new_n4299_ = new_n4296_ & new_n4298_;
  assign n1332 = ~new_n4295_ | ~new_n4299_;
  assign new_n4301_ = ~pencrypt_0_ & n_n2350;
  assign new_n4302_ = ~new_n1200_ & new_n4301_;
  assign new_n4303_ = ~pstart_0_ & new_n4302_;
  assign new_n4304_ = n_n2443 & n_n2350;
  assign new_n4305_ = ~pencrypt_0_ & new_n4304_;
  assign new_n4306_ = new_n1200_ & new_n4305_;
  assign new_n4307_ = ~pstart_0_ & new_n4306_;
  assign new_n4308_ = pkey_3_ & pencrypt_0_;
  assign new_n4309_ = pstart_0_ & new_n4308_;
  assign new_n4310_ = ~pencrypt_0_ & n_n2443;
  assign new_n4311_ = ~new_n1200_ & new_n4310_;
  assign new_n4312_ = ~pstart_0_ & new_n4311_;
  assign new_n4313_ = ~pencrypt_0_ & pkey_11_;
  assign new_n4314_ = pstart_0_ & new_n4313_;
  assign new_n4315_ = ~n_n2350 & ~new_n1220_;
  assign new_n4316_ = pencrypt_0_ & new_n4315_;
  assign new_n4317_ = n_n2443 & new_n4316_;
  assign new_n4318_ = ~pstart_0_ & new_n4317_;
  assign new_n4319_ = n_n2350 & new_n1220_;
  assign new_n4320_ = pencrypt_0_ & new_n4319_;
  assign new_n4321_ = n_n2443 & new_n4320_;
  assign new_n4322_ = ~pstart_0_ & new_n4321_;
  assign new_n4323_ = ~n_n2443 & ~n_n2350;
  assign new_n4324_ = ~pencrypt_0_ & new_n4323_;
  assign new_n4325_ = new_n1200_ & new_n4324_;
  assign new_n4326_ = ~pstart_0_ & new_n4325_;
  assign new_n4327_ = n_n2350 & ~new_n1220_;
  assign new_n4328_ = pencrypt_0_ & new_n4327_;
  assign new_n4329_ = ~n_n2443 & new_n4328_;
  assign new_n4330_ = ~pstart_0_ & new_n4329_;
  assign new_n4331_ = ~new_n4326_ & ~new_n4330_;
  assign new_n4332_ = ~new_n4318_ & ~new_n4322_;
  assign new_n4333_ = new_n4331_ & new_n4332_;
  assign new_n4334_ = ~new_n4312_ & ~new_n4314_;
  assign new_n4335_ = ~new_n4303_ & ~new_n4307_;
  assign new_n4336_ = ~new_n4309_ & new_n4335_;
  assign new_n4337_ = new_n4334_ & new_n4336_;
  assign n1337 = ~new_n4333_ | ~new_n4337_;
  assign new_n4339_ = new_n1200_ & new_n3160_;
  assign new_n4340_ = ~pstart_0_ & new_n4339_;
  assign new_n4341_ = ~new_n1200_ & new_n3155_;
  assign new_n4342_ = ~pstart_0_ & new_n4341_;
  assign new_n4343_ = pkey_218_ & pencrypt_0_;
  assign new_n4344_ = pstart_0_ & new_n4343_;
  assign new_n4345_ = new_n1200_ & new_n3151_;
  assign new_n4346_ = ~pstart_0_ & new_n4345_;
  assign new_n4347_ = pkey_226_ & ~pencrypt_0_;
  assign new_n4348_ = pstart_0_ & new_n4347_;
  assign new_n4349_ = n_n2380 & new_n1220_;
  assign new_n4350_ = pencrypt_0_ & new_n4349_;
  assign new_n4351_ = ~n_n2284 & new_n4350_;
  assign new_n4352_ = ~pstart_0_ & new_n4351_;
  assign new_n4353_ = ~n_n2380 & new_n1220_;
  assign new_n4354_ = pencrypt_0_ & new_n4353_;
  assign new_n4355_ = n_n2284 & new_n4354_;
  assign new_n4356_ = ~pstart_0_ & new_n4355_;
  assign new_n4357_ = ~new_n1200_ & new_n3174_;
  assign new_n4358_ = ~pstart_0_ & new_n4357_;
  assign new_n4359_ = n_n2380 & ~new_n1220_;
  assign new_n4360_ = pencrypt_0_ & new_n4359_;
  assign new_n4361_ = n_n2284 & new_n4360_;
  assign new_n4362_ = ~pstart_0_ & new_n4361_;
  assign new_n4363_ = ~new_n4358_ & ~new_n4362_;
  assign new_n4364_ = ~new_n4352_ & ~new_n4356_;
  assign new_n4365_ = new_n4363_ & new_n4364_;
  assign new_n4366_ = ~new_n4346_ & ~new_n4348_;
  assign new_n4367_ = ~new_n4340_ & ~new_n4342_;
  assign new_n4368_ = ~new_n4344_ & new_n4367_;
  assign new_n4369_ = new_n4366_ & new_n4368_;
  assign n1342 = ~new_n4365_ | ~new_n4369_;
  assign new_n4371_ = ~pencrypt_0_ & n_n2770;
  assign new_n4372_ = ~new_n1200_ & new_n4371_;
  assign new_n4373_ = ~pstart_0_ & new_n4372_;
  assign new_n4374_ = n_n2397 & n_n2770;
  assign new_n4375_ = ~pencrypt_0_ & new_n4374_;
  assign new_n4376_ = new_n1200_ & new_n4375_;
  assign new_n4377_ = ~pstart_0_ & new_n4376_;
  assign new_n4378_ = pkey_147_ & pencrypt_0_;
  assign new_n4379_ = pstart_0_ & new_n4378_;
  assign new_n4380_ = ~pencrypt_0_ & n_n2397;
  assign new_n4381_ = ~new_n1200_ & new_n4380_;
  assign new_n4382_ = ~pstart_0_ & new_n4381_;
  assign new_n4383_ = pkey_155_ & ~pencrypt_0_;
  assign new_n4384_ = pstart_0_ & new_n4383_;
  assign new_n4385_ = ~n_n2770 & ~new_n1220_;
  assign new_n4386_ = pencrypt_0_ & new_n4385_;
  assign new_n4387_ = n_n2397 & new_n4386_;
  assign new_n4388_ = ~pstart_0_ & new_n4387_;
  assign new_n4389_ = n_n2770 & new_n1220_;
  assign new_n4390_ = pencrypt_0_ & new_n4389_;
  assign new_n4391_ = n_n2397 & new_n4390_;
  assign new_n4392_ = ~pstart_0_ & new_n4391_;
  assign new_n4393_ = ~n_n2397 & ~n_n2770;
  assign new_n4394_ = ~pencrypt_0_ & new_n4393_;
  assign new_n4395_ = new_n1200_ & new_n4394_;
  assign new_n4396_ = ~pstart_0_ & new_n4395_;
  assign new_n4397_ = n_n2770 & ~new_n1220_;
  assign new_n4398_ = pencrypt_0_ & new_n4397_;
  assign new_n4399_ = ~n_n2397 & new_n4398_;
  assign new_n4400_ = ~pstart_0_ & new_n4399_;
  assign new_n4401_ = ~new_n4396_ & ~new_n4400_;
  assign new_n4402_ = ~new_n4388_ & ~new_n4392_;
  assign new_n4403_ = new_n4401_ & new_n4402_;
  assign new_n4404_ = ~new_n4382_ & ~new_n4384_;
  assign new_n4405_ = ~new_n4373_ & ~new_n4377_;
  assign new_n4406_ = ~new_n4379_ & new_n4405_;
  assign new_n4407_ = new_n4404_ & new_n4406_;
  assign n1347 = ~new_n4403_ | ~new_n4407_;
  assign new_n4409_ = ~pencrypt_0_ & n_n2310;
  assign new_n4410_ = ~new_n1200_ & new_n4409_;
  assign new_n4411_ = ~pstart_0_ & new_n4410_;
  assign new_n4412_ = n_n2405 & n_n2310;
  assign new_n4413_ = ~pencrypt_0_ & new_n4412_;
  assign new_n4414_ = new_n1200_ & new_n4413_;
  assign new_n4415_ = ~pstart_0_ & new_n4414_;
  assign new_n4416_ = pencrypt_0_ & pkey_188_;
  assign new_n4417_ = pstart_0_ & new_n4416_;
  assign new_n4418_ = ~pencrypt_0_ & n_n2405;
  assign new_n4419_ = ~new_n1200_ & new_n4418_;
  assign new_n4420_ = ~pstart_0_ & new_n4419_;
  assign new_n4421_ = pkey_133_ & ~pencrypt_0_;
  assign new_n4422_ = pstart_0_ & new_n4421_;
  assign new_n4423_ = ~n_n2310 & ~new_n1220_;
  assign new_n4424_ = pencrypt_0_ & new_n4423_;
  assign new_n4425_ = n_n2405 & new_n4424_;
  assign new_n4426_ = ~pstart_0_ & new_n4425_;
  assign new_n4427_ = n_n2310 & new_n1220_;
  assign new_n4428_ = pencrypt_0_ & new_n4427_;
  assign new_n4429_ = n_n2405 & new_n4428_;
  assign new_n4430_ = ~pstart_0_ & new_n4429_;
  assign new_n4431_ = ~n_n2405 & ~n_n2310;
  assign new_n4432_ = ~pencrypt_0_ & new_n4431_;
  assign new_n4433_ = new_n1200_ & new_n4432_;
  assign new_n4434_ = ~pstart_0_ & new_n4433_;
  assign new_n4435_ = n_n2310 & ~new_n1220_;
  assign new_n4436_ = pencrypt_0_ & new_n4435_;
  assign new_n4437_ = ~n_n2405 & new_n4436_;
  assign new_n4438_ = ~pstart_0_ & new_n4437_;
  assign new_n4439_ = ~new_n4434_ & ~new_n4438_;
  assign new_n4440_ = ~new_n4426_ & ~new_n4430_;
  assign new_n4441_ = new_n4439_ & new_n4440_;
  assign new_n4442_ = ~new_n4420_ & ~new_n4422_;
  assign new_n4443_ = ~new_n4411_ & ~new_n4415_;
  assign new_n4444_ = ~new_n4417_ & new_n4443_;
  assign new_n4445_ = new_n4442_ & new_n4444_;
  assign n1352 = ~new_n4441_ | ~new_n4445_;
  assign new_n4447_ = ~pencrypt_0_ & n_n2318;
  assign new_n4448_ = ~new_n1200_ & new_n4447_;
  assign new_n4449_ = ~pstart_0_ & new_n4448_;
  assign new_n4450_ = n_n2921 & n_n2318;
  assign new_n4451_ = ~pencrypt_0_ & new_n4450_;
  assign new_n4452_ = new_n1200_ & new_n4451_;
  assign new_n4453_ = ~pstart_0_ & new_n4452_;
  assign new_n4454_ = pkey_134_ & pencrypt_0_;
  assign new_n4455_ = pstart_0_ & new_n4454_;
  assign new_n4456_ = ~pencrypt_0_ & n_n2921;
  assign new_n4457_ = ~new_n1200_ & new_n4456_;
  assign new_n4458_ = ~pstart_0_ & new_n4457_;
  assign new_n4459_ = pkey_142_ & ~pencrypt_0_;
  assign new_n4460_ = pstart_0_ & new_n4459_;
  assign new_n4461_ = ~n_n2318 & ~new_n1220_;
  assign new_n4462_ = pencrypt_0_ & new_n4461_;
  assign new_n4463_ = n_n2921 & new_n4462_;
  assign new_n4464_ = ~pstart_0_ & new_n4463_;
  assign new_n4465_ = n_n2318 & new_n1220_;
  assign new_n4466_ = pencrypt_0_ & new_n4465_;
  assign new_n4467_ = n_n2921 & new_n4466_;
  assign new_n4468_ = ~pstart_0_ & new_n4467_;
  assign new_n4469_ = ~n_n2921 & ~n_n2318;
  assign new_n4470_ = ~pencrypt_0_ & new_n4469_;
  assign new_n4471_ = new_n1200_ & new_n4470_;
  assign new_n4472_ = ~pstart_0_ & new_n4471_;
  assign new_n4473_ = n_n2318 & ~new_n1220_;
  assign new_n4474_ = pencrypt_0_ & new_n4473_;
  assign new_n4475_ = ~n_n2921 & new_n4474_;
  assign new_n4476_ = ~pstart_0_ & new_n4475_;
  assign new_n4477_ = ~new_n4472_ & ~new_n4476_;
  assign new_n4478_ = ~new_n4464_ & ~new_n4468_;
  assign new_n4479_ = new_n4477_ & new_n4478_;
  assign new_n4480_ = ~new_n4458_ & ~new_n4460_;
  assign new_n4481_ = ~new_n4449_ & ~new_n4453_;
  assign new_n4482_ = ~new_n4455_ & new_n4481_;
  assign new_n4483_ = new_n4480_ & new_n4482_;
  assign n1357 = ~new_n4479_ | ~new_n4483_;
  assign new_n4485_ = ~pencrypt_0_ & n_n2327;
  assign new_n4486_ = ~new_n1200_ & new_n4485_;
  assign new_n4487_ = ~pstart_0_ & new_n4486_;
  assign new_n4488_ = n_n2931 & n_n2327;
  assign new_n4489_ = ~pencrypt_0_ & new_n4488_;
  assign new_n4490_ = new_n1200_ & new_n4489_;
  assign new_n4491_ = ~pstart_0_ & new_n4490_;
  assign new_n4492_ = pencrypt_0_ & pkey_75_;
  assign new_n4493_ = pstart_0_ & new_n4492_;
  assign new_n4494_ = ~pencrypt_0_ & n_n2931;
  assign new_n4495_ = ~new_n1200_ & new_n4494_;
  assign new_n4496_ = ~pstart_0_ & new_n4495_;
  assign new_n4497_ = ~pencrypt_0_ & pkey_83_;
  assign new_n4498_ = pstart_0_ & new_n4497_;
  assign new_n4499_ = ~n_n2327 & ~new_n1220_;
  assign new_n4500_ = pencrypt_0_ & new_n4499_;
  assign new_n4501_ = n_n2931 & new_n4500_;
  assign new_n4502_ = ~pstart_0_ & new_n4501_;
  assign new_n4503_ = n_n2327 & new_n1220_;
  assign new_n4504_ = pencrypt_0_ & new_n4503_;
  assign new_n4505_ = n_n2931 & new_n4504_;
  assign new_n4506_ = ~pstart_0_ & new_n4505_;
  assign new_n4507_ = ~n_n2931 & ~n_n2327;
  assign new_n4508_ = ~pencrypt_0_ & new_n4507_;
  assign new_n4509_ = new_n1200_ & new_n4508_;
  assign new_n4510_ = ~pstart_0_ & new_n4509_;
  assign new_n4511_ = n_n2327 & ~new_n1220_;
  assign new_n4512_ = pencrypt_0_ & new_n4511_;
  assign new_n4513_ = ~n_n2931 & new_n4512_;
  assign new_n4514_ = ~pstart_0_ & new_n4513_;
  assign new_n4515_ = ~new_n4510_ & ~new_n4514_;
  assign new_n4516_ = ~new_n4502_ & ~new_n4506_;
  assign new_n4517_ = new_n4515_ & new_n4516_;
  assign new_n4518_ = ~new_n4496_ & ~new_n4498_;
  assign new_n4519_ = ~new_n4487_ & ~new_n4491_;
  assign new_n4520_ = ~new_n4493_ & new_n4519_;
  assign new_n4521_ = new_n4518_ & new_n4520_;
  assign n1362 = ~new_n4517_ | ~new_n4521_;
  assign new_n4523_ = ~pencrypt_0_ & n_n2821;
  assign new_n4524_ = ~new_n1200_ & new_n4523_;
  assign new_n4525_ = ~pstart_0_ & new_n4524_;
  assign new_n4526_ = n_n2434 & n_n2821;
  assign new_n4527_ = ~pencrypt_0_ & new_n4526_;
  assign new_n4528_ = new_n1200_ & new_n4527_;
  assign new_n4529_ = ~pstart_0_ & new_n4528_;
  assign new_n4530_ = pkey_117_ & pencrypt_0_;
  assign new_n4531_ = pstart_0_ & new_n4530_;
  assign new_n4532_ = ~pencrypt_0_ & n_n2434;
  assign new_n4533_ = ~new_n1200_ & new_n4532_;
  assign new_n4534_ = ~pstart_0_ & new_n4533_;
  assign new_n4535_ = pkey_125_ & ~pencrypt_0_;
  assign new_n4536_ = pstart_0_ & new_n4535_;
  assign new_n4537_ = ~n_n2821 & ~new_n1220_;
  assign new_n4538_ = pencrypt_0_ & new_n4537_;
  assign new_n4539_ = n_n2434 & new_n4538_;
  assign new_n4540_ = ~pstart_0_ & new_n4539_;
  assign new_n4541_ = n_n2821 & new_n1220_;
  assign new_n4542_ = pencrypt_0_ & new_n4541_;
  assign new_n4543_ = n_n2434 & new_n4542_;
  assign new_n4544_ = ~pstart_0_ & new_n4543_;
  assign new_n4545_ = ~n_n2434 & ~n_n2821;
  assign new_n4546_ = ~pencrypt_0_ & new_n4545_;
  assign new_n4547_ = new_n1200_ & new_n4546_;
  assign new_n4548_ = ~pstart_0_ & new_n4547_;
  assign new_n4549_ = n_n2821 & ~new_n1220_;
  assign new_n4550_ = pencrypt_0_ & new_n4549_;
  assign new_n4551_ = ~n_n2434 & new_n4550_;
  assign new_n4552_ = ~pstart_0_ & new_n4551_;
  assign new_n4553_ = ~new_n4548_ & ~new_n4552_;
  assign new_n4554_ = ~new_n4540_ & ~new_n4544_;
  assign new_n4555_ = new_n4553_ & new_n4554_;
  assign new_n4556_ = ~new_n4534_ & ~new_n4536_;
  assign new_n4557_ = ~new_n4525_ & ~new_n4529_;
  assign new_n4558_ = ~new_n4531_ & new_n4557_;
  assign new_n4559_ = new_n4556_ & new_n4558_;
  assign n1367 = ~new_n4555_ | ~new_n4559_;
  assign new_n4561_ = ~pencrypt_0_ & n_n2349;
  assign new_n4562_ = ~new_n1200_ & new_n4561_;
  assign new_n4563_ = ~pstart_0_ & new_n4562_;
  assign new_n4564_ = n_n2442 & n_n2349;
  assign new_n4565_ = ~pencrypt_0_ & new_n4564_;
  assign new_n4566_ = new_n1200_ & new_n4565_;
  assign new_n4567_ = ~pstart_0_ & new_n4566_;
  assign new_n4568_ = pkey_126_ & pencrypt_0_;
  assign new_n4569_ = pstart_0_ & new_n4568_;
  assign new_n4570_ = ~pencrypt_0_ & n_n2442;
  assign new_n4571_ = ~new_n1200_ & new_n4570_;
  assign new_n4572_ = ~pstart_0_ & new_n4571_;
  assign new_n4573_ = pkey_3_ & ~pencrypt_0_;
  assign new_n4574_ = pstart_0_ & new_n4573_;
  assign new_n4575_ = ~n_n2349 & ~new_n1220_;
  assign new_n4576_ = pencrypt_0_ & new_n4575_;
  assign new_n4577_ = n_n2442 & new_n4576_;
  assign new_n4578_ = ~pstart_0_ & new_n4577_;
  assign new_n4579_ = n_n2349 & new_n1220_;
  assign new_n4580_ = pencrypt_0_ & new_n4579_;
  assign new_n4581_ = n_n2442 & new_n4580_;
  assign new_n4582_ = ~pstart_0_ & new_n4581_;
  assign new_n4583_ = ~n_n2442 & ~n_n2349;
  assign new_n4584_ = ~pencrypt_0_ & new_n4583_;
  assign new_n4585_ = new_n1200_ & new_n4584_;
  assign new_n4586_ = ~pstart_0_ & new_n4585_;
  assign new_n4587_ = n_n2349 & ~new_n1220_;
  assign new_n4588_ = pencrypt_0_ & new_n4587_;
  assign new_n4589_ = ~n_n2442 & new_n4588_;
  assign new_n4590_ = ~pstart_0_ & new_n4589_;
  assign new_n4591_ = ~new_n4586_ & ~new_n4590_;
  assign new_n4592_ = ~new_n4578_ & ~new_n4582_;
  assign new_n4593_ = new_n4591_ & new_n4592_;
  assign new_n4594_ = ~new_n4572_ & ~new_n4574_;
  assign new_n4595_ = ~new_n4563_ & ~new_n4567_;
  assign new_n4596_ = ~new_n4569_ & new_n4595_;
  assign new_n4597_ = new_n4594_ & new_n4596_;
  assign n1372 = ~new_n4593_ | ~new_n4597_;
  assign new_n4599_ = new_n1200_ & new_n3122_;
  assign new_n4600_ = ~pstart_0_ & new_n4599_;
  assign new_n4601_ = ~new_n1200_ & new_n3117_;
  assign new_n4602_ = ~pstart_0_ & new_n4601_;
  assign new_n4603_ = pkey_227_ & pencrypt_0_;
  assign new_n4604_ = pstart_0_ & new_n4603_;
  assign new_n4605_ = new_n1200_ & new_n3113_;
  assign new_n4606_ = ~pstart_0_ & new_n4605_;
  assign new_n4607_ = pkey_235_ & ~pencrypt_0_;
  assign new_n4608_ = pstart_0_ & new_n4607_;
  assign new_n4609_ = n_n2374 & new_n1220_;
  assign new_n4610_ = pencrypt_0_ & new_n4609_;
  assign new_n4611_ = ~n_n2279 & new_n4610_;
  assign new_n4612_ = ~pstart_0_ & new_n4611_;
  assign new_n4613_ = ~n_n2374 & new_n1220_;
  assign new_n4614_ = pencrypt_0_ & new_n4613_;
  assign new_n4615_ = n_n2279 & new_n4614_;
  assign new_n4616_ = ~pstart_0_ & new_n4615_;
  assign new_n4617_ = ~new_n1200_ & new_n3136_;
  assign new_n4618_ = ~pstart_0_ & new_n4617_;
  assign new_n4619_ = n_n2374 & ~new_n1220_;
  assign new_n4620_ = pencrypt_0_ & new_n4619_;
  assign new_n4621_ = n_n2279 & new_n4620_;
  assign new_n4622_ = ~pstart_0_ & new_n4621_;
  assign new_n4623_ = ~new_n4618_ & ~new_n4622_;
  assign new_n4624_ = ~new_n4612_ & ~new_n4616_;
  assign new_n4625_ = new_n4623_ & new_n4624_;
  assign new_n4626_ = ~new_n4606_ & ~new_n4608_;
  assign new_n4627_ = ~new_n4600_ & ~new_n4602_;
  assign new_n4628_ = ~new_n4604_ & new_n4627_;
  assign new_n4629_ = new_n4626_ & new_n4628_;
  assign n1377 = ~new_n4625_ | ~new_n4629_;
  assign new_n4631_ = new_n1200_ & new_n3520_;
  assign new_n4632_ = ~pstart_0_ & new_n4631_;
  assign new_n4633_ = ~new_n1200_ & new_n3515_;
  assign new_n4634_ = ~pstart_0_ & new_n4633_;
  assign new_n4635_ = pencrypt_0_ & pkey_24_;
  assign new_n4636_ = pstart_0_ & new_n4635_;
  assign new_n4637_ = new_n1200_ & new_n3511_;
  assign new_n4638_ = ~pstart_0_ & new_n4637_;
  assign new_n4639_ = ~pencrypt_0_ & pkey_32_;
  assign new_n4640_ = pstart_0_ & new_n4639_;
  assign new_n4641_ = n_n2462 & new_n1220_;
  assign new_n4642_ = pencrypt_0_ & new_n4641_;
  assign new_n4643_ = ~n_n2369 & new_n4642_;
  assign new_n4644_ = ~pstart_0_ & new_n4643_;
  assign new_n4645_ = ~n_n2462 & new_n1220_;
  assign new_n4646_ = pencrypt_0_ & new_n4645_;
  assign new_n4647_ = n_n2369 & new_n4646_;
  assign new_n4648_ = ~pstart_0_ & new_n4647_;
  assign new_n4649_ = ~new_n1200_ & new_n3534_;
  assign new_n4650_ = ~pstart_0_ & new_n4649_;
  assign new_n4651_ = n_n2462 & ~new_n1220_;
  assign new_n4652_ = pencrypt_0_ & new_n4651_;
  assign new_n4653_ = n_n2369 & new_n4652_;
  assign new_n4654_ = ~pstart_0_ & new_n4653_;
  assign new_n4655_ = ~new_n4650_ & ~new_n4654_;
  assign new_n4656_ = ~new_n4644_ & ~new_n4648_;
  assign new_n4657_ = new_n4655_ & new_n4656_;
  assign new_n4658_ = ~new_n4638_ & ~new_n4640_;
  assign new_n4659_ = ~new_n4632_ & ~new_n4634_;
  assign new_n4660_ = ~new_n4636_ & new_n4659_;
  assign new_n4661_ = new_n4658_ & new_n4660_;
  assign n1382 = ~new_n4657_ | ~new_n4661_;
  assign new_n4663_ = ~new_n1200_ & new_n4082_;
  assign new_n4664_ = ~pstart_0_ & new_n4663_;
  assign new_n4665_ = new_n1200_ & new_n4077_;
  assign new_n4666_ = ~pstart_0_ & new_n4665_;
  assign new_n4667_ = pkey_212_ & pencrypt_0_;
  assign new_n4668_ = pstart_0_ & new_n4667_;
  assign new_n4669_ = ~new_n1200_ & new_n4073_;
  assign new_n4670_ = ~pstart_0_ & new_n4669_;
  assign new_n4671_ = pkey_220_ & ~pencrypt_0_;
  assign new_n4672_ = pstart_0_ & new_n4671_;
  assign new_n4673_ = ~n_n2283 & ~new_n1220_;
  assign new_n4674_ = pencrypt_0_ & new_n4673_;
  assign new_n4675_ = n_n2379 & new_n4674_;
  assign new_n4676_ = ~pstart_0_ & new_n4675_;
  assign new_n4677_ = n_n2283 & new_n1220_;
  assign new_n4678_ = pencrypt_0_ & new_n4677_;
  assign new_n4679_ = n_n2379 & new_n4678_;
  assign new_n4680_ = ~pstart_0_ & new_n4679_;
  assign new_n4681_ = new_n1200_ & new_n4096_;
  assign new_n4682_ = ~pstart_0_ & new_n4681_;
  assign new_n4683_ = n_n2283 & ~new_n1220_;
  assign new_n4684_ = pencrypt_0_ & new_n4683_;
  assign new_n4685_ = ~n_n2379 & new_n4684_;
  assign new_n4686_ = ~pstart_0_ & new_n4685_;
  assign new_n4687_ = ~new_n4682_ & ~new_n4686_;
  assign new_n4688_ = ~new_n4676_ & ~new_n4680_;
  assign new_n4689_ = new_n4687_ & new_n4688_;
  assign new_n4690_ = ~new_n4670_ & ~new_n4672_;
  assign new_n4691_ = ~new_n4664_ & ~new_n4666_;
  assign new_n4692_ = ~new_n4668_ & new_n4691_;
  assign new_n4693_ = new_n4690_ & new_n4692_;
  assign n1387 = ~new_n4689_ | ~new_n4693_;
  assign new_n4695_ = ~pencrypt_0_ & n_n2304;
  assign new_n4696_ = ~new_n1200_ & new_n4695_;
  assign new_n4697_ = ~pstart_0_ & new_n4696_;
  assign new_n4698_ = n_n2398 & n_n2304;
  assign new_n4699_ = ~pencrypt_0_ & new_n4698_;
  assign new_n4700_ = new_n1200_ & new_n4699_;
  assign new_n4701_ = ~pstart_0_ & new_n4700_;
  assign new_n4702_ = pkey_155_ & pencrypt_0_;
  assign new_n4703_ = pstart_0_ & new_n4702_;
  assign new_n4704_ = ~pencrypt_0_ & n_n2398;
  assign new_n4705_ = ~new_n1200_ & new_n4704_;
  assign new_n4706_ = ~pstart_0_ & new_n4705_;
  assign new_n4707_ = pkey_132_ & ~pencrypt_0_;
  assign new_n4708_ = pstart_0_ & new_n4707_;
  assign new_n4709_ = ~n_n2304 & ~new_n1220_;
  assign new_n4710_ = pencrypt_0_ & new_n4709_;
  assign new_n4711_ = n_n2398 & new_n4710_;
  assign new_n4712_ = ~pstart_0_ & new_n4711_;
  assign new_n4713_ = n_n2304 & new_n1220_;
  assign new_n4714_ = pencrypt_0_ & new_n4713_;
  assign new_n4715_ = n_n2398 & new_n4714_;
  assign new_n4716_ = ~pstart_0_ & new_n4715_;
  assign new_n4717_ = ~n_n2398 & ~n_n2304;
  assign new_n4718_ = ~pencrypt_0_ & new_n4717_;
  assign new_n4719_ = new_n1200_ & new_n4718_;
  assign new_n4720_ = ~pstart_0_ & new_n4719_;
  assign new_n4721_ = n_n2304 & ~new_n1220_;
  assign new_n4722_ = pencrypt_0_ & new_n4721_;
  assign new_n4723_ = ~n_n2398 & new_n4722_;
  assign new_n4724_ = ~pstart_0_ & new_n4723_;
  assign new_n4725_ = ~new_n4720_ & ~new_n4724_;
  assign new_n4726_ = ~new_n4712_ & ~new_n4716_;
  assign new_n4727_ = new_n4725_ & new_n4726_;
  assign new_n4728_ = ~new_n4706_ & ~new_n4708_;
  assign new_n4729_ = ~new_n4697_ & ~new_n4701_;
  assign new_n4730_ = ~new_n4703_ & new_n4729_;
  assign new_n4731_ = new_n4728_ & new_n4730_;
  assign n1392 = ~new_n4727_ | ~new_n4731_;
  assign new_n4733_ = ~pencrypt_0_ & n_n2313;
  assign new_n4734_ = ~new_n1200_ & new_n4733_;
  assign new_n4735_ = ~pstart_0_ & new_n4734_;
  assign new_n4736_ = n_n2408 & n_n2313;
  assign new_n4737_ = ~pencrypt_0_ & new_n4736_;
  assign new_n4738_ = new_n1200_ & new_n4737_;
  assign new_n4739_ = ~pstart_0_ & new_n4738_;
  assign new_n4740_ = pkey_149_ & pencrypt_0_;
  assign new_n4741_ = pstart_0_ & new_n4740_;
  assign new_n4742_ = ~pencrypt_0_ & n_n2408;
  assign new_n4743_ = ~new_n1200_ & new_n4742_;
  assign new_n4744_ = ~pstart_0_ & new_n4743_;
  assign new_n4745_ = pkey_157_ & ~pencrypt_0_;
  assign new_n4746_ = pstart_0_ & new_n4745_;
  assign new_n4747_ = ~n_n2313 & ~new_n1220_;
  assign new_n4748_ = pencrypt_0_ & new_n4747_;
  assign new_n4749_ = n_n2408 & new_n4748_;
  assign new_n4750_ = ~pstart_0_ & new_n4749_;
  assign new_n4751_ = n_n2313 & new_n1220_;
  assign new_n4752_ = pencrypt_0_ & new_n4751_;
  assign new_n4753_ = n_n2408 & new_n4752_;
  assign new_n4754_ = ~pstart_0_ & new_n4753_;
  assign new_n4755_ = ~n_n2408 & ~n_n2313;
  assign new_n4756_ = ~pencrypt_0_ & new_n4755_;
  assign new_n4757_ = new_n1200_ & new_n4756_;
  assign new_n4758_ = ~pstart_0_ & new_n4757_;
  assign new_n4759_ = n_n2313 & ~new_n1220_;
  assign new_n4760_ = pencrypt_0_ & new_n4759_;
  assign new_n4761_ = ~n_n2408 & new_n4760_;
  assign new_n4762_ = ~pstart_0_ & new_n4761_;
  assign new_n4763_ = ~new_n4758_ & ~new_n4762_;
  assign new_n4764_ = ~new_n4750_ & ~new_n4754_;
  assign new_n4765_ = new_n4763_ & new_n4764_;
  assign new_n4766_ = ~new_n4744_ & ~new_n4746_;
  assign new_n4767_ = ~new_n4735_ & ~new_n4739_;
  assign new_n4768_ = ~new_n4741_ & new_n4767_;
  assign new_n4769_ = new_n4766_ & new_n4768_;
  assign n1397 = ~new_n4765_ | ~new_n4769_;
  assign new_n4771_ = ~pencrypt_0_ & n_n2323;
  assign new_n4772_ = ~new_n1200_ & new_n4771_;
  assign new_n4773_ = ~pstart_0_ & new_n4772_;
  assign new_n4774_ = n_n2417 & n_n2323;
  assign new_n4775_ = ~pencrypt_0_ & new_n4774_;
  assign new_n4776_ = new_n1200_ & new_n4775_;
  assign new_n4777_ = ~pstart_0_ & new_n4776_;
  assign new_n4778_ = pencrypt_0_ & pkey_174_;
  assign new_n4779_ = pstart_0_ & new_n4778_;
  assign new_n4780_ = ~pencrypt_0_ & n_n2417;
  assign new_n4781_ = ~new_n1200_ & new_n4780_;
  assign new_n4782_ = ~pstart_0_ & new_n4781_;
  assign new_n4783_ = pkey_182_ & ~pencrypt_0_;
  assign new_n4784_ = pstart_0_ & new_n4783_;
  assign new_n4785_ = ~n_n2323 & ~new_n1220_;
  assign new_n4786_ = pencrypt_0_ & new_n4785_;
  assign new_n4787_ = n_n2417 & new_n4786_;
  assign new_n4788_ = ~pstart_0_ & new_n4787_;
  assign new_n4789_ = n_n2323 & new_n1220_;
  assign new_n4790_ = pencrypt_0_ & new_n4789_;
  assign new_n4791_ = n_n2417 & new_n4790_;
  assign new_n4792_ = ~pstart_0_ & new_n4791_;
  assign new_n4793_ = ~n_n2417 & ~n_n2323;
  assign new_n4794_ = ~pencrypt_0_ & new_n4793_;
  assign new_n4795_ = new_n1200_ & new_n4794_;
  assign new_n4796_ = ~pstart_0_ & new_n4795_;
  assign new_n4797_ = n_n2323 & ~new_n1220_;
  assign new_n4798_ = pencrypt_0_ & new_n4797_;
  assign new_n4799_ = ~n_n2417 & new_n4798_;
  assign new_n4800_ = ~pstart_0_ & new_n4799_;
  assign new_n4801_ = ~new_n4796_ & ~new_n4800_;
  assign new_n4802_ = ~new_n4788_ & ~new_n4792_;
  assign new_n4803_ = new_n4801_ & new_n4802_;
  assign new_n4804_ = ~new_n4782_ & ~new_n4784_;
  assign new_n4805_ = ~new_n4773_ & ~new_n4777_;
  assign new_n4806_ = ~new_n4779_ & new_n4805_;
  assign new_n4807_ = new_n4804_ & new_n4806_;
  assign n1402 = ~new_n4803_ | ~new_n4807_;
  assign new_n4809_ = ~pencrypt_0_ & n_n2332;
  assign new_n4810_ = ~new_n1200_ & new_n4809_;
  assign new_n4811_ = ~pstart_0_ & new_n4810_;
  assign new_n4812_ = n_n2427 & n_n2332;
  assign new_n4813_ = ~pencrypt_0_ & new_n4812_;
  assign new_n4814_ = new_n1200_ & new_n4813_;
  assign new_n4815_ = ~pstart_0_ & new_n4814_;
  assign new_n4816_ = pencrypt_0_ & pkey_100_;
  assign new_n4817_ = pstart_0_ & new_n4816_;
  assign new_n4818_ = ~pencrypt_0_ & n_n2427;
  assign new_n4819_ = ~new_n1200_ & new_n4818_;
  assign new_n4820_ = ~pstart_0_ & new_n4819_;
  assign new_n4821_ = ~n_n2332 & ~new_n1220_;
  assign new_n4822_ = pencrypt_0_ & new_n4821_;
  assign new_n4823_ = n_n2427 & new_n4822_;
  assign new_n4824_ = ~pstart_0_ & new_n4823_;
  assign new_n4825_ = n_n2332 & new_n1220_;
  assign new_n4826_ = pencrypt_0_ & new_n4825_;
  assign new_n4827_ = n_n2427 & new_n4826_;
  assign new_n4828_ = ~pstart_0_ & new_n4827_;
  assign new_n4829_ = ~n_n2427 & ~n_n2332;
  assign new_n4830_ = ~pencrypt_0_ & new_n4829_;
  assign new_n4831_ = new_n1200_ & new_n4830_;
  assign new_n4832_ = ~pstart_0_ & new_n4831_;
  assign new_n4833_ = n_n2332 & ~new_n1220_;
  assign new_n4834_ = pencrypt_0_ & new_n4833_;
  assign new_n4835_ = ~n_n2427 & new_n4834_;
  assign new_n4836_ = ~pstart_0_ & new_n4835_;
  assign new_n4837_ = ~new_n4832_ & ~new_n4836_;
  assign new_n4838_ = ~new_n4824_ & ~new_n4828_;
  assign new_n4839_ = new_n4837_ & new_n4838_;
  assign new_n4840_ = ~new_n2056_ & ~new_n4820_;
  assign new_n4841_ = ~new_n4811_ & ~new_n4815_;
  assign new_n4842_ = ~new_n4817_ & new_n4841_;
  assign new_n4843_ = new_n4840_ & new_n4842_;
  assign n1407 = ~new_n4839_ | ~new_n4843_;
  assign new_n4845_ = ~pencrypt_0_ & n_n2334;
  assign new_n4846_ = ~new_n1200_ & new_n4845_;
  assign new_n4847_ = ~pstart_0_ & new_n4846_;
  assign new_n4848_ = n_n2430 & n_n2334;
  assign new_n4849_ = ~pencrypt_0_ & new_n4848_;
  assign new_n4850_ = new_n1200_ & new_n4849_;
  assign new_n4851_ = ~pstart_0_ & new_n4850_;
  assign new_n4852_ = pkey_124_ & pencrypt_0_;
  assign new_n4853_ = pstart_0_ & new_n4852_;
  assign new_n4854_ = ~pencrypt_0_ & n_n2430;
  assign new_n4855_ = ~new_n1200_ & new_n4854_;
  assign new_n4856_ = ~pstart_0_ & new_n4855_;
  assign new_n4857_ = pkey_69_ & ~pencrypt_0_;
  assign new_n4858_ = pstart_0_ & new_n4857_;
  assign new_n4859_ = ~n_n2334 & ~new_n1220_;
  assign new_n4860_ = pencrypt_0_ & new_n4859_;
  assign new_n4861_ = n_n2430 & new_n4860_;
  assign new_n4862_ = ~pstart_0_ & new_n4861_;
  assign new_n4863_ = n_n2334 & new_n1220_;
  assign new_n4864_ = pencrypt_0_ & new_n4863_;
  assign new_n4865_ = n_n2430 & new_n4864_;
  assign new_n4866_ = ~pstart_0_ & new_n4865_;
  assign new_n4867_ = ~n_n2430 & ~n_n2334;
  assign new_n4868_ = ~pencrypt_0_ & new_n4867_;
  assign new_n4869_ = new_n1200_ & new_n4868_;
  assign new_n4870_ = ~pstart_0_ & new_n4869_;
  assign new_n4871_ = n_n2334 & ~new_n1220_;
  assign new_n4872_ = pencrypt_0_ & new_n4871_;
  assign new_n4873_ = ~n_n2430 & new_n4872_;
  assign new_n4874_ = ~pstart_0_ & new_n4873_;
  assign new_n4875_ = ~new_n4870_ & ~new_n4874_;
  assign new_n4876_ = ~new_n4862_ & ~new_n4866_;
  assign new_n4877_ = new_n4875_ & new_n4876_;
  assign new_n4878_ = ~new_n4856_ & ~new_n4858_;
  assign new_n4879_ = ~new_n4847_ & ~new_n4851_;
  assign new_n4880_ = ~new_n4853_ & new_n4879_;
  assign new_n4881_ = new_n4878_ & new_n4880_;
  assign n1412 = ~new_n4877_ | ~new_n4881_;
  assign new_n4883_ = ~pencrypt_0_ & n_n2344;
  assign new_n4884_ = ~new_n1200_ & new_n4883_;
  assign new_n4885_ = ~pstart_0_ & new_n4884_;
  assign new_n4886_ = n_n2437 & n_n2344;
  assign new_n4887_ = ~pencrypt_0_ & new_n4886_;
  assign new_n4888_ = new_n1200_ & new_n4887_;
  assign new_n4889_ = ~pstart_0_ & new_n4888_;
  assign new_n4890_ = pkey_86_ & pencrypt_0_;
  assign new_n4891_ = pstart_0_ & new_n4890_;
  assign new_n4892_ = ~pencrypt_0_ & n_n2437;
  assign new_n4893_ = ~new_n1200_ & new_n4892_;
  assign new_n4894_ = ~pstart_0_ & new_n4893_;
  assign new_n4895_ = pkey_94_ & ~pencrypt_0_;
  assign new_n4896_ = pstart_0_ & new_n4895_;
  assign new_n4897_ = ~n_n2344 & ~new_n1220_;
  assign new_n4898_ = pencrypt_0_ & new_n4897_;
  assign new_n4899_ = n_n2437 & new_n4898_;
  assign new_n4900_ = ~pstart_0_ & new_n4899_;
  assign new_n4901_ = n_n2344 & new_n1220_;
  assign new_n4902_ = pencrypt_0_ & new_n4901_;
  assign new_n4903_ = n_n2437 & new_n4902_;
  assign new_n4904_ = ~pstart_0_ & new_n4903_;
  assign new_n4905_ = ~n_n2437 & ~n_n2344;
  assign new_n4906_ = ~pencrypt_0_ & new_n4905_;
  assign new_n4907_ = new_n1200_ & new_n4906_;
  assign new_n4908_ = ~pstart_0_ & new_n4907_;
  assign new_n4909_ = n_n2344 & ~new_n1220_;
  assign new_n4910_ = pencrypt_0_ & new_n4909_;
  assign new_n4911_ = ~n_n2437 & new_n4910_;
  assign new_n4912_ = ~pstart_0_ & new_n4911_;
  assign new_n4913_ = ~new_n4908_ & ~new_n4912_;
  assign new_n4914_ = ~new_n4900_ & ~new_n4904_;
  assign new_n4915_ = new_n4913_ & new_n4914_;
  assign new_n4916_ = ~new_n4894_ & ~new_n4896_;
  assign new_n4917_ = ~new_n4885_ & ~new_n4889_;
  assign new_n4918_ = ~new_n4891_ & new_n4917_;
  assign new_n4919_ = new_n4916_ & new_n4918_;
  assign n1417 = ~new_n4915_ | ~new_n4919_;
  assign new_n4921_ = ~pencrypt_0_ & n_n2357;
  assign new_n4922_ = ~new_n1200_ & new_n4921_;
  assign new_n4923_ = ~pstart_0_ & new_n4922_;
  assign new_n4924_ = n_n2452 & n_n2357;
  assign new_n4925_ = ~pencrypt_0_ & new_n4924_;
  assign new_n4926_ = new_n1200_ & new_n4925_;
  assign new_n4927_ = ~pstart_0_ & new_n4926_;
  assign new_n4928_ = pkey_52_ & pencrypt_0_;
  assign new_n4929_ = pstart_0_ & new_n4928_;
  assign new_n4930_ = ~pencrypt_0_ & n_n2452;
  assign new_n4931_ = ~new_n1200_ & new_n4930_;
  assign new_n4932_ = ~pstart_0_ & new_n4931_;
  assign new_n4933_ = pkey_60_ & ~pencrypt_0_;
  assign new_n4934_ = pstart_0_ & new_n4933_;
  assign new_n4935_ = ~n_n2357 & ~new_n1220_;
  assign new_n4936_ = pencrypt_0_ & new_n4935_;
  assign new_n4937_ = n_n2452 & new_n4936_;
  assign new_n4938_ = ~pstart_0_ & new_n4937_;
  assign new_n4939_ = n_n2357 & new_n1220_;
  assign new_n4940_ = pencrypt_0_ & new_n4939_;
  assign new_n4941_ = n_n2452 & new_n4940_;
  assign new_n4942_ = ~pstart_0_ & new_n4941_;
  assign new_n4943_ = ~n_n2452 & ~n_n2357;
  assign new_n4944_ = ~pencrypt_0_ & new_n4943_;
  assign new_n4945_ = new_n1200_ & new_n4944_;
  assign new_n4946_ = ~pstart_0_ & new_n4945_;
  assign new_n4947_ = n_n2357 & ~new_n1220_;
  assign new_n4948_ = pencrypt_0_ & new_n4947_;
  assign new_n4949_ = ~n_n2452 & new_n4948_;
  assign new_n4950_ = ~pstart_0_ & new_n4949_;
  assign new_n4951_ = ~new_n4946_ & ~new_n4950_;
  assign new_n4952_ = ~new_n4938_ & ~new_n4942_;
  assign new_n4953_ = new_n4951_ & new_n4952_;
  assign new_n4954_ = ~new_n4932_ & ~new_n4934_;
  assign new_n4955_ = ~new_n4923_ & ~new_n4927_;
  assign new_n4956_ = ~new_n4929_ & new_n4955_;
  assign new_n4957_ = new_n4954_ & new_n4956_;
  assign n1422 = ~new_n4953_ | ~new_n4957_;
  assign new_n4959_ = ~new_n1200_ & new_n1824_;
  assign new_n4960_ = ~pstart_0_ & new_n4959_;
  assign new_n4961_ = new_n1200_ & new_n1819_;
  assign new_n4962_ = ~pstart_0_ & new_n4961_;
  assign new_n4963_ = pencrypt_0_ & pkey_14_;
  assign new_n4964_ = pstart_0_ & new_n4963_;
  assign new_n4965_ = ~new_n1200_ & new_n1815_;
  assign new_n4966_ = ~pstart_0_ & new_n4965_;
  assign new_n4967_ = ~pencrypt_0_ & pkey_22_;
  assign new_n4968_ = pstart_0_ & new_n4967_;
  assign new_n4969_ = ~n_n2367 & ~new_n1220_;
  assign new_n4970_ = pencrypt_0_ & new_n4969_;
  assign new_n4971_ = n_n2460 & new_n4970_;
  assign new_n4972_ = ~pstart_0_ & new_n4971_;
  assign new_n4973_ = n_n2367 & new_n1220_;
  assign new_n4974_ = pencrypt_0_ & new_n4973_;
  assign new_n4975_ = n_n2460 & new_n4974_;
  assign new_n4976_ = ~pstart_0_ & new_n4975_;
  assign new_n4977_ = new_n1200_ & new_n1838_;
  assign new_n4978_ = ~pstart_0_ & new_n4977_;
  assign new_n4979_ = n_n2367 & ~new_n1220_;
  assign new_n4980_ = pencrypt_0_ & new_n4979_;
  assign new_n4981_ = ~n_n2460 & new_n4980_;
  assign new_n4982_ = ~pstart_0_ & new_n4981_;
  assign new_n4983_ = ~new_n4978_ & ~new_n4982_;
  assign new_n4984_ = ~new_n4972_ & ~new_n4976_;
  assign new_n4985_ = new_n4983_ & new_n4984_;
  assign new_n4986_ = ~new_n4966_ & ~new_n4968_;
  assign new_n4987_ = ~new_n4960_ & ~new_n4962_;
  assign new_n4988_ = ~new_n4964_ & new_n4987_;
  assign new_n4989_ = new_n4986_ & new_n4988_;
  assign n1427 = ~new_n4985_ | ~new_n4989_;
  assign new_n4991_ = new_n1200_ & new_n1558_;
  assign new_n4992_ = ~pstart_0_ & new_n4991_;
  assign new_n4993_ = ~new_n1200_ & new_n1553_;
  assign new_n4994_ = ~pstart_0_ & new_n4993_;
  assign new_n4995_ = pkey_235_ & pencrypt_0_;
  assign new_n4996_ = pstart_0_ & new_n4995_;
  assign new_n4997_ = new_n1200_ & new_n1549_;
  assign new_n4998_ = ~pstart_0_ & new_n4997_;
  assign new_n4999_ = pkey_243_ & ~pencrypt_0_;
  assign new_n5000_ = pstart_0_ & new_n4999_;
  assign new_n5001_ = n_n2865 & new_n1220_;
  assign new_n5002_ = pencrypt_0_ & new_n5001_;
  assign new_n5003_ = ~n_n2280 & new_n5002_;
  assign new_n5004_ = ~pstart_0_ & new_n5003_;
  assign new_n5005_ = ~n_n2865 & new_n1220_;
  assign new_n5006_ = pencrypt_0_ & new_n5005_;
  assign new_n5007_ = n_n2280 & new_n5006_;
  assign new_n5008_ = ~pstart_0_ & new_n5007_;
  assign new_n5009_ = ~new_n1200_ & new_n1572_1_;
  assign new_n5010_ = ~pstart_0_ & new_n5009_;
  assign new_n5011_ = n_n2865 & ~new_n1220_;
  assign new_n5012_ = pencrypt_0_ & new_n5011_;
  assign new_n5013_ = n_n2280 & new_n5012_;
  assign new_n5014_ = ~pstart_0_ & new_n5013_;
  assign new_n5015_ = ~new_n5010_ & ~new_n5014_;
  assign new_n5016_ = ~new_n5004_ & ~new_n5008_;
  assign new_n5017_ = new_n5015_ & new_n5016_;
  assign new_n5018_ = ~new_n4998_ & ~new_n5000_;
  assign new_n5019_ = ~new_n4992_ & ~new_n4994_;
  assign new_n5020_ = ~new_n4996_ & new_n5019_;
  assign new_n5021_ = new_n5018_ & new_n5020_;
  assign n1432 = ~new_n5017_ | ~new_n5021_;
  assign new_n5023_ = new_n1200_ & new_n2760_;
  assign new_n5024_ = ~pstart_0_ & new_n5023_;
  assign new_n5025_ = ~new_n1200_ & new_n2755_;
  assign new_n5026_ = ~pstart_0_ & new_n5025_;
  assign new_n5027_ = pencrypt_0_ & pkey_32_;
  assign new_n5028_ = pstart_0_ & new_n5027_;
  assign new_n5029_ = new_n1200_ & new_n2751_;
  assign new_n5030_ = ~pstart_0_ & new_n5029_;
  assign new_n5031_ = ~pencrypt_0_ & pkey_40_;
  assign new_n5032_ = pstart_0_ & new_n5031_;
  assign new_n5033_ = n_n2463 & new_n1220_;
  assign new_n5034_ = pencrypt_0_ & new_n5033_;
  assign new_n5035_ = ~n_n2370 & new_n5034_;
  assign new_n5036_ = ~pstart_0_ & new_n5035_;
  assign new_n5037_ = ~n_n2463 & new_n1220_;
  assign new_n5038_ = pencrypt_0_ & new_n5037_;
  assign new_n5039_ = n_n2370 & new_n5038_;
  assign new_n5040_ = ~pstart_0_ & new_n5039_;
  assign new_n5041_ = ~new_n1200_ & new_n2774_;
  assign new_n5042_ = ~pstart_0_ & new_n5041_;
  assign new_n5043_ = n_n2463 & ~new_n1220_;
  assign new_n5044_ = pencrypt_0_ & new_n5043_;
  assign new_n5045_ = n_n2370 & new_n5044_;
  assign new_n5046_ = ~pstart_0_ & new_n5045_;
  assign new_n5047_ = ~new_n5042_ & ~new_n5046_;
  assign new_n5048_ = ~new_n5036_ & ~new_n5040_;
  assign new_n5049_ = new_n5047_ & new_n5048_;
  assign new_n5050_ = ~new_n5030_ & ~new_n5032_;
  assign new_n5051_ = ~new_n5024_ & ~new_n5026_;
  assign new_n5052_ = ~new_n5028_ & new_n5051_;
  assign new_n5053_ = new_n5050_ & new_n5052_;
  assign n1437 = ~new_n5049_ | ~new_n5053_;
  assign new_n5055_ = ~new_n1200_ & new_n3818_;
  assign new_n5056_ = ~pstart_0_ & new_n5055_;
  assign new_n5057_ = new_n1200_ & new_n3813_;
  assign new_n5058_ = ~pstart_0_ & new_n5057_;
  assign new_n5059_ = pencrypt_0_ & pkey_204_;
  assign new_n5060_ = pstart_0_ & new_n5059_;
  assign new_n5061_ = ~new_n1200_ & new_n3809_;
  assign new_n5062_ = ~pstart_0_ & new_n5061_;
  assign new_n5063_ = pkey_212_ & ~pencrypt_0_;
  assign new_n5064_ = pstart_0_ & new_n5063_;
  assign new_n5065_ = ~n_n2741 & ~new_n1220_;
  assign new_n5066_ = pencrypt_0_ & new_n5065_;
  assign new_n5067_ = n_n2378 & new_n5066_;
  assign new_n5068_ = ~pstart_0_ & new_n5067_;
  assign new_n5069_ = n_n2741 & new_n1220_;
  assign new_n5070_ = pencrypt_0_ & new_n5069_;
  assign new_n5071_ = n_n2378 & new_n5070_;
  assign new_n5072_ = ~pstart_0_ & new_n5071_;
  assign new_n5073_ = new_n1200_ & new_n3832_;
  assign new_n5074_ = ~pstart_0_ & new_n5073_;
  assign new_n5075_ = n_n2741 & ~new_n1220_;
  assign new_n5076_ = pencrypt_0_ & new_n5075_;
  assign new_n5077_ = ~n_n2378 & new_n5076_;
  assign new_n5078_ = ~pstart_0_ & new_n5077_;
  assign new_n5079_ = ~new_n5074_ & ~new_n5078_;
  assign new_n5080_ = ~new_n5068_ & ~new_n5072_;
  assign new_n5081_ = new_n5079_ & new_n5080_;
  assign new_n5082_ = ~new_n5062_ & ~new_n5064_;
  assign new_n5083_ = ~new_n5056_ & ~new_n5058_;
  assign new_n5084_ = ~new_n5060_ & new_n5083_;
  assign new_n5085_ = new_n5082_ & new_n5084_;
  assign n1442 = ~new_n5081_ | ~new_n5085_;
  assign new_n5087_ = ~pencrypt_0_ & n_n2305;
  assign new_n5088_ = ~new_n1200_ & new_n5087_;
  assign new_n5089_ = ~pstart_0_ & new_n5088_;
  assign new_n5090_ = n_n2399 & n_n2305;
  assign new_n5091_ = ~pencrypt_0_ & new_n5090_;
  assign new_n5092_ = new_n1200_ & new_n5091_;
  assign new_n5093_ = ~pstart_0_ & new_n5092_;
  assign new_n5094_ = pkey_132_ & pencrypt_0_;
  assign new_n5095_ = pstart_0_ & new_n5094_;
  assign new_n5096_ = ~pencrypt_0_ & n_n2399;
  assign new_n5097_ = ~new_n1200_ & new_n5096_;
  assign new_n5098_ = ~pstart_0_ & new_n5097_;
  assign new_n5099_ = pkey_140_ & ~pencrypt_0_;
  assign new_n5100_ = pstart_0_ & new_n5099_;
  assign new_n5101_ = ~n_n2305 & ~new_n1220_;
  assign new_n5102_ = pencrypt_0_ & new_n5101_;
  assign new_n5103_ = n_n2399 & new_n5102_;
  assign new_n5104_ = ~pstart_0_ & new_n5103_;
  assign new_n5105_ = n_n2305 & new_n1220_;
  assign new_n5106_ = pencrypt_0_ & new_n5105_;
  assign new_n5107_ = n_n2399 & new_n5106_;
  assign new_n5108_ = ~pstart_0_ & new_n5107_;
  assign new_n5109_ = ~n_n2399 & ~n_n2305;
  assign new_n5110_ = ~pencrypt_0_ & new_n5109_;
  assign new_n5111_ = new_n1200_ & new_n5110_;
  assign new_n5112_ = ~pstart_0_ & new_n5111_;
  assign new_n5113_ = n_n2305 & ~new_n1220_;
  assign new_n5114_ = pencrypt_0_ & new_n5113_;
  assign new_n5115_ = ~n_n2399 & new_n5114_;
  assign new_n5116_ = ~pstart_0_ & new_n5115_;
  assign new_n5117_ = ~new_n5112_ & ~new_n5116_;
  assign new_n5118_ = ~new_n5104_ & ~new_n5108_;
  assign new_n5119_ = new_n5117_ & new_n5118_;
  assign new_n5120_ = ~new_n5098_ & ~new_n5100_;
  assign new_n5121_ = ~new_n5089_ & ~new_n5093_;
  assign new_n5122_ = ~new_n5095_ & new_n5121_;
  assign new_n5123_ = new_n5120_ & new_n5122_;
  assign n1447 = ~new_n5119_ | ~new_n5123_;
  assign new_n5125_ = ~pencrypt_0_ & n_n2312;
  assign new_n5126_ = ~new_n1200_ & new_n5125_;
  assign new_n5127_ = ~pstart_0_ & new_n5126_;
  assign new_n5128_ = n_n2407 & n_n2312;
  assign new_n5129_ = ~pencrypt_0_ & new_n5128_;
  assign new_n5130_ = new_n1200_ & new_n5129_;
  assign new_n5131_ = ~pstart_0_ & new_n5130_;
  assign new_n5132_ = pkey_141_ & pencrypt_0_;
  assign new_n5133_ = pstart_0_ & new_n5132_;
  assign new_n5134_ = ~pencrypt_0_ & n_n2407;
  assign new_n5135_ = ~new_n1200_ & new_n5134_;
  assign new_n5136_ = ~pstart_0_ & new_n5135_;
  assign new_n5137_ = pkey_149_ & ~pencrypt_0_;
  assign new_n5138_ = pstart_0_ & new_n5137_;
  assign new_n5139_ = ~n_n2312 & ~new_n1220_;
  assign new_n5140_ = pencrypt_0_ & new_n5139_;
  assign new_n5141_ = n_n2407 & new_n5140_;
  assign new_n5142_ = ~pstart_0_ & new_n5141_;
  assign new_n5143_ = n_n2312 & new_n1220_;
  assign new_n5144_ = pencrypt_0_ & new_n5143_;
  assign new_n5145_ = n_n2407 & new_n5144_;
  assign new_n5146_ = ~pstart_0_ & new_n5145_;
  assign new_n5147_ = ~n_n2407 & ~n_n2312;
  assign new_n5148_ = ~pencrypt_0_ & new_n5147_;
  assign new_n5149_ = new_n1200_ & new_n5148_;
  assign new_n5150_ = ~pstart_0_ & new_n5149_;
  assign new_n5151_ = n_n2312 & ~new_n1220_;
  assign new_n5152_ = pencrypt_0_ & new_n5151_;
  assign new_n5153_ = ~n_n2407 & new_n5152_;
  assign new_n5154_ = ~pstart_0_ & new_n5153_;
  assign new_n5155_ = ~new_n5150_ & ~new_n5154_;
  assign new_n5156_ = ~new_n5142_ & ~new_n5146_;
  assign new_n5157_ = new_n5155_ & new_n5156_;
  assign new_n5158_ = ~new_n5136_ & ~new_n5138_;
  assign new_n5159_ = ~new_n5127_ & ~new_n5131_;
  assign new_n5160_ = ~new_n5133_ & new_n5159_;
  assign new_n5161_ = new_n5158_ & new_n5160_;
  assign n1452 = ~new_n5157_ | ~new_n5161_;
  assign new_n5163_ = ~pencrypt_0_ & n_n2324;
  assign new_n5164_ = ~new_n1200_ & new_n5163_;
  assign new_n5165_ = ~pstart_0_ & new_n5164_;
  assign new_n5166_ = n_n2418 & n_n2324;
  assign new_n5167_ = ~pencrypt_0_ & new_n5166_;
  assign new_n5168_ = new_n1200_ & new_n5167_;
  assign new_n5169_ = ~pstart_0_ & new_n5168_;
  assign new_n5170_ = pkey_182_ & pencrypt_0_;
  assign new_n5171_ = pstart_0_ & new_n5170_;
  assign new_n5172_ = ~pencrypt_0_ & n_n2418;
  assign new_n5173_ = ~new_n1200_ & new_n5172_;
  assign new_n5174_ = ~pstart_0_ & new_n5173_;
  assign new_n5175_ = ~pencrypt_0_ & pkey_190_;
  assign new_n5176_ = pstart_0_ & new_n5175_;
  assign new_n5177_ = ~n_n2324 & ~new_n1220_;
  assign new_n5178_ = pencrypt_0_ & new_n5177_;
  assign new_n5179_ = n_n2418 & new_n5178_;
  assign new_n5180_ = ~pstart_0_ & new_n5179_;
  assign new_n5181_ = n_n2324 & new_n1220_;
  assign new_n5182_ = pencrypt_0_ & new_n5181_;
  assign new_n5183_ = n_n2418 & new_n5182_;
  assign new_n5184_ = ~pstart_0_ & new_n5183_;
  assign new_n5185_ = ~n_n2418 & ~n_n2324;
  assign new_n5186_ = ~pencrypt_0_ & new_n5185_;
  assign new_n5187_ = new_n1200_ & new_n5186_;
  assign new_n5188_ = ~pstart_0_ & new_n5187_;
  assign new_n5189_ = n_n2324 & ~new_n1220_;
  assign new_n5190_ = pencrypt_0_ & new_n5189_;
  assign new_n5191_ = ~n_n2418 & new_n5190_;
  assign new_n5192_ = ~pstart_0_ & new_n5191_;
  assign new_n5193_ = ~new_n5188_ & ~new_n5192_;
  assign new_n5194_ = ~new_n5180_ & ~new_n5184_;
  assign new_n5195_ = new_n5193_ & new_n5194_;
  assign new_n5196_ = ~new_n5174_ & ~new_n5176_;
  assign new_n5197_ = ~new_n5165_ & ~new_n5169_;
  assign new_n5198_ = ~new_n5171_ & new_n5197_;
  assign new_n5199_ = new_n5196_ & new_n5198_;
  assign n1457 = ~new_n5195_ | ~new_n5199_;
  assign new_n5201_ = ~pencrypt_0_ & n_n2331;
  assign new_n5202_ = ~new_n1200_ & new_n5201_;
  assign new_n5203_ = ~pstart_0_ & new_n5202_;
  assign new_n5204_ = n_n2426 & n_n2331;
  assign new_n5205_ = ~pencrypt_0_ & new_n5204_;
  assign new_n5206_ = new_n1200_ & new_n5205_;
  assign new_n5207_ = ~pstart_0_ & new_n5206_;
  assign new_n5208_ = pkey_92_ & pencrypt_0_;
  assign new_n5209_ = pstart_0_ & new_n5208_;
  assign new_n5210_ = ~pencrypt_0_ & n_n2426;
  assign new_n5211_ = ~new_n1200_ & new_n5210_;
  assign new_n5212_ = ~pstart_0_ & new_n5211_;
  assign new_n5213_ = ~pencrypt_0_ & pkey_100_;
  assign new_n5214_ = pstart_0_ & new_n5213_;
  assign new_n5215_ = ~n_n2331 & ~new_n1220_;
  assign new_n5216_ = pencrypt_0_ & new_n5215_;
  assign new_n5217_ = n_n2426 & new_n5216_;
  assign new_n5218_ = ~pstart_0_ & new_n5217_;
  assign new_n5219_ = n_n2331 & new_n1220_;
  assign new_n5220_ = pencrypt_0_ & new_n5219_;
  assign new_n5221_ = n_n2426 & new_n5220_;
  assign new_n5222_ = ~pstart_0_ & new_n5221_;
  assign new_n5223_ = ~n_n2426 & ~n_n2331;
  assign new_n5224_ = ~pencrypt_0_ & new_n5223_;
  assign new_n5225_ = new_n1200_ & new_n5224_;
  assign new_n5226_ = ~pstart_0_ & new_n5225_;
  assign new_n5227_ = n_n2331 & ~new_n1220_;
  assign new_n5228_ = pencrypt_0_ & new_n5227_;
  assign new_n5229_ = ~n_n2426 & new_n5228_;
  assign new_n5230_ = ~pstart_0_ & new_n5229_;
  assign new_n5231_ = ~new_n5226_ & ~new_n5230_;
  assign new_n5232_ = ~new_n5218_ & ~new_n5222_;
  assign new_n5233_ = new_n5231_ & new_n5232_;
  assign new_n5234_ = ~new_n5212_ & ~new_n5214_;
  assign new_n5235_ = ~new_n5203_ & ~new_n5207_;
  assign new_n5236_ = ~new_n5209_ & new_n5235_;
  assign new_n5237_ = new_n5234_ & new_n5236_;
  assign n1462 = ~new_n5233_ | ~new_n5237_;
  assign new_n5239_ = ~pencrypt_0_ & n_n2335;
  assign new_n5240_ = ~new_n1200_ & new_n5239_;
  assign new_n5241_ = ~pstart_0_ & new_n5240_;
  assign new_n5242_ = n_n2943 & n_n2335;
  assign new_n5243_ = ~pencrypt_0_ & new_n5242_;
  assign new_n5244_ = new_n1200_ & new_n5243_;
  assign new_n5245_ = ~pstart_0_ & new_n5244_;
  assign new_n5246_ = pkey_69_ & pencrypt_0_;
  assign new_n5247_ = pstart_0_ & new_n5246_;
  assign new_n5248_ = ~pencrypt_0_ & n_n2943;
  assign new_n5249_ = ~new_n1200_ & new_n5248_;
  assign new_n5250_ = ~pstart_0_ & new_n5249_;
  assign new_n5251_ = pkey_77_ & ~pencrypt_0_;
  assign new_n5252_ = pstart_0_ & new_n5251_;
  assign new_n5253_ = ~n_n2335 & ~new_n1220_;
  assign new_n5254_ = pencrypt_0_ & new_n5253_;
  assign new_n5255_ = n_n2943 & new_n5254_;
  assign new_n5256_ = ~pstart_0_ & new_n5255_;
  assign new_n5257_ = n_n2335 & new_n1220_;
  assign new_n5258_ = pencrypt_0_ & new_n5257_;
  assign new_n5259_ = n_n2943 & new_n5258_;
  assign new_n5260_ = ~pstart_0_ & new_n5259_;
  assign new_n5261_ = ~n_n2943 & ~n_n2335;
  assign new_n5262_ = ~pencrypt_0_ & new_n5261_;
  assign new_n5263_ = new_n1200_ & new_n5262_;
  assign new_n5264_ = ~pstart_0_ & new_n5263_;
  assign new_n5265_ = n_n2335 & ~new_n1220_;
  assign new_n5266_ = pencrypt_0_ & new_n5265_;
  assign new_n5267_ = ~n_n2943 & new_n5266_;
  assign new_n5268_ = ~pstart_0_ & new_n5267_;
  assign new_n5269_ = ~new_n5264_ & ~new_n5268_;
  assign new_n5270_ = ~new_n5256_ & ~new_n5260_;
  assign new_n5271_ = new_n5269_ & new_n5270_;
  assign new_n5272_ = ~new_n5250_ & ~new_n5252_;
  assign new_n5273_ = ~new_n5241_ & ~new_n5245_;
  assign new_n5274_ = ~new_n5247_ & new_n5273_;
  assign new_n5275_ = new_n5272_ & new_n5274_;
  assign n1467 = ~new_n5271_ | ~new_n5275_;
  assign new_n5277_ = ~pencrypt_0_ & n_n2343;
  assign new_n5278_ = ~new_n1200_ & new_n5277_;
  assign new_n5279_ = ~pstart_0_ & new_n5278_;
  assign new_n5280_ = n_n2436 & n_n2343;
  assign new_n5281_ = ~pencrypt_0_ & new_n5280_;
  assign new_n5282_ = new_n1200_ & new_n5281_;
  assign new_n5283_ = ~pstart_0_ & new_n5282_;
  assign new_n5284_ = pkey_78_ & pencrypt_0_;
  assign new_n5285_ = pstart_0_ & new_n5284_;
  assign new_n5286_ = ~pencrypt_0_ & n_n2436;
  assign new_n5287_ = ~new_n1200_ & new_n5286_;
  assign new_n5288_ = ~pstart_0_ & new_n5287_;
  assign new_n5289_ = pkey_86_ & ~pencrypt_0_;
  assign new_n5290_ = pstart_0_ & new_n5289_;
  assign new_n5291_ = ~n_n2343 & ~new_n1220_;
  assign new_n5292_ = pencrypt_0_ & new_n5291_;
  assign new_n5293_ = n_n2436 & new_n5292_;
  assign new_n5294_ = ~pstart_0_ & new_n5293_;
  assign new_n5295_ = n_n2343 & new_n1220_;
  assign new_n5296_ = pencrypt_0_ & new_n5295_;
  assign new_n5297_ = n_n2436 & new_n5296_;
  assign new_n5298_ = ~pstart_0_ & new_n5297_;
  assign new_n5299_ = ~n_n2436 & ~n_n2343;
  assign new_n5300_ = ~pencrypt_0_ & new_n5299_;
  assign new_n5301_ = new_n1200_ & new_n5300_;
  assign new_n5302_ = ~pstart_0_ & new_n5301_;
  assign new_n5303_ = n_n2343 & ~new_n1220_;
  assign new_n5304_ = pencrypt_0_ & new_n5303_;
  assign new_n5305_ = ~n_n2436 & new_n5304_;
  assign new_n5306_ = ~pstart_0_ & new_n5305_;
  assign new_n5307_ = ~new_n5302_ & ~new_n5306_;
  assign new_n5308_ = ~new_n5294_ & ~new_n5298_;
  assign new_n5309_ = new_n5307_ & new_n5308_;
  assign new_n5310_ = ~new_n5288_ & ~new_n5290_;
  assign new_n5311_ = ~new_n5279_ & ~new_n5283_;
  assign new_n5312_ = ~new_n5285_ & new_n5311_;
  assign new_n5313_ = new_n5310_ & new_n5312_;
  assign n1472 = ~new_n5309_ | ~new_n5313_;
  assign new_n5315_ = ~pencrypt_0_ & n_n2358;
  assign new_n5316_ = ~new_n1200_ & new_n5315_;
  assign new_n5317_ = ~pstart_0_ & new_n5316_;
  assign new_n5318_ = n_n2453 & n_n2358;
  assign new_n5319_ = ~pencrypt_0_ & new_n5318_;
  assign new_n5320_ = new_n1200_ & new_n5319_;
  assign new_n5321_ = ~pstart_0_ & new_n5320_;
  assign new_n5322_ = pkey_60_ & pencrypt_0_;
  assign new_n5323_ = pstart_0_ & new_n5322_;
  assign new_n5324_ = ~pencrypt_0_ & n_n2453;
  assign new_n5325_ = ~new_n1200_ & new_n5324_;
  assign new_n5326_ = ~pstart_0_ & new_n5325_;
  assign new_n5327_ = pkey_5_ & ~pencrypt_0_;
  assign new_n5328_ = pstart_0_ & new_n5327_;
  assign new_n5329_ = ~n_n2358 & ~new_n1220_;
  assign new_n5330_ = pencrypt_0_ & new_n5329_;
  assign new_n5331_ = n_n2453 & new_n5330_;
  assign new_n5332_ = ~pstart_0_ & new_n5331_;
  assign new_n5333_ = n_n2358 & new_n1220_;
  assign new_n5334_ = pencrypt_0_ & new_n5333_;
  assign new_n5335_ = n_n2453 & new_n5334_;
  assign new_n5336_ = ~pstart_0_ & new_n5335_;
  assign new_n5337_ = ~n_n2453 & ~n_n2358;
  assign new_n5338_ = ~pencrypt_0_ & new_n5337_;
  assign new_n5339_ = new_n1200_ & new_n5338_;
  assign new_n5340_ = ~pstart_0_ & new_n5339_;
  assign new_n5341_ = n_n2358 & ~new_n1220_;
  assign new_n5342_ = pencrypt_0_ & new_n5341_;
  assign new_n5343_ = ~n_n2453 & new_n5342_;
  assign new_n5344_ = ~pstart_0_ & new_n5343_;
  assign new_n5345_ = ~new_n5340_ & ~new_n5344_;
  assign new_n5346_ = ~new_n5332_ & ~new_n5336_;
  assign new_n5347_ = new_n5345_ & new_n5346_;
  assign new_n5348_ = ~new_n5326_ & ~new_n5328_;
  assign new_n5349_ = ~new_n5317_ & ~new_n5321_;
  assign new_n5350_ = ~new_n5323_ & new_n5349_;
  assign new_n5351_ = new_n5348_ & new_n5350_;
  assign n1477 = ~new_n5347_ | ~new_n5351_;
  assign new_n5353_ = ~new_n1200_ & new_n1520_;
  assign new_n5354_ = ~pstart_0_ & new_n5353_;
  assign new_n5355_ = new_n1200_ & new_n1515_;
  assign new_n5356_ = ~pstart_0_ & new_n5355_;
  assign new_n5357_ = pkey_6_ & pencrypt_0_;
  assign new_n5358_ = pstart_0_ & new_n5357_;
  assign new_n5359_ = ~new_n1200_ & new_n1511_;
  assign new_n5360_ = ~pstart_0_ & new_n5359_;
  assign new_n5361_ = ~pencrypt_0_ & pkey_14_;
  assign new_n5362_ = pstart_0_ & new_n5361_;
  assign new_n5363_ = ~n_n2366 & ~new_n1220_;
  assign new_n5364_ = pencrypt_0_ & new_n5363_;
  assign new_n5365_ = n_n2986 & new_n5364_;
  assign new_n5366_ = ~pstart_0_ & new_n5365_;
  assign new_n5367_ = n_n2366 & new_n1220_;
  assign new_n5368_ = pencrypt_0_ & new_n5367_;
  assign new_n5369_ = n_n2986 & new_n5368_;
  assign new_n5370_ = ~pstart_0_ & new_n5369_;
  assign new_n5371_ = new_n1200_ & new_n1534_;
  assign new_n5372_ = ~pstart_0_ & new_n5371_;
  assign new_n5373_ = n_n2366 & ~new_n1220_;
  assign new_n5374_ = pencrypt_0_ & new_n5373_;
  assign new_n5375_ = ~n_n2986 & new_n5374_;
  assign new_n5376_ = ~pstart_0_ & new_n5375_;
  assign new_n5377_ = ~new_n5372_ & ~new_n5376_;
  assign new_n5378_ = ~new_n5366_ & ~new_n5370_;
  assign new_n5379_ = new_n5377_ & new_n5378_;
  assign new_n5380_ = ~new_n5360_ & ~new_n5362_;
  assign new_n5381_ = ~new_n5354_ & ~new_n5356_;
  assign new_n5382_ = ~new_n5358_ & new_n5381_;
  assign new_n5383_ = new_n5380_ & new_n5382_;
  assign n1482 = ~new_n5379_ | ~new_n5383_;
  assign new_n5385_ = new_n1200_ & new_n1254_;
  assign new_n5386_ = ~pstart_0_ & new_n5385_;
  assign new_n5387_ = ~new_n1200_ & new_n1249_;
  assign new_n5388_ = ~pstart_0_ & new_n5387_;
  assign new_n5389_ = pkey_243_ & pencrypt_0_;
  assign new_n5390_ = pstart_0_ & new_n5389_;
  assign new_n5391_ = new_n1200_ & new_n1245_;
  assign new_n5392_ = ~pstart_0_ & new_n5391_;
  assign new_n5393_ = pkey_251_ & ~pencrypt_0_;
  assign new_n5394_ = pstart_0_ & new_n5393_;
  assign new_n5395_ = n_n2375 & new_n1220_;
  assign new_n5396_ = pencrypt_0_ & new_n5395_;
  assign new_n5397_ = ~n_n2737 & new_n5396_;
  assign new_n5398_ = ~pstart_0_ & new_n5397_;
  assign new_n5399_ = ~n_n2375 & new_n1220_;
  assign new_n5400_ = pencrypt_0_ & new_n5399_;
  assign new_n5401_ = n_n2737 & new_n5400_;
  assign new_n5402_ = ~pstart_0_ & new_n5401_;
  assign new_n5403_ = ~new_n1200_ & new_n1268_;
  assign new_n5404_ = ~pstart_0_ & new_n5403_;
  assign new_n5405_ = n_n2375 & ~new_n1220_;
  assign new_n5406_ = pencrypt_0_ & new_n5405_;
  assign new_n5407_ = n_n2737 & new_n5406_;
  assign new_n5408_ = ~pstart_0_ & new_n5407_;
  assign new_n5409_ = ~new_n5404_ & ~new_n5408_;
  assign new_n5410_ = ~new_n5398_ & ~new_n5402_;
  assign new_n5411_ = new_n5409_ & new_n5410_;
  assign new_n5412_ = ~new_n5392_ & ~new_n5394_;
  assign new_n5413_ = ~new_n5386_ & ~new_n5388_;
  assign new_n5414_ = ~new_n5390_ & new_n5413_;
  assign new_n5415_ = new_n5412_ & new_n5414_;
  assign n1487 = ~new_n5411_ | ~new_n5415_;
  assign new_n5417_ = ~pencrypt_0_ & n_n2290;
  assign new_n5418_ = ~new_n1200_ & new_n5417_;
  assign new_n5419_ = ~pstart_0_ & new_n5418_;
  assign new_n5420_ = n_n2385 & n_n2290;
  assign new_n5421_ = ~pencrypt_0_ & new_n5420_;
  assign new_n5422_ = new_n1200_ & new_n5421_;
  assign new_n5423_ = ~pstart_0_ & new_n5422_;
  assign new_n5424_ = pkey_221_ & pencrypt_0_;
  assign new_n5425_ = pstart_0_ & new_n5424_;
  assign new_n5426_ = ~pencrypt_0_ & n_n2385;
  assign new_n5427_ = ~new_n1200_ & new_n5426_;
  assign new_n5428_ = ~pstart_0_ & new_n5427_;
  assign new_n5429_ = pkey_229_ & ~pencrypt_0_;
  assign new_n5430_ = pstart_0_ & new_n5429_;
  assign new_n5431_ = ~n_n2290 & ~new_n1220_;
  assign new_n5432_ = pencrypt_0_ & new_n5431_;
  assign new_n5433_ = n_n2385 & new_n5432_;
  assign new_n5434_ = ~pstart_0_ & new_n5433_;
  assign new_n5435_ = n_n2290 & new_n1220_;
  assign new_n5436_ = pencrypt_0_ & new_n5435_;
  assign new_n5437_ = n_n2385 & new_n5436_;
  assign new_n5438_ = ~pstart_0_ & new_n5437_;
  assign new_n5439_ = ~n_n2385 & ~n_n2290;
  assign new_n5440_ = ~pencrypt_0_ & new_n5439_;
  assign new_n5441_ = new_n1200_ & new_n5440_;
  assign new_n5442_ = ~pstart_0_ & new_n5441_;
  assign new_n5443_ = n_n2290 & ~new_n1220_;
  assign new_n5444_ = pencrypt_0_ & new_n5443_;
  assign new_n5445_ = ~n_n2385 & new_n5444_;
  assign new_n5446_ = ~pstart_0_ & new_n5445_;
  assign new_n5447_ = ~new_n5442_ & ~new_n5446_;
  assign new_n5448_ = ~new_n5434_ & ~new_n5438_;
  assign new_n5449_ = new_n5447_ & new_n5448_;
  assign new_n5450_ = ~new_n5428_ & ~new_n5430_;
  assign new_n5451_ = ~new_n5419_ & ~new_n5423_;
  assign new_n5452_ = ~new_n5425_ & new_n5451_;
  assign new_n5453_ = new_n5450_ & new_n5452_;
  assign n1492 = ~new_n5449_ | ~new_n5453_;
  assign new_n5455_ = ~pencrypt_0_ & n_n2300;
  assign new_n5456_ = ~new_n1200_ & new_n5455_;
  assign new_n5457_ = ~pstart_0_ & new_n5456_;
  assign new_n5458_ = n_n2394 & n_n2300;
  assign new_n5459_ = ~pencrypt_0_ & new_n5458_;
  assign new_n5460_ = new_n1200_ & new_n5459_;
  assign new_n5461_ = ~pstart_0_ & new_n5460_;
  assign new_n5462_ = pkey_246_ & pencrypt_0_;
  assign new_n5463_ = pstart_0_ & new_n5462_;
  assign new_n5464_ = ~pencrypt_0_ & n_n2394;
  assign new_n5465_ = ~new_n1200_ & new_n5464_;
  assign new_n5466_ = ~pstart_0_ & new_n5465_;
  assign new_n5467_ = pkey_254_ & ~pencrypt_0_;
  assign new_n5468_ = pstart_0_ & new_n5467_;
  assign new_n5469_ = ~n_n2300 & ~new_n1220_;
  assign new_n5470_ = pencrypt_0_ & new_n5469_;
  assign new_n5471_ = n_n2394 & new_n5470_;
  assign new_n5472_ = ~pstart_0_ & new_n5471_;
  assign new_n5473_ = n_n2300 & new_n1220_;
  assign new_n5474_ = pencrypt_0_ & new_n5473_;
  assign new_n5475_ = n_n2394 & new_n5474_;
  assign new_n5476_ = ~pstart_0_ & new_n5475_;
  assign new_n5477_ = ~n_n2394 & ~n_n2300;
  assign new_n5478_ = ~pencrypt_0_ & new_n5477_;
  assign new_n5479_ = new_n1200_ & new_n5478_;
  assign new_n5480_ = ~pstart_0_ & new_n5479_;
  assign new_n5481_ = n_n2300 & ~new_n1220_;
  assign new_n5482_ = pencrypt_0_ & new_n5481_;
  assign new_n5483_ = ~n_n2394 & new_n5482_;
  assign new_n5484_ = ~pstart_0_ & new_n5483_;
  assign new_n5485_ = ~new_n5480_ & ~new_n5484_;
  assign new_n5486_ = ~new_n5472_ & ~new_n5476_;
  assign new_n5487_ = new_n5485_ & new_n5486_;
  assign new_n5488_ = ~new_n5466_ & ~new_n5468_;
  assign new_n5489_ = ~new_n5457_ & ~new_n5461_;
  assign new_n5490_ = ~new_n5463_ & new_n5489_;
  assign new_n5491_ = new_n5488_ & new_n5490_;
  assign n1497 = ~new_n5487_ | ~new_n5491_;
  assign new_n5493_ = ~pencrypt_0_ & n_n2774;
  assign new_n5494_ = ~new_n1200_ & new_n5493_;
  assign new_n5495_ = ~pstart_0_ & new_n5494_;
  assign new_n5496_ = n_n2400 & n_n2774;
  assign new_n5497_ = ~pencrypt_0_ & new_n5496_;
  assign new_n5498_ = new_n1200_ & new_n5497_;
  assign new_n5499_ = ~pstart_0_ & new_n5498_;
  assign new_n5500_ = pkey_140_ & pencrypt_0_;
  assign new_n5501_ = pstart_0_ & new_n5500_;
  assign new_n5502_ = ~pencrypt_0_ & n_n2400;
  assign new_n5503_ = ~new_n1200_ & new_n5502_;
  assign new_n5504_ = ~pstart_0_ & new_n5503_;
  assign new_n5505_ = pkey_148_ & ~pencrypt_0_;
  assign new_n5506_ = pstart_0_ & new_n5505_;
  assign new_n5507_ = ~n_n2774 & ~new_n1220_;
  assign new_n5508_ = pencrypt_0_ & new_n5507_;
  assign new_n5509_ = n_n2400 & new_n5508_;
  assign new_n5510_ = ~pstart_0_ & new_n5509_;
  assign new_n5511_ = n_n2774 & new_n1220_;
  assign new_n5512_ = pencrypt_0_ & new_n5511_;
  assign new_n5513_ = n_n2400 & new_n5512_;
  assign new_n5514_ = ~pstart_0_ & new_n5513_;
  assign new_n5515_ = ~n_n2400 & ~n_n2774;
  assign new_n5516_ = ~pencrypt_0_ & new_n5515_;
  assign new_n5517_ = new_n1200_ & new_n5516_;
  assign new_n5518_ = ~pstart_0_ & new_n5517_;
  assign new_n5519_ = n_n2774 & ~new_n1220_;
  assign new_n5520_ = pencrypt_0_ & new_n5519_;
  assign new_n5521_ = ~n_n2400 & new_n5520_;
  assign new_n5522_ = ~pstart_0_ & new_n5521_;
  assign new_n5523_ = ~new_n5518_ & ~new_n5522_;
  assign new_n5524_ = ~new_n5510_ & ~new_n5514_;
  assign new_n5525_ = new_n5523_ & new_n5524_;
  assign new_n5526_ = ~new_n5504_ & ~new_n5506_;
  assign new_n5527_ = ~new_n5495_ & ~new_n5499_;
  assign new_n5528_ = ~new_n5501_ & new_n5527_;
  assign new_n5529_ = new_n5526_ & new_n5528_;
  assign n1502 = ~new_n5525_ | ~new_n5529_;
  assign new_n5531_ = ~pencrypt_0_ & n_n2315;
  assign new_n5532_ = ~new_n1200_ & new_n5531_;
  assign new_n5533_ = ~pstart_0_ & new_n5532_;
  assign new_n5534_ = n_n2410 & n_n2315;
  assign new_n5535_ = ~pencrypt_0_ & new_n5534_;
  assign new_n5536_ = new_n1200_ & new_n5535_;
  assign new_n5537_ = ~pstart_0_ & new_n5536_;
  assign new_n5538_ = pkey_165_ & pencrypt_0_;
  assign new_n5539_ = pstart_0_ & new_n5538_;
  assign new_n5540_ = ~pencrypt_0_ & n_n2410;
  assign new_n5541_ = ~new_n1200_ & new_n5540_;
  assign new_n5542_ = ~pstart_0_ & new_n5541_;
  assign new_n5543_ = ~pencrypt_0_ & pkey_173_;
  assign new_n5544_ = pstart_0_ & new_n5543_;
  assign new_n5545_ = ~n_n2315 & ~new_n1220_;
  assign new_n5546_ = pencrypt_0_ & new_n5545_;
  assign new_n5547_ = n_n2410 & new_n5546_;
  assign new_n5548_ = ~pstart_0_ & new_n5547_;
  assign new_n5549_ = n_n2315 & new_n1220_;
  assign new_n5550_ = pencrypt_0_ & new_n5549_;
  assign new_n5551_ = n_n2410 & new_n5550_;
  assign new_n5552_ = ~pstart_0_ & new_n5551_;
  assign new_n5553_ = ~n_n2410 & ~n_n2315;
  assign new_n5554_ = ~pencrypt_0_ & new_n5553_;
  assign new_n5555_ = new_n1200_ & new_n5554_;
  assign new_n5556_ = ~pstart_0_ & new_n5555_;
  assign new_n5557_ = n_n2315 & ~new_n1220_;
  assign new_n5558_ = pencrypt_0_ & new_n5557_;
  assign new_n5559_ = ~n_n2410 & new_n5558_;
  assign new_n5560_ = ~pstart_0_ & new_n5559_;
  assign new_n5561_ = ~new_n5556_ & ~new_n5560_;
  assign new_n5562_ = ~new_n5548_ & ~new_n5552_;
  assign new_n5563_ = new_n5561_ & new_n5562_;
  assign new_n5564_ = ~new_n5542_ & ~new_n5544_;
  assign new_n5565_ = ~new_n5533_ & ~new_n5537_;
  assign new_n5566_ = ~new_n5539_ & new_n5565_;
  assign new_n5567_ = new_n5564_ & new_n5566_;
  assign n1507 = ~new_n5563_ | ~new_n5567_;
  assign new_n5569_ = ~pencrypt_0_ & n_n2321;
  assign new_n5570_ = ~new_n1200_ & new_n5569_;
  assign new_n5571_ = ~pstart_0_ & new_n5570_;
  assign new_n5572_ = n_n2415 & n_n2321;
  assign new_n5573_ = ~pencrypt_0_ & new_n5572_;
  assign new_n5574_ = new_n1200_ & new_n5573_;
  assign new_n5575_ = ~pstart_0_ & new_n5574_;
  assign new_n5576_ = pkey_158_ & pencrypt_0_;
  assign new_n5577_ = pstart_0_ & new_n5576_;
  assign new_n5578_ = ~pencrypt_0_ & n_n2415;
  assign new_n5579_ = ~new_n1200_ & new_n5578_;
  assign new_n5580_ = ~pstart_0_ & new_n5579_;
  assign new_n5581_ = pkey_166_ & ~pencrypt_0_;
  assign new_n5582_ = pstart_0_ & new_n5581_;
  assign new_n5583_ = ~n_n2321 & ~new_n1220_;
  assign new_n5584_ = pencrypt_0_ & new_n5583_;
  assign new_n5585_ = n_n2415 & new_n5584_;
  assign new_n5586_ = ~pstart_0_ & new_n5585_;
  assign new_n5587_ = n_n2321 & new_n1220_;
  assign new_n5588_ = pencrypt_0_ & new_n5587_;
  assign new_n5589_ = n_n2415 & new_n5588_;
  assign new_n5590_ = ~pstart_0_ & new_n5589_;
  assign new_n5591_ = ~n_n2415 & ~n_n2321;
  assign new_n5592_ = ~pencrypt_0_ & new_n5591_;
  assign new_n5593_ = new_n1200_ & new_n5592_;
  assign new_n5594_ = ~pstart_0_ & new_n5593_;
  assign new_n5595_ = n_n2321 & ~new_n1220_;
  assign new_n5596_ = pencrypt_0_ & new_n5595_;
  assign new_n5597_ = ~n_n2415 & new_n5596_;
  assign new_n5598_ = ~pstart_0_ & new_n5597_;
  assign new_n5599_ = ~new_n5594_ & ~new_n5598_;
  assign new_n5600_ = ~new_n5586_ & ~new_n5590_;
  assign new_n5601_ = new_n5599_ & new_n5600_;
  assign new_n5602_ = ~new_n5580_ & ~new_n5582_;
  assign new_n5603_ = ~new_n5571_ & ~new_n5575_;
  assign new_n5604_ = ~new_n5577_ & new_n5603_;
  assign new_n5605_ = new_n5602_ & new_n5604_;
  assign n1512 = ~new_n5601_ | ~new_n5605_;
  assign new_n5607_ = ~pencrypt_0_ & n_n2330;
  assign new_n5608_ = ~new_n1200_ & new_n5607_;
  assign new_n5609_ = ~pstart_0_ & new_n5608_;
  assign new_n5610_ = n_n2425 & n_n2330;
  assign new_n5611_ = ~pencrypt_0_ & new_n5610_;
  assign new_n5612_ = new_n1200_ & new_n5611_;
  assign new_n5613_ = ~pstart_0_ & new_n5612_;
  assign new_n5614_ = pencrypt_0_ & pkey_84_;
  assign new_n5615_ = pstart_0_ & new_n5614_;
  assign new_n5616_ = ~pencrypt_0_ & n_n2425;
  assign new_n5617_ = ~new_n1200_ & new_n5616_;
  assign new_n5618_ = ~pstart_0_ & new_n5617_;
  assign new_n5619_ = pkey_92_ & ~pencrypt_0_;
  assign new_n5620_ = pstart_0_ & new_n5619_;
  assign new_n5621_ = ~n_n2330 & ~new_n1220_;
  assign new_n5622_ = pencrypt_0_ & new_n5621_;
  assign new_n5623_ = n_n2425 & new_n5622_;
  assign new_n5624_ = ~pstart_0_ & new_n5623_;
  assign new_n5625_ = n_n2330 & new_n1220_;
  assign new_n5626_ = pencrypt_0_ & new_n5625_;
  assign new_n5627_ = n_n2425 & new_n5626_;
  assign new_n5628_ = ~pstart_0_ & new_n5627_;
  assign new_n5629_ = ~n_n2425 & ~n_n2330;
  assign new_n5630_ = ~pencrypt_0_ & new_n5629_;
  assign new_n5631_ = new_n1200_ & new_n5630_;
  assign new_n5632_ = ~pstart_0_ & new_n5631_;
  assign new_n5633_ = n_n2330 & ~new_n1220_;
  assign new_n5634_ = pencrypt_0_ & new_n5633_;
  assign new_n5635_ = ~n_n2425 & new_n5634_;
  assign new_n5636_ = ~pstart_0_ & new_n5635_;
  assign new_n5637_ = ~new_n5632_ & ~new_n5636_;
  assign new_n5638_ = ~new_n5624_ & ~new_n5628_;
  assign new_n5639_ = new_n5637_ & new_n5638_;
  assign new_n5640_ = ~new_n5618_ & ~new_n5620_;
  assign new_n5641_ = ~new_n5609_ & ~new_n5613_;
  assign new_n5642_ = ~new_n5615_ & new_n5641_;
  assign new_n5643_ = new_n5640_ & new_n5642_;
  assign n1517 = ~new_n5639_ | ~new_n5643_;
  assign new_n5645_ = ~pencrypt_0_ & n_n2336;
  assign new_n5646_ = ~new_n1200_ & new_n5645_;
  assign new_n5647_ = ~pstart_0_ & new_n5646_;
  assign new_n5648_ = n_n2945 & n_n2336;
  assign new_n5649_ = ~pencrypt_0_ & new_n5648_;
  assign new_n5650_ = new_n1200_ & new_n5649_;
  assign new_n5651_ = ~pstart_0_ & new_n5650_;
  assign new_n5652_ = pkey_77_ & pencrypt_0_;
  assign new_n5653_ = pstart_0_ & new_n5652_;
  assign new_n5654_ = ~pencrypt_0_ & n_n2945;
  assign new_n5655_ = ~new_n1200_ & new_n5654_;
  assign new_n5656_ = ~pstart_0_ & new_n5655_;
  assign new_n5657_ = pkey_85_ & ~pencrypt_0_;
  assign new_n5658_ = pstart_0_ & new_n5657_;
  assign new_n5659_ = ~n_n2336 & ~new_n1220_;
  assign new_n5660_ = pencrypt_0_ & new_n5659_;
  assign new_n5661_ = n_n2945 & new_n5660_;
  assign new_n5662_ = ~pstart_0_ & new_n5661_;
  assign new_n5663_ = n_n2336 & new_n1220_;
  assign new_n5664_ = pencrypt_0_ & new_n5663_;
  assign new_n5665_ = n_n2945 & new_n5664_;
  assign new_n5666_ = ~pstart_0_ & new_n5665_;
  assign new_n5667_ = ~n_n2945 & ~n_n2336;
  assign new_n5668_ = ~pencrypt_0_ & new_n5667_;
  assign new_n5669_ = new_n1200_ & new_n5668_;
  assign new_n5670_ = ~pstart_0_ & new_n5669_;
  assign new_n5671_ = n_n2336 & ~new_n1220_;
  assign new_n5672_ = pencrypt_0_ & new_n5671_;
  assign new_n5673_ = ~n_n2945 & new_n5672_;
  assign new_n5674_ = ~pstart_0_ & new_n5673_;
  assign new_n5675_ = ~new_n5670_ & ~new_n5674_;
  assign new_n5676_ = ~new_n5662_ & ~new_n5666_;
  assign new_n5677_ = new_n5675_ & new_n5676_;
  assign new_n5678_ = ~new_n5656_ & ~new_n5658_;
  assign new_n5679_ = ~new_n5647_ & ~new_n5651_;
  assign new_n5680_ = ~new_n5653_ & new_n5679_;
  assign new_n5681_ = new_n5678_ & new_n5680_;
  assign n1522 = ~new_n5677_ | ~new_n5681_;
  assign new_n5683_ = ~pencrypt_0_ & n_n2346;
  assign new_n5684_ = ~new_n1200_ & new_n5683_;
  assign new_n5685_ = ~pstart_0_ & new_n5684_;
  assign new_n5686_ = n_n2439 & n_n2346;
  assign new_n5687_ = ~pencrypt_0_ & new_n5686_;
  assign new_n5688_ = new_n1200_ & new_n5687_;
  assign new_n5689_ = ~pstart_0_ & new_n5688_;
  assign new_n5690_ = pencrypt_0_ & pkey_102_;
  assign new_n5691_ = pstart_0_ & new_n5690_;
  assign new_n5692_ = ~pencrypt_0_ & n_n2439;
  assign new_n5693_ = ~new_n1200_ & new_n5692_;
  assign new_n5694_ = ~pstart_0_ & new_n5693_;
  assign new_n5695_ = pkey_110_ & ~pencrypt_0_;
  assign new_n5696_ = pstart_0_ & new_n5695_;
  assign new_n5697_ = ~n_n2346 & ~new_n1220_;
  assign new_n5698_ = pencrypt_0_ & new_n5697_;
  assign new_n5699_ = n_n2439 & new_n5698_;
  assign new_n5700_ = ~pstart_0_ & new_n5699_;
  assign new_n5701_ = n_n2346 & new_n1220_;
  assign new_n5702_ = pencrypt_0_ & new_n5701_;
  assign new_n5703_ = n_n2439 & new_n5702_;
  assign new_n5704_ = ~pstart_0_ & new_n5703_;
  assign new_n5705_ = ~n_n2439 & ~n_n2346;
  assign new_n5706_ = ~pencrypt_0_ & new_n5705_;
  assign new_n5707_ = new_n1200_ & new_n5706_;
  assign new_n5708_ = ~pstart_0_ & new_n5707_;
  assign new_n5709_ = n_n2346 & ~new_n1220_;
  assign new_n5710_ = pencrypt_0_ & new_n5709_;
  assign new_n5711_ = ~n_n2439 & new_n5710_;
  assign new_n5712_ = ~pstart_0_ & new_n5711_;
  assign new_n5713_ = ~new_n5708_ & ~new_n5712_;
  assign new_n5714_ = ~new_n5700_ & ~new_n5704_;
  assign new_n5715_ = new_n5713_ & new_n5714_;
  assign new_n5716_ = ~new_n5694_ & ~new_n5696_;
  assign new_n5717_ = ~new_n5685_ & ~new_n5689_;
  assign new_n5718_ = ~new_n5691_ & new_n5717_;
  assign new_n5719_ = new_n5716_ & new_n5718_;
  assign n1527 = ~new_n5715_ | ~new_n5719_;
  assign new_n5721_ = ~pencrypt_0_ & n_n2359;
  assign new_n5722_ = ~new_n1200_ & new_n5721_;
  assign new_n5723_ = ~pstart_0_ & new_n5722_;
  assign new_n5724_ = n_n2976 & n_n2359;
  assign new_n5725_ = ~pencrypt_0_ & new_n5724_;
  assign new_n5726_ = new_n1200_ & new_n5725_;
  assign new_n5727_ = ~pstart_0_ & new_n5726_;
  assign new_n5728_ = pkey_5_ & pencrypt_0_;
  assign new_n5729_ = pstart_0_ & new_n5728_;
  assign new_n5730_ = ~pencrypt_0_ & n_n2976;
  assign new_n5731_ = ~new_n1200_ & new_n5730_;
  assign new_n5732_ = ~pstart_0_ & new_n5731_;
  assign new_n5733_ = ~pencrypt_0_ & pkey_13_;
  assign new_n5734_ = pstart_0_ & new_n5733_;
  assign new_n5735_ = ~n_n2359 & ~new_n1220_;
  assign new_n5736_ = pencrypt_0_ & new_n5735_;
  assign new_n5737_ = n_n2976 & new_n5736_;
  assign new_n5738_ = ~pstart_0_ & new_n5737_;
  assign new_n5739_ = n_n2359 & new_n1220_;
  assign new_n5740_ = pencrypt_0_ & new_n5739_;
  assign new_n5741_ = n_n2976 & new_n5740_;
  assign new_n5742_ = ~pstart_0_ & new_n5741_;
  assign new_n5743_ = ~n_n2976 & ~n_n2359;
  assign new_n5744_ = ~pencrypt_0_ & new_n5743_;
  assign new_n5745_ = new_n1200_ & new_n5744_;
  assign new_n5746_ = ~pstart_0_ & new_n5745_;
  assign new_n5747_ = n_n2359 & ~new_n1220_;
  assign new_n5748_ = pencrypt_0_ & new_n5747_;
  assign new_n5749_ = ~n_n2976 & new_n5748_;
  assign new_n5750_ = ~pstart_0_ & new_n5749_;
  assign new_n5751_ = ~new_n5746_ & ~new_n5750_;
  assign new_n5752_ = ~new_n5738_ & ~new_n5742_;
  assign new_n5753_ = new_n5751_ & new_n5752_;
  assign new_n5754_ = ~new_n5732_ & ~new_n5734_;
  assign new_n5755_ = ~new_n5723_ & ~new_n5727_;
  assign new_n5756_ = ~new_n5729_ & new_n5755_;
  assign new_n5757_ = new_n5754_ & new_n5756_;
  assign n1532 = ~new_n5753_ | ~new_n5757_;
  assign new_n5759_ = new_n1200_ & new_n2198_;
  assign new_n5760_ = ~pstart_0_ & new_n5759_;
  assign new_n5761_ = ~new_n1200_ & new_n2193_;
  assign new_n5762_ = ~pstart_0_ & new_n5761_;
  assign new_n5763_ = pkey_251_ & pencrypt_0_;
  assign new_n5764_ = pstart_0_ & new_n5763_;
  assign new_n5765_ = new_n1200_ & new_n2189_;
  assign new_n5766_ = ~pstart_0_ & new_n5765_;
  assign new_n5767_ = pkey_194_ & ~pencrypt_0_;
  assign new_n5768_ = pstart_0_ & new_n5767_;
  assign new_n5769_ = n_n2376 & new_n1220_;
  assign new_n5770_ = pencrypt_0_ & new_n5769_;
  assign new_n5771_ = ~n_n2281 & new_n5770_;
  assign new_n5772_ = ~pstart_0_ & new_n5771_;
  assign new_n5773_ = ~n_n2376 & new_n1220_;
  assign new_n5774_ = pencrypt_0_ & new_n5773_;
  assign new_n5775_ = n_n2281 & new_n5774_;
  assign new_n5776_ = ~pstart_0_ & new_n5775_;
  assign new_n5777_ = ~new_n1200_ & new_n2212_;
  assign new_n5778_ = ~pstart_0_ & new_n5777_;
  assign new_n5779_ = n_n2376 & ~new_n1220_;
  assign new_n5780_ = pencrypt_0_ & new_n5779_;
  assign new_n5781_ = n_n2281 & new_n5780_;
  assign new_n5782_ = ~pstart_0_ & new_n5781_;
  assign new_n5783_ = ~new_n5778_ & ~new_n5782_;
  assign new_n5784_ = ~new_n5772_ & ~new_n5776_;
  assign new_n5785_ = new_n5783_ & new_n5784_;
  assign new_n5786_ = ~new_n5766_ & ~new_n5768_;
  assign new_n5787_ = ~new_n5760_ & ~new_n5762_;
  assign new_n5788_ = ~new_n5764_ & new_n5787_;
  assign new_n5789_ = new_n5786_ & new_n5788_;
  assign n1537 = ~new_n5785_ | ~new_n5789_;
  assign new_n5791_ = ~pencrypt_0_ & n_n2291;
  assign new_n5792_ = ~new_n1200_ & new_n5791_;
  assign new_n5793_ = ~pstart_0_ & new_n5792_;
  assign new_n5794_ = n_n2386 & n_n2291;
  assign new_n5795_ = ~pencrypt_0_ & new_n5794_;
  assign new_n5796_ = new_n1200_ & new_n5795_;
  assign new_n5797_ = ~pstart_0_ & new_n5796_;
  assign new_n5798_ = pkey_229_ & pencrypt_0_;
  assign new_n5799_ = pstart_0_ & new_n5798_;
  assign new_n5800_ = ~pencrypt_0_ & n_n2386;
  assign new_n5801_ = ~new_n1200_ & new_n5800_;
  assign new_n5802_ = ~pstart_0_ & new_n5801_;
  assign new_n5803_ = pkey_237_ & ~pencrypt_0_;
  assign new_n5804_ = pstart_0_ & new_n5803_;
  assign new_n5805_ = ~n_n2291 & ~new_n1220_;
  assign new_n5806_ = pencrypt_0_ & new_n5805_;
  assign new_n5807_ = n_n2386 & new_n5806_;
  assign new_n5808_ = ~pstart_0_ & new_n5807_;
  assign new_n5809_ = n_n2291 & new_n1220_;
  assign new_n5810_ = pencrypt_0_ & new_n5809_;
  assign new_n5811_ = n_n2386 & new_n5810_;
  assign new_n5812_ = ~pstart_0_ & new_n5811_;
  assign new_n5813_ = ~n_n2386 & ~n_n2291;
  assign new_n5814_ = ~pencrypt_0_ & new_n5813_;
  assign new_n5815_ = new_n1200_ & new_n5814_;
  assign new_n5816_ = ~pstart_0_ & new_n5815_;
  assign new_n5817_ = n_n2291 & ~new_n1220_;
  assign new_n5818_ = pencrypt_0_ & new_n5817_;
  assign new_n5819_ = ~n_n2386 & new_n5818_;
  assign new_n5820_ = ~pstart_0_ & new_n5819_;
  assign new_n5821_ = ~new_n5816_ & ~new_n5820_;
  assign new_n5822_ = ~new_n5808_ & ~new_n5812_;
  assign new_n5823_ = new_n5821_ & new_n5822_;
  assign new_n5824_ = ~new_n5802_ & ~new_n5804_;
  assign new_n5825_ = ~new_n5793_ & ~new_n5797_;
  assign new_n5826_ = ~new_n5799_ & new_n5825_;
  assign new_n5827_ = new_n5824_ & new_n5826_;
  assign n1542 = ~new_n5823_ | ~new_n5827_;
  assign new_n5829_ = ~pencrypt_0_ & n_n2299;
  assign new_n5830_ = ~new_n1200_ & new_n5829_;
  assign new_n5831_ = ~pstart_0_ & new_n5830_;
  assign new_n5832_ = n_n2393 & n_n2299;
  assign new_n5833_ = ~pencrypt_0_ & new_n5832_;
  assign new_n5834_ = new_n1200_ & new_n5833_;
  assign new_n5835_ = ~pstart_0_ & new_n5834_;
  assign new_n5836_ = pkey_238_ & pencrypt_0_;
  assign new_n5837_ = pstart_0_ & new_n5836_;
  assign new_n5838_ = ~pencrypt_0_ & n_n2393;
  assign new_n5839_ = ~new_n1200_ & new_n5838_;
  assign new_n5840_ = ~pstart_0_ & new_n5839_;
  assign new_n5841_ = pkey_246_ & ~pencrypt_0_;
  assign new_n5842_ = pstart_0_ & new_n5841_;
  assign new_n5843_ = ~n_n2299 & ~new_n1220_;
  assign new_n5844_ = pencrypt_0_ & new_n5843_;
  assign new_n5845_ = n_n2393 & new_n5844_;
  assign new_n5846_ = ~pstart_0_ & new_n5845_;
  assign new_n5847_ = n_n2299 & new_n1220_;
  assign new_n5848_ = pencrypt_0_ & new_n5847_;
  assign new_n5849_ = n_n2393 & new_n5848_;
  assign new_n5850_ = ~pstart_0_ & new_n5849_;
  assign new_n5851_ = ~n_n2393 & ~n_n2299;
  assign new_n5852_ = ~pencrypt_0_ & new_n5851_;
  assign new_n5853_ = new_n1200_ & new_n5852_;
  assign new_n5854_ = ~pstart_0_ & new_n5853_;
  assign new_n5855_ = n_n2299 & ~new_n1220_;
  assign new_n5856_ = pencrypt_0_ & new_n5855_;
  assign new_n5857_ = ~n_n2393 & new_n5856_;
  assign new_n5858_ = ~pstart_0_ & new_n5857_;
  assign new_n5859_ = ~new_n5854_ & ~new_n5858_;
  assign new_n5860_ = ~new_n5846_ & ~new_n5850_;
  assign new_n5861_ = new_n5859_ & new_n5860_;
  assign new_n5862_ = ~new_n5840_ & ~new_n5842_;
  assign new_n5863_ = ~new_n5831_ & ~new_n5835_;
  assign new_n5864_ = ~new_n5837_ & new_n5863_;
  assign new_n5865_ = new_n5862_ & new_n5864_;
  assign n1547 = ~new_n5861_ | ~new_n5865_;
  assign new_n5867_ = ~pencrypt_0_ & n_n2306;
  assign new_n5868_ = ~new_n1200_ & new_n5867_;
  assign new_n5869_ = ~pstart_0_ & new_n5868_;
  assign new_n5870_ = n_n2401 & n_n2306;
  assign new_n5871_ = ~pencrypt_0_ & new_n5870_;
  assign new_n5872_ = new_n1200_ & new_n5871_;
  assign new_n5873_ = ~pstart_0_ & new_n5872_;
  assign new_n5874_ = pkey_148_ & pencrypt_0_;
  assign new_n5875_ = pstart_0_ & new_n5874_;
  assign new_n5876_ = ~pencrypt_0_ & n_n2401;
  assign new_n5877_ = ~new_n1200_ & new_n5876_;
  assign new_n5878_ = ~pstart_0_ & new_n5877_;
  assign new_n5879_ = pkey_156_ & ~pencrypt_0_;
  assign new_n5880_ = pstart_0_ & new_n5879_;
  assign new_n5881_ = ~n_n2306 & ~new_n1220_;
  assign new_n5882_ = pencrypt_0_ & new_n5881_;
  assign new_n5883_ = n_n2401 & new_n5882_;
  assign new_n5884_ = ~pstart_0_ & new_n5883_;
  assign new_n5885_ = n_n2306 & new_n1220_;
  assign new_n5886_ = pencrypt_0_ & new_n5885_;
  assign new_n5887_ = n_n2401 & new_n5886_;
  assign new_n5888_ = ~pstart_0_ & new_n5887_;
  assign new_n5889_ = ~n_n2401 & ~n_n2306;
  assign new_n5890_ = ~pencrypt_0_ & new_n5889_;
  assign new_n5891_ = new_n1200_ & new_n5890_;
  assign new_n5892_ = ~pstart_0_ & new_n5891_;
  assign new_n5893_ = n_n2306 & ~new_n1220_;
  assign new_n5894_ = pencrypt_0_ & new_n5893_;
  assign new_n5895_ = ~n_n2401 & new_n5894_;
  assign new_n5896_ = ~pstart_0_ & new_n5895_;
  assign new_n5897_ = ~new_n5892_ & ~new_n5896_;
  assign new_n5898_ = ~new_n5884_ & ~new_n5888_;
  assign new_n5899_ = new_n5897_ & new_n5898_;
  assign new_n5900_ = ~new_n5878_ & ~new_n5880_;
  assign new_n5901_ = ~new_n5869_ & ~new_n5873_;
  assign new_n5902_ = ~new_n5875_ & new_n5901_;
  assign new_n5903_ = new_n5900_ & new_n5902_;
  assign n1552 = ~new_n5899_ | ~new_n5903_;
  assign new_n5905_ = ~pencrypt_0_ & n_n2314;
  assign new_n5906_ = ~new_n1200_ & new_n5905_;
  assign new_n5907_ = ~pstart_0_ & new_n5906_;
  assign new_n5908_ = n_n2409 & n_n2314;
  assign new_n5909_ = ~pencrypt_0_ & new_n5908_;
  assign new_n5910_ = new_n1200_ & new_n5909_;
  assign new_n5911_ = ~pstart_0_ & new_n5910_;
  assign new_n5912_ = pkey_157_ & pencrypt_0_;
  assign new_n5913_ = pstart_0_ & new_n5912_;
  assign new_n5914_ = ~pencrypt_0_ & n_n2409;
  assign new_n5915_ = ~new_n1200_ & new_n5914_;
  assign new_n5916_ = ~pstart_0_ & new_n5915_;
  assign new_n5917_ = pkey_165_ & ~pencrypt_0_;
  assign new_n5918_ = pstart_0_ & new_n5917_;
  assign new_n5919_ = ~n_n2314 & ~new_n1220_;
  assign new_n5920_ = pencrypt_0_ & new_n5919_;
  assign new_n5921_ = n_n2409 & new_n5920_;
  assign new_n5922_ = ~pstart_0_ & new_n5921_;
  assign new_n5923_ = n_n2314 & new_n1220_;
  assign new_n5924_ = pencrypt_0_ & new_n5923_;
  assign new_n5925_ = n_n2409 & new_n5924_;
  assign new_n5926_ = ~pstart_0_ & new_n5925_;
  assign new_n5927_ = ~n_n2409 & ~n_n2314;
  assign new_n5928_ = ~pencrypt_0_ & new_n5927_;
  assign new_n5929_ = new_n1200_ & new_n5928_;
  assign new_n5930_ = ~pstart_0_ & new_n5929_;
  assign new_n5931_ = n_n2314 & ~new_n1220_;
  assign new_n5932_ = pencrypt_0_ & new_n5931_;
  assign new_n5933_ = ~n_n2409 & new_n5932_;
  assign new_n5934_ = ~pstart_0_ & new_n5933_;
  assign new_n5935_ = ~new_n5930_ & ~new_n5934_;
  assign new_n5936_ = ~new_n5922_ & ~new_n5926_;
  assign new_n5937_ = new_n5935_ & new_n5936_;
  assign new_n5938_ = ~new_n5916_ & ~new_n5918_;
  assign new_n5939_ = ~new_n5907_ & ~new_n5911_;
  assign new_n5940_ = ~new_n5913_ & new_n5939_;
  assign new_n5941_ = new_n5938_ & new_n5940_;
  assign n1557 = ~new_n5937_ | ~new_n5941_;
  assign new_n5943_ = ~pencrypt_0_ & n_n2322;
  assign new_n5944_ = ~new_n1200_ & new_n5943_;
  assign new_n5945_ = ~pstart_0_ & new_n5944_;
  assign new_n5946_ = n_n2416 & n_n2322;
  assign new_n5947_ = ~pencrypt_0_ & new_n5946_;
  assign new_n5948_ = new_n1200_ & new_n5947_;
  assign new_n5949_ = ~pstart_0_ & new_n5948_;
  assign new_n5950_ = pkey_166_ & pencrypt_0_;
  assign new_n5951_ = pstart_0_ & new_n5950_;
  assign new_n5952_ = ~pencrypt_0_ & n_n2416;
  assign new_n5953_ = ~new_n1200_ & new_n5952_;
  assign new_n5954_ = ~pstart_0_ & new_n5953_;
  assign new_n5955_ = ~pencrypt_0_ & pkey_174_;
  assign new_n5956_ = pstart_0_ & new_n5955_;
  assign new_n5957_ = ~n_n2322 & ~new_n1220_;
  assign new_n5958_ = pencrypt_0_ & new_n5957_;
  assign new_n5959_ = n_n2416 & new_n5958_;
  assign new_n5960_ = ~pstart_0_ & new_n5959_;
  assign new_n5961_ = n_n2322 & new_n1220_;
  assign new_n5962_ = pencrypt_0_ & new_n5961_;
  assign new_n5963_ = n_n2416 & new_n5962_;
  assign new_n5964_ = ~pstart_0_ & new_n5963_;
  assign new_n5965_ = ~n_n2416 & ~n_n2322;
  assign new_n5966_ = ~pencrypt_0_ & new_n5965_;
  assign new_n5967_ = new_n1200_ & new_n5966_;
  assign new_n5968_ = ~pstart_0_ & new_n5967_;
  assign new_n5969_ = n_n2322 & ~new_n1220_;
  assign new_n5970_ = pencrypt_0_ & new_n5969_;
  assign new_n5971_ = ~n_n2416 & new_n5970_;
  assign new_n5972_ = ~pstart_0_ & new_n5971_;
  assign new_n5973_ = ~new_n5968_ & ~new_n5972_;
  assign new_n5974_ = ~new_n5960_ & ~new_n5964_;
  assign new_n5975_ = new_n5973_ & new_n5974_;
  assign new_n5976_ = ~new_n5954_ & ~new_n5956_;
  assign new_n5977_ = ~new_n5945_ & ~new_n5949_;
  assign new_n5978_ = ~new_n5951_ & new_n5977_;
  assign new_n5979_ = new_n5976_ & new_n5978_;
  assign n1562 = ~new_n5975_ | ~new_n5979_;
  assign new_n5981_ = ~pencrypt_0_ & n_n2806;
  assign new_n5982_ = ~new_n1200_ & new_n5981_;
  assign new_n5983_ = ~pstart_0_ & new_n5982_;
  assign new_n5984_ = n_n2424 & n_n2806;
  assign new_n5985_ = ~pencrypt_0_ & new_n5984_;
  assign new_n5986_ = new_n1200_ & new_n5985_;
  assign new_n5987_ = ~pstart_0_ & new_n5986_;
  assign new_n5988_ = pkey_76_ & pencrypt_0_;
  assign new_n5989_ = pstart_0_ & new_n5988_;
  assign new_n5990_ = ~pencrypt_0_ & n_n2424;
  assign new_n5991_ = ~new_n1200_ & new_n5990_;
  assign new_n5992_ = ~pstart_0_ & new_n5991_;
  assign new_n5993_ = ~pencrypt_0_ & pkey_84_;
  assign new_n5994_ = pstart_0_ & new_n5993_;
  assign new_n5995_ = ~n_n2806 & ~new_n1220_;
  assign new_n5996_ = pencrypt_0_ & new_n5995_;
  assign new_n5997_ = n_n2424 & new_n5996_;
  assign new_n5998_ = ~pstart_0_ & new_n5997_;
  assign new_n5999_ = n_n2806 & new_n1220_;
  assign new_n6000_ = pencrypt_0_ & new_n5999_;
  assign new_n6001_ = n_n2424 & new_n6000_;
  assign new_n6002_ = ~pstart_0_ & new_n6001_;
  assign new_n6003_ = ~n_n2424 & ~n_n2806;
  assign new_n6004_ = ~pencrypt_0_ & new_n6003_;
  assign new_n6005_ = new_n1200_ & new_n6004_;
  assign new_n6006_ = ~pstart_0_ & new_n6005_;
  assign new_n6007_ = n_n2806 & ~new_n1220_;
  assign new_n6008_ = pencrypt_0_ & new_n6007_;
  assign new_n6009_ = ~n_n2424 & new_n6008_;
  assign new_n6010_ = ~pstart_0_ & new_n6009_;
  assign new_n6011_ = ~new_n6006_ & ~new_n6010_;
  assign new_n6012_ = ~new_n5998_ & ~new_n6002_;
  assign new_n6013_ = new_n6011_ & new_n6012_;
  assign new_n6014_ = ~new_n5992_ & ~new_n5994_;
  assign new_n6015_ = ~new_n5983_ & ~new_n5987_;
  assign new_n6016_ = ~new_n5989_ & new_n6015_;
  assign new_n6017_ = new_n6014_ & new_n6016_;
  assign n1567 = ~new_n6013_ | ~new_n6017_;
  assign new_n6019_ = ~pencrypt_0_ & n_n2337;
  assign new_n6020_ = ~new_n1200_ & new_n6019_;
  assign new_n6021_ = ~pstart_0_ & new_n6020_;
  assign new_n6022_ = n_n2431 & n_n2337;
  assign new_n6023_ = ~pencrypt_0_ & new_n6022_;
  assign new_n6024_ = new_n1200_ & new_n6023_;
  assign new_n6025_ = ~pstart_0_ & new_n6024_;
  assign new_n6026_ = pkey_85_ & pencrypt_0_;
  assign new_n6027_ = pstart_0_ & new_n6026_;
  assign new_n6028_ = ~pencrypt_0_ & n_n2431;
  assign new_n6029_ = ~new_n1200_ & new_n6028_;
  assign new_n6030_ = ~pstart_0_ & new_n6029_;
  assign new_n6031_ = pkey_93_ & ~pencrypt_0_;
  assign new_n6032_ = pstart_0_ & new_n6031_;
  assign new_n6033_ = ~n_n2337 & ~new_n1220_;
  assign new_n6034_ = pencrypt_0_ & new_n6033_;
  assign new_n6035_ = n_n2431 & new_n6034_;
  assign new_n6036_ = ~pstart_0_ & new_n6035_;
  assign new_n6037_ = n_n2337 & new_n1220_;
  assign new_n6038_ = pencrypt_0_ & new_n6037_;
  assign new_n6039_ = n_n2431 & new_n6038_;
  assign new_n6040_ = ~pstart_0_ & new_n6039_;
  assign new_n6041_ = ~n_n2431 & ~n_n2337;
  assign new_n6042_ = ~pencrypt_0_ & new_n6041_;
  assign new_n6043_ = new_n1200_ & new_n6042_;
  assign new_n6044_ = ~pstart_0_ & new_n6043_;
  assign new_n6045_ = n_n2337 & ~new_n1220_;
  assign new_n6046_ = pencrypt_0_ & new_n6045_;
  assign new_n6047_ = ~n_n2431 & new_n6046_;
  assign new_n6048_ = ~pstart_0_ & new_n6047_;
  assign new_n6049_ = ~new_n6044_ & ~new_n6048_;
  assign new_n6050_ = ~new_n6036_ & ~new_n6040_;
  assign new_n6051_ = new_n6049_ & new_n6050_;
  assign new_n6052_ = ~new_n6030_ & ~new_n6032_;
  assign new_n6053_ = ~new_n6021_ & ~new_n6025_;
  assign new_n6054_ = ~new_n6027_ & new_n6053_;
  assign new_n6055_ = new_n6052_ & new_n6054_;
  assign n1572 = ~new_n6051_ | ~new_n6055_;
  assign new_n6057_ = ~pencrypt_0_ & n_n2345;
  assign new_n6058_ = ~new_n1200_ & new_n6057_;
  assign new_n6059_ = ~pstart_0_ & new_n6058_;
  assign new_n6060_ = n_n2438 & n_n2345;
  assign new_n6061_ = ~pencrypt_0_ & new_n6060_;
  assign new_n6062_ = new_n1200_ & new_n6061_;
  assign new_n6063_ = ~pstart_0_ & new_n6062_;
  assign new_n6064_ = pkey_94_ & pencrypt_0_;
  assign new_n6065_ = pstart_0_ & new_n6064_;
  assign new_n6066_ = ~pencrypt_0_ & n_n2438;
  assign new_n6067_ = ~new_n1200_ & new_n6066_;
  assign new_n6068_ = ~pstart_0_ & new_n6067_;
  assign new_n6069_ = ~pencrypt_0_ & pkey_102_;
  assign new_n6070_ = pstart_0_ & new_n6069_;
  assign new_n6071_ = ~n_n2345 & ~new_n1220_;
  assign new_n6072_ = pencrypt_0_ & new_n6071_;
  assign new_n6073_ = n_n2438 & new_n6072_;
  assign new_n6074_ = ~pstart_0_ & new_n6073_;
  assign new_n6075_ = n_n2345 & new_n1220_;
  assign new_n6076_ = pencrypt_0_ & new_n6075_;
  assign new_n6077_ = n_n2438 & new_n6076_;
  assign new_n6078_ = ~pstart_0_ & new_n6077_;
  assign new_n6079_ = ~n_n2438 & ~n_n2345;
  assign new_n6080_ = ~pencrypt_0_ & new_n6079_;
  assign new_n6081_ = new_n1200_ & new_n6080_;
  assign new_n6082_ = ~pstart_0_ & new_n6081_;
  assign new_n6083_ = n_n2345 & ~new_n1220_;
  assign new_n6084_ = pencrypt_0_ & new_n6083_;
  assign new_n6085_ = ~n_n2438 & new_n6084_;
  assign new_n6086_ = ~pstart_0_ & new_n6085_;
  assign new_n6087_ = ~new_n6082_ & ~new_n6086_;
  assign new_n6088_ = ~new_n6074_ & ~new_n6078_;
  assign new_n6089_ = new_n6087_ & new_n6088_;
  assign new_n6090_ = ~new_n6068_ & ~new_n6070_;
  assign new_n6091_ = ~new_n6059_ & ~new_n6063_;
  assign new_n6092_ = ~new_n6065_ & new_n6091_;
  assign new_n6093_ = new_n6090_ & new_n6092_;
  assign n1577 = ~new_n6089_ | ~new_n6093_;
  assign new_n6095_ = ~new_n1200_ & new_n2160_;
  assign new_n6096_ = ~pstart_0_ & new_n6095_;
  assign new_n6097_ = new_n1200_ & new_n2155_;
  assign new_n6098_ = ~pstart_0_ & new_n6097_;
  assign new_n6099_ = pencrypt_0_ & pkey_22_;
  assign new_n6100_ = pstart_0_ & new_n6099_;
  assign new_n6101_ = ~new_n1200_ & new_n2151_;
  assign new_n6102_ = ~pstart_0_ & new_n6101_;
  assign new_n6103_ = ~pencrypt_0_ & pkey_30_;
  assign new_n6104_ = pstart_0_ & new_n6103_;
  assign new_n6105_ = ~n_n2368 & ~new_n1220_;
  assign new_n6106_ = pencrypt_0_ & new_n6105_;
  assign new_n6107_ = n_n2461 & new_n6106_;
  assign new_n6108_ = ~pstart_0_ & new_n6107_;
  assign new_n6109_ = n_n2368 & new_n1220_;
  assign new_n6110_ = pencrypt_0_ & new_n6109_;
  assign new_n6111_ = n_n2461 & new_n6110_;
  assign new_n6112_ = ~pstart_0_ & new_n6111_;
  assign new_n6113_ = new_n1200_ & new_n2174_;
  assign new_n6114_ = ~pstart_0_ & new_n6113_;
  assign new_n6115_ = n_n2368 & ~new_n1220_;
  assign new_n6116_ = pencrypt_0_ & new_n6115_;
  assign new_n6117_ = ~n_n2461 & new_n6116_;
  assign new_n6118_ = ~pstart_0_ & new_n6117_;
  assign new_n6119_ = ~new_n6114_ & ~new_n6118_;
  assign new_n6120_ = ~new_n6108_ & ~new_n6112_;
  assign new_n6121_ = new_n6119_ & new_n6120_;
  assign new_n6122_ = ~new_n6102_ & ~new_n6104_;
  assign new_n6123_ = ~new_n6096_ & ~new_n6098_;
  assign new_n6124_ = ~new_n6100_ & new_n6123_;
  assign new_n6125_ = new_n6122_ & new_n6124_;
  assign n1582 = ~new_n6121_ | ~new_n6125_;
  assign new_n6127_ = new_n1200_ & new_n3666_;
  assign new_n6128_ = ~pstart_0_ & new_n6127_;
  assign new_n6129_ = ~new_n1200_ & new_n3661_;
  assign new_n6130_ = ~pstart_0_ & new_n6129_;
  assign new_n6131_ = pkey_136_ & pencrypt_0_;
  assign new_n6132_ = pstart_0_ & new_n6131_;
  assign new_n6133_ = new_n1200_ & new_n3657_;
  assign new_n6134_ = ~pstart_0_ & new_n6133_;
  assign new_n6135_ = pkey_144_ & ~pencrypt_0_;
  assign new_n6136_ = pstart_0_ & new_n6135_;
  assign new_n6137_ = n_n2413 & new_n1220_;
  assign new_n6138_ = pencrypt_0_ & new_n6137_;
  assign new_n6139_ = ~n_n2319 & new_n6138_;
  assign new_n6140_ = ~pstart_0_ & new_n6139_;
  assign new_n6141_ = ~n_n2413 & new_n1220_;
  assign new_n6142_ = pencrypt_0_ & new_n6141_;
  assign new_n6143_ = n_n2319 & new_n6142_;
  assign new_n6144_ = ~pstart_0_ & new_n6143_;
  assign new_n6145_ = ~new_n1200_ & new_n3680_;
  assign new_n6146_ = ~pstart_0_ & new_n6145_;
  assign new_n6147_ = n_n2413 & ~new_n1220_;
  assign new_n6148_ = pencrypt_0_ & new_n6147_;
  assign new_n6149_ = n_n2319 & new_n6148_;
  assign new_n6150_ = ~pstart_0_ & new_n6149_;
  assign new_n6151_ = ~new_n6146_ & ~new_n6150_;
  assign new_n6152_ = ~new_n6140_ & ~new_n6144_;
  assign new_n6153_ = new_n6151_ & new_n6152_;
  assign new_n6154_ = ~new_n6134_ & ~new_n6136_;
  assign new_n6155_ = ~new_n6128_ & ~new_n6130_;
  assign new_n6156_ = ~new_n6132_ & new_n6155_;
  assign new_n6157_ = new_n6154_ & new_n6156_;
  assign n1587 = ~new_n6153_ | ~new_n6157_;
  assign new_n6159_ = new_n1200_ & new_n3704_;
  assign new_n6160_ = ~pstart_0_ & new_n6159_;
  assign new_n6161_ = ~new_n1200_ & new_n3699_;
  assign new_n6162_ = ~pstart_0_ & new_n6161_;
  assign new_n6163_ = pkey_66_ & pencrypt_0_;
  assign new_n6164_ = pstart_0_ & new_n6163_;
  assign new_n6165_ = new_n1200_ & new_n3695_;
  assign new_n6166_ = ~pstart_0_ & new_n6165_;
  assign new_n6167_ = pkey_74_ & ~pencrypt_0_;
  assign new_n6168_ = pstart_0_ & new_n6167_;
  assign new_n6169_ = n_n2423 & new_n1220_;
  assign new_n6170_ = pencrypt_0_ & new_n6169_;
  assign new_n6171_ = ~n_n2329 & new_n6170_;
  assign new_n6172_ = ~pstart_0_ & new_n6171_;
  assign new_n6173_ = ~n_n2423 & new_n1220_;
  assign new_n6174_ = pencrypt_0_ & new_n6173_;
  assign new_n6175_ = n_n2329 & new_n6174_;
  assign new_n6176_ = ~pstart_0_ & new_n6175_;
  assign new_n6177_ = ~new_n1200_ & new_n3718_;
  assign new_n6178_ = ~pstart_0_ & new_n6177_;
  assign new_n6179_ = n_n2423 & ~new_n1220_;
  assign new_n6180_ = pencrypt_0_ & new_n6179_;
  assign new_n6181_ = n_n2329 & new_n6180_;
  assign new_n6182_ = ~pstart_0_ & new_n6181_;
  assign new_n6183_ = ~new_n6178_ & ~new_n6182_;
  assign new_n6184_ = ~new_n6172_ & ~new_n6176_;
  assign new_n6185_ = new_n6183_ & new_n6184_;
  assign new_n6186_ = ~new_n6166_ & ~new_n6168_;
  assign new_n6187_ = ~new_n6160_ & ~new_n6162_;
  assign new_n6188_ = ~new_n6164_ & new_n6187_;
  assign new_n6189_ = new_n6186_ & new_n6188_;
  assign n1592 = ~new_n6185_ | ~new_n6189_;
  assign new_n6191_ = new_n1200_ & new_n3742_;
  assign new_n6192_ = ~pstart_0_ & new_n6191_;
  assign new_n6193_ = ~new_n1200_ & new_n3737_;
  assign new_n6194_ = ~pstart_0_ & new_n6193_;
  assign new_n6195_ = pkey_89_ & pencrypt_0_;
  assign new_n6196_ = pstart_0_ & new_n6195_;
  assign new_n6197_ = new_n1200_ & new_n3733_;
  assign new_n6198_ = ~pstart_0_ & new_n6197_;
  assign new_n6199_ = pkey_97_ & ~pencrypt_0_;
  assign new_n6200_ = pstart_0_ & new_n6199_;
  assign new_n6201_ = n_n2432 & new_n1220_;
  assign new_n6202_ = pencrypt_0_ & new_n6201_;
  assign new_n6203_ = ~n_n2338 & new_n6202_;
  assign new_n6204_ = ~pstart_0_ & new_n6203_;
  assign new_n6205_ = ~n_n2432 & new_n1220_;
  assign new_n6206_ = pencrypt_0_ & new_n6205_;
  assign new_n6207_ = n_n2338 & new_n6206_;
  assign new_n6208_ = ~pstart_0_ & new_n6207_;
  assign new_n6209_ = ~new_n1200_ & new_n3756_;
  assign new_n6210_ = ~pstart_0_ & new_n6209_;
  assign new_n6211_ = n_n2432 & ~new_n1220_;
  assign new_n6212_ = pencrypt_0_ & new_n6211_;
  assign new_n6213_ = n_n2338 & new_n6212_;
  assign new_n6214_ = ~pstart_0_ & new_n6213_;
  assign new_n6215_ = ~new_n6210_ & ~new_n6214_;
  assign new_n6216_ = ~new_n6204_ & ~new_n6208_;
  assign new_n6217_ = new_n6215_ & new_n6216_;
  assign new_n6218_ = ~new_n6198_ & ~new_n6200_;
  assign new_n6219_ = ~new_n6192_ & ~new_n6194_;
  assign new_n6220_ = ~new_n6196_ & new_n6219_;
  assign new_n6221_ = new_n6218_ & new_n6220_;
  assign n1597 = ~new_n6217_ | ~new_n6221_;
  assign new_n6223_ = new_n1200_ & new_n3780_;
  assign new_n6224_ = ~pstart_0_ & new_n6223_;
  assign new_n6225_ = ~new_n1200_ & new_n3775_;
  assign new_n6226_ = ~pstart_0_ & new_n6225_;
  assign new_n6227_ = pkey_112_ & pencrypt_0_;
  assign new_n6228_ = pstart_0_ & new_n6227_;
  assign new_n6229_ = new_n1200_ & new_n3771_;
  assign new_n6230_ = ~pstart_0_ & new_n6229_;
  assign new_n6231_ = pkey_120_ & ~pencrypt_0_;
  assign new_n6232_ = pstart_0_ & new_n6231_;
  assign new_n6233_ = n_n2441 & new_n1220_;
  assign new_n6234_ = pencrypt_0_ & new_n6233_;
  assign new_n6235_ = ~n_n2348 & new_n6234_;
  assign new_n6236_ = ~pstart_0_ & new_n6235_;
  assign new_n6237_ = ~n_n2441 & new_n1220_;
  assign new_n6238_ = pencrypt_0_ & new_n6237_;
  assign new_n6239_ = n_n2348 & new_n6238_;
  assign new_n6240_ = ~pstart_0_ & new_n6239_;
  assign new_n6241_ = ~new_n1200_ & new_n3794_;
  assign new_n6242_ = ~pstart_0_ & new_n6241_;
  assign new_n6243_ = n_n2441 & ~new_n1220_;
  assign new_n6244_ = pencrypt_0_ & new_n6243_;
  assign new_n6245_ = n_n2348 & new_n6244_;
  assign new_n6246_ = ~pstart_0_ & new_n6245_;
  assign new_n6247_ = ~new_n6242_ & ~new_n6246_;
  assign new_n6248_ = ~new_n6236_ & ~new_n6240_;
  assign new_n6249_ = new_n6247_ & new_n6248_;
  assign new_n6250_ = ~new_n6230_ & ~new_n6232_;
  assign new_n6251_ = ~new_n6224_ & ~new_n6226_;
  assign new_n6252_ = ~new_n6228_ & new_n6251_;
  assign new_n6253_ = new_n6250_ & new_n6252_;
  assign n1602 = ~new_n6249_ | ~new_n6253_;
  assign new_n6255_ = new_n1200_ & new_n2386_;
  assign new_n6256_ = ~pstart_0_ & new_n6255_;
  assign new_n6257_ = ~new_n1200_ & new_n2383_;
  assign new_n6258_ = ~pstart_0_ & new_n6257_;
  assign new_n6259_ = pencrypt_0_ & pkey_42_;
  assign new_n6260_ = pstart_0_ & new_n6259_;
  assign new_n6261_ = new_n1200_ & new_n2379_;
  assign new_n6262_ = ~pstart_0_ & new_n6261_;
  assign new_n6263_ = pkey_50_ & ~pencrypt_0_;
  assign new_n6264_ = pstart_0_ & new_n6263_;
  assign new_n6265_ = n_n2451 & new_n1220_;
  assign new_n6266_ = pencrypt_0_ & new_n6265_;
  assign new_n6267_ = ~n_n2843 & new_n6266_;
  assign new_n6268_ = ~pstart_0_ & new_n6267_;
  assign new_n6269_ = ~n_n2451 & new_n1220_;
  assign new_n6270_ = pencrypt_0_ & new_n6269_;
  assign new_n6271_ = n_n2843 & new_n6270_;
  assign new_n6272_ = ~pstart_0_ & new_n6271_;
  assign new_n6273_ = ~new_n1200_ & new_n2400_;
  assign new_n6274_ = ~pstart_0_ & new_n6273_;
  assign new_n6275_ = n_n2451 & ~new_n1220_;
  assign new_n6276_ = pencrypt_0_ & new_n6275_;
  assign new_n6277_ = n_n2843 & new_n6276_;
  assign new_n6278_ = ~pstart_0_ & new_n6277_;
  assign new_n6279_ = ~new_n6274_ & ~new_n6278_;
  assign new_n6280_ = ~new_n6268_ & ~new_n6272_;
  assign new_n6281_ = new_n6279_ & new_n6280_;
  assign new_n6282_ = ~new_n6262_ & ~new_n6264_;
  assign new_n6283_ = ~new_n6256_ & ~new_n6258_;
  assign new_n6284_ = ~new_n6260_ & new_n6283_;
  assign new_n6285_ = new_n6282_ & new_n6284_;
  assign n1607 = ~new_n6281_ | ~new_n6285_;
  assign new_n6287_ = new_n1200_ & new_n3930_;
  assign new_n6288_ = ~pstart_0_ & new_n6287_;
  assign new_n6289_ = ~new_n1200_ & new_n3925_;
  assign new_n6290_ = ~pstart_0_ & new_n6289_;
  assign new_n6291_ = pkey_144_ & pencrypt_0_;
  assign new_n6292_ = pstart_0_ & new_n6291_;
  assign new_n6293_ = new_n1200_ & new_n3921_;
  assign new_n6294_ = ~pstart_0_ & new_n6293_;
  assign new_n6295_ = pkey_152_ & ~pencrypt_0_;
  assign new_n6296_ = pstart_0_ & new_n6295_;
  assign new_n6297_ = n_n2414 & new_n1220_;
  assign new_n6298_ = pencrypt_0_ & new_n6297_;
  assign new_n6299_ = ~n_n2320 & new_n6298_;
  assign new_n6300_ = ~pstart_0_ & new_n6299_;
  assign new_n6301_ = ~n_n2414 & new_n1220_;
  assign new_n6302_ = pencrypt_0_ & new_n6301_;
  assign new_n6303_ = n_n2320 & new_n6302_;
  assign new_n6304_ = ~pstart_0_ & new_n6303_;
  assign new_n6305_ = ~new_n1200_ & new_n3944_;
  assign new_n6306_ = ~pstart_0_ & new_n6305_;
  assign new_n6307_ = n_n2414 & ~new_n1220_;
  assign new_n6308_ = pencrypt_0_ & new_n6307_;
  assign new_n6309_ = n_n2320 & new_n6308_;
  assign new_n6310_ = ~pstart_0_ & new_n6309_;
  assign new_n6311_ = ~new_n6306_ & ~new_n6310_;
  assign new_n6312_ = ~new_n6300_ & ~new_n6304_;
  assign new_n6313_ = new_n6311_ & new_n6312_;
  assign new_n6314_ = ~new_n6294_ & ~new_n6296_;
  assign new_n6315_ = ~new_n6288_ & ~new_n6290_;
  assign new_n6316_ = ~new_n6292_ & new_n6315_;
  assign new_n6317_ = new_n6314_ & new_n6316_;
  assign n1612 = ~new_n6313_ | ~new_n6317_;
  assign new_n6319_ = new_n1200_ & new_n3968_;
  assign new_n6320_ = ~pstart_0_ & new_n6319_;
  assign new_n6321_ = ~new_n1200_ & new_n3963_;
  assign new_n6322_ = ~pstart_0_ & new_n6321_;
  assign new_n6323_ = pkey_123_ & pencrypt_0_;
  assign new_n6324_ = pstart_0_ & new_n6323_;
  assign new_n6325_ = new_n1200_ & new_n3959_;
  assign new_n6326_ = ~pstart_0_ & new_n6325_;
  assign new_n6327_ = pkey_66_ & ~pencrypt_0_;
  assign new_n6328_ = pstart_0_ & new_n6327_;
  assign new_n6329_ = n_n2422 & new_n1220_;
  assign new_n6330_ = pencrypt_0_ & new_n6329_;
  assign new_n6331_ = ~n_n2328 & new_n6330_;
  assign new_n6332_ = ~pstart_0_ & new_n6331_;
  assign new_n6333_ = ~n_n2422 & new_n1220_;
  assign new_n6334_ = pencrypt_0_ & new_n6333_;
  assign new_n6335_ = n_n2328 & new_n6334_;
  assign new_n6336_ = ~pstart_0_ & new_n6335_;
  assign new_n6337_ = ~new_n1200_ & new_n3982_;
  assign new_n6338_ = ~pstart_0_ & new_n6337_;
  assign new_n6339_ = n_n2422 & ~new_n1220_;
  assign new_n6340_ = pencrypt_0_ & new_n6339_;
  assign new_n6341_ = n_n2328 & new_n6340_;
  assign new_n6342_ = ~pstart_0_ & new_n6341_;
  assign new_n6343_ = ~new_n6338_ & ~new_n6342_;
  assign new_n6344_ = ~new_n6332_ & ~new_n6336_;
  assign new_n6345_ = new_n6343_ & new_n6344_;
  assign new_n6346_ = ~new_n6326_ & ~new_n6328_;
  assign new_n6347_ = ~new_n6320_ & ~new_n6322_;
  assign new_n6348_ = ~new_n6324_ & new_n6347_;
  assign new_n6349_ = new_n6346_ & new_n6348_;
  assign n1617 = ~new_n6345_ | ~new_n6349_;
  assign new_n6351_ = new_n1200_ & new_n4006_;
  assign new_n6352_ = ~pstart_0_ & new_n6351_;
  assign new_n6353_ = ~new_n1200_ & new_n4001_;
  assign new_n6354_ = ~pstart_0_ & new_n6353_;
  assign new_n6355_ = pkey_97_ & pencrypt_0_;
  assign new_n6356_ = pstart_0_ & new_n6355_;
  assign new_n6357_ = new_n1200_ & new_n3997_;
  assign new_n6358_ = ~pstart_0_ & new_n6357_;
  assign new_n6359_ = ~pencrypt_0_ & pkey_105_;
  assign new_n6360_ = pstart_0_ & new_n6359_;
  assign new_n6361_ = n_n2433 & new_n1220_;
  assign new_n6362_ = pencrypt_0_ & new_n6361_;
  assign new_n6363_ = ~n_n2339 & new_n6362_;
  assign new_n6364_ = ~pstart_0_ & new_n6363_;
  assign new_n6365_ = ~n_n2433 & new_n1220_;
  assign new_n6366_ = pencrypt_0_ & new_n6365_;
  assign new_n6367_ = n_n2339 & new_n6366_;
  assign new_n6368_ = ~pstart_0_ & new_n6367_;
  assign new_n6369_ = ~new_n1200_ & new_n4020_;
  assign new_n6370_ = ~pstart_0_ & new_n6369_;
  assign new_n6371_ = n_n2433 & ~new_n1220_;
  assign new_n6372_ = pencrypt_0_ & new_n6371_;
  assign new_n6373_ = n_n2339 & new_n6372_;
  assign new_n6374_ = ~pstart_0_ & new_n6373_;
  assign new_n6375_ = ~new_n6370_ & ~new_n6374_;
  assign new_n6376_ = ~new_n6364_ & ~new_n6368_;
  assign new_n6377_ = new_n6375_ & new_n6376_;
  assign new_n6378_ = ~new_n6358_ & ~new_n6360_;
  assign new_n6379_ = ~new_n6352_ & ~new_n6354_;
  assign new_n6380_ = ~new_n6356_ & new_n6379_;
  assign new_n6381_ = new_n6378_ & new_n6380_;
  assign n1622 = ~new_n6377_ | ~new_n6381_;
  assign new_n6383_ = new_n1200_ & new_n4044_;
  assign new_n6384_ = ~pstart_0_ & new_n6383_;
  assign new_n6385_ = ~new_n1200_ & new_n4039_;
  assign new_n6386_ = ~pstart_0_ & new_n6385_;
  assign new_n6387_ = pkey_104_ & pencrypt_0_;
  assign new_n6388_ = pstart_0_ & new_n6387_;
  assign new_n6389_ = new_n1200_ & new_n4035_;
  assign new_n6390_ = ~pstart_0_ & new_n6389_;
  assign new_n6391_ = pkey_112_ & ~pencrypt_0_;
  assign new_n6392_ = pstart_0_ & new_n6391_;
  assign new_n6393_ = n_n2440 & new_n1220_;
  assign new_n6394_ = pencrypt_0_ & new_n6393_;
  assign new_n6395_ = ~n_n2347 & new_n6394_;
  assign new_n6396_ = ~pstart_0_ & new_n6395_;
  assign new_n6397_ = ~n_n2440 & new_n1220_;
  assign new_n6398_ = pencrypt_0_ & new_n6397_;
  assign new_n6399_ = n_n2347 & new_n6398_;
  assign new_n6400_ = ~pstart_0_ & new_n6399_;
  assign new_n6401_ = ~new_n1200_ & new_n4058_;
  assign new_n6402_ = ~pstart_0_ & new_n6401_;
  assign new_n6403_ = n_n2440 & ~new_n1220_;
  assign new_n6404_ = pencrypt_0_ & new_n6403_;
  assign new_n6405_ = n_n2347 & new_n6404_;
  assign new_n6406_ = ~pstart_0_ & new_n6405_;
  assign new_n6407_ = ~new_n6402_ & ~new_n6406_;
  assign new_n6408_ = ~new_n6396_ & ~new_n6400_;
  assign new_n6409_ = new_n6407_ & new_n6408_;
  assign new_n6410_ = ~new_n6390_ & ~new_n6392_;
  assign new_n6411_ = ~new_n6384_ & ~new_n6386_;
  assign new_n6412_ = ~new_n6388_ & new_n6411_;
  assign new_n6413_ = new_n6410_ & new_n6412_;
  assign n1627 = ~new_n6409_ | ~new_n6413_;
  assign new_n6415_ = new_n1200_ & new_n4930_;
  assign new_n6416_ = ~pstart_0_ & new_n6415_;
  assign new_n6417_ = ~new_n1200_ & new_n4925_;
  assign new_n6418_ = ~pstart_0_ & new_n6417_;
  assign new_n6419_ = pkey_50_ & pencrypt_0_;
  assign new_n6420_ = pstart_0_ & new_n6419_;
  assign new_n6421_ = new_n1200_ & new_n4921_;
  assign new_n6422_ = ~pstart_0_ & new_n6421_;
  assign new_n6423_ = pkey_58_ & ~pencrypt_0_;
  assign new_n6424_ = pstart_0_ & new_n6423_;
  assign new_n6425_ = n_n2452 & new_n1220_;
  assign new_n6426_ = pencrypt_0_ & new_n6425_;
  assign new_n6427_ = ~n_n2357 & new_n6426_;
  assign new_n6428_ = ~pstart_0_ & new_n6427_;
  assign new_n6429_ = ~n_n2452 & new_n1220_;
  assign new_n6430_ = pencrypt_0_ & new_n6429_;
  assign new_n6431_ = n_n2357 & new_n6430_;
  assign new_n6432_ = ~pstart_0_ & new_n6431_;
  assign new_n6433_ = ~new_n1200_ & new_n4944_;
  assign new_n6434_ = ~pstart_0_ & new_n6433_;
  assign new_n6435_ = n_n2452 & ~new_n1220_;
  assign new_n6436_ = pencrypt_0_ & new_n6435_;
  assign new_n6437_ = n_n2357 & new_n6436_;
  assign new_n6438_ = ~pstart_0_ & new_n6437_;
  assign new_n6439_ = ~new_n6434_ & ~new_n6438_;
  assign new_n6440_ = ~new_n6428_ & ~new_n6432_;
  assign new_n6441_ = new_n6439_ & new_n6440_;
  assign new_n6442_ = ~new_n6422_ & ~new_n6424_;
  assign new_n6443_ = ~new_n6416_ & ~new_n6418_;
  assign new_n6444_ = ~new_n6420_ & new_n6443_;
  assign new_n6445_ = new_n6442_ & new_n6444_;
  assign n1632 = ~new_n6441_ | ~new_n6445_;
  assign new_n6447_ = new_n1200_ & new_n5578_;
  assign new_n6448_ = ~pstart_0_ & new_n6447_;
  assign new_n6449_ = ~new_n1200_ & new_n5573_;
  assign new_n6450_ = ~pstart_0_ & new_n6449_;
  assign new_n6451_ = pkey_152_ & pencrypt_0_;
  assign new_n6452_ = pstart_0_ & new_n6451_;
  assign new_n6453_ = new_n1200_ & new_n5569_;
  assign new_n6454_ = ~pstart_0_ & new_n6453_;
  assign new_n6455_ = pkey_160_ & ~pencrypt_0_;
  assign new_n6456_ = pstart_0_ & new_n6455_;
  assign new_n6457_ = n_n2415 & new_n1220_;
  assign new_n6458_ = pencrypt_0_ & new_n6457_;
  assign new_n6459_ = ~n_n2321 & new_n6458_;
  assign new_n6460_ = ~pstart_0_ & new_n6459_;
  assign new_n6461_ = ~n_n2415 & new_n1220_;
  assign new_n6462_ = pencrypt_0_ & new_n6461_;
  assign new_n6463_ = n_n2321 & new_n6462_;
  assign new_n6464_ = ~pstart_0_ & new_n6463_;
  assign new_n6465_ = ~new_n1200_ & new_n5592_;
  assign new_n6466_ = ~pstart_0_ & new_n6465_;
  assign new_n6467_ = n_n2415 & ~new_n1220_;
  assign new_n6468_ = pencrypt_0_ & new_n6467_;
  assign new_n6469_ = n_n2321 & new_n6468_;
  assign new_n6470_ = ~pstart_0_ & new_n6469_;
  assign new_n6471_ = ~new_n6466_ & ~new_n6470_;
  assign new_n6472_ = ~new_n6460_ & ~new_n6464_;
  assign new_n6473_ = new_n6471_ & new_n6472_;
  assign new_n6474_ = ~new_n6454_ & ~new_n6456_;
  assign new_n6475_ = ~new_n6448_ & ~new_n6450_;
  assign new_n6476_ = ~new_n6452_ & new_n6475_;
  assign new_n6477_ = new_n6474_ & new_n6476_;
  assign n1637 = ~new_n6473_ | ~new_n6477_;
  assign new_n6479_ = new_n1200_ & new_n5616_;
  assign new_n6480_ = ~pstart_0_ & new_n6479_;
  assign new_n6481_ = ~new_n1200_ & new_n5611_;
  assign new_n6482_ = ~pstart_0_ & new_n6481_;
  assign new_n6483_ = pencrypt_0_ & pkey_82_;
  assign new_n6484_ = pstart_0_ & new_n6483_;
  assign new_n6485_ = new_n1200_ & new_n5607_;
  assign new_n6486_ = ~pstart_0_ & new_n6485_;
  assign new_n6487_ = ~pencrypt_0_ & pkey_90_;
  assign new_n6488_ = pstart_0_ & new_n6487_;
  assign new_n6489_ = n_n2425 & new_n1220_;
  assign new_n6490_ = pencrypt_0_ & new_n6489_;
  assign new_n6491_ = ~n_n2330 & new_n6490_;
  assign new_n6492_ = ~pstart_0_ & new_n6491_;
  assign new_n6493_ = ~n_n2425 & new_n1220_;
  assign new_n6494_ = pencrypt_0_ & new_n6493_;
  assign new_n6495_ = n_n2330 & new_n6494_;
  assign new_n6496_ = ~pstart_0_ & new_n6495_;
  assign new_n6497_ = ~new_n1200_ & new_n5630_;
  assign new_n6498_ = ~pstart_0_ & new_n6497_;
  assign new_n6499_ = n_n2425 & ~new_n1220_;
  assign new_n6500_ = pencrypt_0_ & new_n6499_;
  assign new_n6501_ = n_n2330 & new_n6500_;
  assign new_n6502_ = ~pstart_0_ & new_n6501_;
  assign new_n6503_ = ~new_n6498_ & ~new_n6502_;
  assign new_n6504_ = ~new_n6492_ & ~new_n6496_;
  assign new_n6505_ = new_n6503_ & new_n6504_;
  assign new_n6506_ = ~new_n6486_ & ~new_n6488_;
  assign new_n6507_ = ~new_n6480_ & ~new_n6482_;
  assign new_n6508_ = ~new_n6484_ & new_n6507_;
  assign new_n6509_ = new_n6506_ & new_n6508_;
  assign n1642 = ~new_n6505_ | ~new_n6509_;
  assign new_n6511_ = new_n1200_ & new_n5654_;
  assign new_n6512_ = ~pstart_0_ & new_n6511_;
  assign new_n6513_ = ~new_n1200_ & new_n5649_;
  assign new_n6514_ = ~pstart_0_ & new_n6513_;
  assign new_n6515_ = pencrypt_0_ & pkey_73_;
  assign new_n6516_ = pstart_0_ & new_n6515_;
  assign new_n6517_ = new_n1200_ & new_n5645_;
  assign new_n6518_ = ~pstart_0_ & new_n6517_;
  assign new_n6519_ = pkey_81_ & ~pencrypt_0_;
  assign new_n6520_ = pstart_0_ & new_n6519_;
  assign new_n6521_ = n_n2945 & new_n1220_;
  assign new_n6522_ = pencrypt_0_ & new_n6521_;
  assign new_n6523_ = ~n_n2336 & new_n6522_;
  assign new_n6524_ = ~pstart_0_ & new_n6523_;
  assign new_n6525_ = ~n_n2945 & new_n1220_;
  assign new_n6526_ = pencrypt_0_ & new_n6525_;
  assign new_n6527_ = n_n2336 & new_n6526_;
  assign new_n6528_ = ~pstart_0_ & new_n6527_;
  assign new_n6529_ = ~new_n1200_ & new_n5668_;
  assign new_n6530_ = ~pstart_0_ & new_n6529_;
  assign new_n6531_ = n_n2945 & ~new_n1220_;
  assign new_n6532_ = pencrypt_0_ & new_n6531_;
  assign new_n6533_ = n_n2336 & new_n6532_;
  assign new_n6534_ = ~pstart_0_ & new_n6533_;
  assign new_n6535_ = ~new_n6530_ & ~new_n6534_;
  assign new_n6536_ = ~new_n6524_ & ~new_n6528_;
  assign new_n6537_ = new_n6535_ & new_n6536_;
  assign new_n6538_ = ~new_n6518_ & ~new_n6520_;
  assign new_n6539_ = ~new_n6512_ & ~new_n6514_;
  assign new_n6540_ = ~new_n6516_ & new_n6539_;
  assign new_n6541_ = new_n6538_ & new_n6540_;
  assign n1647 = ~new_n6537_ | ~new_n6541_;
  assign new_n6543_ = new_n1200_ & new_n5692_;
  assign new_n6544_ = ~pstart_0_ & new_n6543_;
  assign new_n6545_ = ~new_n1200_ & new_n5687_;
  assign new_n6546_ = ~pstart_0_ & new_n6545_;
  assign new_n6547_ = pkey_96_ & pencrypt_0_;
  assign new_n6548_ = pstart_0_ & new_n6547_;
  assign new_n6549_ = new_n1200_ & new_n5683_;
  assign new_n6550_ = ~pstart_0_ & new_n6549_;
  assign new_n6551_ = pkey_104_ & ~pencrypt_0_;
  assign new_n6552_ = pstart_0_ & new_n6551_;
  assign new_n6553_ = n_n2439 & new_n1220_;
  assign new_n6554_ = pencrypt_0_ & new_n6553_;
  assign new_n6555_ = ~n_n2346 & new_n6554_;
  assign new_n6556_ = ~pstart_0_ & new_n6555_;
  assign new_n6557_ = ~n_n2439 & new_n1220_;
  assign new_n6558_ = pencrypt_0_ & new_n6557_;
  assign new_n6559_ = n_n2346 & new_n6558_;
  assign new_n6560_ = ~pstart_0_ & new_n6559_;
  assign new_n6561_ = ~new_n1200_ & new_n5706_;
  assign new_n6562_ = ~pstart_0_ & new_n6561_;
  assign new_n6563_ = n_n2439 & ~new_n1220_;
  assign new_n6564_ = pencrypt_0_ & new_n6563_;
  assign new_n6565_ = n_n2346 & new_n6564_;
  assign new_n6566_ = ~pstart_0_ & new_n6565_;
  assign new_n6567_ = ~new_n6562_ & ~new_n6566_;
  assign new_n6568_ = ~new_n6556_ & ~new_n6560_;
  assign new_n6569_ = new_n6567_ & new_n6568_;
  assign new_n6570_ = ~new_n6550_ & ~new_n6552_;
  assign new_n6571_ = ~new_n6544_ & ~new_n6546_;
  assign new_n6572_ = ~new_n6548_ & new_n6571_;
  assign new_n6573_ = new_n6570_ & new_n6572_;
  assign n1652 = ~new_n6569_ | ~new_n6573_;
  assign new_n6575_ = new_n1200_ & new_n5324_;
  assign new_n6576_ = ~pstart_0_ & new_n6575_;
  assign new_n6577_ = ~new_n1200_ & new_n5319_;
  assign new_n6578_ = ~pstart_0_ & new_n6577_;
  assign new_n6579_ = pkey_58_ & pencrypt_0_;
  assign new_n6580_ = pstart_0_ & new_n6579_;
  assign new_n6581_ = new_n1200_ & new_n5315_;
  assign new_n6582_ = ~pstart_0_ & new_n6581_;
  assign new_n6583_ = pkey_1_ & ~pencrypt_0_;
  assign new_n6584_ = pstart_0_ & new_n6583_;
  assign new_n6585_ = n_n2453 & new_n1220_;
  assign new_n6586_ = pencrypt_0_ & new_n6585_;
  assign new_n6587_ = ~n_n2358 & new_n6586_;
  assign new_n6588_ = ~pstart_0_ & new_n6587_;
  assign new_n6589_ = ~n_n2453 & new_n1220_;
  assign new_n6590_ = pencrypt_0_ & new_n6589_;
  assign new_n6591_ = n_n2358 & new_n6590_;
  assign new_n6592_ = ~pstart_0_ & new_n6591_;
  assign new_n6593_ = ~new_n1200_ & new_n5338_;
  assign new_n6594_ = ~pstart_0_ & new_n6593_;
  assign new_n6595_ = n_n2453 & ~new_n1220_;
  assign new_n6596_ = pencrypt_0_ & new_n6595_;
  assign new_n6597_ = n_n2358 & new_n6596_;
  assign new_n6598_ = ~pstart_0_ & new_n6597_;
  assign new_n6599_ = ~new_n6594_ & ~new_n6598_;
  assign new_n6600_ = ~new_n6588_ & ~new_n6592_;
  assign new_n6601_ = new_n6599_ & new_n6600_;
  assign new_n6602_ = ~new_n6582_ & ~new_n6584_;
  assign new_n6603_ = ~new_n6576_ & ~new_n6578_;
  assign new_n6604_ = ~new_n6580_ & new_n6603_;
  assign new_n6605_ = new_n6602_ & new_n6604_;
  assign n1657 = ~new_n6601_ | ~new_n6605_;
  assign new_n6607_ = new_n1200_ & new_n3338_;
  assign new_n6608_ = ~pstart_0_ & new_n6607_;
  assign new_n6609_ = ~new_n1200_ & new_n3333_;
  assign new_n6610_ = ~pstart_0_ & new_n6609_;
  assign new_n6611_ = pkey_56_ & pencrypt_0_;
  assign new_n6612_ = pstart_0_ & new_n6611_;
  assign new_n6613_ = new_n1200_ & new_n3329_;
  assign new_n6614_ = ~pstart_0_ & new_n6613_;
  assign new_n6615_ = pkey_227_ & ~pencrypt_0_;
  assign new_n6616_ = pstart_0_ & new_n6615_;
  assign new_n6617_ = n_n2373 & new_n1220_;
  assign new_n6618_ = pencrypt_0_ & new_n6617_;
  assign new_n6619_ = ~n_n2278 & new_n6618_;
  assign new_n6620_ = ~pstart_0_ & new_n6619_;
  assign new_n6621_ = ~n_n2373 & new_n1220_;
  assign new_n6622_ = pencrypt_0_ & new_n6621_;
  assign new_n6623_ = n_n2278 & new_n6622_;
  assign new_n6624_ = ~pstart_0_ & new_n6623_;
  assign new_n6625_ = ~new_n1200_ & new_n3352_;
  assign new_n6626_ = ~pstart_0_ & new_n6625_;
  assign new_n6627_ = n_n2373 & ~new_n1220_;
  assign new_n6628_ = pencrypt_0_ & new_n6627_;
  assign new_n6629_ = n_n2278 & new_n6628_;
  assign new_n6630_ = ~pstart_0_ & new_n6629_;
  assign new_n6631_ = ~new_n6626_ & ~new_n6630_;
  assign new_n6632_ = ~new_n6620_ & ~new_n6624_;
  assign new_n6633_ = new_n6631_ & new_n6632_;
  assign new_n6634_ = ~new_n6614_ & ~new_n6616_;
  assign new_n6635_ = ~new_n6608_ & ~new_n6610_;
  assign new_n6636_ = ~new_n6612_ & new_n6635_;
  assign new_n6637_ = new_n6634_ & new_n6636_;
  assign n1662 = ~new_n6633_ | ~new_n6637_;
  assign new_n6639_ = new_n1200_ & new_n5952_;
  assign new_n6640_ = ~pstart_0_ & new_n6639_;
  assign new_n6641_ = ~new_n1200_ & new_n5947_;
  assign new_n6642_ = ~pstart_0_ & new_n6641_;
  assign new_n6643_ = pkey_160_ & pencrypt_0_;
  assign new_n6644_ = pstart_0_ & new_n6643_;
  assign new_n6645_ = new_n1200_ & new_n5943_;
  assign new_n6646_ = ~pstart_0_ & new_n6645_;
  assign new_n6647_ = pkey_168_ & ~pencrypt_0_;
  assign new_n6648_ = pstart_0_ & new_n6647_;
  assign new_n6649_ = n_n2416 & new_n1220_;
  assign new_n6650_ = pencrypt_0_ & new_n6649_;
  assign new_n6651_ = ~n_n2322 & new_n6650_;
  assign new_n6652_ = ~pstart_0_ & new_n6651_;
  assign new_n6653_ = ~n_n2416 & new_n1220_;
  assign new_n6654_ = pencrypt_0_ & new_n6653_;
  assign new_n6655_ = n_n2322 & new_n6654_;
  assign new_n6656_ = ~pstart_0_ & new_n6655_;
  assign new_n6657_ = ~new_n1200_ & new_n5966_;
  assign new_n6658_ = ~pstart_0_ & new_n6657_;
  assign new_n6659_ = n_n2416 & ~new_n1220_;
  assign new_n6660_ = pencrypt_0_ & new_n6659_;
  assign new_n6661_ = n_n2322 & new_n6660_;
  assign new_n6662_ = ~pstart_0_ & new_n6661_;
  assign new_n6663_ = ~new_n6658_ & ~new_n6662_;
  assign new_n6664_ = ~new_n6652_ & ~new_n6656_;
  assign new_n6665_ = new_n6663_ & new_n6664_;
  assign new_n6666_ = ~new_n6646_ & ~new_n6648_;
  assign new_n6667_ = ~new_n6640_ & ~new_n6642_;
  assign new_n6668_ = ~new_n6644_ & new_n6667_;
  assign new_n6669_ = new_n6666_ & new_n6668_;
  assign n1667 = ~new_n6665_ | ~new_n6669_;
  assign new_n6671_ = new_n1200_ & new_n5990_;
  assign new_n6672_ = ~pstart_0_ & new_n6671_;
  assign new_n6673_ = ~new_n1200_ & new_n5985_;
  assign new_n6674_ = ~pstart_0_ & new_n6673_;
  assign new_n6675_ = pkey_74_ & pencrypt_0_;
  assign new_n6676_ = pstart_0_ & new_n6675_;
  assign new_n6677_ = new_n1200_ & new_n5981_;
  assign new_n6678_ = ~pstart_0_ & new_n6677_;
  assign new_n6679_ = ~pencrypt_0_ & pkey_82_;
  assign new_n6680_ = pstart_0_ & new_n6679_;
  assign new_n6681_ = n_n2424 & new_n1220_;
  assign new_n6682_ = pencrypt_0_ & new_n6681_;
  assign new_n6683_ = ~n_n2806 & new_n6682_;
  assign new_n6684_ = ~pstart_0_ & new_n6683_;
  assign new_n6685_ = ~n_n2424 & new_n1220_;
  assign new_n6686_ = pencrypt_0_ & new_n6685_;
  assign new_n6687_ = n_n2806 & new_n6686_;
  assign new_n6688_ = ~pstart_0_ & new_n6687_;
  assign new_n6689_ = ~new_n1200_ & new_n6004_;
  assign new_n6690_ = ~pstart_0_ & new_n6689_;
  assign new_n6691_ = n_n2424 & ~new_n1220_;
  assign new_n6692_ = pencrypt_0_ & new_n6691_;
  assign new_n6693_ = n_n2806 & new_n6692_;
  assign new_n6694_ = ~pstart_0_ & new_n6693_;
  assign new_n6695_ = ~new_n6690_ & ~new_n6694_;
  assign new_n6696_ = ~new_n6684_ & ~new_n6688_;
  assign new_n6697_ = new_n6695_ & new_n6696_;
  assign new_n6698_ = ~new_n6678_ & ~new_n6680_;
  assign new_n6699_ = ~new_n6672_ & ~new_n6674_;
  assign new_n6700_ = ~new_n6676_ & new_n6699_;
  assign new_n6701_ = new_n6698_ & new_n6700_;
  assign n1672 = ~new_n6697_ | ~new_n6701_;
  assign new_n6703_ = new_n1200_ & new_n6028_;
  assign new_n6704_ = ~pstart_0_ & new_n6703_;
  assign new_n6705_ = ~new_n1200_ & new_n6023_;
  assign new_n6706_ = ~pstart_0_ & new_n6705_;
  assign new_n6707_ = pkey_81_ & pencrypt_0_;
  assign new_n6708_ = pstart_0_ & new_n6707_;
  assign new_n6709_ = new_n1200_ & new_n6019_;
  assign new_n6710_ = ~pstart_0_ & new_n6709_;
  assign new_n6711_ = pkey_89_ & ~pencrypt_0_;
  assign new_n6712_ = pstart_0_ & new_n6711_;
  assign new_n6713_ = n_n2431 & new_n1220_;
  assign new_n6714_ = pencrypt_0_ & new_n6713_;
  assign new_n6715_ = ~n_n2337 & new_n6714_;
  assign new_n6716_ = ~pstart_0_ & new_n6715_;
  assign new_n6717_ = ~n_n2431 & new_n1220_;
  assign new_n6718_ = pencrypt_0_ & new_n6717_;
  assign new_n6719_ = n_n2337 & new_n6718_;
  assign new_n6720_ = ~pstart_0_ & new_n6719_;
  assign new_n6721_ = ~new_n1200_ & new_n6042_;
  assign new_n6722_ = ~pstart_0_ & new_n6721_;
  assign new_n6723_ = n_n2431 & ~new_n1220_;
  assign new_n6724_ = pencrypt_0_ & new_n6723_;
  assign new_n6725_ = n_n2337 & new_n6724_;
  assign new_n6726_ = ~pstart_0_ & new_n6725_;
  assign new_n6727_ = ~new_n6722_ & ~new_n6726_;
  assign new_n6728_ = ~new_n6716_ & ~new_n6720_;
  assign new_n6729_ = new_n6727_ & new_n6728_;
  assign new_n6730_ = ~new_n6710_ & ~new_n6712_;
  assign new_n6731_ = ~new_n6704_ & ~new_n6706_;
  assign new_n6732_ = ~new_n6708_ & new_n6731_;
  assign new_n6733_ = new_n6730_ & new_n6732_;
  assign n1677 = ~new_n6729_ | ~new_n6733_;
  assign new_n6735_ = new_n1200_ & new_n6066_;
  assign new_n6736_ = ~pstart_0_ & new_n6735_;
  assign new_n6737_ = ~new_n1200_ & new_n6061_;
  assign new_n6738_ = ~pstart_0_ & new_n6737_;
  assign new_n6739_ = pkey_88_ & pencrypt_0_;
  assign new_n6740_ = pstart_0_ & new_n6739_;
  assign new_n6741_ = new_n1200_ & new_n6057_;
  assign new_n6742_ = ~pstart_0_ & new_n6741_;
  assign new_n6743_ = pkey_96_ & ~pencrypt_0_;
  assign new_n6744_ = pstart_0_ & new_n6743_;
  assign new_n6745_ = n_n2438 & new_n1220_;
  assign new_n6746_ = pencrypt_0_ & new_n6745_;
  assign new_n6747_ = ~n_n2345 & new_n6746_;
  assign new_n6748_ = ~pstart_0_ & new_n6747_;
  assign new_n6749_ = ~n_n2438 & new_n1220_;
  assign new_n6750_ = pencrypt_0_ & new_n6749_;
  assign new_n6751_ = n_n2345 & new_n6750_;
  assign new_n6752_ = ~pstart_0_ & new_n6751_;
  assign new_n6753_ = ~new_n1200_ & new_n6080_;
  assign new_n6754_ = ~pstart_0_ & new_n6753_;
  assign new_n6755_ = n_n2438 & ~new_n1220_;
  assign new_n6756_ = pencrypt_0_ & new_n6755_;
  assign new_n6757_ = n_n2345 & new_n6756_;
  assign new_n6758_ = ~pstart_0_ & new_n6757_;
  assign new_n6759_ = ~new_n6754_ & ~new_n6758_;
  assign new_n6760_ = ~new_n6748_ & ~new_n6752_;
  assign new_n6761_ = new_n6759_ & new_n6760_;
  assign new_n6762_ = ~new_n6742_ & ~new_n6744_;
  assign new_n6763_ = ~new_n6736_ & ~new_n6738_;
  assign new_n6764_ = ~new_n6740_ & new_n6763_;
  assign new_n6765_ = new_n6762_ & new_n6764_;
  assign n1682 = ~new_n6761_ | ~new_n6765_;
  assign new_n6767_ = new_n1200_ & new_n5730_;
  assign new_n6768_ = ~pstart_0_ & new_n6767_;
  assign new_n6769_ = ~new_n1200_ & new_n5725_;
  assign new_n6770_ = ~pstart_0_ & new_n6769_;
  assign new_n6771_ = pkey_1_ & pencrypt_0_;
  assign new_n6772_ = pstart_0_ & new_n6771_;
  assign new_n6773_ = new_n1200_ & new_n5721_;
  assign new_n6774_ = ~pstart_0_ & new_n6773_;
  assign new_n6775_ = pkey_9_ & ~pencrypt_0_;
  assign new_n6776_ = pstart_0_ & new_n6775_;
  assign new_n6777_ = n_n2976 & new_n1220_;
  assign new_n6778_ = pencrypt_0_ & new_n6777_;
  assign new_n6779_ = ~n_n2359 & new_n6778_;
  assign new_n6780_ = ~pstart_0_ & new_n6779_;
  assign new_n6781_ = ~n_n2976 & new_n1220_;
  assign new_n6782_ = pencrypt_0_ & new_n6781_;
  assign new_n6783_ = n_n2359 & new_n6782_;
  assign new_n6784_ = ~pstart_0_ & new_n6783_;
  assign new_n6785_ = ~new_n1200_ & new_n5744_;
  assign new_n6786_ = ~pstart_0_ & new_n6785_;
  assign new_n6787_ = n_n2976 & ~new_n1220_;
  assign new_n6788_ = pencrypt_0_ & new_n6787_;
  assign new_n6789_ = n_n2359 & new_n6788_;
  assign new_n6790_ = ~pstart_0_ & new_n6789_;
  assign new_n6791_ = ~new_n6786_ & ~new_n6790_;
  assign new_n6792_ = ~new_n6780_ & ~new_n6784_;
  assign new_n6793_ = new_n6791_ & new_n6792_;
  assign new_n6794_ = ~new_n6774_ & ~new_n6776_;
  assign new_n6795_ = ~new_n6768_ & ~new_n6770_;
  assign new_n6796_ = ~new_n6772_ & new_n6795_;
  assign new_n6797_ = new_n6794_ & new_n6796_;
  assign n1687 = ~new_n6793_ | ~new_n6797_;
  assign new_n6799_ = new_n1200_ & new_n2570_;
  assign new_n6800_ = ~pstart_0_ & new_n6799_;
  assign new_n6801_ = ~new_n1200_ & new_n2565_;
  assign new_n6802_ = ~pstart_0_ & new_n6801_;
  assign new_n6803_ = pkey_234_ & pencrypt_0_;
  assign new_n6804_ = pstart_0_ & new_n6803_;
  assign new_n6805_ = new_n1200_ & new_n2561_;
  assign new_n6806_ = ~pstart_0_ & new_n6805_;
  assign new_n6807_ = pkey_242_ & ~pencrypt_0_;
  assign new_n6808_ = pstart_0_ & new_n6807_;
  assign new_n6809_ = n_n2382 & new_n1220_;
  assign new_n6810_ = pencrypt_0_ & new_n6809_;
  assign new_n6811_ = ~n_n2746 & new_n6810_;
  assign new_n6812_ = ~pstart_0_ & new_n6811_;
  assign new_n6813_ = ~n_n2382 & new_n1220_;
  assign new_n6814_ = pencrypt_0_ & new_n6813_;
  assign new_n6815_ = n_n2746 & new_n6814_;
  assign new_n6816_ = ~pstart_0_ & new_n6815_;
  assign new_n6817_ = ~new_n1200_ & new_n2584_;
  assign new_n6818_ = ~pstart_0_ & new_n6817_;
  assign new_n6819_ = n_n2382 & ~new_n1220_;
  assign new_n6820_ = pencrypt_0_ & new_n6819_;
  assign new_n6821_ = n_n2746 & new_n6820_;
  assign new_n6822_ = ~pstart_0_ & new_n6821_;
  assign new_n6823_ = ~new_n6818_ & ~new_n6822_;
  assign new_n6824_ = ~new_n6812_ & ~new_n6816_;
  assign new_n6825_ = new_n6823_ & new_n6824_;
  assign new_n6826_ = ~new_n6806_ & ~new_n6808_;
  assign new_n6827_ = ~new_n6800_ & ~new_n6802_;
  assign new_n6828_ = ~new_n6804_ & new_n6827_;
  assign new_n6829_ = new_n6826_ & new_n6828_;
  assign n1692 = ~new_n6825_ | ~new_n6829_;
  assign new_n6831_ = new_n1200_ & new_n2608_;
  assign new_n6832_ = ~pstart_0_ & new_n6831_;
  assign new_n6833_ = ~new_n1200_ & new_n2603_;
  assign new_n6834_ = ~pstart_0_ & new_n6833_;
  assign new_n6835_ = pencrypt_0_ & pkey_192_;
  assign new_n6836_ = pstart_0_ & new_n6835_;
  assign new_n6837_ = new_n1200_ & new_n2599_;
  assign new_n6838_ = ~pstart_0_ & new_n6837_;
  assign new_n6839_ = ~pencrypt_0_ & pkey_200_;
  assign new_n6840_ = pstart_0_ & new_n6839_;
  assign new_n6841_ = n_n2889 & new_n1220_;
  assign new_n6842_ = pencrypt_0_ & new_n6841_;
  assign new_n6843_ = ~n_n2294 & new_n6842_;
  assign new_n6844_ = ~pstart_0_ & new_n6843_;
  assign new_n6845_ = ~n_n2889 & new_n1220_;
  assign new_n6846_ = pencrypt_0_ & new_n6845_;
  assign new_n6847_ = n_n2294 & new_n6846_;
  assign new_n6848_ = ~pstart_0_ & new_n6847_;
  assign new_n6849_ = ~new_n1200_ & new_n2622_;
  assign new_n6850_ = ~pstart_0_ & new_n6849_;
  assign new_n6851_ = n_n2889 & ~new_n1220_;
  assign new_n6852_ = pencrypt_0_ & new_n6851_;
  assign new_n6853_ = n_n2294 & new_n6852_;
  assign new_n6854_ = ~pstart_0_ & new_n6853_;
  assign new_n6855_ = ~new_n6850_ & ~new_n6854_;
  assign new_n6856_ = ~new_n6844_ & ~new_n6848_;
  assign new_n6857_ = new_n6855_ & new_n6856_;
  assign new_n6858_ = ~new_n6838_ & ~new_n6840_;
  assign new_n6859_ = ~new_n6832_ & ~new_n6834_;
  assign new_n6860_ = ~new_n6836_ & new_n6859_;
  assign new_n6861_ = new_n6858_ & new_n6860_;
  assign n1697 = ~new_n6857_ | ~new_n6861_;
  assign new_n6863_ = new_n1200_ & new_n4704_;
  assign new_n6864_ = ~pstart_0_ & new_n6863_;
  assign new_n6865_ = ~new_n1200_ & new_n4699_;
  assign new_n6866_ = ~pstart_0_ & new_n6865_;
  assign new_n6867_ = pencrypt_0_ & pkey_187_;
  assign new_n6868_ = pstart_0_ & new_n6867_;
  assign new_n6869_ = new_n1200_ & new_n4695_;
  assign new_n6870_ = ~pstart_0_ & new_n6869_;
  assign new_n6871_ = pkey_130_ & ~pencrypt_0_;
  assign new_n6872_ = pstart_0_ & new_n6871_;
  assign new_n6873_ = n_n2398 & new_n1220_;
  assign new_n6874_ = pencrypt_0_ & new_n6873_;
  assign new_n6875_ = ~n_n2304 & new_n6874_;
  assign new_n6876_ = ~pstart_0_ & new_n6875_;
  assign new_n6877_ = ~n_n2398 & new_n1220_;
  assign new_n6878_ = pencrypt_0_ & new_n6877_;
  assign new_n6879_ = n_n2304 & new_n6878_;
  assign new_n6880_ = ~pstart_0_ & new_n6879_;
  assign new_n6881_ = ~new_n1200_ & new_n4718_;
  assign new_n6882_ = ~pstart_0_ & new_n6881_;
  assign new_n6883_ = n_n2398 & ~new_n1220_;
  assign new_n6884_ = pencrypt_0_ & new_n6883_;
  assign new_n6885_ = n_n2304 & new_n6884_;
  assign new_n6886_ = ~pstart_0_ & new_n6885_;
  assign new_n6887_ = ~new_n6882_ & ~new_n6886_;
  assign new_n6888_ = ~new_n6876_ & ~new_n6880_;
  assign new_n6889_ = new_n6887_ & new_n6888_;
  assign new_n6890_ = ~new_n6870_ & ~new_n6872_;
  assign new_n6891_ = ~new_n6864_ & ~new_n6866_;
  assign new_n6892_ = ~new_n6868_ & new_n6891_;
  assign new_n6893_ = new_n6890_ & new_n6892_;
  assign n1702 = ~new_n6889_ | ~new_n6893_;
  assign new_n6895_ = new_n1200_ & new_n4742_;
  assign new_n6896_ = ~pstart_0_ & new_n6895_;
  assign new_n6897_ = ~new_n1200_ & new_n4737_;
  assign new_n6898_ = ~pstart_0_ & new_n6897_;
  assign new_n6899_ = pkey_145_ & pencrypt_0_;
  assign new_n6900_ = pstart_0_ & new_n6899_;
  assign new_n6901_ = new_n1200_ & new_n4733_;
  assign new_n6902_ = ~pstart_0_ & new_n6901_;
  assign new_n6903_ = pkey_153_ & ~pencrypt_0_;
  assign new_n6904_ = pstart_0_ & new_n6903_;
  assign new_n6905_ = n_n2408 & new_n1220_;
  assign new_n6906_ = pencrypt_0_ & new_n6905_;
  assign new_n6907_ = ~n_n2313 & new_n6906_;
  assign new_n6908_ = ~pstart_0_ & new_n6907_;
  assign new_n6909_ = ~n_n2408 & new_n1220_;
  assign new_n6910_ = pencrypt_0_ & new_n6909_;
  assign new_n6911_ = n_n2313 & new_n6910_;
  assign new_n6912_ = ~pstart_0_ & new_n6911_;
  assign new_n6913_ = ~new_n1200_ & new_n4756_;
  assign new_n6914_ = ~pstart_0_ & new_n6913_;
  assign new_n6915_ = n_n2408 & ~new_n1220_;
  assign new_n6916_ = pencrypt_0_ & new_n6915_;
  assign new_n6917_ = n_n2313 & new_n6916_;
  assign new_n6918_ = ~pstart_0_ & new_n6917_;
  assign new_n6919_ = ~new_n6914_ & ~new_n6918_;
  assign new_n6920_ = ~new_n6908_ & ~new_n6912_;
  assign new_n6921_ = new_n6919_ & new_n6920_;
  assign new_n6922_ = ~new_n6902_ & ~new_n6904_;
  assign new_n6923_ = ~new_n6896_ & ~new_n6898_;
  assign new_n6924_ = ~new_n6900_ & new_n6923_;
  assign new_n6925_ = new_n6922_ & new_n6924_;
  assign n1707 = ~new_n6921_ | ~new_n6925_;
  assign new_n6927_ = new_n1200_ & new_n2722_;
  assign new_n6928_ = ~pstart_0_ & new_n6927_;
  assign new_n6929_ = ~new_n1200_ & new_n2717_;
  assign new_n6930_ = ~pstart_0_ & new_n6929_;
  assign new_n6931_ = pkey_9_ & pencrypt_0_;
  assign new_n6932_ = pstart_0_ & new_n6931_;
  assign new_n6933_ = new_n1200_ & new_n2713_;
  assign new_n6934_ = ~pstart_0_ & new_n6933_;
  assign new_n6935_ = pkey_17_ & ~pencrypt_0_;
  assign new_n6936_ = pstart_0_ & new_n6935_;
  assign new_n6937_ = n_n2454 & new_n1220_;
  assign new_n6938_ = pencrypt_0_ & new_n6937_;
  assign new_n6939_ = ~n_n2360 & new_n6938_;
  assign new_n6940_ = ~pstart_0_ & new_n6939_;
  assign new_n6941_ = ~n_n2454 & new_n1220_;
  assign new_n6942_ = pencrypt_0_ & new_n6941_;
  assign new_n6943_ = n_n2360 & new_n6942_;
  assign new_n6944_ = ~pstart_0_ & new_n6943_;
  assign new_n6945_ = ~new_n1200_ & new_n2736_;
  assign new_n6946_ = ~pstart_0_ & new_n6945_;
  assign new_n6947_ = n_n2454 & ~new_n1220_;
  assign new_n6948_ = pencrypt_0_ & new_n6947_;
  assign new_n6949_ = n_n2360 & new_n6948_;
  assign new_n6950_ = ~pstart_0_ & new_n6949_;
  assign new_n6951_ = ~new_n6946_ & ~new_n6950_;
  assign new_n6952_ = ~new_n6940_ & ~new_n6944_;
  assign new_n6953_ = new_n6951_ & new_n6952_;
  assign new_n6954_ = ~new_n6934_ & ~new_n6936_;
  assign new_n6955_ = ~new_n6928_ & ~new_n6930_;
  assign new_n6956_ = ~new_n6932_ & new_n6955_;
  assign new_n6957_ = new_n6954_ & new_n6956_;
  assign n1712 = ~new_n6953_ | ~new_n6957_;
  assign new_n6959_ = new_n1200_ & new_n2868_;
  assign new_n6960_ = ~pstart_0_ & new_n6959_;
  assign new_n6961_ = ~new_n1200_ & new_n2863_;
  assign new_n6962_ = ~pstart_0_ & new_n6961_;
  assign new_n6963_ = pkey_242_ & pencrypt_0_;
  assign new_n6964_ = pstart_0_ & new_n6963_;
  assign new_n6965_ = new_n1200_ & new_n2859_;
  assign new_n6966_ = ~pstart_0_ & new_n6965_;
  assign new_n6967_ = pkey_250_ & ~pencrypt_0_;
  assign new_n6968_ = pstart_0_ & new_n6967_;
  assign new_n6969_ = n_n2383 & new_n1220_;
  assign new_n6970_ = pencrypt_0_ & new_n6969_;
  assign new_n6971_ = ~n_n2286 & new_n6970_;
  assign new_n6972_ = ~pstart_0_ & new_n6971_;
  assign new_n6973_ = ~n_n2383 & new_n1220_;
  assign new_n6974_ = pencrypt_0_ & new_n6973_;
  assign new_n6975_ = n_n2286 & new_n6974_;
  assign new_n6976_ = ~pstart_0_ & new_n6975_;
  assign new_n6977_ = ~new_n1200_ & new_n2882_;
  assign new_n6978_ = ~pstart_0_ & new_n6977_;
  assign new_n6979_ = n_n2383 & ~new_n1220_;
  assign new_n6980_ = pencrypt_0_ & new_n6979_;
  assign new_n6981_ = n_n2286 & new_n6980_;
  assign new_n6982_ = ~pstart_0_ & new_n6981_;
  assign new_n6983_ = ~new_n6978_ & ~new_n6982_;
  assign new_n6984_ = ~new_n6972_ & ~new_n6976_;
  assign new_n6985_ = new_n6983_ & new_n6984_;
  assign new_n6986_ = ~new_n6966_ & ~new_n6968_;
  assign new_n6987_ = ~new_n6960_ & ~new_n6962_;
  assign new_n6988_ = ~new_n6964_ & new_n6987_;
  assign new_n6989_ = new_n6986_ & new_n6988_;
  assign n1717 = ~new_n6985_ | ~new_n6989_;
  assign new_n6991_ = new_n1200_ & new_n2906_;
  assign new_n6992_ = ~pstart_0_ & new_n6991_;
  assign new_n6993_ = ~new_n1200_ & new_n2901_;
  assign new_n6994_ = ~pstart_0_ & new_n6993_;
  assign new_n6995_ = pkey_249_ & pencrypt_0_;
  assign new_n6996_ = pstart_0_ & new_n6995_;
  assign new_n6997_ = new_n1200_ & new_n2897_;
  assign new_n6998_ = ~pstart_0_ & new_n6997_;
  assign new_n6999_ = ~pencrypt_0_ & pkey_192_;
  assign new_n7000_ = pstart_0_ & new_n6999_;
  assign new_n7001_ = n_n2388 & new_n1220_;
  assign new_n7002_ = pencrypt_0_ & new_n7001_;
  assign new_n7003_ = ~n_n2293 & new_n7002_;
  assign new_n7004_ = ~pstart_0_ & new_n7003_;
  assign new_n7005_ = ~n_n2388 & new_n1220_;
  assign new_n7006_ = pencrypt_0_ & new_n7005_;
  assign new_n7007_ = n_n2293 & new_n7006_;
  assign new_n7008_ = ~pstart_0_ & new_n7007_;
  assign new_n7009_ = ~new_n1200_ & new_n2920_;
  assign new_n7010_ = ~pstart_0_ & new_n7009_;
  assign new_n7011_ = n_n2388 & ~new_n1220_;
  assign new_n7012_ = pencrypt_0_ & new_n7011_;
  assign new_n7013_ = n_n2293 & new_n7012_;
  assign new_n7014_ = ~pstart_0_ & new_n7013_;
  assign new_n7015_ = ~new_n7010_ & ~new_n7014_;
  assign new_n7016_ = ~new_n7004_ & ~new_n7008_;
  assign new_n7017_ = new_n7015_ & new_n7016_;
  assign new_n7018_ = ~new_n6998_ & ~new_n7000_;
  assign new_n7019_ = ~new_n6992_ & ~new_n6994_;
  assign new_n7020_ = ~new_n6996_ & new_n7019_;
  assign new_n7021_ = new_n7018_ & new_n7020_;
  assign n1722 = ~new_n7017_ | ~new_n7021_;
  assign new_n7023_ = new_n1200_ & new_n5096_;
  assign new_n7024_ = ~pstart_0_ & new_n7023_;
  assign new_n7025_ = ~new_n1200_ & new_n5091_;
  assign new_n7026_ = ~pstart_0_ & new_n7025_;
  assign new_n7027_ = pkey_130_ & pencrypt_0_;
  assign new_n7028_ = pstart_0_ & new_n7027_;
  assign new_n7029_ = new_n1200_ & new_n5087_;
  assign new_n7030_ = ~pstart_0_ & new_n7029_;
  assign new_n7031_ = pkey_138_ & ~pencrypt_0_;
  assign new_n7032_ = pstart_0_ & new_n7031_;
  assign new_n7033_ = n_n2399 & new_n1220_;
  assign new_n7034_ = pencrypt_0_ & new_n7033_;
  assign new_n7035_ = ~n_n2305 & new_n7034_;
  assign new_n7036_ = ~pstart_0_ & new_n7035_;
  assign new_n7037_ = ~n_n2399 & new_n1220_;
  assign new_n7038_ = pencrypt_0_ & new_n7037_;
  assign new_n7039_ = n_n2305 & new_n7038_;
  assign new_n7040_ = ~pstart_0_ & new_n7039_;
  assign new_n7041_ = ~new_n1200_ & new_n5110_;
  assign new_n7042_ = ~pstart_0_ & new_n7041_;
  assign new_n7043_ = n_n2399 & ~new_n1220_;
  assign new_n7044_ = pencrypt_0_ & new_n7043_;
  assign new_n7045_ = n_n2305 & new_n7044_;
  assign new_n7046_ = ~pstart_0_ & new_n7045_;
  assign new_n7047_ = ~new_n7042_ & ~new_n7046_;
  assign new_n7048_ = ~new_n7036_ & ~new_n7040_;
  assign new_n7049_ = new_n7047_ & new_n7048_;
  assign new_n7050_ = ~new_n7030_ & ~new_n7032_;
  assign new_n7051_ = ~new_n7024_ & ~new_n7026_;
  assign new_n7052_ = ~new_n7028_ & new_n7051_;
  assign new_n7053_ = new_n7050_ & new_n7052_;
  assign n1727 = ~new_n7049_ | ~new_n7053_;
  assign new_n7055_ = new_n1200_ & new_n5134_;
  assign new_n7056_ = ~pstart_0_ & new_n7055_;
  assign new_n7057_ = ~new_n1200_ & new_n5129_;
  assign new_n7058_ = ~pstart_0_ & new_n7057_;
  assign new_n7059_ = pkey_137_ & pencrypt_0_;
  assign new_n7060_ = pstart_0_ & new_n7059_;
  assign new_n7061_ = new_n1200_ & new_n5125_;
  assign new_n7062_ = ~pstart_0_ & new_n7061_;
  assign new_n7063_ = pkey_145_ & ~pencrypt_0_;
  assign new_n7064_ = pstart_0_ & new_n7063_;
  assign new_n7065_ = n_n2407 & new_n1220_;
  assign new_n7066_ = pencrypt_0_ & new_n7065_;
  assign new_n7067_ = ~n_n2312 & new_n7066_;
  assign new_n7068_ = ~pstart_0_ & new_n7067_;
  assign new_n7069_ = ~n_n2407 & new_n1220_;
  assign new_n7070_ = pencrypt_0_ & new_n7069_;
  assign new_n7071_ = n_n2312 & new_n7070_;
  assign new_n7072_ = ~pstart_0_ & new_n7071_;
  assign new_n7073_ = ~new_n1200_ & new_n5148_;
  assign new_n7074_ = ~pstart_0_ & new_n7073_;
  assign new_n7075_ = n_n2407 & ~new_n1220_;
  assign new_n7076_ = pencrypt_0_ & new_n7075_;
  assign new_n7077_ = n_n2312 & new_n7076_;
  assign new_n7078_ = ~pstart_0_ & new_n7077_;
  assign new_n7079_ = ~new_n7074_ & ~new_n7078_;
  assign new_n7080_ = ~new_n7068_ & ~new_n7072_;
  assign new_n7081_ = new_n7079_ & new_n7080_;
  assign new_n7082_ = ~new_n7062_ & ~new_n7064_;
  assign new_n7083_ = ~new_n7056_ & ~new_n7058_;
  assign new_n7084_ = ~new_n7060_ & new_n7083_;
  assign new_n7085_ = new_n7082_ & new_n7084_;
  assign n1732 = ~new_n7081_ | ~new_n7085_;
  assign new_n7087_ = new_n1200_ & new_n3482_;
  assign new_n7088_ = ~pstart_0_ & new_n7087_;
  assign new_n7089_ = ~new_n1200_ & new_n3477_;
  assign new_n7090_ = ~pstart_0_ & new_n7089_;
  assign new_n7091_ = pkey_17_ & pencrypt_0_;
  assign new_n7092_ = pstart_0_ & new_n7091_;
  assign new_n7093_ = new_n1200_ & new_n3473_;
  assign new_n7094_ = ~pstart_0_ & new_n7093_;
  assign new_n7095_ = ~pencrypt_0_ & pkey_25_;
  assign new_n7096_ = pstart_0_ & new_n7095_;
  assign new_n7097_ = n_n2455 & new_n1220_;
  assign new_n7098_ = pencrypt_0_ & new_n7097_;
  assign new_n7099_ = ~n_n2361 & new_n7098_;
  assign new_n7100_ = ~pstart_0_ & new_n7099_;
  assign new_n7101_ = ~n_n2455 & new_n1220_;
  assign new_n7102_ = pencrypt_0_ & new_n7101_;
  assign new_n7103_ = n_n2361 & new_n7102_;
  assign new_n7104_ = ~pstart_0_ & new_n7103_;
  assign new_n7105_ = ~new_n1200_ & new_n3496_;
  assign new_n7106_ = ~pstart_0_ & new_n7105_;
  assign new_n7107_ = n_n2455 & ~new_n1220_;
  assign new_n7108_ = pencrypt_0_ & new_n7107_;
  assign new_n7109_ = n_n2361 & new_n7108_;
  assign new_n7110_ = ~pstart_0_ & new_n7109_;
  assign new_n7111_ = ~new_n7106_ & ~new_n7110_;
  assign new_n7112_ = ~new_n7100_ & ~new_n7104_;
  assign new_n7113_ = new_n7111_ & new_n7112_;
  assign new_n7114_ = ~new_n7094_ & ~new_n7096_;
  assign new_n7115_ = ~new_n7088_ & ~new_n7090_;
  assign new_n7116_ = ~new_n7092_ & new_n7115_;
  assign new_n7117_ = new_n7114_ & new_n7116_;
  assign n1737 = ~new_n7113_ | ~new_n7117_;
  assign new_n7119_ = new_n1200_ & new_n1900_;
  assign new_n7120_ = ~pstart_0_ & new_n7119_;
  assign new_n7121_ = ~new_n1200_ & new_n1895_;
  assign new_n7122_ = ~pstart_0_ & new_n7121_;
  assign new_n7123_ = pkey_250_ & pencrypt_0_;
  assign new_n7124_ = pstart_0_ & new_n7123_;
  assign new_n7125_ = new_n1200_ & new_n1891_;
  assign new_n7126_ = ~pstart_0_ & new_n7125_;
  assign new_n7127_ = pkey_193_ & ~pencrypt_0_;
  assign new_n7128_ = pstart_0_ & new_n7127_;
  assign new_n7129_ = n_n2384 & new_n1220_;
  assign new_n7130_ = pencrypt_0_ & new_n7129_;
  assign new_n7131_ = ~n_n2749 & new_n7130_;
  assign new_n7132_ = ~pstart_0_ & new_n7131_;
  assign new_n7133_ = ~n_n2384 & new_n1220_;
  assign new_n7134_ = pencrypt_0_ & new_n7133_;
  assign new_n7135_ = n_n2749 & new_n7134_;
  assign new_n7136_ = ~pstart_0_ & new_n7135_;
  assign new_n7137_ = ~new_n1200_ & new_n1914_;
  assign new_n7138_ = ~pstart_0_ & new_n7137_;
  assign new_n7139_ = n_n2384 & ~new_n1220_;
  assign new_n7140_ = pencrypt_0_ & new_n7139_;
  assign new_n7141_ = n_n2749 & new_n7140_;
  assign new_n7142_ = ~pstart_0_ & new_n7141_;
  assign new_n7143_ = ~new_n7138_ & ~new_n7142_;
  assign new_n7144_ = ~new_n7132_ & ~new_n7136_;
  assign new_n7145_ = new_n7143_ & new_n7144_;
  assign new_n7146_ = ~new_n7126_ & ~new_n7128_;
  assign new_n7147_ = ~new_n7120_ & ~new_n7122_;
  assign new_n7148_ = ~new_n7124_ & new_n7147_;
  assign new_n7149_ = new_n7146_ & new_n7148_;
  assign n1742 = ~new_n7145_ | ~new_n7149_;
  assign new_n7151_ = new_n1200_ & new_n1938_;
  assign new_n7152_ = ~pstart_0_ & new_n7151_;
  assign new_n7153_ = ~new_n1200_ & new_n1933_;
  assign new_n7154_ = ~pstart_0_ & new_n7153_;
  assign new_n7155_ = pkey_208_ & pencrypt_0_;
  assign new_n7156_ = pstart_0_ & new_n7155_;
  assign new_n7157_ = new_n1200_ & new_n1929_;
  assign new_n7158_ = ~pstart_0_ & new_n7157_;
  assign new_n7159_ = pkey_216_ & ~pencrypt_0_;
  assign new_n7160_ = pstart_0_ & new_n7159_;
  assign new_n7161_ = n_n2390 & new_n1220_;
  assign new_n7162_ = pencrypt_0_ & new_n7161_;
  assign new_n7163_ = ~n_n2296 & new_n7162_;
  assign new_n7164_ = ~pstart_0_ & new_n7163_;
  assign new_n7165_ = ~n_n2390 & new_n1220_;
  assign new_n7166_ = pencrypt_0_ & new_n7165_;
  assign new_n7167_ = n_n2296 & new_n7166_;
  assign new_n7168_ = ~pstart_0_ & new_n7167_;
  assign new_n7169_ = ~new_n1200_ & new_n1952_1_;
  assign new_n7170_ = ~pstart_0_ & new_n7169_;
  assign new_n7171_ = n_n2390 & ~new_n1220_;
  assign new_n7172_ = pencrypt_0_ & new_n7171_;
  assign new_n7173_ = n_n2296 & new_n7172_;
  assign new_n7174_ = ~pstart_0_ & new_n7173_;
  assign new_n7175_ = ~new_n7170_ & ~new_n7174_;
  assign new_n7176_ = ~new_n7164_ & ~new_n7168_;
  assign new_n7177_ = new_n7175_ & new_n7176_;
  assign new_n7178_ = ~new_n7158_ & ~new_n7160_;
  assign new_n7179_ = ~new_n7152_ & ~new_n7154_;
  assign new_n7180_ = ~new_n7156_ & new_n7179_;
  assign new_n7181_ = new_n7178_ & new_n7180_;
  assign n1747 = ~new_n7177_ | ~new_n7181_;
  assign new_n7183_ = new_n1200_ & new_n4120_;
  assign new_n7184_ = ~pstart_0_ & new_n7183_;
  assign new_n7185_ = ~new_n1200_ & new_n4115_;
  assign new_n7186_ = ~pstart_0_ & new_n7185_;
  assign new_n7187_ = pkey_171_ & pencrypt_0_;
  assign new_n7188_ = pstart_0_ & new_n7187_;
  assign new_n7189_ = new_n1200_ & new_n4111_;
  assign new_n7190_ = ~pstart_0_ & new_n7189_;
  assign new_n7191_ = ~pencrypt_0_ & pkey_179_;
  assign new_n7192_ = pstart_0_ & new_n7191_;
  assign new_n7193_ = n_n2899 & new_n1220_;
  assign new_n7194_ = pencrypt_0_ & new_n7193_;
  assign new_n7195_ = ~n_n2303 & new_n7194_;
  assign new_n7196_ = ~pstart_0_ & new_n7195_;
  assign new_n7197_ = ~n_n2899 & new_n1220_;
  assign new_n7198_ = pencrypt_0_ & new_n7197_;
  assign new_n7199_ = n_n2303 & new_n7198_;
  assign new_n7200_ = ~pstart_0_ & new_n7199_;
  assign new_n7201_ = ~new_n1200_ & new_n4134_;
  assign new_n7202_ = ~pstart_0_ & new_n7201_;
  assign new_n7203_ = n_n2899 & ~new_n1220_;
  assign new_n7204_ = pencrypt_0_ & new_n7203_;
  assign new_n7205_ = n_n2303 & new_n7204_;
  assign new_n7206_ = ~pstart_0_ & new_n7205_;
  assign new_n7207_ = ~new_n7202_ & ~new_n7206_;
  assign new_n7208_ = ~new_n7196_ & ~new_n7200_;
  assign new_n7209_ = new_n7207_ & new_n7208_;
  assign new_n7210_ = ~new_n7190_ & ~new_n7192_;
  assign new_n7211_ = ~new_n7184_ & ~new_n7186_;
  assign new_n7212_ = ~new_n7188_ & new_n7211_;
  assign new_n7213_ = new_n7210_ & new_n7212_;
  assign n1752 = ~new_n7209_ | ~new_n7213_;
  assign new_n7215_ = new_n1200_ & new_n4158_;
  assign new_n7216_ = ~pstart_0_ & new_n7215_;
  assign new_n7217_ = ~new_n1200_ & new_n4153_;
  assign new_n7218_ = ~pstart_0_ & new_n7217_;
  assign new_n7219_ = pkey_129_ & pencrypt_0_;
  assign new_n7220_ = pstart_0_ & new_n7219_;
  assign new_n7221_ = new_n1200_ & new_n4149_;
  assign new_n7222_ = ~pstart_0_ & new_n7221_;
  assign new_n7223_ = pkey_137_ & ~pencrypt_0_;
  assign new_n7224_ = pstart_0_ & new_n7223_;
  assign new_n7225_ = n_n2406 & new_n1220_;
  assign new_n7226_ = pencrypt_0_ & new_n7225_;
  assign new_n7227_ = ~n_n2311 & new_n7226_;
  assign new_n7228_ = ~pstart_0_ & new_n7227_;
  assign new_n7229_ = ~n_n2406 & new_n1220_;
  assign new_n7230_ = pencrypt_0_ & new_n7229_;
  assign new_n7231_ = n_n2311 & new_n7230_;
  assign new_n7232_ = ~pstart_0_ & new_n7231_;
  assign new_n7233_ = ~new_n1200_ & new_n4172_;
  assign new_n7234_ = ~pstart_0_ & new_n7233_;
  assign new_n7235_ = n_n2406 & ~new_n1220_;
  assign new_n7236_ = pencrypt_0_ & new_n7235_;
  assign new_n7237_ = n_n2311 & new_n7236_;
  assign new_n7238_ = ~pstart_0_ & new_n7237_;
  assign new_n7239_ = ~new_n7234_ & ~new_n7238_;
  assign new_n7240_ = ~new_n7228_ & ~new_n7232_;
  assign new_n7241_ = new_n7239_ & new_n7240_;
  assign new_n7242_ = ~new_n7222_ & ~new_n7224_;
  assign new_n7243_ = ~new_n7216_ & ~new_n7218_;
  assign new_n7244_ = ~new_n7220_ & new_n7243_;
  assign new_n7245_ = new_n7242_ & new_n7244_;
  assign n1757 = ~new_n7241_ | ~new_n7245_;
  assign new_n7247_ = new_n1200_ & new_n2236_;
  assign new_n7248_ = ~pstart_0_ & new_n7247_;
  assign new_n7249_ = ~new_n1200_ & new_n2231_;
  assign new_n7250_ = ~pstart_0_ & new_n7249_;
  assign new_n7251_ = pkey_193_ & pencrypt_0_;
  assign new_n7252_ = pstart_0_ & new_n7251_;
  assign new_n7253_ = new_n1200_ & new_n2227_;
  assign new_n7254_ = ~pstart_0_ & new_n7253_;
  assign new_n7255_ = ~pencrypt_0_ & pkey_201_;
  assign new_n7256_ = pstart_0_ & new_n7255_;
  assign new_n7257_ = n_n2877 & new_n1220_;
  assign new_n7258_ = pencrypt_0_ & new_n7257_;
  assign new_n7259_ = ~n_n2287 & new_n7258_;
  assign new_n7260_ = ~pstart_0_ & new_n7259_;
  assign new_n7261_ = ~n_n2877 & new_n1220_;
  assign new_n7262_ = pencrypt_0_ & new_n7261_;
  assign new_n7263_ = n_n2287 & new_n7262_;
  assign new_n7264_ = ~pstart_0_ & new_n7263_;
  assign new_n7265_ = ~new_n1200_ & new_n2250_;
  assign new_n7266_ = ~pstart_0_ & new_n7265_;
  assign new_n7267_ = n_n2877 & ~new_n1220_;
  assign new_n7268_ = pencrypt_0_ & new_n7267_;
  assign new_n7269_ = n_n2287 & new_n7268_;
  assign new_n7270_ = ~pstart_0_ & new_n7269_;
  assign new_n7271_ = ~new_n7266_ & ~new_n7270_;
  assign new_n7272_ = ~new_n7260_ & ~new_n7264_;
  assign new_n7273_ = new_n7271_ & new_n7272_;
  assign new_n7274_ = ~new_n7254_ & ~new_n7256_;
  assign new_n7275_ = ~new_n7248_ & ~new_n7250_;
  assign new_n7276_ = ~new_n7252_ & new_n7275_;
  assign new_n7277_ = new_n7274_ & new_n7276_;
  assign n1762 = ~new_n7273_ | ~new_n7277_;
  assign new_n7279_ = new_n1200_ & new_n2274_;
  assign new_n7280_ = ~pstart_0_ & new_n7279_;
  assign new_n7281_ = ~new_n1200_ & new_n2269_;
  assign new_n7282_ = ~pstart_0_ & new_n7281_;
  assign new_n7283_ = pencrypt_0_ & pkey_200_;
  assign new_n7284_ = pstart_0_ & new_n7283_;
  assign new_n7285_ = new_n1200_ & new_n2265_;
  assign new_n7286_ = ~pstart_0_ & new_n7285_;
  assign new_n7287_ = pkey_208_ & ~pencrypt_0_;
  assign new_n7288_ = pstart_0_ & new_n7287_;
  assign new_n7289_ = n_n2389 & new_n1220_;
  assign new_n7290_ = pencrypt_0_ & new_n7289_;
  assign new_n7291_ = ~n_n2295 & new_n7290_;
  assign new_n7292_ = ~pstart_0_ & new_n7291_;
  assign new_n7293_ = ~n_n2389 & new_n1220_;
  assign new_n7294_ = pencrypt_0_ & new_n7293_;
  assign new_n7295_ = n_n2295 & new_n7294_;
  assign new_n7296_ = ~pstart_0_ & new_n7295_;
  assign new_n7297_ = ~new_n1200_ & new_n2288_;
  assign new_n7298_ = ~pstart_0_ & new_n7297_;
  assign new_n7299_ = n_n2389 & ~new_n1220_;
  assign new_n7300_ = pencrypt_0_ & new_n7299_;
  assign new_n7301_ = n_n2295 & new_n7300_;
  assign new_n7302_ = ~pstart_0_ & new_n7301_;
  assign new_n7303_ = ~new_n7298_ & ~new_n7302_;
  assign new_n7304_ = ~new_n7292_ & ~new_n7296_;
  assign new_n7305_ = new_n7303_ & new_n7304_;
  assign new_n7306_ = ~new_n7286_ & ~new_n7288_;
  assign new_n7307_ = ~new_n7280_ & ~new_n7282_;
  assign new_n7308_ = ~new_n7284_ & new_n7307_;
  assign new_n7309_ = new_n7306_ & new_n7308_;
  assign n1767 = ~new_n7305_ | ~new_n7309_;
  assign new_n7311_ = new_n1200_ & new_n4380_;
  assign new_n7312_ = ~pstart_0_ & new_n7311_;
  assign new_n7313_ = ~new_n1200_ & new_n4375_;
  assign new_n7314_ = ~pstart_0_ & new_n7313_;
  assign new_n7315_ = pencrypt_0_ & pkey_179_;
  assign new_n7316_ = pstart_0_ & new_n7315_;
  assign new_n7317_ = new_n1200_ & new_n4371_;
  assign new_n7318_ = ~pstart_0_ & new_n7317_;
  assign new_n7319_ = ~pencrypt_0_ & pkey_187_;
  assign new_n7320_ = pstart_0_ & new_n7319_;
  assign new_n7321_ = n_n2397 & new_n1220_;
  assign new_n7322_ = pencrypt_0_ & new_n7321_;
  assign new_n7323_ = ~n_n2770 & new_n7322_;
  assign new_n7324_ = ~pstart_0_ & new_n7323_;
  assign new_n7325_ = ~n_n2397 & new_n1220_;
  assign new_n7326_ = pencrypt_0_ & new_n7325_;
  assign new_n7327_ = n_n2770 & new_n7326_;
  assign new_n7328_ = ~pstart_0_ & new_n7327_;
  assign new_n7329_ = ~new_n1200_ & new_n4394_;
  assign new_n7330_ = ~pstart_0_ & new_n7329_;
  assign new_n7331_ = n_n2397 & ~new_n1220_;
  assign new_n7332_ = pencrypt_0_ & new_n7331_;
  assign new_n7333_ = n_n2770 & new_n7332_;
  assign new_n7334_ = ~pstart_0_ & new_n7333_;
  assign new_n7335_ = ~new_n7330_ & ~new_n7334_;
  assign new_n7336_ = ~new_n7324_ & ~new_n7328_;
  assign new_n7337_ = new_n7335_ & new_n7336_;
  assign new_n7338_ = ~new_n7318_ & ~new_n7320_;
  assign new_n7339_ = ~new_n7312_ & ~new_n7314_;
  assign new_n7340_ = ~new_n7316_ & new_n7339_;
  assign new_n7341_ = new_n7338_ & new_n7340_;
  assign n1772 = ~new_n7337_ | ~new_n7341_;
  assign new_n7343_ = new_n1200_ & new_n4418_;
  assign new_n7344_ = ~pstart_0_ & new_n7343_;
  assign new_n7345_ = ~new_n1200_ & new_n4413_;
  assign new_n7346_ = ~pstart_0_ & new_n7345_;
  assign new_n7347_ = pencrypt_0_ & pkey_186_;
  assign new_n7348_ = pstart_0_ & new_n7347_;
  assign new_n7349_ = new_n1200_ & new_n4409_;
  assign new_n7350_ = ~pstart_0_ & new_n7349_;
  assign new_n7351_ = pkey_129_ & ~pencrypt_0_;
  assign new_n7352_ = pstart_0_ & new_n7351_;
  assign new_n7353_ = n_n2405 & new_n1220_;
  assign new_n7354_ = pencrypt_0_ & new_n7353_;
  assign new_n7355_ = ~n_n2310 & new_n7354_;
  assign new_n7356_ = ~pstart_0_ & new_n7355_;
  assign new_n7357_ = ~n_n2405 & new_n1220_;
  assign new_n7358_ = pencrypt_0_ & new_n7357_;
  assign new_n7359_ = n_n2310 & new_n7358_;
  assign new_n7360_ = ~pstart_0_ & new_n7359_;
  assign new_n7361_ = ~new_n1200_ & new_n4432_;
  assign new_n7362_ = ~pstart_0_ & new_n7361_;
  assign new_n7363_ = n_n2405 & ~new_n1220_;
  assign new_n7364_ = pencrypt_0_ & new_n7363_;
  assign new_n7365_ = n_n2310 & new_n7364_;
  assign new_n7366_ = ~pstart_0_ & new_n7365_;
  assign new_n7367_ = ~new_n7362_ & ~new_n7366_;
  assign new_n7368_ = ~new_n7356_ & ~new_n7360_;
  assign new_n7369_ = new_n7367_ & new_n7368_;
  assign new_n7370_ = ~new_n7350_ & ~new_n7352_;
  assign new_n7371_ = ~new_n7344_ & ~new_n7346_;
  assign new_n7372_ = ~new_n7348_ & new_n7371_;
  assign new_n7373_ = new_n7370_ & new_n7372_;
  assign n1777 = ~new_n7369_ | ~new_n7373_;
  assign new_n7375_ = new_n1200_ & new_n1292_1_;
  assign new_n7376_ = ~pstart_0_ & new_n7375_;
  assign new_n7377_ = ~new_n1200_ & new_n1287_1_;
  assign new_n7378_ = ~pstart_0_ & new_n7377_;
  assign new_n7379_ = pencrypt_0_ & pkey_201_;
  assign new_n7380_ = pstart_0_ & new_n7379_;
  assign new_n7381_ = new_n1200_ & new_n1283_;
  assign new_n7382_ = ~pstart_0_ & new_n7381_;
  assign new_n7383_ = pkey_209_ & ~pencrypt_0_;
  assign new_n7384_ = pstart_0_ & new_n7383_;
  assign new_n7385_ = n_n2879 & new_n1220_;
  assign new_n7386_ = pencrypt_0_ & new_n7385_;
  assign new_n7387_ = ~n_n2288 & new_n7386_;
  assign new_n7388_ = ~pstart_0_ & new_n7387_;
  assign new_n7389_ = ~n_n2879 & new_n1220_;
  assign new_n7390_ = pencrypt_0_ & new_n7389_;
  assign new_n7391_ = n_n2288 & new_n7390_;
  assign new_n7392_ = ~pstart_0_ & new_n7391_;
  assign new_n7393_ = ~new_n1200_ & new_n1306_;
  assign new_n7394_ = ~pstart_0_ & new_n7393_;
  assign new_n7395_ = n_n2879 & ~new_n1220_;
  assign new_n7396_ = pencrypt_0_ & new_n7395_;
  assign new_n7397_ = n_n2288 & new_n7396_;
  assign new_n7398_ = ~pstart_0_ & new_n7397_;
  assign new_n7399_ = ~new_n7394_ & ~new_n7398_;
  assign new_n7400_ = ~new_n7388_ & ~new_n7392_;
  assign new_n7401_ = new_n7399_ & new_n7400_;
  assign new_n7402_ = ~new_n7382_ & ~new_n7384_;
  assign new_n7403_ = ~new_n7376_ & ~new_n7378_;
  assign new_n7404_ = ~new_n7380_ & new_n7403_;
  assign new_n7405_ = new_n7402_ & new_n7404_;
  assign n1782 = ~new_n7401_ | ~new_n7405_;
  assign new_n7407_ = new_n1200_ & new_n1330_;
  assign new_n7408_ = ~pstart_0_ & new_n7407_;
  assign new_n7409_ = ~new_n1200_ & new_n1325_;
  assign new_n7410_ = ~pstart_0_ & new_n7409_;
  assign new_n7411_ = pkey_224_ & pencrypt_0_;
  assign new_n7412_ = pstart_0_ & new_n7411_;
  assign new_n7413_ = new_n1200_ & new_n1321_;
  assign new_n7414_ = ~pstart_0_ & new_n7413_;
  assign new_n7415_ = pkey_232_ & ~pencrypt_0_;
  assign new_n7416_ = pstart_0_ & new_n7415_;
  assign new_n7417_ = n_n2392 & new_n1220_;
  assign new_n7418_ = pencrypt_0_ & new_n7417_;
  assign new_n7419_ = ~n_n2298 & new_n7418_;
  assign new_n7420_ = ~pstart_0_ & new_n7419_;
  assign new_n7421_ = ~n_n2392 & new_n1220_;
  assign new_n7422_ = pencrypt_0_ & new_n7421_;
  assign new_n7423_ = n_n2298 & new_n7422_;
  assign new_n7424_ = ~pstart_0_ & new_n7423_;
  assign new_n7425_ = ~new_n1200_ & new_n1344_;
  assign new_n7426_ = ~pstart_0_ & new_n7425_;
  assign new_n7427_ = n_n2392 & ~new_n1220_;
  assign new_n7428_ = pencrypt_0_ & new_n7427_;
  assign new_n7429_ = n_n2298 & new_n7428_;
  assign new_n7430_ = ~pstart_0_ & new_n7429_;
  assign new_n7431_ = ~new_n7426_ & ~new_n7430_;
  assign new_n7432_ = ~new_n7420_ & ~new_n7424_;
  assign new_n7433_ = new_n7431_ & new_n7432_;
  assign new_n7434_ = ~new_n7414_ & ~new_n7416_;
  assign new_n7435_ = ~new_n7408_ & ~new_n7410_;
  assign new_n7436_ = ~new_n7412_ & new_n7435_;
  assign new_n7437_ = new_n7434_ & new_n7436_;
  assign n1787 = ~new_n7433_ | ~new_n7437_;
  assign new_n7439_ = new_n1200_ & new_n1368_;
  assign new_n7440_ = ~pstart_0_ & new_n7439_;
  assign new_n7441_ = ~new_n1200_ & new_n1363_;
  assign new_n7442_ = ~pstart_0_ & new_n7441_;
  assign new_n7443_ = pkey_154_ & pencrypt_0_;
  assign new_n7444_ = pstart_0_ & new_n7443_;
  assign new_n7445_ = new_n1200_ & new_n1359_;
  assign new_n7446_ = ~pstart_0_ & new_n7445_;
  assign new_n7447_ = pkey_162_ & ~pencrypt_0_;
  assign new_n7448_ = pstart_0_ & new_n7447_;
  assign new_n7449_ = n_n2402 & new_n1220_;
  assign new_n7450_ = pencrypt_0_ & new_n7449_;
  assign new_n7451_ = ~n_n2307 & new_n7450_;
  assign new_n7452_ = ~pstart_0_ & new_n7451_;
  assign new_n7453_ = ~n_n2402 & new_n1220_;
  assign new_n7454_ = pencrypt_0_ & new_n7453_;
  assign new_n7455_ = n_n2307 & new_n7454_;
  assign new_n7456_ = ~pstart_0_ & new_n7455_;
  assign new_n7457_ = ~new_n1200_ & new_n1382_1_;
  assign new_n7458_ = ~pstart_0_ & new_n7457_;
  assign new_n7459_ = n_n2402 & ~new_n1220_;
  assign new_n7460_ = pencrypt_0_ & new_n7459_;
  assign new_n7461_ = n_n2307 & new_n7460_;
  assign new_n7462_ = ~pstart_0_ & new_n7461_;
  assign new_n7463_ = ~new_n7458_ & ~new_n7462_;
  assign new_n7464_ = ~new_n7452_ & ~new_n7456_;
  assign new_n7465_ = new_n7463_ & new_n7464_;
  assign new_n7466_ = ~new_n7446_ & ~new_n7448_;
  assign new_n7467_ = ~new_n7440_ & ~new_n7442_;
  assign new_n7468_ = ~new_n7444_ & new_n7467_;
  assign new_n7469_ = new_n7466_ & new_n7468_;
  assign n1792 = ~new_n7465_ | ~new_n7469_;
  assign new_n7471_ = new_n1200_ & new_n1406_;
  assign new_n7472_ = ~pstart_0_ & new_n7471_;
  assign new_n7473_ = ~new_n1200_ & new_n1401_;
  assign new_n7474_ = ~pstart_0_ & new_n7473_;
  assign new_n7475_ = pencrypt_0_ & pkey_177_;
  assign new_n7476_ = pstart_0_ & new_n7475_;
  assign new_n7477_ = new_n1200_ & new_n1397_1_;
  assign new_n7478_ = ~pstart_0_ & new_n7477_;
  assign new_n7479_ = ~pencrypt_0_ & pkey_185_;
  assign new_n7480_ = pstart_0_ & new_n7479_;
  assign new_n7481_ = n_n2411 & new_n1220_;
  assign new_n7482_ = pencrypt_0_ & new_n7481_;
  assign new_n7483_ = ~n_n2789 & new_n7482_;
  assign new_n7484_ = ~pstart_0_ & new_n7483_;
  assign new_n7485_ = ~n_n2411 & new_n1220_;
  assign new_n7486_ = pencrypt_0_ & new_n7485_;
  assign new_n7487_ = n_n2789 & new_n7486_;
  assign new_n7488_ = ~pstart_0_ & new_n7487_;
  assign new_n7489_ = ~new_n1200_ & new_n1420_;
  assign new_n7490_ = ~pstart_0_ & new_n7489_;
  assign new_n7491_ = n_n2411 & ~new_n1220_;
  assign new_n7492_ = pencrypt_0_ & new_n7491_;
  assign new_n7493_ = n_n2789 & new_n7492_;
  assign new_n7494_ = ~pstart_0_ & new_n7493_;
  assign new_n7495_ = ~new_n7490_ & ~new_n7494_;
  assign new_n7496_ = ~new_n7484_ & ~new_n7488_;
  assign new_n7497_ = new_n7495_ & new_n7496_;
  assign new_n7498_ = ~new_n7478_ & ~new_n7480_;
  assign new_n7499_ = ~new_n7472_ & ~new_n7474_;
  assign new_n7500_ = ~new_n7476_ & new_n7499_;
  assign new_n7501_ = new_n7498_ & new_n7500_;
  assign n1797 = ~new_n7497_ | ~new_n7501_;
  assign new_n7503_ = new_n1200_ & new_n4494_;
  assign new_n7504_ = ~pstart_0_ & new_n7503_;
  assign new_n7505_ = ~new_n1200_ & new_n4489_;
  assign new_n7506_ = ~pstart_0_ & new_n7505_;
  assign new_n7507_ = pkey_107_ & pencrypt_0_;
  assign new_n7508_ = pstart_0_ & new_n7507_;
  assign new_n7509_ = new_n1200_ & new_n4485_;
  assign new_n7510_ = ~pstart_0_ & new_n7509_;
  assign new_n7511_ = pkey_115_ & ~pencrypt_0_;
  assign new_n7512_ = pstart_0_ & new_n7511_;
  assign new_n7513_ = n_n2931 & new_n1220_;
  assign new_n7514_ = pencrypt_0_ & new_n7513_;
  assign new_n7515_ = ~n_n2327 & new_n7514_;
  assign new_n7516_ = ~pstart_0_ & new_n7515_;
  assign new_n7517_ = ~n_n2931 & new_n1220_;
  assign new_n7518_ = pencrypt_0_ & new_n7517_;
  assign new_n7519_ = n_n2327 & new_n7518_;
  assign new_n7520_ = ~pstart_0_ & new_n7519_;
  assign new_n7521_ = ~new_n1200_ & new_n4508_;
  assign new_n7522_ = ~pstart_0_ & new_n7521_;
  assign new_n7523_ = n_n2931 & ~new_n1220_;
  assign new_n7524_ = pencrypt_0_ & new_n7523_;
  assign new_n7525_ = n_n2327 & new_n7524_;
  assign new_n7526_ = ~pstart_0_ & new_n7525_;
  assign new_n7527_ = ~new_n7522_ & ~new_n7526_;
  assign new_n7528_ = ~new_n7516_ & ~new_n7520_;
  assign new_n7529_ = new_n7527_ & new_n7528_;
  assign new_n7530_ = ~new_n7510_ & ~new_n7512_;
  assign new_n7531_ = ~new_n7504_ & ~new_n7506_;
  assign new_n7532_ = ~new_n7508_ & new_n7531_;
  assign new_n7533_ = new_n7530_ & new_n7532_;
  assign n1802 = ~new_n7529_ | ~new_n7533_;
  assign new_n7535_ = new_n1200_ & new_n5248_;
  assign new_n7536_ = ~pstart_0_ & new_n7535_;
  assign new_n7537_ = ~new_n1200_ & new_n5243_;
  assign new_n7538_ = ~pstart_0_ & new_n7537_;
  assign new_n7539_ = pencrypt_0_ & pkey_65_;
  assign new_n7540_ = pstart_0_ & new_n7539_;
  assign new_n7541_ = new_n1200_ & new_n5239_;
  assign new_n7542_ = ~pstart_0_ & new_n7541_;
  assign new_n7543_ = ~pencrypt_0_ & pkey_73_;
  assign new_n7544_ = pstart_0_ & new_n7543_;
  assign new_n7545_ = n_n2943 & new_n1220_;
  assign new_n7546_ = pencrypt_0_ & new_n7545_;
  assign new_n7547_ = ~n_n2335 & new_n7546_;
  assign new_n7548_ = ~pstart_0_ & new_n7547_;
  assign new_n7549_ = ~n_n2943 & new_n1220_;
  assign new_n7550_ = pencrypt_0_ & new_n7549_;
  assign new_n7551_ = n_n2335 & new_n7550_;
  assign new_n7552_ = ~pstart_0_ & new_n7551_;
  assign new_n7553_ = ~new_n1200_ & new_n5262_;
  assign new_n7554_ = ~pstart_0_ & new_n7553_;
  assign new_n7555_ = n_n2943 & ~new_n1220_;
  assign new_n7556_ = pencrypt_0_ & new_n7555_;
  assign new_n7557_ = n_n2335 & new_n7556_;
  assign new_n7558_ = ~pstart_0_ & new_n7557_;
  assign new_n7559_ = ~new_n7554_ & ~new_n7558_;
  assign new_n7560_ = ~new_n7548_ & ~new_n7552_;
  assign new_n7561_ = new_n7559_ & new_n7560_;
  assign new_n7562_ = ~new_n7542_ & ~new_n7544_;
  assign new_n7563_ = ~new_n7536_ & ~new_n7538_;
  assign new_n7564_ = ~new_n7540_ & new_n7563_;
  assign new_n7565_ = new_n7562_ & new_n7564_;
  assign n1807 = ~new_n7561_ | ~new_n7565_;
  assign new_n7567_ = new_n1200_ & new_n1596_;
  assign new_n7568_ = ~pstart_0_ & new_n7567_;
  assign new_n7569_ = ~new_n1200_ & new_n1591_;
  assign new_n7570_ = ~pstart_0_ & new_n7569_;
  assign new_n7571_ = pkey_209_ & pencrypt_0_;
  assign new_n7572_ = pstart_0_ & new_n7571_;
  assign new_n7573_ = new_n1200_ & new_n1587_1_;
  assign new_n7574_ = ~pstart_0_ & new_n7573_;
  assign new_n7575_ = pkey_217_ & ~pencrypt_0_;
  assign new_n7576_ = pstart_0_ & new_n7575_;
  assign new_n7577_ = n_n2881 & new_n1220_;
  assign new_n7578_ = pencrypt_0_ & new_n7577_;
  assign new_n7579_ = ~n_n2289 & new_n7578_;
  assign new_n7580_ = ~pstart_0_ & new_n7579_;
  assign new_n7581_ = ~n_n2881 & new_n1220_;
  assign new_n7582_ = pencrypt_0_ & new_n7581_;
  assign new_n7583_ = n_n2289 & new_n7582_;
  assign new_n7584_ = ~pstart_0_ & new_n7583_;
  assign new_n7585_ = ~new_n1200_ & new_n1610_;
  assign new_n7586_ = ~pstart_0_ & new_n7585_;
  assign new_n7587_ = n_n2881 & ~new_n1220_;
  assign new_n7588_ = pencrypt_0_ & new_n7587_;
  assign new_n7589_ = n_n2289 & new_n7588_;
  assign new_n7590_ = ~pstart_0_ & new_n7589_;
  assign new_n7591_ = ~new_n7586_ & ~new_n7590_;
  assign new_n7592_ = ~new_n7580_ & ~new_n7584_;
  assign new_n7593_ = new_n7591_ & new_n7592_;
  assign new_n7594_ = ~new_n7574_ & ~new_n7576_;
  assign new_n7595_ = ~new_n7568_ & ~new_n7570_;
  assign new_n7596_ = ~new_n7572_ & new_n7595_;
  assign new_n7597_ = new_n7594_ & new_n7596_;
  assign n1812 = ~new_n7593_ | ~new_n7597_;
  assign new_n7599_ = new_n1200_ & new_n1634_;
  assign new_n7600_ = ~pstart_0_ & new_n7599_;
  assign new_n7601_ = ~new_n1200_ & new_n1629_;
  assign new_n7602_ = ~pstart_0_ & new_n7601_;
  assign new_n7603_ = pkey_216_ & pencrypt_0_;
  assign new_n7604_ = pstart_0_ & new_n7603_;
  assign new_n7605_ = new_n1200_ & new_n1625_;
  assign new_n7606_ = ~pstart_0_ & new_n7605_;
  assign new_n7607_ = pkey_224_ & ~pencrypt_0_;
  assign new_n7608_ = pstart_0_ & new_n7607_;
  assign new_n7609_ = n_n2391 & new_n1220_;
  assign new_n7610_ = pencrypt_0_ & new_n7609_;
  assign new_n7611_ = ~n_n2297 & new_n7610_;
  assign new_n7612_ = ~pstart_0_ & new_n7611_;
  assign new_n7613_ = ~n_n2391 & new_n1220_;
  assign new_n7614_ = pencrypt_0_ & new_n7613_;
  assign new_n7615_ = n_n2297 & new_n7614_;
  assign new_n7616_ = ~pstart_0_ & new_n7615_;
  assign new_n7617_ = ~new_n1200_ & new_n1648_;
  assign new_n7618_ = ~pstart_0_ & new_n7617_;
  assign new_n7619_ = n_n2391 & ~new_n1220_;
  assign new_n7620_ = pencrypt_0_ & new_n7619_;
  assign new_n7621_ = n_n2297 & new_n7620_;
  assign new_n7622_ = ~pstart_0_ & new_n7621_;
  assign new_n7623_ = ~new_n7618_ & ~new_n7622_;
  assign new_n7624_ = ~new_n7612_ & ~new_n7616_;
  assign new_n7625_ = new_n7623_ & new_n7624_;
  assign new_n7626_ = ~new_n7606_ & ~new_n7608_;
  assign new_n7627_ = ~new_n7600_ & ~new_n7602_;
  assign new_n7628_ = ~new_n7604_ & new_n7627_;
  assign new_n7629_ = new_n7626_ & new_n7628_;
  assign n1817 = ~new_n7625_ | ~new_n7629_;
  assign new_n7631_ = new_n1200_ & new_n1672_1_;
  assign new_n7632_ = ~pstart_0_ & new_n7631_;
  assign new_n7633_ = ~new_n1200_ & new_n1667_1_;
  assign new_n7634_ = ~pstart_0_ & new_n7633_;
  assign new_n7635_ = pkey_162_ & pencrypt_0_;
  assign new_n7636_ = pstart_0_ & new_n7635_;
  assign new_n7637_ = new_n1200_ & new_n1663_;
  assign new_n7638_ = ~pstart_0_ & new_n7637_;
  assign new_n7639_ = ~pencrypt_0_ & pkey_170_;
  assign new_n7640_ = pstart_0_ & new_n7639_;
  assign new_n7641_ = n_n2403 & new_n1220_;
  assign new_n7642_ = pencrypt_0_ & new_n7641_;
  assign new_n7643_ = ~n_n2308 & new_n7642_;
  assign new_n7644_ = ~pstart_0_ & new_n7643_;
  assign new_n7645_ = ~n_n2403 & new_n1220_;
  assign new_n7646_ = pencrypt_0_ & new_n7645_;
  assign new_n7647_ = n_n2308 & new_n7646_;
  assign new_n7648_ = ~pstart_0_ & new_n7647_;
  assign new_n7649_ = ~new_n1200_ & new_n1686_;
  assign new_n7650_ = ~pstart_0_ & new_n7649_;
  assign new_n7651_ = n_n2403 & ~new_n1220_;
  assign new_n7652_ = pencrypt_0_ & new_n7651_;
  assign new_n7653_ = n_n2308 & new_n7652_;
  assign new_n7654_ = ~pstart_0_ & new_n7653_;
  assign new_n7655_ = ~new_n7650_ & ~new_n7654_;
  assign new_n7656_ = ~new_n7644_ & ~new_n7648_;
  assign new_n7657_ = new_n7655_ & new_n7656_;
  assign new_n7658_ = ~new_n7638_ & ~new_n7640_;
  assign new_n7659_ = ~new_n7632_ & ~new_n7634_;
  assign new_n7660_ = ~new_n7636_ & new_n7659_;
  assign new_n7661_ = new_n7658_ & new_n7660_;
  assign n1822 = ~new_n7657_ | ~new_n7661_;
  assign new_n7663_ = new_n1200_ & new_n1710_;
  assign new_n7664_ = ~pstart_0_ & new_n7663_;
  assign new_n7665_ = ~new_n1200_ & new_n1705_;
  assign new_n7666_ = ~pstart_0_ & new_n7665_;
  assign new_n7667_ = pkey_169_ & pencrypt_0_;
  assign new_n7668_ = pstart_0_ & new_n7667_;
  assign new_n7669_ = new_n1200_ & new_n1701_;
  assign new_n7670_ = ~pstart_0_ & new_n7669_;
  assign new_n7671_ = ~pencrypt_0_ & pkey_177_;
  assign new_n7672_ = pstart_0_ & new_n7671_;
  assign new_n7673_ = n_n2917 & new_n1220_;
  assign new_n7674_ = pencrypt_0_ & new_n7673_;
  assign new_n7675_ = ~n_n2316 & new_n7674_;
  assign new_n7676_ = ~pstart_0_ & new_n7675_;
  assign new_n7677_ = ~n_n2917 & new_n1220_;
  assign new_n7678_ = pencrypt_0_ & new_n7677_;
  assign new_n7679_ = n_n2316 & new_n7678_;
  assign new_n7680_ = ~pstart_0_ & new_n7679_;
  assign new_n7681_ = ~new_n1200_ & new_n1724_;
  assign new_n7682_ = ~pstart_0_ & new_n7681_;
  assign new_n7683_ = n_n2917 & ~new_n1220_;
  assign new_n7684_ = pencrypt_0_ & new_n7683_;
  assign new_n7685_ = n_n2316 & new_n7684_;
  assign new_n7686_ = ~pstart_0_ & new_n7685_;
  assign new_n7687_ = ~new_n7682_ & ~new_n7686_;
  assign new_n7688_ = ~new_n7676_ & ~new_n7680_;
  assign new_n7689_ = new_n7687_ & new_n7688_;
  assign new_n7690_ = ~new_n7670_ & ~new_n7672_;
  assign new_n7691_ = ~new_n7664_ & ~new_n7666_;
  assign new_n7692_ = ~new_n7668_ & new_n7691_;
  assign new_n7693_ = new_n7690_ & new_n7692_;
  assign n1827 = ~new_n7689_ | ~new_n7693_;
  assign new_n7695_ = new_n1200_ & new_n4234_;
  assign new_n7696_ = ~pstart_0_ & new_n7695_;
  assign new_n7697_ = ~new_n1200_ & new_n4229_;
  assign new_n7698_ = ~pstart_0_ & new_n7697_;
  assign new_n7699_ = pkey_115_ & pencrypt_0_;
  assign new_n7700_ = pstart_0_ & new_n7699_;
  assign new_n7701_ = new_n1200_ & new_n4225_;
  assign new_n7702_ = ~pstart_0_ & new_n7701_;
  assign new_n7703_ = pkey_123_ & ~pencrypt_0_;
  assign new_n7704_ = pstart_0_ & new_n7703_;
  assign new_n7705_ = n_n2421 & new_n1220_;
  assign new_n7706_ = pencrypt_0_ & new_n7705_;
  assign new_n7707_ = ~n_n2802 & new_n7706_;
  assign new_n7708_ = ~pstart_0_ & new_n7707_;
  assign new_n7709_ = ~n_n2421 & new_n1220_;
  assign new_n7710_ = pencrypt_0_ & new_n7709_;
  assign new_n7711_ = n_n2802 & new_n7710_;
  assign new_n7712_ = ~pstart_0_ & new_n7711_;
  assign new_n7713_ = ~new_n1200_ & new_n4248_;
  assign new_n7714_ = ~pstart_0_ & new_n7713_;
  assign new_n7715_ = n_n2421 & ~new_n1220_;
  assign new_n7716_ = pencrypt_0_ & new_n7715_;
  assign new_n7717_ = n_n2802 & new_n7716_;
  assign new_n7718_ = ~pstart_0_ & new_n7717_;
  assign new_n7719_ = ~new_n7714_ & ~new_n7718_;
  assign new_n7720_ = ~new_n7708_ & ~new_n7712_;
  assign new_n7721_ = new_n7719_ & new_n7720_;
  assign new_n7722_ = ~new_n7702_ & ~new_n7704_;
  assign new_n7723_ = ~new_n7696_ & ~new_n7698_;
  assign new_n7724_ = ~new_n7700_ & new_n7723_;
  assign new_n7725_ = new_n7722_ & new_n7724_;
  assign n1832 = ~new_n7721_ | ~new_n7725_;
  assign new_n7727_ = new_n1200_ & new_n4854_;
  assign new_n7728_ = ~pstart_0_ & new_n7727_;
  assign new_n7729_ = ~new_n1200_ & new_n4849_;
  assign new_n7730_ = ~pstart_0_ & new_n7729_;
  assign new_n7731_ = pkey_122_ & pencrypt_0_;
  assign new_n7732_ = pstart_0_ & new_n7731_;
  assign new_n7733_ = new_n1200_ & new_n4845_;
  assign new_n7734_ = ~pstart_0_ & new_n7733_;
  assign new_n7735_ = ~pencrypt_0_ & pkey_65_;
  assign new_n7736_ = pstart_0_ & new_n7735_;
  assign new_n7737_ = n_n2430 & new_n1220_;
  assign new_n7738_ = pencrypt_0_ & new_n7737_;
  assign new_n7739_ = ~n_n2334 & new_n7738_;
  assign new_n7740_ = ~pstart_0_ & new_n7739_;
  assign new_n7741_ = ~n_n2430 & new_n1220_;
  assign new_n7742_ = pencrypt_0_ & new_n7741_;
  assign new_n7743_ = n_n2334 & new_n7742_;
  assign new_n7744_ = ~pstart_0_ & new_n7743_;
  assign new_n7745_ = ~new_n1200_ & new_n4868_;
  assign new_n7746_ = ~pstart_0_ & new_n7745_;
  assign new_n7747_ = n_n2430 & ~new_n1220_;
  assign new_n7748_ = pencrypt_0_ & new_n7747_;
  assign new_n7749_ = n_n2334 & new_n7748_;
  assign new_n7750_ = ~pstart_0_ & new_n7749_;
  assign new_n7751_ = ~new_n7746_ & ~new_n7750_;
  assign new_n7752_ = ~new_n7740_ & ~new_n7744_;
  assign new_n7753_ = new_n7751_ & new_n7752_;
  assign new_n7754_ = ~new_n7734_ & ~new_n7736_;
  assign new_n7755_ = ~new_n7728_ & ~new_n7730_;
  assign new_n7756_ = ~new_n7732_ & new_n7755_;
  assign new_n7757_ = new_n7754_ & new_n7756_;
  assign n1837 = ~new_n7753_ | ~new_n7757_;
  assign new_n7759_ = new_n1200_ & new_n5426_;
  assign new_n7760_ = ~pstart_0_ & new_n7759_;
  assign new_n7761_ = ~new_n1200_ & new_n5421_;
  assign new_n7762_ = ~pstart_0_ & new_n7761_;
  assign new_n7763_ = pkey_217_ & pencrypt_0_;
  assign new_n7764_ = pstart_0_ & new_n7763_;
  assign new_n7765_ = new_n1200_ & new_n5417_;
  assign new_n7766_ = ~pstart_0_ & new_n7765_;
  assign new_n7767_ = pkey_225_ & ~pencrypt_0_;
  assign new_n7768_ = pstart_0_ & new_n7767_;
  assign new_n7769_ = n_n2385 & new_n1220_;
  assign new_n7770_ = pencrypt_0_ & new_n7769_;
  assign new_n7771_ = ~n_n2290 & new_n7770_;
  assign new_n7772_ = ~pstart_0_ & new_n7771_;
  assign new_n7773_ = ~n_n2385 & new_n1220_;
  assign new_n7774_ = pencrypt_0_ & new_n7773_;
  assign new_n7775_ = n_n2290 & new_n7774_;
  assign new_n7776_ = ~pstart_0_ & new_n7775_;
  assign new_n7777_ = ~new_n1200_ & new_n5440_;
  assign new_n7778_ = ~pstart_0_ & new_n7777_;
  assign new_n7779_ = n_n2385 & ~new_n1220_;
  assign new_n7780_ = pencrypt_0_ & new_n7779_;
  assign new_n7781_ = n_n2290 & new_n7780_;
  assign new_n7782_ = ~pstart_0_ & new_n7781_;
  assign new_n7783_ = ~new_n7778_ & ~new_n7782_;
  assign new_n7784_ = ~new_n7772_ & ~new_n7776_;
  assign new_n7785_ = new_n7783_ & new_n7784_;
  assign new_n7786_ = ~new_n7766_ & ~new_n7768_;
  assign new_n7787_ = ~new_n7760_ & ~new_n7762_;
  assign new_n7788_ = ~new_n7764_ & new_n7787_;
  assign new_n7789_ = new_n7786_ & new_n7788_;
  assign n1842 = ~new_n7785_ | ~new_n7789_;
  assign new_n7791_ = new_n1200_ & new_n5464_;
  assign new_n7792_ = ~pstart_0_ & new_n7791_;
  assign new_n7793_ = ~new_n1200_ & new_n5459_;
  assign new_n7794_ = ~pstart_0_ & new_n7793_;
  assign new_n7795_ = pkey_240_ & pencrypt_0_;
  assign new_n7796_ = pstart_0_ & new_n7795_;
  assign new_n7797_ = new_n1200_ & new_n5455_;
  assign new_n7798_ = ~pstart_0_ & new_n7797_;
  assign new_n7799_ = pkey_248_ & ~pencrypt_0_;
  assign new_n7800_ = pstart_0_ & new_n7799_;
  assign new_n7801_ = n_n2394 & new_n1220_;
  assign new_n7802_ = pencrypt_0_ & new_n7801_;
  assign new_n7803_ = ~n_n2300 & new_n7802_;
  assign new_n7804_ = ~pstart_0_ & new_n7803_;
  assign new_n7805_ = ~n_n2394 & new_n1220_;
  assign new_n7806_ = pencrypt_0_ & new_n7805_;
  assign new_n7807_ = n_n2300 & new_n7806_;
  assign new_n7808_ = ~pstart_0_ & new_n7807_;
  assign new_n7809_ = ~new_n1200_ & new_n5478_;
  assign new_n7810_ = ~pstart_0_ & new_n7809_;
  assign new_n7811_ = n_n2394 & ~new_n1220_;
  assign new_n7812_ = pencrypt_0_ & new_n7811_;
  assign new_n7813_ = n_n2300 & new_n7812_;
  assign new_n7814_ = ~pstart_0_ & new_n7813_;
  assign new_n7815_ = ~new_n7810_ & ~new_n7814_;
  assign new_n7816_ = ~new_n7804_ & ~new_n7808_;
  assign new_n7817_ = new_n7815_ & new_n7816_;
  assign new_n7818_ = ~new_n7798_ & ~new_n7800_;
  assign new_n7819_ = ~new_n7792_ & ~new_n7794_;
  assign new_n7820_ = ~new_n7796_ & new_n7819_;
  assign new_n7821_ = new_n7818_ & new_n7820_;
  assign n1847 = ~new_n7817_ | ~new_n7821_;
  assign new_n7823_ = new_n1200_ & new_n5502_;
  assign new_n7824_ = ~pstart_0_ & new_n7823_;
  assign new_n7825_ = ~new_n1200_ & new_n5497_;
  assign new_n7826_ = ~pstart_0_ & new_n7825_;
  assign new_n7827_ = pkey_138_ & pencrypt_0_;
  assign new_n7828_ = pstart_0_ & new_n7827_;
  assign new_n7829_ = new_n1200_ & new_n5493_;
  assign new_n7830_ = ~pstart_0_ & new_n7829_;
  assign new_n7831_ = pkey_146_ & ~pencrypt_0_;
  assign new_n7832_ = pstart_0_ & new_n7831_;
  assign new_n7833_ = n_n2400 & new_n1220_;
  assign new_n7834_ = pencrypt_0_ & new_n7833_;
  assign new_n7835_ = ~n_n2774 & new_n7834_;
  assign new_n7836_ = ~pstart_0_ & new_n7835_;
  assign new_n7837_ = ~n_n2400 & new_n1220_;
  assign new_n7838_ = pencrypt_0_ & new_n7837_;
  assign new_n7839_ = n_n2774 & new_n7838_;
  assign new_n7840_ = ~pstart_0_ & new_n7839_;
  assign new_n7841_ = ~new_n1200_ & new_n5516_;
  assign new_n7842_ = ~pstart_0_ & new_n7841_;
  assign new_n7843_ = n_n2400 & ~new_n1220_;
  assign new_n7844_ = pencrypt_0_ & new_n7843_;
  assign new_n7845_ = n_n2774 & new_n7844_;
  assign new_n7846_ = ~pstart_0_ & new_n7845_;
  assign new_n7847_ = ~new_n7842_ & ~new_n7846_;
  assign new_n7848_ = ~new_n7836_ & ~new_n7840_;
  assign new_n7849_ = new_n7847_ & new_n7848_;
  assign new_n7850_ = ~new_n7830_ & ~new_n7832_;
  assign new_n7851_ = ~new_n7824_ & ~new_n7826_;
  assign new_n7852_ = ~new_n7828_ & new_n7851_;
  assign new_n7853_ = new_n7850_ & new_n7852_;
  assign n1852 = ~new_n7849_ | ~new_n7853_;
  assign new_n7855_ = new_n1200_ & new_n5540_;
  assign new_n7856_ = ~pstart_0_ & new_n7855_;
  assign new_n7857_ = ~new_n1200_ & new_n5535_;
  assign new_n7858_ = ~pstart_0_ & new_n7857_;
  assign new_n7859_ = pkey_161_ & pencrypt_0_;
  assign new_n7860_ = pstart_0_ & new_n7859_;
  assign new_n7861_ = new_n1200_ & new_n5531_;
  assign new_n7862_ = ~pstart_0_ & new_n7861_;
  assign new_n7863_ = pkey_169_ & ~pencrypt_0_;
  assign new_n7864_ = pstart_0_ & new_n7863_;
  assign new_n7865_ = n_n2410 & new_n1220_;
  assign new_n7866_ = pencrypt_0_ & new_n7865_;
  assign new_n7867_ = ~n_n2315 & new_n7866_;
  assign new_n7868_ = ~pstart_0_ & new_n7867_;
  assign new_n7869_ = ~n_n2410 & new_n1220_;
  assign new_n7870_ = pencrypt_0_ & new_n7869_;
  assign new_n7871_ = n_n2315 & new_n7870_;
  assign new_n7872_ = ~pstart_0_ & new_n7871_;
  assign new_n7873_ = ~new_n1200_ & new_n5554_;
  assign new_n7874_ = ~pstart_0_ & new_n7873_;
  assign new_n7875_ = n_n2410 & ~new_n1220_;
  assign new_n7876_ = pencrypt_0_ & new_n7875_;
  assign new_n7877_ = n_n2315 & new_n7876_;
  assign new_n7878_ = ~pstart_0_ & new_n7877_;
  assign new_n7879_ = ~new_n7874_ & ~new_n7878_;
  assign new_n7880_ = ~new_n7868_ & ~new_n7872_;
  assign new_n7881_ = new_n7879_ & new_n7880_;
  assign new_n7882_ = ~new_n7862_ & ~new_n7864_;
  assign new_n7883_ = ~new_n7856_ & ~new_n7858_;
  assign new_n7884_ = ~new_n7860_ & new_n7883_;
  assign new_n7885_ = new_n7882_ & new_n7884_;
  assign n1857 = ~new_n7881_ | ~new_n7885_;
  assign new_n7887_ = new_n1200_ & new_n5286_;
  assign new_n7888_ = ~pstart_0_ & new_n7887_;
  assign new_n7889_ = ~new_n1200_ & new_n5281_;
  assign new_n7890_ = ~pstart_0_ & new_n7889_;
  assign new_n7891_ = pencrypt_0_ & pkey_72_;
  assign new_n7892_ = pstart_0_ & new_n7891_;
  assign new_n7893_ = new_n1200_ & new_n5277_;
  assign new_n7894_ = ~pstart_0_ & new_n7893_;
  assign new_n7895_ = pkey_80_ & ~pencrypt_0_;
  assign new_n7896_ = pstart_0_ & new_n7895_;
  assign new_n7897_ = n_n2436 & new_n1220_;
  assign new_n7898_ = pencrypt_0_ & new_n7897_;
  assign new_n7899_ = ~n_n2343 & new_n7898_;
  assign new_n7900_ = ~pstart_0_ & new_n7899_;
  assign new_n7901_ = ~n_n2436 & new_n1220_;
  assign new_n7902_ = pencrypt_0_ & new_n7901_;
  assign new_n7903_ = n_n2343 & new_n7902_;
  assign new_n7904_ = ~pstart_0_ & new_n7903_;
  assign new_n7905_ = ~new_n1200_ & new_n5300_;
  assign new_n7906_ = ~pstart_0_ & new_n7905_;
  assign new_n7907_ = n_n2436 & ~new_n1220_;
  assign new_n7908_ = pencrypt_0_ & new_n7907_;
  assign new_n7909_ = n_n2343 & new_n7908_;
  assign new_n7910_ = ~pstart_0_ & new_n7909_;
  assign new_n7911_ = ~new_n7906_ & ~new_n7910_;
  assign new_n7912_ = ~new_n7900_ & ~new_n7904_;
  assign new_n7913_ = new_n7911_ & new_n7912_;
  assign new_n7914_ = ~new_n7894_ & ~new_n7896_;
  assign new_n7915_ = ~new_n7888_ & ~new_n7890_;
  assign new_n7916_ = ~new_n7892_ & new_n7915_;
  assign new_n7917_ = new_n7914_ & new_n7916_;
  assign n1862 = ~new_n7913_ | ~new_n7917_;
  assign new_n7919_ = new_n1200_ & new_n3236_;
  assign new_n7920_ = ~pstart_0_ & new_n7919_;
  assign new_n7921_ = ~new_n1200_ & new_n3231_;
  assign new_n7922_ = ~pstart_0_ & new_n7921_;
  assign new_n7923_ = pkey_2_ & pencrypt_0_;
  assign new_n7924_ = pstart_0_ & new_n7923_;
  assign new_n7925_ = new_n1200_ & new_n3227_;
  assign new_n7926_ = ~pstart_0_ & new_n7925_;
  assign new_n7927_ = ~pencrypt_0_ & pkey_10_;
  assign new_n7928_ = pstart_0_ & new_n7927_;
  assign new_n7929_ = n_n2446 & new_n1220_;
  assign new_n7930_ = pencrypt_0_ & new_n7929_;
  assign new_n7931_ = ~n_n2353 & new_n7930_;
  assign new_n7932_ = ~pstart_0_ & new_n7931_;
  assign new_n7933_ = ~n_n2446 & new_n1220_;
  assign new_n7934_ = pencrypt_0_ & new_n7933_;
  assign new_n7935_ = n_n2353 & new_n7934_;
  assign new_n7936_ = ~pstart_0_ & new_n7935_;
  assign new_n7937_ = ~new_n1200_ & new_n3250_;
  assign new_n7938_ = ~pstart_0_ & new_n7937_;
  assign new_n7939_ = n_n2446 & ~new_n1220_;
  assign new_n7940_ = pencrypt_0_ & new_n7939_;
  assign new_n7941_ = n_n2353 & new_n7940_;
  assign new_n7942_ = ~pstart_0_ & new_n7941_;
  assign new_n7943_ = ~new_n7938_ & ~new_n7942_;
  assign new_n7944_ = ~new_n7932_ & ~new_n7936_;
  assign new_n7945_ = new_n7943_ & new_n7944_;
  assign new_n7946_ = ~new_n7926_ & ~new_n7928_;
  assign new_n7947_ = ~new_n7920_ & ~new_n7922_;
  assign new_n7948_ = ~new_n7924_ & new_n7947_;
  assign new_n7949_ = new_n7946_ & new_n7948_;
  assign n1867 = ~new_n7945_ | ~new_n7949_;
  assign new_n7951_ = new_n1200_ & new_n5800_;
  assign new_n7952_ = ~pstart_0_ & new_n7951_;
  assign new_n7953_ = ~new_n1200_ & new_n5795_;
  assign new_n7954_ = ~pstart_0_ & new_n7953_;
  assign new_n7955_ = pkey_225_ & pencrypt_0_;
  assign new_n7956_ = pstart_0_ & new_n7955_;
  assign new_n7957_ = new_n1200_ & new_n5791_;
  assign new_n7958_ = ~pstart_0_ & new_n7957_;
  assign new_n7959_ = pkey_233_ & ~pencrypt_0_;
  assign new_n7960_ = pstart_0_ & new_n7959_;
  assign new_n7961_ = n_n2386 & new_n1220_;
  assign new_n7962_ = pencrypt_0_ & new_n7961_;
  assign new_n7963_ = ~n_n2291 & new_n7962_;
  assign new_n7964_ = ~pstart_0_ & new_n7963_;
  assign new_n7965_ = ~n_n2386 & new_n1220_;
  assign new_n7966_ = pencrypt_0_ & new_n7965_;
  assign new_n7967_ = n_n2291 & new_n7966_;
  assign new_n7968_ = ~pstart_0_ & new_n7967_;
  assign new_n7969_ = ~new_n1200_ & new_n5814_;
  assign new_n7970_ = ~pstart_0_ & new_n7969_;
  assign new_n7971_ = n_n2386 & ~new_n1220_;
  assign new_n7972_ = pencrypt_0_ & new_n7971_;
  assign new_n7973_ = n_n2291 & new_n7972_;
  assign new_n7974_ = ~pstart_0_ & new_n7973_;
  assign new_n7975_ = ~new_n7970_ & ~new_n7974_;
  assign new_n7976_ = ~new_n7964_ & ~new_n7968_;
  assign new_n7977_ = new_n7975_ & new_n7976_;
  assign new_n7978_ = ~new_n7958_ & ~new_n7960_;
  assign new_n7979_ = ~new_n7952_ & ~new_n7954_;
  assign new_n7980_ = ~new_n7956_ & new_n7979_;
  assign new_n7981_ = new_n7978_ & new_n7980_;
  assign n1872 = ~new_n7977_ | ~new_n7981_;
  assign new_n7983_ = new_n1200_ & new_n5838_;
  assign new_n7984_ = ~pstart_0_ & new_n7983_;
  assign new_n7985_ = ~new_n1200_ & new_n5833_;
  assign new_n7986_ = ~pstart_0_ & new_n7985_;
  assign new_n7987_ = pkey_232_ & pencrypt_0_;
  assign new_n7988_ = pstart_0_ & new_n7987_;
  assign new_n7989_ = new_n1200_ & new_n5829_;
  assign new_n7990_ = ~pstart_0_ & new_n7989_;
  assign new_n7991_ = pkey_240_ & ~pencrypt_0_;
  assign new_n7992_ = pstart_0_ & new_n7991_;
  assign new_n7993_ = n_n2393 & new_n1220_;
  assign new_n7994_ = pencrypt_0_ & new_n7993_;
  assign new_n7995_ = ~n_n2299 & new_n7994_;
  assign new_n7996_ = ~pstart_0_ & new_n7995_;
  assign new_n7997_ = ~n_n2393 & new_n1220_;
  assign new_n7998_ = pencrypt_0_ & new_n7997_;
  assign new_n7999_ = n_n2299 & new_n7998_;
  assign new_n8000_ = ~pstart_0_ & new_n7999_;
  assign new_n8001_ = ~new_n1200_ & new_n5852_;
  assign new_n8002_ = ~pstart_0_ & new_n8001_;
  assign new_n8003_ = n_n2393 & ~new_n1220_;
  assign new_n8004_ = pencrypt_0_ & new_n8003_;
  assign new_n8005_ = n_n2299 & new_n8004_;
  assign new_n8006_ = ~pstart_0_ & new_n8005_;
  assign new_n8007_ = ~new_n8002_ & ~new_n8006_;
  assign new_n8008_ = ~new_n7996_ & ~new_n8000_;
  assign new_n8009_ = new_n8007_ & new_n8008_;
  assign new_n8010_ = ~new_n7990_ & ~new_n7992_;
  assign new_n8011_ = ~new_n7984_ & ~new_n7986_;
  assign new_n8012_ = ~new_n7988_ & new_n8011_;
  assign new_n8013_ = new_n8010_ & new_n8012_;
  assign n1877 = ~new_n8009_ | ~new_n8013_;
  assign new_n8015_ = new_n1200_ & new_n5876_;
  assign new_n8016_ = ~pstart_0_ & new_n8015_;
  assign new_n8017_ = ~new_n1200_ & new_n5871_;
  assign new_n8018_ = ~pstart_0_ & new_n8017_;
  assign new_n8019_ = pkey_146_ & pencrypt_0_;
  assign new_n8020_ = pstart_0_ & new_n8019_;
  assign new_n8021_ = new_n1200_ & new_n5867_;
  assign new_n8022_ = ~pstart_0_ & new_n8021_;
  assign new_n8023_ = pkey_154_ & ~pencrypt_0_;
  assign new_n8024_ = pstart_0_ & new_n8023_;
  assign new_n8025_ = n_n2401 & new_n1220_;
  assign new_n8026_ = pencrypt_0_ & new_n8025_;
  assign new_n8027_ = ~n_n2306 & new_n8026_;
  assign new_n8028_ = ~pstart_0_ & new_n8027_;
  assign new_n8029_ = ~n_n2401 & new_n1220_;
  assign new_n8030_ = pencrypt_0_ & new_n8029_;
  assign new_n8031_ = n_n2306 & new_n8030_;
  assign new_n8032_ = ~pstart_0_ & new_n8031_;
  assign new_n8033_ = ~new_n1200_ & new_n5890_;
  assign new_n8034_ = ~pstart_0_ & new_n8033_;
  assign new_n8035_ = n_n2401 & ~new_n1220_;
  assign new_n8036_ = pencrypt_0_ & new_n8035_;
  assign new_n8037_ = n_n2306 & new_n8036_;
  assign new_n8038_ = ~pstart_0_ & new_n8037_;
  assign new_n8039_ = ~new_n8034_ & ~new_n8038_;
  assign new_n8040_ = ~new_n8028_ & ~new_n8032_;
  assign new_n8041_ = new_n8039_ & new_n8040_;
  assign new_n8042_ = ~new_n8022_ & ~new_n8024_;
  assign new_n8043_ = ~new_n8016_ & ~new_n8018_;
  assign new_n8044_ = ~new_n8020_ & new_n8043_;
  assign new_n8045_ = new_n8042_ & new_n8044_;
  assign n1882 = ~new_n8041_ | ~new_n8045_;
  assign new_n8047_ = new_n1200_ & new_n5914_;
  assign new_n8048_ = ~pstart_0_ & new_n8047_;
  assign new_n8049_ = ~new_n1200_ & new_n5909_;
  assign new_n8050_ = ~pstart_0_ & new_n8049_;
  assign new_n8051_ = pkey_153_ & pencrypt_0_;
  assign new_n8052_ = pstart_0_ & new_n8051_;
  assign new_n8053_ = new_n1200_ & new_n5905_;
  assign new_n8054_ = ~pstart_0_ & new_n8053_;
  assign new_n8055_ = pkey_161_ & ~pencrypt_0_;
  assign new_n8056_ = pstart_0_ & new_n8055_;
  assign new_n8057_ = n_n2409 & new_n1220_;
  assign new_n8058_ = pencrypt_0_ & new_n8057_;
  assign new_n8059_ = ~n_n2314 & new_n8058_;
  assign new_n8060_ = ~pstart_0_ & new_n8059_;
  assign new_n8061_ = ~n_n2409 & new_n1220_;
  assign new_n8062_ = pencrypt_0_ & new_n8061_;
  assign new_n8063_ = n_n2314 & new_n8062_;
  assign new_n8064_ = ~pstart_0_ & new_n8063_;
  assign new_n8065_ = ~new_n1200_ & new_n5928_;
  assign new_n8066_ = ~pstart_0_ & new_n8065_;
  assign new_n8067_ = n_n2409 & ~new_n1220_;
  assign new_n8068_ = pencrypt_0_ & new_n8067_;
  assign new_n8069_ = n_n2314 & new_n8068_;
  assign new_n8070_ = ~pstart_0_ & new_n8069_;
  assign new_n8071_ = ~new_n8066_ & ~new_n8070_;
  assign new_n8072_ = ~new_n8060_ & ~new_n8064_;
  assign new_n8073_ = new_n8071_ & new_n8072_;
  assign new_n8074_ = ~new_n8054_ & ~new_n8056_;
  assign new_n8075_ = ~new_n8048_ & ~new_n8050_;
  assign new_n8076_ = ~new_n8052_ & new_n8075_;
  assign new_n8077_ = new_n8074_ & new_n8076_;
  assign n1887 = ~new_n8073_ | ~new_n8077_;
  assign new_n8079_ = new_n1200_ & new_n4892_;
  assign new_n8080_ = ~pstart_0_ & new_n8079_;
  assign new_n8081_ = ~new_n1200_ & new_n4887_;
  assign new_n8082_ = ~pstart_0_ & new_n8081_;
  assign new_n8083_ = pkey_80_ & pencrypt_0_;
  assign new_n8084_ = pstart_0_ & new_n8083_;
  assign new_n8085_ = new_n1200_ & new_n4883_;
  assign new_n8086_ = ~pstart_0_ & new_n8085_;
  assign new_n8087_ = pkey_88_ & ~pencrypt_0_;
  assign new_n8088_ = pstart_0_ & new_n8087_;
  assign new_n8089_ = n_n2437 & new_n1220_;
  assign new_n8090_ = pencrypt_0_ & new_n8089_;
  assign new_n8091_ = ~n_n2344 & new_n8090_;
  assign new_n8092_ = ~pstart_0_ & new_n8091_;
  assign new_n8093_ = ~n_n2437 & new_n1220_;
  assign new_n8094_ = pencrypt_0_ & new_n8093_;
  assign new_n8095_ = n_n2344 & new_n8094_;
  assign new_n8096_ = ~pstart_0_ & new_n8095_;
  assign new_n8097_ = ~new_n1200_ & new_n4906_;
  assign new_n8098_ = ~pstart_0_ & new_n8097_;
  assign new_n8099_ = n_n2437 & ~new_n1220_;
  assign new_n8100_ = pencrypt_0_ & new_n8099_;
  assign new_n8101_ = n_n2344 & new_n8100_;
  assign new_n8102_ = ~pstart_0_ & new_n8101_;
  assign new_n8103_ = ~new_n8098_ & ~new_n8102_;
  assign new_n8104_ = ~new_n8092_ & ~new_n8096_;
  assign new_n8105_ = new_n8103_ & new_n8104_;
  assign new_n8106_ = ~new_n8086_ & ~new_n8088_;
  assign new_n8107_ = ~new_n8080_ & ~new_n8082_;
  assign new_n8108_ = ~new_n8084_ & new_n8107_;
  assign new_n8109_ = new_n8106_ & new_n8108_;
  assign n1892 = ~new_n8105_ | ~new_n8109_;
  assign new_n8111_ = new_n1200_ & new_n3020_;
  assign new_n8112_ = ~pstart_0_ & new_n8111_;
  assign new_n8113_ = ~new_n1200_ & new_n3015_;
  assign new_n8114_ = ~pstart_0_ & new_n8113_;
  assign new_n8115_ = pkey_59_ & pencrypt_0_;
  assign new_n8116_ = pstart_0_ & new_n8115_;
  assign new_n8117_ = new_n1200_ & new_n3011_;
  assign new_n8118_ = ~pstart_0_ & new_n8117_;
  assign new_n8119_ = pkey_2_ & ~pencrypt_0_;
  assign new_n8120_ = pstart_0_ & new_n8119_;
  assign new_n8121_ = n_n2445 & new_n1220_;
  assign new_n8122_ = pencrypt_0_ & new_n8121_;
  assign new_n8123_ = ~n_n2352 & new_n8122_;
  assign new_n8124_ = ~pstart_0_ & new_n8123_;
  assign new_n8125_ = ~n_n2445 & new_n1220_;
  assign new_n8126_ = pencrypt_0_ & new_n8125_;
  assign new_n8127_ = n_n2352 & new_n8126_;
  assign new_n8128_ = ~pstart_0_ & new_n8127_;
  assign new_n8129_ = ~new_n1200_ & new_n3034_;
  assign new_n8130_ = ~pstart_0_ & new_n8129_;
  assign new_n8131_ = n_n2445 & ~new_n1220_;
  assign new_n8132_ = pencrypt_0_ & new_n8131_;
  assign new_n8133_ = n_n2352 & new_n8132_;
  assign new_n8134_ = ~pstart_0_ & new_n8133_;
  assign new_n8135_ = ~new_n8130_ & ~new_n8134_;
  assign new_n8136_ = ~new_n8124_ & ~new_n8128_;
  assign new_n8137_ = new_n8135_ & new_n8136_;
  assign new_n8138_ = ~new_n8118_ & ~new_n8120_;
  assign new_n8139_ = ~new_n8112_ & ~new_n8114_;
  assign new_n8140_ = ~new_n8116_ & new_n8139_;
  assign new_n8141_ = new_n8138_ & new_n8140_;
  assign n1897 = ~new_n8137_ | ~new_n8141_;
  assign new_n8143_ = new_n1200_ & new_n3406_;
  assign new_n8144_ = ~pstart_0_ & new_n8143_;
  assign new_n8145_ = ~new_n1200_ & new_n3401_;
  assign new_n8146_ = ~pstart_0_ & new_n8145_;
  assign new_n8147_ = pkey_233_ & pencrypt_0_;
  assign new_n8148_ = pstart_0_ & new_n8147_;
  assign new_n8149_ = new_n1200_ & new_n3397_;
  assign new_n8150_ = ~pstart_0_ & new_n8149_;
  assign new_n8151_ = pkey_241_ & ~pencrypt_0_;
  assign new_n8152_ = pstart_0_ & new_n8151_;
  assign new_n8153_ = n_n2885 & new_n1220_;
  assign new_n8154_ = pencrypt_0_ & new_n8153_;
  assign new_n8155_ = ~n_n2292 & new_n8154_;
  assign new_n8156_ = ~pstart_0_ & new_n8155_;
  assign new_n8157_ = ~n_n2885 & new_n1220_;
  assign new_n8158_ = pencrypt_0_ & new_n8157_;
  assign new_n8159_ = n_n2292 & new_n8158_;
  assign new_n8160_ = ~pstart_0_ & new_n8159_;
  assign new_n8161_ = ~new_n1200_ & new_n3420_;
  assign new_n8162_ = ~pstart_0_ & new_n8161_;
  assign new_n8163_ = n_n2885 & ~new_n1220_;
  assign new_n8164_ = pencrypt_0_ & new_n8163_;
  assign new_n8165_ = n_n2292 & new_n8164_;
  assign new_n8166_ = ~pstart_0_ & new_n8165_;
  assign new_n8167_ = ~new_n8162_ & ~new_n8166_;
  assign new_n8168_ = ~new_n8156_ & ~new_n8160_;
  assign new_n8169_ = new_n8167_ & new_n8168_;
  assign new_n8170_ = ~new_n8150_ & ~new_n8152_;
  assign new_n8171_ = ~new_n8144_ & ~new_n8146_;
  assign new_n8172_ = ~new_n8148_ & new_n8171_;
  assign new_n8173_ = new_n8170_ & new_n8172_;
  assign n1902 = ~new_n8169_ | ~new_n8173_;
  assign new_n8175_ = new_n1200_ & new_n3856_;
  assign new_n8176_ = ~pstart_0_ & new_n8175_;
  assign new_n8177_ = ~new_n1200_ & new_n3851_;
  assign new_n8178_ = ~pstart_0_ & new_n8177_;
  assign new_n8179_ = pkey_163_ & pencrypt_0_;
  assign new_n8180_ = pstart_0_ & new_n8179_;
  assign new_n8181_ = new_n1200_ & new_n3847_;
  assign new_n8182_ = ~pstart_0_ & new_n8181_;
  assign new_n8183_ = pkey_171_ & ~pencrypt_0_;
  assign new_n8184_ = pstart_0_ & new_n8183_;
  assign new_n8185_ = n_n2396 & new_n1220_;
  assign new_n8186_ = pencrypt_0_ & new_n8185_;
  assign new_n8187_ = ~n_n2302 & new_n8186_;
  assign new_n8188_ = ~pstart_0_ & new_n8187_;
  assign new_n8189_ = ~n_n2396 & new_n1220_;
  assign new_n8190_ = pencrypt_0_ & new_n8189_;
  assign new_n8191_ = n_n2302 & new_n8190_;
  assign new_n8192_ = ~pstart_0_ & new_n8191_;
  assign new_n8193_ = ~new_n1200_ & new_n3870_;
  assign new_n8194_ = ~pstart_0_ & new_n8193_;
  assign new_n8195_ = n_n2396 & ~new_n1220_;
  assign new_n8196_ = pencrypt_0_ & new_n8195_;
  assign new_n8197_ = n_n2302 & new_n8196_;
  assign new_n8198_ = ~pstart_0_ & new_n8197_;
  assign new_n8199_ = ~new_n8194_ & ~new_n8198_;
  assign new_n8200_ = ~new_n8188_ & ~new_n8192_;
  assign new_n8201_ = new_n8199_ & new_n8200_;
  assign new_n8202_ = ~new_n8182_ & ~new_n8184_;
  assign new_n8203_ = ~new_n8176_ & ~new_n8178_;
  assign new_n8204_ = ~new_n8180_ & new_n8203_;
  assign new_n8205_ = new_n8202_ & new_n8204_;
  assign n1907 = ~new_n8201_ | ~new_n8205_;
  assign new_n8207_ = new_n1200_ & new_n4780_;
  assign new_n8208_ = ~pstart_0_ & new_n8207_;
  assign new_n8209_ = ~new_n1200_ & new_n4775_;
  assign new_n8210_ = ~pstart_0_ & new_n8209_;
  assign new_n8211_ = pkey_168_ & pencrypt_0_;
  assign new_n8212_ = pstart_0_ & new_n8211_;
  assign new_n8213_ = new_n1200_ & new_n4771_;
  assign new_n8214_ = ~pstart_0_ & new_n8213_;
  assign new_n8215_ = ~pencrypt_0_ & pkey_176_;
  assign new_n8216_ = pstart_0_ & new_n8215_;
  assign new_n8217_ = n_n2417 & new_n1220_;
  assign new_n8218_ = pencrypt_0_ & new_n8217_;
  assign new_n8219_ = ~n_n2323 & new_n8218_;
  assign new_n8220_ = ~pstart_0_ & new_n8219_;
  assign new_n8221_ = ~n_n2417 & new_n1220_;
  assign new_n8222_ = pencrypt_0_ & new_n8221_;
  assign new_n8223_ = n_n2323 & new_n8222_;
  assign new_n8224_ = ~pstart_0_ & new_n8223_;
  assign new_n8225_ = ~new_n1200_ & new_n4794_;
  assign new_n8226_ = ~pstart_0_ & new_n8225_;
  assign new_n8227_ = n_n2417 & ~new_n1220_;
  assign new_n8228_ = pencrypt_0_ & new_n8227_;
  assign new_n8229_ = n_n2323 & new_n8228_;
  assign new_n8230_ = ~pstart_0_ & new_n8229_;
  assign new_n8231_ = ~new_n8226_ & ~new_n8230_;
  assign new_n8232_ = ~new_n8220_ & ~new_n8224_;
  assign new_n8233_ = new_n8231_ & new_n8232_;
  assign new_n8234_ = ~new_n8214_ & ~new_n8216_;
  assign new_n8235_ = ~new_n8208_ & ~new_n8210_;
  assign new_n8236_ = ~new_n8212_ & new_n8235_;
  assign new_n8237_ = new_n8234_ & new_n8236_;
  assign n1912 = ~new_n8233_ | ~new_n8237_;
  assign new_n8239_ = new_n1200_ & new_n4818_;
  assign new_n8240_ = ~pstart_0_ & new_n8239_;
  assign new_n8241_ = ~new_n1200_ & new_n4813_;
  assign new_n8242_ = ~pstart_0_ & new_n8241_;
  assign new_n8243_ = pkey_98_ & pencrypt_0_;
  assign new_n8244_ = pstart_0_ & new_n8243_;
  assign new_n8245_ = new_n1200_ & new_n4809_;
  assign new_n8246_ = ~pstart_0_ & new_n8245_;
  assign new_n8247_ = ~pencrypt_0_ & pkey_106_;
  assign new_n8248_ = pstart_0_ & new_n8247_;
  assign new_n8249_ = n_n2427 & new_n1220_;
  assign new_n8250_ = pencrypt_0_ & new_n8249_;
  assign new_n8251_ = ~n_n2332 & new_n8250_;
  assign new_n8252_ = ~pstart_0_ & new_n8251_;
  assign new_n8253_ = ~n_n2427 & new_n1220_;
  assign new_n8254_ = pencrypt_0_ & new_n8253_;
  assign new_n8255_ = n_n2332 & new_n8254_;
  assign new_n8256_ = ~pstart_0_ & new_n8255_;
  assign new_n8257_ = ~new_n1200_ & new_n4830_;
  assign new_n8258_ = ~pstart_0_ & new_n8257_;
  assign new_n8259_ = n_n2427 & ~new_n1220_;
  assign new_n8260_ = pencrypt_0_ & new_n8259_;
  assign new_n8261_ = n_n2332 & new_n8260_;
  assign new_n8262_ = ~pstart_0_ & new_n8261_;
  assign new_n8263_ = ~new_n8258_ & ~new_n8262_;
  assign new_n8264_ = ~new_n8252_ & ~new_n8256_;
  assign new_n8265_ = new_n8263_ & new_n8264_;
  assign new_n8266_ = ~new_n8246_ & ~new_n8248_;
  assign new_n8267_ = ~new_n8240_ & ~new_n8242_;
  assign new_n8268_ = ~new_n8244_ & new_n8267_;
  assign new_n8269_ = new_n8266_ & new_n8268_;
  assign n1917 = ~new_n8265_ | ~new_n8269_;
  assign new_n8271_ = new_n1200_ & new_n2646_;
  assign new_n8272_ = ~pstart_0_ & new_n8271_;
  assign new_n8273_ = ~new_n1200_ & new_n2641_;
  assign new_n8274_ = ~pstart_0_ & new_n8273_;
  assign new_n8275_ = pkey_121_ & pencrypt_0_;
  assign new_n8276_ = pstart_0_ & new_n8275_;
  assign new_n8277_ = new_n1200_ & new_n2637_;
  assign new_n8278_ = ~pstart_0_ & new_n8277_;
  assign new_n8279_ = ~pencrypt_0_ & pkey_64_;
  assign new_n8280_ = pstart_0_ & new_n8279_;
  assign new_n8281_ = n_n2435 & new_n1220_;
  assign new_n8282_ = pencrypt_0_ & new_n8281_;
  assign new_n8283_ = ~n_n2341 & new_n8282_;
  assign new_n8284_ = ~pstart_0_ & new_n8283_;
  assign new_n8285_ = ~n_n2435 & new_n1220_;
  assign new_n8286_ = pencrypt_0_ & new_n8285_;
  assign new_n8287_ = n_n2341 & new_n8286_;
  assign new_n8288_ = ~pstart_0_ & new_n8287_;
  assign new_n8289_ = ~new_n1200_ & new_n2660_;
  assign new_n8290_ = ~pstart_0_ & new_n8289_;
  assign new_n8291_ = n_n2435 & ~new_n1220_;
  assign new_n8292_ = pencrypt_0_ & new_n8291_;
  assign new_n8293_ = n_n2341 & new_n8292_;
  assign new_n8294_ = ~pstart_0_ & new_n8293_;
  assign new_n8295_ = ~new_n8290_ & ~new_n8294_;
  assign new_n8296_ = ~new_n8284_ & ~new_n8288_;
  assign new_n8297_ = new_n8295_ & new_n8296_;
  assign new_n8298_ = ~new_n8278_ & ~new_n8280_;
  assign new_n8299_ = ~new_n8272_ & ~new_n8274_;
  assign new_n8300_ = ~new_n8276_ & new_n8299_;
  assign new_n8301_ = new_n8298_ & new_n8300_;
  assign n1922 = ~new_n8297_ | ~new_n8301_;
  assign new_n8303_ = new_n1200_ & new_n2684_;
  assign new_n8304_ = ~pstart_0_ & new_n8303_;
  assign new_n8305_ = ~new_n1200_ & new_n2679_;
  assign new_n8306_ = ~pstart_0_ & new_n8305_;
  assign new_n8307_ = pkey_51_ & pencrypt_0_;
  assign new_n8308_ = pstart_0_ & new_n8307_;
  assign new_n8309_ = new_n1200_ & new_n2675_;
  assign new_n8310_ = ~pstart_0_ & new_n8309_;
  assign new_n8311_ = pkey_59_ & ~pencrypt_0_;
  assign new_n8312_ = pstart_0_ & new_n8311_;
  assign new_n8313_ = n_n2444 & new_n1220_;
  assign new_n8314_ = pencrypt_0_ & new_n8313_;
  assign new_n8315_ = ~n_n2834 & new_n8314_;
  assign new_n8316_ = ~pstart_0_ & new_n8315_;
  assign new_n8317_ = ~n_n2444 & new_n1220_;
  assign new_n8318_ = pencrypt_0_ & new_n8317_;
  assign new_n8319_ = n_n2834 & new_n8318_;
  assign new_n8320_ = ~pstart_0_ & new_n8319_;
  assign new_n8321_ = ~new_n1200_ & new_n2698_;
  assign new_n8322_ = ~pstart_0_ & new_n8321_;
  assign new_n8323_ = n_n2444 & ~new_n1220_;
  assign new_n8324_ = pencrypt_0_ & new_n8323_;
  assign new_n8325_ = n_n2834 & new_n8324_;
  assign new_n8326_ = ~pstart_0_ & new_n8325_;
  assign new_n8327_ = ~new_n8322_ & ~new_n8326_;
  assign new_n8328_ = ~new_n8316_ & ~new_n8320_;
  assign new_n8329_ = new_n8327_ & new_n8328_;
  assign new_n8330_ = ~new_n8310_ & ~new_n8312_;
  assign new_n8331_ = ~new_n8304_ & ~new_n8306_;
  assign new_n8332_ = ~new_n8308_ & new_n8331_;
  assign new_n8333_ = new_n8330_ & new_n8332_;
  assign n1927 = ~new_n8329_ | ~new_n8333_;
  assign new_n8335_ = new_n1200_ & new_n3444_;
  assign new_n8336_ = ~pstart_0_ & new_n8335_;
  assign new_n8337_ = ~new_n1200_ & new_n3439_;
  assign new_n8338_ = ~pstart_0_ & new_n8337_;
  assign new_n8339_ = pencrypt_0_ & pkey_10_;
  assign new_n8340_ = pstart_0_ & new_n8339_;
  assign new_n8341_ = new_n1200_ & new_n3435_;
  assign new_n8342_ = ~pstart_0_ & new_n8341_;
  assign new_n8343_ = pkey_18_ & ~pencrypt_0_;
  assign new_n8344_ = pstart_0_ & new_n8343_;
  assign new_n8345_ = n_n2447 & new_n1220_;
  assign new_n8346_ = pencrypt_0_ & new_n8345_;
  assign new_n8347_ = ~n_n2838 & new_n8346_;
  assign new_n8348_ = ~pstart_0_ & new_n8347_;
  assign new_n8349_ = ~n_n2447 & new_n1220_;
  assign new_n8350_ = pencrypt_0_ & new_n8349_;
  assign new_n8351_ = n_n2838 & new_n8350_;
  assign new_n8352_ = ~pstart_0_ & new_n8351_;
  assign new_n8353_ = ~new_n1200_ & new_n3458_;
  assign new_n8354_ = ~pstart_0_ & new_n8353_;
  assign new_n8355_ = n_n2447 & ~new_n1220_;
  assign new_n8356_ = pencrypt_0_ & new_n8355_;
  assign new_n8357_ = n_n2838 & new_n8356_;
  assign new_n8358_ = ~pstart_0_ & new_n8357_;
  assign new_n8359_ = ~new_n8354_ & ~new_n8358_;
  assign new_n8360_ = ~new_n8348_ & ~new_n8352_;
  assign new_n8361_ = new_n8359_ & new_n8360_;
  assign new_n8362_ = ~new_n8342_ & ~new_n8344_;
  assign new_n8363_ = ~new_n8336_ & ~new_n8338_;
  assign new_n8364_ = ~new_n8340_ & new_n8363_;
  assign new_n8365_ = new_n8362_ & new_n8364_;
  assign n1932 = ~new_n8361_ | ~new_n8365_;
  assign new_n8367_ = new_n1200_ & new_n3198_;
  assign new_n8368_ = ~pstart_0_ & new_n8367_;
  assign new_n8369_ = ~new_n1200_ & new_n3193_;
  assign new_n8370_ = ~pstart_0_ & new_n8369_;
  assign new_n8371_ = pkey_241_ & pencrypt_0_;
  assign new_n8372_ = pstart_0_ & new_n8371_;
  assign new_n8373_ = new_n1200_ & new_n3189_;
  assign new_n8374_ = ~pstart_0_ & new_n8373_;
  assign new_n8375_ = pkey_249_ & ~pencrypt_0_;
  assign new_n8376_ = pstart_0_ & new_n8375_;
  assign new_n8377_ = n_n2387 & new_n1220_;
  assign new_n8378_ = pencrypt_0_ & new_n8377_;
  assign new_n8379_ = ~n_n2757 & new_n8378_;
  assign new_n8380_ = ~pstart_0_ & new_n8379_;
  assign new_n8381_ = ~n_n2387 & new_n1220_;
  assign new_n8382_ = pencrypt_0_ & new_n8381_;
  assign new_n8383_ = n_n2757 & new_n8382_;
  assign new_n8384_ = ~pstart_0_ & new_n8383_;
  assign new_n8385_ = ~new_n1200_ & new_n3212_;
  assign new_n8386_ = ~pstart_0_ & new_n8385_;
  assign new_n8387_ = n_n2387 & ~new_n1220_;
  assign new_n8388_ = pencrypt_0_ & new_n8387_;
  assign new_n8389_ = n_n2757 & new_n8388_;
  assign new_n8390_ = ~pstart_0_ & new_n8389_;
  assign new_n8391_ = ~new_n8386_ & ~new_n8390_;
  assign new_n8392_ = ~new_n8380_ & ~new_n8384_;
  assign new_n8393_ = new_n8391_ & new_n8392_;
  assign new_n8394_ = ~new_n8374_ & ~new_n8376_;
  assign new_n8395_ = ~new_n8368_ & ~new_n8370_;
  assign new_n8396_ = ~new_n8372_ & new_n8395_;
  assign new_n8397_ = new_n8394_ & new_n8396_;
  assign n1937 = ~new_n8393_ | ~new_n8397_;
  assign new_n8399_ = new_n1200_ & new_n3590_;
  assign new_n8400_ = ~pstart_0_ & new_n8399_;
  assign new_n8401_ = ~new_n1200_ & new_n3585_;
  assign new_n8402_ = ~pstart_0_ & new_n8401_;
  assign new_n8403_ = pkey_248_ & pencrypt_0_;
  assign new_n8404_ = pstart_0_ & new_n8403_;
  assign new_n8405_ = new_n1200_ & new_n3581_;
  assign new_n8406_ = ~pstart_0_ & new_n8405_;
  assign new_n8407_ = pkey_163_ & ~pencrypt_0_;
  assign new_n8408_ = pstart_0_ & new_n8407_;
  assign new_n8409_ = n_n2395 & new_n1220_;
  assign new_n8410_ = pencrypt_0_ & new_n8409_;
  assign new_n8411_ = ~n_n2301 & new_n8410_;
  assign new_n8412_ = ~pstart_0_ & new_n8411_;
  assign new_n8413_ = ~n_n2395 & new_n1220_;
  assign new_n8414_ = pencrypt_0_ & new_n8413_;
  assign new_n8415_ = n_n2301 & new_n8414_;
  assign new_n8416_ = ~pstart_0_ & new_n8415_;
  assign new_n8417_ = ~new_n1200_ & new_n3604_;
  assign new_n8418_ = ~pstart_0_ & new_n8417_;
  assign new_n8419_ = n_n2395 & ~new_n1220_;
  assign new_n8420_ = pencrypt_0_ & new_n8419_;
  assign new_n8421_ = n_n2301 & new_n8420_;
  assign new_n8422_ = ~pstart_0_ & new_n8421_;
  assign new_n8423_ = ~new_n8418_ & ~new_n8422_;
  assign new_n8424_ = ~new_n8412_ & ~new_n8416_;
  assign new_n8425_ = new_n8423_ & new_n8424_;
  assign new_n8426_ = ~new_n8406_ & ~new_n8408_;
  assign new_n8427_ = ~new_n8400_ & ~new_n8402_;
  assign new_n8428_ = ~new_n8404_ & new_n8427_;
  assign new_n8429_ = new_n8426_ & new_n8428_;
  assign n1942 = ~new_n8425_ | ~new_n8429_;
  assign new_n8431_ = new_n1200_ & new_n5172_;
  assign new_n8432_ = ~pstart_0_ & new_n8431_;
  assign new_n8433_ = ~new_n1200_ & new_n5167_;
  assign new_n8434_ = ~pstart_0_ & new_n8433_;
  assign new_n8435_ = pencrypt_0_ & pkey_176_;
  assign new_n8436_ = pstart_0_ & new_n8435_;
  assign new_n8437_ = new_n1200_ & new_n5163_;
  assign new_n8438_ = ~pstart_0_ & new_n8437_;
  assign new_n8439_ = ~pencrypt_0_ & pkey_184_;
  assign new_n8440_ = pstart_0_ & new_n8439_;
  assign new_n8441_ = n_n2418 & new_n1220_;
  assign new_n8442_ = pencrypt_0_ & new_n8441_;
  assign new_n8443_ = ~n_n2324 & new_n8442_;
  assign new_n8444_ = ~pstart_0_ & new_n8443_;
  assign new_n8445_ = ~n_n2418 & new_n1220_;
  assign new_n8446_ = pencrypt_0_ & new_n8445_;
  assign new_n8447_ = n_n2324 & new_n8446_;
  assign new_n8448_ = ~pstart_0_ & new_n8447_;
  assign new_n8449_ = ~new_n1200_ & new_n5186_;
  assign new_n8450_ = ~pstart_0_ & new_n8449_;
  assign new_n8451_ = n_n2418 & ~new_n1220_;
  assign new_n8452_ = pencrypt_0_ & new_n8451_;
  assign new_n8453_ = n_n2324 & new_n8452_;
  assign new_n8454_ = ~pstart_0_ & new_n8453_;
  assign new_n8455_ = ~new_n8450_ & ~new_n8454_;
  assign new_n8456_ = ~new_n8444_ & ~new_n8448_;
  assign new_n8457_ = new_n8455_ & new_n8456_;
  assign new_n8458_ = ~new_n8438_ & ~new_n8440_;
  assign new_n8459_ = ~new_n8432_ & ~new_n8434_;
  assign new_n8460_ = ~new_n8436_ & new_n8459_;
  assign new_n8461_ = new_n8458_ & new_n8460_;
  assign n1947 = ~new_n8457_ | ~new_n8461_;
  assign new_n8463_ = new_n1200_ & new_n5210_;
  assign new_n8464_ = ~pstart_0_ & new_n8463_;
  assign new_n8465_ = ~new_n1200_ & new_n5205_;
  assign new_n8466_ = ~pstart_0_ & new_n8465_;
  assign new_n8467_ = pencrypt_0_ & pkey_90_;
  assign new_n8468_ = pstart_0_ & new_n8467_;
  assign new_n8469_ = new_n1200_ & new_n5201_;
  assign new_n8470_ = ~pstart_0_ & new_n8469_;
  assign new_n8471_ = pkey_98_ & ~pencrypt_0_;
  assign new_n8472_ = pstart_0_ & new_n8471_;
  assign new_n8473_ = n_n2426 & new_n1220_;
  assign new_n8474_ = pencrypt_0_ & new_n8473_;
  assign new_n8475_ = ~n_n2331 & new_n8474_;
  assign new_n8476_ = ~pstart_0_ & new_n8475_;
  assign new_n8477_ = ~n_n2426 & new_n1220_;
  assign new_n8478_ = pencrypt_0_ & new_n8477_;
  assign new_n8479_ = n_n2331 & new_n8478_;
  assign new_n8480_ = ~pstart_0_ & new_n8479_;
  assign new_n8481_ = ~new_n1200_ & new_n5224_;
  assign new_n8482_ = ~pstart_0_ & new_n8481_;
  assign new_n8483_ = n_n2426 & ~new_n1220_;
  assign new_n8484_ = pencrypt_0_ & new_n8483_;
  assign new_n8485_ = n_n2331 & new_n8484_;
  assign new_n8486_ = ~pstart_0_ & new_n8485_;
  assign new_n8487_ = ~new_n8482_ & ~new_n8486_;
  assign new_n8488_ = ~new_n8476_ & ~new_n8480_;
  assign new_n8489_ = new_n8487_ & new_n8488_;
  assign new_n8490_ = ~new_n8470_ & ~new_n8472_;
  assign new_n8491_ = ~new_n8464_ & ~new_n8466_;
  assign new_n8492_ = ~new_n8468_ & new_n8491_;
  assign new_n8493_ = new_n8490_ & new_n8492_;
  assign n1952 = ~new_n8489_ | ~new_n8493_;
  assign new_n8495_ = new_n1200_ & new_n2944_;
  assign new_n8496_ = ~pstart_0_ & new_n8495_;
  assign new_n8497_ = ~new_n1200_ & new_n2939_;
  assign new_n8498_ = ~pstart_0_ & new_n8497_;
  assign new_n8499_ = pencrypt_0_ & pkey_64_;
  assign new_n8500_ = pstart_0_ & new_n8499_;
  assign new_n8501_ = new_n1200_ & new_n2935_;
  assign new_n8502_ = ~pstart_0_ & new_n8501_;
  assign new_n8503_ = ~pencrypt_0_ & pkey_72_;
  assign new_n8504_ = pstart_0_ & new_n8503_;
  assign new_n8505_ = n_n2954 & new_n1220_;
  assign new_n8506_ = pencrypt_0_ & new_n8505_;
  assign new_n8507_ = ~n_n2342 & new_n8506_;
  assign new_n8508_ = ~pstart_0_ & new_n8507_;
  assign new_n8509_ = ~n_n2954 & new_n1220_;
  assign new_n8510_ = pencrypt_0_ & new_n8509_;
  assign new_n8511_ = n_n2342 & new_n8510_;
  assign new_n8512_ = ~pstart_0_ & new_n8511_;
  assign new_n8513_ = ~new_n1200_ & new_n2958_;
  assign new_n8514_ = ~pstart_0_ & new_n8513_;
  assign new_n8515_ = n_n2954 & ~new_n1220_;
  assign new_n8516_ = pencrypt_0_ & new_n8515_;
  assign new_n8517_ = n_n2342 & new_n8516_;
  assign new_n8518_ = ~pstart_0_ & new_n8517_;
  assign new_n8519_ = ~new_n8514_ & ~new_n8518_;
  assign new_n8520_ = ~new_n8508_ & ~new_n8512_;
  assign new_n8521_ = new_n8519_ & new_n8520_;
  assign new_n8522_ = ~new_n8502_ & ~new_n8504_;
  assign new_n8523_ = ~new_n8496_ & ~new_n8498_;
  assign new_n8524_ = ~new_n8500_ & new_n8523_;
  assign new_n8525_ = new_n8522_ & new_n8524_;
  assign n1957 = ~new_n8521_ | ~new_n8525_;
  assign new_n8527_ = new_n1200_ & new_n2982_;
  assign new_n8528_ = ~pstart_0_ & new_n8527_;
  assign new_n8529_ = ~new_n1200_ & new_n2977_;
  assign new_n8530_ = ~pstart_0_ & new_n8529_;
  assign new_n8531_ = pencrypt_0_ & pkey_43_;
  assign new_n8532_ = pstart_0_ & new_n8531_;
  assign new_n8533_ = new_n1200_ & new_n2973_;
  assign new_n8534_ = ~pstart_0_ & new_n8533_;
  assign new_n8535_ = pkey_51_ & ~pencrypt_0_;
  assign new_n8536_ = pstart_0_ & new_n8535_;
  assign new_n8537_ = n_n2964 & new_n1220_;
  assign new_n8538_ = pencrypt_0_ & new_n8537_;
  assign new_n8539_ = ~n_n2351 & new_n8538_;
  assign new_n8540_ = ~pstart_0_ & new_n8539_;
  assign new_n8541_ = ~n_n2964 & new_n1220_;
  assign new_n8542_ = pencrypt_0_ & new_n8541_;
  assign new_n8543_ = n_n2351 & new_n8542_;
  assign new_n8544_ = ~pstart_0_ & new_n8543_;
  assign new_n8545_ = ~new_n1200_ & new_n2996_;
  assign new_n8546_ = ~pstart_0_ & new_n8545_;
  assign new_n8547_ = n_n2964 & ~new_n1220_;
  assign new_n8548_ = pencrypt_0_ & new_n8547_;
  assign new_n8549_ = n_n2351 & new_n8548_;
  assign new_n8550_ = ~pstart_0_ & new_n8549_;
  assign new_n8551_ = ~new_n8546_ & ~new_n8550_;
  assign new_n8552_ = ~new_n8540_ & ~new_n8544_;
  assign new_n8553_ = new_n8551_ & new_n8552_;
  assign new_n8554_ = ~new_n8534_ & ~new_n8536_;
  assign new_n8555_ = ~new_n8528_ & ~new_n8530_;
  assign new_n8556_ = ~new_n8532_ & new_n8555_;
  assign new_n8557_ = new_n8554_ & new_n8556_;
  assign n1962 = ~new_n8553_ | ~new_n8557_;
  assign new_n8559_ = new_n1200_ & new_n1444_;
  assign new_n8560_ = ~pstart_0_ & new_n8559_;
  assign new_n8561_ = ~new_n1200_ & new_n1439_;
  assign new_n8562_ = ~pstart_0_ & new_n8561_;
  assign new_n8563_ = pkey_18_ & pencrypt_0_;
  assign new_n8564_ = pstart_0_ & new_n8563_;
  assign new_n8565_ = new_n1200_ & new_n1435_;
  assign new_n8566_ = ~pstart_0_ & new_n8565_;
  assign new_n8567_ = pkey_26_ & ~pencrypt_0_;
  assign new_n8568_ = pstart_0_ & new_n8567_;
  assign new_n8569_ = n_n2448 & new_n1220_;
  assign new_n8570_ = pencrypt_0_ & new_n8569_;
  assign new_n8571_ = ~n_n2354 & new_n8570_;
  assign new_n8572_ = ~pstart_0_ & new_n8571_;
  assign new_n8573_ = ~n_n2448 & new_n1220_;
  assign new_n8574_ = pencrypt_0_ & new_n8573_;
  assign new_n8575_ = n_n2354 & new_n8574_;
  assign new_n8576_ = ~pstart_0_ & new_n8575_;
  assign new_n8577_ = ~new_n1200_ & new_n1458_;
  assign new_n8578_ = ~pstart_0_ & new_n8577_;
  assign new_n8579_ = n_n2448 & ~new_n1220_;
  assign new_n8580_ = pencrypt_0_ & new_n8579_;
  assign new_n8581_ = n_n2354 & new_n8580_;
  assign new_n8582_ = ~pstart_0_ & new_n8581_;
  assign new_n8583_ = ~new_n8578_ & ~new_n8582_;
  assign new_n8584_ = ~new_n8572_ & ~new_n8576_;
  assign new_n8585_ = new_n8583_ & new_n8584_;
  assign new_n8586_ = ~new_n8566_ & ~new_n8568_;
  assign new_n8587_ = ~new_n8560_ & ~new_n8562_;
  assign new_n8588_ = ~new_n8564_ & new_n8587_;
  assign new_n8589_ = new_n8586_ & new_n8588_;
  assign n1967 = ~new_n8585_ | ~new_n8589_;
  assign new_n8591_ = new_n1200_ & new_n3892_;
  assign new_n8592_ = ~pstart_0_ & new_n8591_;
  assign new_n8593_ = ~new_n1200_ & new_n3889_;
  assign new_n8594_ = ~pstart_0_ & new_n8593_;
  assign new_n8595_ = pencrypt_0_ & pkey_170_;
  assign new_n8596_ = pstart_0_ & new_n8595_;
  assign new_n8597_ = new_n1200_ & new_n3885_;
  assign new_n8598_ = ~pstart_0_ & new_n8597_;
  assign new_n8599_ = ~pencrypt_0_ & pkey_178_;
  assign new_n8600_ = pstart_0_ & new_n8599_;
  assign new_n8601_ = n_n2404 & new_n1220_;
  assign new_n8602_ = pencrypt_0_ & new_n8601_;
  assign new_n8603_ = ~n_n2779 & new_n8602_;
  assign new_n8604_ = ~pstart_0_ & new_n8603_;
  assign new_n8605_ = ~n_n2404 & new_n1220_;
  assign new_n8606_ = pencrypt_0_ & new_n8605_;
  assign new_n8607_ = n_n2779 & new_n8606_;
  assign new_n8608_ = ~pstart_0_ & new_n8607_;
  assign new_n8609_ = ~new_n1200_ & new_n3906_;
  assign new_n8610_ = ~pstart_0_ & new_n8609_;
  assign new_n8611_ = n_n2404 & ~new_n1220_;
  assign new_n8612_ = pencrypt_0_ & new_n8611_;
  assign new_n8613_ = n_n2779 & new_n8612_;
  assign new_n8614_ = ~pstart_0_ & new_n8613_;
  assign new_n8615_ = ~new_n8610_ & ~new_n8614_;
  assign new_n8616_ = ~new_n8604_ & ~new_n8608_;
  assign new_n8617_ = new_n8615_ & new_n8616_;
  assign new_n8618_ = ~new_n8598_ & ~new_n8600_;
  assign new_n8619_ = ~new_n8592_ & ~new_n8594_;
  assign new_n8620_ = ~new_n8596_ & new_n8619_;
  assign new_n8621_ = new_n8618_ & new_n8620_;
  assign n1972 = ~new_n8617_ | ~new_n8621_;
  assign new_n8623_ = new_n1200_ & new_n4456_;
  assign new_n8624_ = ~pstart_0_ & new_n8623_;
  assign new_n8625_ = ~new_n1200_ & new_n4451_;
  assign new_n8626_ = ~pstart_0_ & new_n8625_;
  assign new_n8627_ = pkey_128_ & pencrypt_0_;
  assign new_n8628_ = pstart_0_ & new_n8627_;
  assign new_n8629_ = new_n1200_ & new_n4447_;
  assign new_n8630_ = ~pstart_0_ & new_n8629_;
  assign new_n8631_ = pkey_136_ & ~pencrypt_0_;
  assign new_n8632_ = pstart_0_ & new_n8631_;
  assign new_n8633_ = n_n2921 & new_n1220_;
  assign new_n8634_ = pencrypt_0_ & new_n8633_;
  assign new_n8635_ = ~n_n2318 & new_n8634_;
  assign new_n8636_ = ~pstart_0_ & new_n8635_;
  assign new_n8637_ = ~n_n2921 & new_n1220_;
  assign new_n8638_ = pencrypt_0_ & new_n8637_;
  assign new_n8639_ = n_n2318 & new_n8638_;
  assign new_n8640_ = ~pstart_0_ & new_n8639_;
  assign new_n8641_ = ~new_n1200_ & new_n4470_;
  assign new_n8642_ = ~pstart_0_ & new_n8641_;
  assign new_n8643_ = n_n2921 & ~new_n1220_;
  assign new_n8644_ = pencrypt_0_ & new_n8643_;
  assign new_n8645_ = n_n2318 & new_n8644_;
  assign new_n8646_ = ~pstart_0_ & new_n8645_;
  assign new_n8647_ = ~new_n8642_ & ~new_n8646_;
  assign new_n8648_ = ~new_n8636_ & ~new_n8640_;
  assign new_n8649_ = new_n8647_ & new_n8648_;
  assign new_n8650_ = ~new_n8630_ & ~new_n8632_;
  assign new_n8651_ = ~new_n8624_ & ~new_n8626_;
  assign new_n8652_ = ~new_n8628_ & new_n8651_;
  assign new_n8653_ = new_n8650_ & new_n8652_;
  assign n1977 = ~new_n8649_ | ~new_n8653_;
  assign new_n8655_ = new_n1200_ & new_n1976_;
  assign new_n8656_ = ~pstart_0_ & new_n8655_;
  assign new_n8657_ = ~new_n1200_ & new_n1971_;
  assign new_n8658_ = ~pstart_0_ & new_n8657_;
  assign new_n8659_ = pencrypt_0_ & pkey_184_;
  assign new_n8660_ = pstart_0_ & new_n8659_;
  assign new_n8661_ = new_n1200_ & new_n1967_1_;
  assign new_n8662_ = ~pstart_0_ & new_n8661_;
  assign new_n8663_ = pkey_99_ & ~pencrypt_0_;
  assign new_n8664_ = pstart_0_ & new_n8663_;
  assign new_n8665_ = n_n2419 & new_n1220_;
  assign new_n8666_ = pencrypt_0_ & new_n8665_;
  assign new_n8667_ = ~n_n2325 & new_n8666_;
  assign new_n8668_ = ~pstart_0_ & new_n8667_;
  assign new_n8669_ = ~n_n2419 & new_n1220_;
  assign new_n8670_ = pencrypt_0_ & new_n8669_;
  assign new_n8671_ = n_n2325 & new_n8670_;
  assign new_n8672_ = ~pstart_0_ & new_n8671_;
  assign new_n8673_ = ~new_n1200_ & new_n1990_;
  assign new_n8674_ = ~pstart_0_ & new_n8673_;
  assign new_n8675_ = n_n2419 & ~new_n1220_;
  assign new_n8676_ = pencrypt_0_ & new_n8675_;
  assign new_n8677_ = n_n2325 & new_n8676_;
  assign new_n8678_ = ~pstart_0_ & new_n8677_;
  assign new_n8679_ = ~new_n8674_ & ~new_n8678_;
  assign new_n8680_ = ~new_n8668_ & ~new_n8672_;
  assign new_n8681_ = new_n8679_ & new_n8680_;
  assign new_n8682_ = ~new_n8662_ & ~new_n8664_;
  assign new_n8683_ = ~new_n8656_ & ~new_n8658_;
  assign new_n8684_ = ~new_n8660_ & new_n8683_;
  assign new_n8685_ = new_n8682_ & new_n8684_;
  assign n1982 = ~new_n8681_ | ~new_n8685_;
  assign new_n8687_ = new_n1200_ & new_n2014_;
  assign new_n8688_ = ~pstart_0_ & new_n8687_;
  assign new_n8689_ = ~new_n1200_ & new_n2009_;
  assign new_n8690_ = ~pstart_0_ & new_n8689_;
  assign new_n8691_ = pkey_114_ & pencrypt_0_;
  assign new_n8692_ = pstart_0_ & new_n8691_;
  assign new_n8693_ = new_n1200_ & new_n2005_;
  assign new_n8694_ = ~pstart_0_ & new_n8693_;
  assign new_n8695_ = pkey_122_ & ~pencrypt_0_;
  assign new_n8696_ = pstart_0_ & new_n8695_;
  assign new_n8697_ = n_n2429 & new_n1220_;
  assign new_n8698_ = pencrypt_0_ & new_n8697_;
  assign new_n8699_ = ~n_n2333 & new_n8698_;
  assign new_n8700_ = ~pstart_0_ & new_n8699_;
  assign new_n8701_ = ~n_n2429 & new_n1220_;
  assign new_n8702_ = pencrypt_0_ & new_n8701_;
  assign new_n8703_ = n_n2333 & new_n8702_;
  assign new_n8704_ = ~pstart_0_ & new_n8703_;
  assign new_n8705_ = ~new_n1200_ & new_n2028_;
  assign new_n8706_ = ~pstart_0_ & new_n8705_;
  assign new_n8707_ = n_n2429 & ~new_n1220_;
  assign new_n8708_ = pencrypt_0_ & new_n8707_;
  assign new_n8709_ = n_n2333 & new_n8708_;
  assign new_n8710_ = ~pstart_0_ & new_n8709_;
  assign new_n8711_ = ~new_n8706_ & ~new_n8710_;
  assign new_n8712_ = ~new_n8700_ & ~new_n8704_;
  assign new_n8713_ = new_n8711_ & new_n8712_;
  assign new_n8714_ = ~new_n8694_ & ~new_n8696_;
  assign new_n8715_ = ~new_n8688_ & ~new_n8690_;
  assign new_n8716_ = ~new_n8692_ & new_n8715_;
  assign new_n8717_ = new_n8714_ & new_n8716_;
  assign n1987 = ~new_n8713_ | ~new_n8717_;
  assign new_n8719_ = new_n1200_ & new_n4272_;
  assign new_n8720_ = ~pstart_0_ & new_n8719_;
  assign new_n8721_ = ~new_n1200_ & new_n4267_;
  assign new_n8722_ = ~pstart_0_ & new_n8721_;
  assign new_n8723_ = pencrypt_0_ & pkey_105_;
  assign new_n8724_ = pstart_0_ & new_n8723_;
  assign new_n8725_ = new_n1200_ & new_n4263_;
  assign new_n8726_ = ~pstart_0_ & new_n8725_;
  assign new_n8727_ = pkey_113_ & ~pencrypt_0_;
  assign new_n8728_ = pstart_0_ & new_n8727_;
  assign new_n8729_ = n_n2950 & new_n1220_;
  assign new_n8730_ = pencrypt_0_ & new_n8729_;
  assign new_n8731_ = ~n_n2340 & new_n8730_;
  assign new_n8732_ = ~pstart_0_ & new_n8731_;
  assign new_n8733_ = ~n_n2950 & new_n1220_;
  assign new_n8734_ = pencrypt_0_ & new_n8733_;
  assign new_n8735_ = n_n2340 & new_n8734_;
  assign new_n8736_ = ~pstart_0_ & new_n8735_;
  assign new_n8737_ = ~new_n1200_ & new_n4286_;
  assign new_n8738_ = ~pstart_0_ & new_n8737_;
  assign new_n8739_ = n_n2950 & ~new_n1220_;
  assign new_n8740_ = pencrypt_0_ & new_n8739_;
  assign new_n8741_ = n_n2340 & new_n8740_;
  assign new_n8742_ = ~pstart_0_ & new_n8741_;
  assign new_n8743_ = ~new_n8738_ & ~new_n8742_;
  assign new_n8744_ = ~new_n8732_ & ~new_n8736_;
  assign new_n8745_ = new_n8743_ & new_n8744_;
  assign new_n8746_ = ~new_n8726_ & ~new_n8728_;
  assign new_n8747_ = ~new_n8720_ & ~new_n8722_;
  assign new_n8748_ = ~new_n8724_ & new_n8747_;
  assign new_n8749_ = new_n8746_ & new_n8748_;
  assign n1992 = ~new_n8745_ | ~new_n8749_;
  assign new_n8751_ = new_n1200_ & new_n4310_;
  assign new_n8752_ = ~pstart_0_ & new_n8751_;
  assign new_n8753_ = ~new_n1200_ & new_n4305_;
  assign new_n8754_ = ~pstart_0_ & new_n8753_;
  assign new_n8755_ = pencrypt_0_ & pkey_35_;
  assign new_n8756_ = pstart_0_ & new_n8755_;
  assign new_n8757_ = new_n1200_ & new_n4301_;
  assign new_n8758_ = ~pstart_0_ & new_n8757_;
  assign new_n8759_ = ~pencrypt_0_ & pkey_43_;
  assign new_n8760_ = pstart_0_ & new_n8759_;
  assign new_n8761_ = n_n2443 & new_n1220_;
  assign new_n8762_ = pencrypt_0_ & new_n8761_;
  assign new_n8763_ = ~n_n2350 & new_n8762_;
  assign new_n8764_ = ~pstart_0_ & new_n8763_;
  assign new_n8765_ = ~n_n2443 & new_n1220_;
  assign new_n8766_ = pencrypt_0_ & new_n8765_;
  assign new_n8767_ = n_n2350 & new_n8766_;
  assign new_n8768_ = ~pstart_0_ & new_n8767_;
  assign new_n8769_ = ~new_n1200_ & new_n4324_;
  assign new_n8770_ = ~pstart_0_ & new_n8769_;
  assign new_n8771_ = n_n2443 & ~new_n1220_;
  assign new_n8772_ = pencrypt_0_ & new_n8771_;
  assign new_n8773_ = n_n2350 & new_n8772_;
  assign new_n8774_ = ~pstart_0_ & new_n8773_;
  assign new_n8775_ = ~new_n8770_ & ~new_n8774_;
  assign new_n8776_ = ~new_n8764_ & ~new_n8768_;
  assign new_n8777_ = new_n8775_ & new_n8776_;
  assign new_n8778_ = ~new_n8758_ & ~new_n8760_;
  assign new_n8779_ = ~new_n8752_ & ~new_n8754_;
  assign new_n8780_ = ~new_n8756_ & new_n8779_;
  assign new_n8781_ = new_n8778_ & new_n8780_;
  assign n1997 = ~new_n8777_ | ~new_n8781_;
  assign new_n8783_ = new_n1200_ & new_n1748_;
  assign new_n8784_ = ~pstart_0_ & new_n8783_;
  assign new_n8785_ = ~new_n1200_ & new_n1743_;
  assign new_n8786_ = ~pstart_0_ & new_n8785_;
  assign new_n8787_ = pkey_26_ & pencrypt_0_;
  assign new_n8788_ = pstart_0_ & new_n8787_;
  assign new_n8789_ = new_n1200_ & new_n1739_;
  assign new_n8790_ = ~pstart_0_ & new_n8789_;
  assign new_n8791_ = ~pencrypt_0_ & pkey_34_;
  assign new_n8792_ = pstart_0_ & new_n8791_;
  assign new_n8793_ = n_n2449 & new_n1220_;
  assign new_n8794_ = pencrypt_0_ & new_n8793_;
  assign new_n8795_ = ~n_n2355 & new_n8794_;
  assign new_n8796_ = ~pstart_0_ & new_n8795_;
  assign new_n8797_ = ~n_n2449 & new_n1220_;
  assign new_n8798_ = pencrypt_0_ & new_n8797_;
  assign new_n8799_ = n_n2355 & new_n8798_;
  assign new_n8800_ = ~pstart_0_ & new_n8799_;
  assign new_n8801_ = ~new_n1200_ & new_n1762_1_;
  assign new_n8802_ = ~pstart_0_ & new_n8801_;
  assign new_n8803_ = n_n2449 & ~new_n1220_;
  assign new_n8804_ = pencrypt_0_ & new_n8803_;
  assign new_n8805_ = n_n2355 & new_n8804_;
  assign new_n8806_ = ~pstart_0_ & new_n8805_;
  assign new_n8807_ = ~new_n8802_ & ~new_n8806_;
  assign new_n8808_ = ~new_n8796_ & ~new_n8800_;
  assign new_n8809_ = new_n8807_ & new_n8808_;
  assign new_n8810_ = ~new_n8790_ & ~new_n8792_;
  assign new_n8811_ = ~new_n8784_ & ~new_n8786_;
  assign new_n8812_ = ~new_n8788_ & new_n8811_;
  assign new_n8813_ = new_n8810_ & new_n8812_;
  assign n2002 = ~new_n8809_ | ~new_n8813_;
  assign new_n8815_ = new_n1200_ & new_n3628_;
  assign new_n8816_ = ~pstart_0_ & new_n8815_;
  assign new_n8817_ = ~new_n1200_ & new_n3623_;
  assign new_n8818_ = ~pstart_0_ & new_n8817_;
  assign new_n8819_ = pencrypt_0_ & pkey_178_;
  assign new_n8820_ = pstart_0_ & new_n8819_;
  assign new_n8821_ = new_n1200_ & new_n3619_;
  assign new_n8822_ = ~pstart_0_ & new_n8821_;
  assign new_n8823_ = ~pencrypt_0_ & pkey_186_;
  assign new_n8824_ = pstart_0_ & new_n8823_;
  assign new_n8825_ = n_n2909 & new_n1220_;
  assign new_n8826_ = pencrypt_0_ & new_n8825_;
  assign new_n8827_ = ~n_n2309 & new_n8826_;
  assign new_n8828_ = ~pstart_0_ & new_n8827_;
  assign new_n8829_ = ~n_n2909 & new_n1220_;
  assign new_n8830_ = pencrypt_0_ & new_n8829_;
  assign new_n8831_ = n_n2309 & new_n8830_;
  assign new_n8832_ = ~pstart_0_ & new_n8831_;
  assign new_n8833_ = ~new_n1200_ & new_n3642_;
  assign new_n8834_ = ~pstart_0_ & new_n8833_;
  assign new_n8835_ = n_n2909 & ~new_n1220_;
  assign new_n8836_ = pencrypt_0_ & new_n8835_;
  assign new_n8837_ = n_n2309 & new_n8836_;
  assign new_n8838_ = ~pstart_0_ & new_n8837_;
  assign new_n8839_ = ~new_n8834_ & ~new_n8838_;
  assign new_n8840_ = ~new_n8828_ & ~new_n8832_;
  assign new_n8841_ = new_n8839_ & new_n8840_;
  assign new_n8842_ = ~new_n8822_ & ~new_n8824_;
  assign new_n8843_ = ~new_n8816_ & ~new_n8818_;
  assign new_n8844_ = ~new_n8820_ & new_n8843_;
  assign new_n8845_ = new_n8842_ & new_n8844_;
  assign n2007 = ~new_n8841_ | ~new_n8845_;
  assign new_n8847_ = new_n1200_ & new_n4196_;
  assign new_n8848_ = ~pstart_0_ & new_n8847_;
  assign new_n8849_ = ~new_n1200_ & new_n4191_;
  assign new_n8850_ = ~pstart_0_ & new_n8849_;
  assign new_n8851_ = pencrypt_0_ & pkey_185_;
  assign new_n8852_ = pstart_0_ & new_n8851_;
  assign new_n8853_ = new_n1200_ & new_n4187_;
  assign new_n8854_ = ~pstart_0_ & new_n8853_;
  assign new_n8855_ = pkey_128_ & ~pencrypt_0_;
  assign new_n8856_ = pstart_0_ & new_n8855_;
  assign new_n8857_ = n_n2412 & new_n1220_;
  assign new_n8858_ = pencrypt_0_ & new_n8857_;
  assign new_n8859_ = ~n_n2317 & new_n8858_;
  assign new_n8860_ = ~pstart_0_ & new_n8859_;
  assign new_n8861_ = ~n_n2412 & new_n1220_;
  assign new_n8862_ = pencrypt_0_ & new_n8861_;
  assign new_n8863_ = n_n2317 & new_n8862_;
  assign new_n8864_ = ~pstart_0_ & new_n8863_;
  assign new_n8865_ = ~new_n1200_ & new_n4210_;
  assign new_n8866_ = ~pstart_0_ & new_n8865_;
  assign new_n8867_ = n_n2412 & ~new_n1220_;
  assign new_n8868_ = pencrypt_0_ & new_n8867_;
  assign new_n8869_ = n_n2317 & new_n8868_;
  assign new_n8870_ = ~pstart_0_ & new_n8869_;
  assign new_n8871_ = ~new_n8866_ & ~new_n8870_;
  assign new_n8872_ = ~new_n8860_ & ~new_n8864_;
  assign new_n8873_ = new_n8871_ & new_n8872_;
  assign new_n8874_ = ~new_n8854_ & ~new_n8856_;
  assign new_n8875_ = ~new_n8848_ & ~new_n8850_;
  assign new_n8876_ = ~new_n8852_ & new_n8875_;
  assign new_n8877_ = new_n8874_ & new_n8876_;
  assign n2012 = ~new_n8873_ | ~new_n8877_;
  assign new_n8879_ = new_n1200_ & new_n2312_;
  assign new_n8880_ = ~pstart_0_ & new_n8879_;
  assign new_n8881_ = ~new_n1200_ & new_n2307_;
  assign new_n8882_ = ~pstart_0_ & new_n8881_;
  assign new_n8883_ = pkey_99_ & pencrypt_0_;
  assign new_n8884_ = pstart_0_ & new_n8883_;
  assign new_n8885_ = new_n1200_ & new_n2303_;
  assign new_n8886_ = ~pstart_0_ & new_n8885_;
  assign new_n8887_ = pkey_107_ & ~pencrypt_0_;
  assign new_n8888_ = pstart_0_ & new_n8887_;
  assign new_n8889_ = n_n2420 & new_n1220_;
  assign new_n8890_ = pencrypt_0_ & new_n8889_;
  assign new_n8891_ = ~n_n2326 & new_n8890_;
  assign new_n8892_ = ~pstart_0_ & new_n8891_;
  assign new_n8893_ = ~n_n2420 & new_n1220_;
  assign new_n8894_ = pencrypt_0_ & new_n8893_;
  assign new_n8895_ = n_n2326 & new_n8894_;
  assign new_n8896_ = ~pstart_0_ & new_n8895_;
  assign new_n8897_ = ~new_n1200_ & new_n2326_;
  assign new_n8898_ = ~pstart_0_ & new_n8897_;
  assign new_n8899_ = n_n2420 & ~new_n1220_;
  assign new_n8900_ = pencrypt_0_ & new_n8899_;
  assign new_n8901_ = n_n2326 & new_n8900_;
  assign new_n8902_ = ~pstart_0_ & new_n8901_;
  assign new_n8903_ = ~new_n8898_ & ~new_n8902_;
  assign new_n8904_ = ~new_n8892_ & ~new_n8896_;
  assign new_n8905_ = new_n8903_ & new_n8904_;
  assign new_n8906_ = ~new_n8886_ & ~new_n8888_;
  assign new_n8907_ = ~new_n8880_ & ~new_n8882_;
  assign new_n8908_ = ~new_n8884_ & new_n8907_;
  assign new_n8909_ = new_n8906_ & new_n8908_;
  assign n2017 = ~new_n8905_ | ~new_n8909_;
  assign new_n8911_ = new_n1200_ & new_n2350_;
  assign new_n8912_ = ~pstart_0_ & new_n8911_;
  assign new_n8913_ = ~new_n1200_ & new_n2345_;
  assign new_n8914_ = ~pstart_0_ & new_n8913_;
  assign new_n8915_ = pencrypt_0_ & pkey_106_;
  assign new_n8916_ = pstart_0_ & new_n8915_;
  assign new_n8917_ = new_n1200_ & new_n2341_;
  assign new_n8918_ = ~pstart_0_ & new_n8917_;
  assign new_n8919_ = pkey_114_ & ~pencrypt_0_;
  assign new_n8920_ = pstart_0_ & new_n8919_;
  assign new_n8921_ = n_n2428 & new_n1220_;
  assign new_n8922_ = pencrypt_0_ & new_n8921_;
  assign new_n8923_ = ~n_n2811 & new_n8922_;
  assign new_n8924_ = ~pstart_0_ & new_n8923_;
  assign new_n8925_ = ~n_n2428 & new_n1220_;
  assign new_n8926_ = pencrypt_0_ & new_n8925_;
  assign new_n8927_ = n_n2811 & new_n8926_;
  assign new_n8928_ = ~pstart_0_ & new_n8927_;
  assign new_n8929_ = ~new_n1200_ & new_n2364_;
  assign new_n8930_ = ~pstart_0_ & new_n8929_;
  assign new_n8931_ = n_n2428 & ~new_n1220_;
  assign new_n8932_ = pencrypt_0_ & new_n8931_;
  assign new_n8933_ = n_n2811 & new_n8932_;
  assign new_n8934_ = ~pstart_0_ & new_n8933_;
  assign new_n8935_ = ~new_n8930_ & ~new_n8934_;
  assign new_n8936_ = ~new_n8924_ & ~new_n8928_;
  assign new_n8937_ = new_n8935_ & new_n8936_;
  assign new_n8938_ = ~new_n8918_ & ~new_n8920_;
  assign new_n8939_ = ~new_n8912_ & ~new_n8914_;
  assign new_n8940_ = ~new_n8916_ & new_n8939_;
  assign new_n8941_ = new_n8938_ & new_n8940_;
  assign n2022 = ~new_n8937_ | ~new_n8941_;
  assign new_n8943_ = new_n1200_ & new_n4532_;
  assign new_n8944_ = ~pstart_0_ & new_n8943_;
  assign new_n8945_ = ~new_n1200_ & new_n4527_;
  assign new_n8946_ = ~pstart_0_ & new_n8945_;
  assign new_n8947_ = pkey_113_ & pencrypt_0_;
  assign new_n8948_ = pstart_0_ & new_n8947_;
  assign new_n8949_ = new_n1200_ & new_n4523_;
  assign new_n8950_ = ~pstart_0_ & new_n8949_;
  assign new_n8951_ = pkey_121_ & ~pencrypt_0_;
  assign new_n8952_ = pstart_0_ & new_n8951_;
  assign new_n8953_ = n_n2434 & new_n1220_;
  assign new_n8954_ = pencrypt_0_ & new_n8953_;
  assign new_n8955_ = ~n_n2821 & new_n8954_;
  assign new_n8956_ = ~pstart_0_ & new_n8955_;
  assign new_n8957_ = ~n_n2434 & new_n1220_;
  assign new_n8958_ = pencrypt_0_ & new_n8957_;
  assign new_n8959_ = n_n2821 & new_n8958_;
  assign new_n8960_ = ~pstart_0_ & new_n8959_;
  assign new_n8961_ = ~new_n1200_ & new_n4546_;
  assign new_n8962_ = ~pstart_0_ & new_n8961_;
  assign new_n8963_ = n_n2434 & ~new_n1220_;
  assign new_n8964_ = pencrypt_0_ & new_n8963_;
  assign new_n8965_ = n_n2821 & new_n8964_;
  assign new_n8966_ = ~pstart_0_ & new_n8965_;
  assign new_n8967_ = ~new_n8962_ & ~new_n8966_;
  assign new_n8968_ = ~new_n8956_ & ~new_n8960_;
  assign new_n8969_ = new_n8967_ & new_n8968_;
  assign new_n8970_ = ~new_n8950_ & ~new_n8952_;
  assign new_n8971_ = ~new_n8944_ & ~new_n8946_;
  assign new_n8972_ = ~new_n8948_ & new_n8971_;
  assign new_n8973_ = new_n8970_ & new_n8972_;
  assign n2027 = ~new_n8969_ | ~new_n8973_;
  assign new_n8975_ = new_n1200_ & new_n4570_;
  assign new_n8976_ = ~pstart_0_ & new_n8975_;
  assign new_n8977_ = ~new_n1200_ & new_n4565_;
  assign new_n8978_ = ~pstart_0_ & new_n8977_;
  assign new_n8979_ = pkey_120_ & pencrypt_0_;
  assign new_n8980_ = pstart_0_ & new_n8979_;
  assign new_n8981_ = new_n1200_ & new_n4561_;
  assign new_n8982_ = ~pstart_0_ & new_n8981_;
  assign new_n8983_ = ~pencrypt_0_ & pkey_35_;
  assign new_n8984_ = pstart_0_ & new_n8983_;
  assign new_n8985_ = n_n2442 & new_n1220_;
  assign new_n8986_ = pencrypt_0_ & new_n8985_;
  assign new_n8987_ = ~n_n2349 & new_n8986_;
  assign new_n8988_ = ~pstart_0_ & new_n8987_;
  assign new_n8989_ = ~n_n2442 & new_n1220_;
  assign new_n8990_ = pencrypt_0_ & new_n8989_;
  assign new_n8991_ = n_n2349 & new_n8990_;
  assign new_n8992_ = ~pstart_0_ & new_n8991_;
  assign new_n8993_ = ~new_n1200_ & new_n4584_;
  assign new_n8994_ = ~pstart_0_ & new_n8993_;
  assign new_n8995_ = n_n2442 & ~new_n1220_;
  assign new_n8996_ = pencrypt_0_ & new_n8995_;
  assign new_n8997_ = n_n2349 & new_n8996_;
  assign new_n8998_ = ~pstart_0_ & new_n8997_;
  assign new_n8999_ = ~new_n8994_ & ~new_n8998_;
  assign new_n9000_ = ~new_n8988_ & ~new_n8992_;
  assign new_n9001_ = new_n8999_ & new_n9000_;
  assign new_n9002_ = ~new_n8982_ & ~new_n8984_;
  assign new_n9003_ = ~new_n8976_ & ~new_n8978_;
  assign new_n9004_ = ~new_n8980_ & new_n9003_;
  assign new_n9005_ = new_n9002_ & new_n9004_;
  assign n2032 = ~new_n9001_ | ~new_n9005_;
  assign new_n9007_ = new_n1200_ & new_n2052_;
  assign new_n9008_ = ~pstart_0_ & new_n9007_;
  assign new_n9009_ = ~new_n1200_ & new_n2047_;
  assign new_n9010_ = ~pstart_0_ & new_n9009_;
  assign new_n9011_ = pencrypt_0_ & pkey_34_;
  assign new_n9012_ = pstart_0_ & new_n9011_;
  assign new_n9013_ = new_n1200_ & new_n2043_;
  assign new_n9014_ = ~pstart_0_ & new_n9013_;
  assign new_n9015_ = ~pencrypt_0_ & pkey_42_;
  assign new_n9016_ = pstart_0_ & new_n9015_;
  assign new_n9017_ = n_n2450 & new_n1220_;
  assign new_n9018_ = pencrypt_0_ & new_n9017_;
  assign new_n9019_ = ~n_n2356 & new_n9018_;
  assign new_n9020_ = ~pstart_0_ & new_n9019_;
  assign new_n9021_ = ~n_n2450 & new_n1220_;
  assign new_n9022_ = pencrypt_0_ & new_n9021_;
  assign new_n9023_ = n_n2356 & new_n9022_;
  assign new_n9024_ = ~pstart_0_ & new_n9023_;
  assign new_n9025_ = ~new_n1200_ & new_n2066_;
  assign new_n9026_ = ~pstart_0_ & new_n9025_;
  assign new_n9027_ = n_n2450 & ~new_n1220_;
  assign new_n9028_ = pencrypt_0_ & new_n9027_;
  assign new_n9029_ = n_n2356 & new_n9028_;
  assign new_n9030_ = ~pstart_0_ & new_n9029_;
  assign new_n9031_ = ~new_n9026_ & ~new_n9030_;
  assign new_n9032_ = ~new_n9020_ & ~new_n9024_;
  assign new_n9033_ = new_n9031_ & new_n9032_;
  assign new_n9034_ = ~new_n9014_ & ~new_n9016_;
  assign new_n9035_ = ~new_n9008_ & ~new_n9010_;
  assign new_n9036_ = ~new_n9012_ & new_n9035_;
  assign new_n9037_ = new_n9034_ & new_n9036_;
  assign n2037 = ~new_n9033_ | ~new_n9037_;
  assign pksi_50_ = n_n2315;
  assign pksi_61_ = n_n2308;
  assign pksi_72_ = n_n2288;
  assign pksi_83_ = n_n2292;
  assign pksi_94_ = n_n2289;
  assign pksi_102_ = n_n2464;
  assign pksi_115_ = n_n2454;
  assign pksi_128_ = n_n2423;
  assign pksi_51_ = n_n2304;
  assign pksi_60_ = n_n2305;
  assign pksi_73_ = n_n2286;
  assign pksi_82_ = n_n2283;
  assign pksi_95_ = n_n2299;
  assign pksi_101_ = n_n2443;
  assign pksi_116_ = n_n2447;
  assign pksi_127_ = n_n2432;
  assign pksi_52_ = n_n2324;
  assign pksi_63_ = n_n2321;
  assign pksi_70_ = n_n2313;
  assign pksi_81_ = n_n2295;
  assign pksi_96_ = n_n2455;
  assign pksi_100_ = n_n2450;
  assign pksi_113_ = n_n2444;
  assign pksi_53_ = n_n2320;
  assign pksi_62_ = n_n2314;
  assign pksi_71_ = n_n2323;
  assign pksi_80_ = n_n2287;
  assign pksi_97_ = n_n2445;
  assign pksi_114_ = n_n2451;
  assign pksi_129_ = n_n2429;
  assign pksi_54_ = n_n2322;
  assign pksi_65_ = n_n2317;
  assign pksi_76_ = n_n2300;
  assign pksi_87_ = n_n2297;
  assign pksi_90_ = n_n2280;
  assign pksi_119_ = n_n2462;
  assign pksi_124_ = n_n2427;
  assign pksi_191_ = n_n2391;
  assign pksi_55_ = n_n2301;
  assign pksi_64_ = n_n2303;
  assign pksi_77_ = n_n2296;
  assign pksi_86_ = n_n2290;
  assign pksi_91_ = n_n2294;
  assign pksi_123_ = n_n2434;
  assign pksi_56_ = n_n2311;
  assign pksi_67_ = n_n2318;
  assign pksi_74_ = n_n2291;
  assign pksi_85_ = n_n2285;
  assign pksi_92_ = n_n2279;
  assign pksi_117_ = n_n2459;
  assign pksi_126_ = n_n2440;
  assign pksi_57_ = n_n2319;
  assign pksi_66_ = n_n2310;
  assign pksi_75_ = n_n2281;
  assign pksi_84_ = n_n2282;
  assign pksi_93_ = n_n2284;
  assign pksi_118_ = n_n2465;
  assign pksi_125_ = n_n2420;
  assign pksi_190_ = n_n2394;
  assign pksi_14_ = n_n2362;
  assign pksi_25_ = n_n2333;
  assign pksi_36_ = n_n2329;
  assign pksi_47_ = n_n2347;
  assign pksi_120_ = n_n2431;
  assign pksi_15_ = n_n2369;
  assign pksi_24_ = n_n2336;
  assign pksi_37_ = n_n2332;
  assign pksi_46_ = n_n2337;
  assign pksi_109_ = n_n2448;
  assign pksi_16_ = n_n2351;
  assign pksi_27_ = n_n2328;
  assign pksi_34_ = n_n2330;
  assign pksi_45_ = n_n2331;
  assign pksi_108_ = n_n2453;
  assign pksi_122_ = n_n2439;
  assign pksi_17_ = n_n2365;
  assign pksi_26_ = n_n2339;
  assign pksi_35_ = n_n2340;
  assign pksi_44_ = n_n2326;
  assign pksi_107_ = n_n2449;
  assign pksi_121_ = n_n2422;
  assign pksi_10_ = n_n2354;
  assign pksi_21_ = n_n2355;
  assign pksi_32_ = n_n2335;
  assign pksi_43_ = n_n2342;
  assign pksi_106_ = n_n2461;
  assign pksi_111_ = n_n2442;
  assign pksi_11_ = n_n2364;
  assign pksi_20_ = n_n2350;
  assign pksi_33_ = n_n2343;
  assign pksi_42_ = n_n2334;
  assign pksi_105_ = n_n2452;
  assign pksi_112_ = n_n2460;
  assign pksi_12_ = n_n2353;
  assign pksi_23_ = n_n2371;
  assign pksi_30_ = n_n2346;
  assign pksi_41_ = n_n2341;
  assign pksi_104_ = n_n2446;
  assign pksi_13_ = n_n2356;
  assign pksi_22_ = n_n2361;
  assign pksi_31_ = n_n2325;
  assign pksi_40_ = n_n2327;
  assign pksi_103_ = n_n2456;
  assign pksi_110_ = n_n2457;
  assign pksi_3_ = n_n2352;
  assign pksi_151_ = n_n2409;
  assign pksi_164_ = n_n2400;
  assign pksi_177_ = n_n2383;
  assign pksi_2_ = n_n2363;
  assign pksi_152_ = n_n2399;
  assign pksi_163_ = n_n2407;
  assign pksi_178_ = n_n2390;
  assign pksi_189_ = n_n2388;
  assign pksi_1_ = n_n2357;
  assign pksi_166_ = n_n2418;
  assign pksi_179_ = n_n2380;
  assign pksi_188_ = n_n2378;
  assign pksi_0_ = n_n2360;
  assign pksi_150_ = n_n2417;
  assign pksi_165_ = n_n2412;
  assign pksi_187_ = n_n2391;
  assign pksi_18_ = n_n2358;
  assign pksi_29_ = n_n2344;
  assign pksi_142_ = n_n2441;
  assign pksi_168_ = n_n2379;
  assign pksi_173_ = n_n2374;
  assign pksi_186_ = n_n2382;
  assign pksi_19_ = n_n2366;
  assign pksi_28_ = n_n2348;
  assign pksi_130_ = n_n2437;
  assign pksi_141_ = n_n2435;
  assign pksi_167_ = n_n2415;
  assign pksi_174_ = n_n2393;
  assign pksi_185_ = n_n2375;
  assign pksi_38_ = n_n2338;
  assign pksi_49_ = n_n2309;
  assign pksi_131_ = n_n2426;
  assign pksi_140_ = n_n2424;
  assign pksi_175_ = n_n2385;
  assign pksi_184_ = n_n2389;
  assign pksi_39_ = n_n2345;
  assign pksi_48_ = n_n2312;
  assign pksi_132_ = n_n2430;
  assign pksi_169_ = n_n2376;
  assign pksi_176_ = n_n2377;
  assign pksi_183_ = n_n2373;
  assign pksi_58_ = n_n2306;
  assign pksi_69_ = n_n2307;
  assign pksi_133_ = n_n2425;
  assign pksi_146_ = n_n2416;
  assign pksi_159_ = n_n2395;
  assign pksi_182_ = n_n2386;
  assign pksi_59_ = n_n2316;
  assign pksi_68_ = n_n2302;
  assign pksi_134_ = n_n2433;
  assign pksi_145_ = n_n2398;
  assign pksi_170_ = n_n2392;
  assign pksi_181_ = n_n2379;
  assign pksi_9_ = n_n2367;
  assign pksi_78_ = n_n2298;
  assign pksi_89_ = n_n2293;
  assign pksi_135_ = n_n2419;
  assign pksi_144_ = n_n2408;
  assign pksi_157_ = n_n2401;
  assign pksi_171_ = n_n2387;
  assign pksi_180_ = n_n2384;
  assign pksi_8_ = n_n2359;
  assign pksi_79_ = n_n2278;
  assign pksi_88_ = n_n2280;
  assign pksi_136_ = n_n2436;
  assign pksi_143_ = n_n2438;
  assign pksi_158_ = n_n2410;
  assign pksi_172_ = n_n2381;
  assign pksi_7_ = n_n2349;
  assign pksi_98_ = n_n2463;
  assign pksi_137_ = n_n2421;
  assign pksi_155_ = n_n2402;
  assign pksi_160_ = n_n2413;
  assign pksi_6_ = n_n2370;
  assign pksi_99_ = n_n2458;
  assign pksi_138_ = n_n2428;
  assign pksi_149_ = n_n2396;
  assign pksi_156_ = n_n2405;
  assign pksi_5_ = n_n2368;
  assign pksi_139_ = n_n2438;
  assign pksi_148_ = n_n2403;
  assign pksi_153_ = n_n2406;
  assign pksi_162_ = n_n2404;
  assign pksi_4_ = n_n2372;
  assign pksi_147_ = n_n2411;
  assign pksi_154_ = n_n2414;
  assign pksi_161_ = n_n2397;
  always @ (posedge clock) begin
    n_n2365 <= n922;
    n_n2375 <= n927;
    n_n2879 <= n932;
    n_n2392 <= n937;
    n_n2402 <= n942;
    n_n2411 <= n947;
    n_n2448 <= n952;
    n_n2982 <= n957;
    n_n2366 <= n962;
    n_n2865 <= n967;
    n_n2881 <= n972;
    n_n2391 <= n977;
    n_n2403 <= n982;
    n_n2917 <= n987;
    n_n2449 <= n992;
    n_n2457 <= n997;
    n_n2367 <= n1002;
    n_n2377 <= n1007;
    n_n2384 <= n1012;
    n_n2390 <= n1017;
    n_n2419 <= n1022;
    n_n2429 <= n1027;
    n_n2450 <= n1032;
    n_n2459 <= n1037;
    n_n2465 <= n1042;
    n_n2368 <= n1047;
    n_n2376 <= n1052;
    n_n2877 <= n1057;
    n_n2389 <= n1062;
    n_n2420 <= n1067;
    n_n2428 <= n1072;
    n_n2451 <= n1077;
    n_n2458 <= n1082;
    n_n2285 <= n1087;
    n_n2362 <= n1092;
    n_n2372 <= n1097;
    n_n2382 <= n1102;
    n_n2889 <= n1107;
    n_n2435 <= n1112;
    n_n2444 <= n1117;
    n_n2454 <= n1122;
    n_n2463 <= n1127;
    n_n2363 <= n1132;
    n_n2371 <= n1137;
    n_n2383 <= n1142;
    n_n2388 <= n1147;
    n_n2954 <= n1152;
    n_n2964 <= n1157;
    n_n2445 <= n1162;
    n_n2464 <= n1167;
    n_n2364 <= n1172;
    n_n2374 <= n1177;
    n_n2380 <= n1182;
    n_n2387 <= n1187;
    n_n2446 <= n1192;
    n_n2456 <= n1197;
    n_n2853 <= n1202;
    n_n2373 <= n1207;
    n_n2381 <= n1212;
    n_n2885 <= n1217;
    n_n2447 <= n1222;
    n_n2455 <= n1227;
    n_n2462 <= n1232;
    n_n2282 <= n1237;
    n_n2395 <= n1242;
    n_n2909 <= n1247;
    n_n2413 <= n1252;
    n_n2423 <= n1257;
    n_n2432 <= n1262;
    n_n2441 <= n1267;
    n_n2741 <= n1272;
    n_n2396 <= n1277;
    n_n2404 <= n1282;
    n_n2414 <= n1287;
    n_n2422 <= n1292;
    n_n2433 <= n1297;
    n_n2440 <= n1302;
    n_n2283 <= n1307;
    n_n2899 <= n1312;
    n_n2406 <= n1317;
    n_n2412 <= n1322;
    n_n2421 <= n1327;
    n_n2950 <= n1332;
    n_n2443 <= n1337;
    n_n2284 <= n1342;
    n_n2397 <= n1347;
    n_n2405 <= n1352;
    n_n2921 <= n1357;
    n_n2931 <= n1362;
    n_n2434 <= n1367;
    n_n2442 <= n1372;
    n_n2279 <= n1377;
    n_n2369 <= n1382;
    n_n2379 <= n1387;
    n_n2398 <= n1392;
    n_n2408 <= n1397;
    n_n2417 <= n1402;
    n_n2427 <= n1407;
    n_n2430 <= n1412;
    n_n2437 <= n1417;
    n_n2452 <= n1422;
    n_n2460 <= n1427;
    n_n2280 <= n1432;
    n_n2370 <= n1437;
    n_n2378 <= n1442;
    n_n2399 <= n1447;
    n_n2407 <= n1452;
    n_n2418 <= n1457;
    n_n2426 <= n1462;
    n_n2943 <= n1467;
    n_n2436 <= n1472;
    n_n2453 <= n1477;
    n_n2986 <= n1482;
    n_n2737 <= n1487;
    n_n2385 <= n1492;
    n_n2394 <= n1497;
    n_n2400 <= n1502;
    n_n2410 <= n1507;
    n_n2415 <= n1512;
    n_n2425 <= n1517;
    n_n2945 <= n1522;
    n_n2439 <= n1527;
    n_n2976 <= n1532;
    n_n2281 <= n1537;
    n_n2386 <= n1542;
    n_n2393 <= n1547;
    n_n2401 <= n1552;
    n_n2409 <= n1557;
    n_n2416 <= n1562;
    n_n2424 <= n1567;
    n_n2431 <= n1572;
    n_n2438 <= n1577;
    n_n2461 <= n1582;
    n_n2319 <= n1587;
    n_n2329 <= n1592;
    n_n2338 <= n1597;
    n_n2348 <= n1602;
    n_n2843 <= n1607;
    n_n2320 <= n1612;
    n_n2328 <= n1617;
    n_n2339 <= n1622;
    n_n2347 <= n1627;
    n_n2357 <= n1632;
    n_n2321 <= n1637;
    n_n2330 <= n1642;
    n_n2336 <= n1647;
    n_n2346 <= n1652;
    n_n2358 <= n1657;
    n_n2278 <= n1662;
    n_n2322 <= n1667;
    n_n2806 <= n1672;
    n_n2337 <= n1677;
    n_n2345 <= n1682;
    n_n2359 <= n1687;
    n_n2746 <= n1692;
    n_n2294 <= n1697;
    n_n2304 <= n1702;
    n_n2313 <= n1707;
    n_n2360 <= n1712;
    n_n2286 <= n1717;
    n_n2293 <= n1722;
    n_n2305 <= n1727;
    n_n2312 <= n1732;
    n_n2361 <= n1737;
    n_n2749 <= n1742;
    n_n2296 <= n1747;
    n_n2303 <= n1752;
    n_n2311 <= n1757;
    n_n2287 <= n1762;
    n_n2295 <= n1767;
    n_n2770 <= n1772;
    n_n2310 <= n1777;
    n_n2288 <= n1782;
    n_n2298 <= n1787;
    n_n2307 <= n1792;
    n_n2789 <= n1797;
    n_n2327 <= n1802;
    n_n2335 <= n1807;
    n_n2289 <= n1812;
    n_n2297 <= n1817;
    n_n2308 <= n1822;
    n_n2316 <= n1827;
    n_n2802 <= n1832;
    n_n2334 <= n1837;
    n_n2290 <= n1842;
    n_n2300 <= n1847;
    n_n2774 <= n1852;
    n_n2315 <= n1857;
    n_n2343 <= n1862;
    n_n2353 <= n1867;
    n_n2291 <= n1872;
    n_n2299 <= n1877;
    n_n2306 <= n1882;
    n_n2314 <= n1887;
    n_n2344 <= n1892;
    n_n2352 <= n1897;
    n_n2292 <= n1902;
    n_n2302 <= n1907;
    n_n2323 <= n1912;
    n_n2332 <= n1917;
    n_n2341 <= n1922;
    n_n2834 <= n1927;
    n_n2838 <= n1932;
    n_n2757 <= n1937;
    n_n2301 <= n1942;
    n_n2324 <= n1947;
    n_n2331 <= n1952;
    n_n2342 <= n1957;
    n_n2351 <= n1962;
    n_n2354 <= n1967;
    n_n2779 <= n1972;
    n_n2318 <= n1977;
    n_n2325 <= n1982;
    n_n2333 <= n1987;
    n_n2340 <= n1992;
    n_n2350 <= n1997;
    n_n2355 <= n2002;
    n_n2309 <= n2007;
    n_n2317 <= n2012;
    n_n2326 <= n2017;
    n_n2811 <= n2022;
    n_n2821 <= n2027;
    n_n2349 <= n2032;
    n_n2356 <= n2037;
  end
endmodule

