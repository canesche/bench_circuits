module top ( clock, 
    ck, g7, g6, g5, g4, g10, g3, g2, g12, g1, g11, g0, g13, g9, g8,
    g535, g546, g537, g548, g547, g539, g549, g551, g530, g552, g542, g532,
    g550, g45  );
  input  clock;
  input  ck, g7, g6, g5, g4, g10, g3, g2, g12, g1, g11, g0, g13, g9, g8;
  output g535, g546, g537, g548, g547, g539, g549, g551, g530, g552, g542,
    g532, g550, g45;
  reg ng38, ng39, ng36, ng35, ng37, ng42, ng43, ng40, ng41, ng30, ng46,
    ng29, ng44, ng45, ng34, ng33, ng32, ng31;
  wire new_n84_, new_n85_1_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_1_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_1_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n100_1_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_1_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_1_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_1_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_1_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_1_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_1_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_1_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_1_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_1_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n518_, new_n520_, new_n521_, new_n523_, new_n524_,
    new_n525_, new_n527_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n563_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n605_, new_n606_, new_n607_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, n60, n65, n70, n75, n80,
    n85, n90, n95, n100, n105, n110, n115, n120, n125, n130, n135, n140,
    n145;
  assign new_n84_ = g10 & ~g8;
  assign new_n85_1_ = ~g7 & ~g5;
  assign new_n86_ = g6 & ~g9;
  assign new_n87_ = ~g3 & new_n84_;
  assign new_n88_ = new_n85_1_ & new_n87_;
  assign new_n89_ = new_n86_ & new_n88_;
  assign new_n90_1_ = g5 & g3;
  assign new_n91_ = g7 & ~g10;
  assign new_n92_ = g8 & ng37;
  assign new_n93_ = new_n90_1_ & new_n92_;
  assign new_n94_ = new_n91_ & new_n93_;
  assign new_n95_1_ = ~new_n89_ & ~new_n94_;
  assign new_n96_ = ~g4 & ~g0;
  assign new_n97_ = g11 & ~new_n95_1_;
  assign new_n98_ = new_n96_ & new_n97_;
  assign new_n99_ = g6 & g4;
  assign new_n100_1_ = g11 & g9;
  assign new_n101_ = g8 & new_n100_1_;
  assign new_n102_ = g7 & g10;
  assign new_n103_ = new_n101_ & new_n102_;
  assign new_n104_ = new_n90_1_ & new_n99_;
  assign new_n105_1_ = new_n103_ & new_n104_;
  assign new_n106_ = g0 & new_n105_1_;
  assign new_n107_ = ~new_n98_ & ~new_n106_;
  assign new_n108_ = g2 & g1;
  assign new_n109_ = ~new_n107_ & new_n108_;
  assign new_n110_1_ = g7 & ~g6;
  assign new_n111_ = ng30 & new_n110_1_;
  assign new_n112_ = ~g10 & ~g11;
  assign new_n113_ = ~g9 & new_n112_;
  assign new_n114_ = g8 & ng31;
  assign new_n115_1_ = ~new_n111_ & new_n113_;
  assign new_n116_ = ~new_n114_ & new_n115_1_;
  assign new_n117_ = ~g6 & ~ng30;
  assign new_n118_ = g10 & g8;
  assign new_n119_ = g9 & ~new_n118_;
  assign new_n120_1_ = g8 & ~ng31;
  assign new_n121_ = ~new_n111_ & ~new_n119_;
  assign new_n122_ = new_n120_1_ & new_n121_;
  assign new_n123_ = g10 & new_n118_;
  assign new_n124_ = g9 & ~new_n123_;
  assign new_n125_1_ = ~g7 & ~g8;
  assign new_n126_ = ~new_n124_ & new_n125_1_;
  assign new_n127_ = ~new_n117_ & ~new_n122_;
  assign new_n128_ = ~new_n126_ & new_n127_;
  assign new_n129_ = g11 & ~new_n128_;
  assign new_n130_1_ = ~new_n84_ & ~new_n120_1_;
  assign new_n131_ = ~g7 & ~g11;
  assign new_n132_ = g9 & ~new_n130_1_;
  assign new_n133_ = new_n131_ & new_n132_;
  assign new_n134_ = g3 & new_n96_;
  assign new_n135_1_ = ~g3 & g0;
  assign new_n136_ = ~g2 & new_n135_1_;
  assign new_n137_ = g5 & ~g1;
  assign new_n138_ = g4 & ~new_n90_1_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_1_ = g2 & ~new_n139_;
  assign new_n141_ = ~g3 & ~new_n140_1_;
  assign new_n142_ = g0 & ~new_n141_;
  assign new_n143_ = ~g4 & ~new_n142_;
  assign new_n144_ = ~new_n136_ & ~new_n143_;
  assign new_n145_1_ = ~g5 & ~new_n144_;
  assign new_n146_ = ~new_n134_ & ~new_n145_1_;
  assign new_n147_ = ~g5 & g4;
  assign new_n148_ = ~new_n146_ & ~new_n147_;
  assign new_n149_ = ~new_n116_ & ~new_n129_;
  assign new_n150_ = ~new_n133_ & ~new_n148_;
  assign new_n151_ = new_n149_ & new_n150_;
  assign new_n152_ = ng46 & new_n151_;
  assign new_n153_ = g12 & ~g13;
  assign new_n154_ = ~new_n152_ & new_n153_;
  assign new_n155_ = new_n109_ & new_n154_;
  assign new_n156_ = g1 & new_n90_1_;
  assign new_n157_ = g8 & new_n155_;
  assign new_n158_ = new_n156_ & new_n157_;
  assign new_n159_ = ng37 & new_n158_;
  assign new_n160_ = ng38 & new_n159_;
  assign new_n161_ = g3 & g1;
  assign new_n162_ = ~g4 & new_n161_;
  assign new_n163_ = g6 & new_n162_;
  assign new_n164_ = g3 & new_n99_;
  assign new_n165_ = ~g1 & new_n164_;
  assign new_n166_ = ~new_n163_ & ~new_n165_;
  assign new_n167_ = new_n84_ & new_n100_1_;
  assign new_n168_ = ~new_n166_ & new_n167_;
  assign new_n169_ = ~g10 & new_n101_;
  assign new_n170_ = new_n165_ & new_n169_;
  assign new_n171_ = ~new_n168_ & ~new_n170_;
  assign new_n172_ = ~g7 & ~new_n171_;
  assign new_n173_ = ~g6 & ~g4;
  assign new_n174_ = g3 & ~g1;
  assign new_n175_ = ~g8 & new_n173_;
  assign new_n176_ = new_n174_ & new_n175_;
  assign new_n177_ = g8 & ~new_n166_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~g9 & new_n91_;
  assign new_n180_ = g11 & new_n179_;
  assign new_n181_ = ~new_n178_ & new_n180_;
  assign new_n182_ = ~new_n172_ & ~new_n181_;
  assign new_n183_ = ~g5 & g2;
  assign new_n184_ = ~new_n182_ & new_n183_;
  assign new_n185_ = g2 & new_n99_;
  assign new_n186_ = ~g10 & g9;
  assign new_n187_ = ~g8 & new_n131_;
  assign new_n188_ = new_n186_ & new_n187_;
  assign new_n189_ = ~new_n103_ & ~new_n188_;
  assign new_n190_ = new_n185_ & ~new_n189_;
  assign new_n191_ = new_n156_ & new_n190_;
  assign new_n192_ = ~new_n184_ & ~new_n191_;
  assign new_n193_ = g4 & g1;
  assign new_n194_ = ~g5 & ~new_n193_;
  assign new_n195_ = g2 & ~new_n194_;
  assign new_n196_ = ~g6 & new_n195_;
  assign new_n197_ = ~g3 & g2;
  assign new_n198_ = g3 & ~g2;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = ~new_n138_ & new_n199_;
  assign new_n201_ = g6 & ~new_n200_;
  assign new_n202_ = ~g3 & new_n147_;
  assign new_n203_ = g3 & ~new_n99_;
  assign new_n204_ = ~new_n173_ & ~new_n203_;
  assign new_n205_ = g5 & ~new_n204_;
  assign new_n206_ = ~new_n201_ & ~new_n202_;
  assign new_n207_ = ~new_n205_ & new_n206_;
  assign new_n208_ = g1 & ~new_n207_;
  assign new_n209_ = g6 & ~g4;
  assign new_n210_ = ~g5 & ~new_n209_;
  assign new_n211_ = g2 & ~g1;
  assign new_n212_ = ~new_n210_ & new_n211_;
  assign new_n213_ = ~new_n196_ & ~new_n208_;
  assign new_n214_ = ~new_n212_ & new_n213_;
  assign new_n215_ = ~new_n101_ & new_n102_;
  assign new_n216_ = ~g7 & g8;
  assign new_n217_ = ng30 & new_n216_;
  assign new_n218_ = g7 & new_n186_;
  assign new_n219_ = ~new_n215_ & ~new_n217_;
  assign new_n220_ = ~new_n218_ & new_n219_;
  assign new_n221_ = ~new_n214_ & ~new_n220_;
  assign new_n222_ = g13 & ~new_n192_;
  assign new_n223_ = ~new_n221_ & new_n222_;
  assign new_n224_ = ~g1 & new_n223_;
  assign new_n225_ = ~g7 & new_n186_;
  assign new_n226_ = ~new_n179_ & ~new_n225_;
  assign new_n227_ = g8 & ~new_n226_;
  assign new_n228_ = new_n147_ & new_n224_;
  assign new_n229_ = new_n227_ & new_n228_;
  assign new_n230_ = g1 & new_n223_;
  assign new_n231_ = ~g5 & ~g4;
  assign new_n232_ = g3 & ng35;
  assign new_n233_ = g11 & new_n232_;
  assign new_n234_ = new_n231_ & new_n233_;
  assign new_n235_ = g5 & new_n188_;
  assign new_n236_ = new_n164_ & new_n235_;
  assign new_n237_ = ~new_n105_1_ & ~new_n234_;
  assign new_n238_ = ~new_n236_ & new_n237_;
  assign new_n239_ = g2 & ~new_n238_;
  assign new_n240_ = new_n186_ & new_n216_;
  assign new_n241_ = ~g7 & g9;
  assign new_n242_ = new_n84_ & new_n241_;
  assign new_n243_ = g8 & new_n179_;
  assign new_n244_ = ~new_n242_ & ~new_n243_;
  assign new_n245_ = ~new_n240_ & new_n244_;
  assign new_n246_ = ~g5 & g11;
  assign new_n247_ = new_n164_ & new_n246_;
  assign new_n248_ = ~g2 & ~new_n245_;
  assign new_n249_ = new_n247_ & new_n248_;
  assign new_n250_ = ~g6 & ng36;
  assign new_n251_ = g5 & new_n99_;
  assign new_n252_ = g11 & ~new_n244_;
  assign new_n253_ = new_n251_ & new_n252_;
  assign new_n254_ = ~new_n250_ & ~new_n253_;
  assign new_n255_ = ~g3 & ~new_n254_;
  assign new_n256_ = ~g2 & new_n255_;
  assign new_n257_ = ~new_n239_ & ~new_n249_;
  assign new_n258_ = ~new_n256_ & new_n257_;
  assign new_n259_ = ng32 & ~new_n220_;
  assign new_n260_ = ~g13 & ~new_n259_;
  assign new_n261_ = ~new_n258_ & new_n260_;
  assign new_n262_ = ~new_n230_ & ~new_n261_;
  assign new_n263_ = ~g5 & ~new_n244_;
  assign new_n264_ = ~g4 & new_n263_;
  assign new_n265_ = ~new_n262_ & new_n264_;
  assign new_n266_ = ~new_n229_ & ~new_n265_;
  assign new_n267_ = g6 & g3;
  assign new_n268_ = ~g12 & ~new_n266_;
  assign new_n269_ = new_n267_ & new_n268_;
  assign new_n270_ = ~new_n160_ & ~new_n269_;
  assign new_n271_ = g2 & g11;
  assign new_n272_ = ~new_n270_ & new_n271_;
  assign new_n273_ = new_n227_ & new_n247_;
  assign new_n274_ = ~g3 & ~ng44;
  assign new_n275_ = ~new_n273_ & ~new_n274_;
  assign new_n276_ = ~g2 & new_n261_;
  assign new_n277_ = ~g12 & new_n276_;
  assign new_n278_ = ~new_n275_ & new_n277_;
  assign g535 = new_n272_ | new_n278_;
  assign new_n280_ = new_n231_ & new_n267_;
  assign new_n281_ = new_n179_ & new_n280_;
  assign new_n282_ = g9 & new_n102_;
  assign new_n283_ = new_n99_ & new_n282_;
  assign new_n284_ = new_n90_1_ & new_n283_;
  assign new_n285_ = ~new_n281_ & ~new_n284_;
  assign new_n286_ = g8 & ~new_n262_;
  assign new_n287_ = ~new_n285_ & new_n286_;
  assign new_n288_ = new_n164_ & new_n263_;
  assign new_n289_ = new_n224_ & new_n288_;
  assign new_n290_ = ~new_n287_ & ~new_n289_;
  assign new_n291_ = ~g12 & ~new_n290_;
  assign new_n292_ = ng38 & new_n86_;
  assign new_n293_ = g0 & new_n283_;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign new_n295_ = new_n158_ & ~new_n294_;
  assign new_n296_ = ~new_n291_ & ~new_n295_;
  assign new_n297_ = new_n271_ & ~new_n296_;
  assign new_n298_ = ~g6 & new_n102_;
  assign new_n299_ = new_n101_ & new_n147_;
  assign new_n300_ = new_n298_ & new_n299_;
  assign new_n301_ = ~g5 & new_n173_;
  assign new_n302_ = new_n112_ & new_n301_;
  assign new_n303_ = g10 & new_n100_1_;
  assign new_n304_ = new_n251_ & new_n303_;
  assign new_n305_ = ~new_n302_ & ~new_n304_;
  assign new_n306_ = new_n125_1_ & ~new_n305_;
  assign new_n307_ = ~new_n300_ & ~new_n306_;
  assign new_n308_ = ~g3 & ~new_n307_;
  assign new_n309_ = g11 & new_n288_;
  assign new_n310_ = ~new_n308_ & ~new_n309_;
  assign new_n311_ = new_n277_ & ~new_n310_;
  assign g537 = new_n297_ | new_n311_;
  assign new_n313_ = g12 & new_n152_;
  assign new_n314_ = ~g13 & new_n313_;
  assign new_n315_ = ~ng42 & new_n314_;
  assign new_n316_ = g7 & ~new_n118_;
  assign new_n317_ = new_n100_1_ & new_n316_;
  assign new_n318_ = ~g9 & new_n102_;
  assign new_n319_ = ~new_n186_ & new_n216_;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign new_n321_ = g11 & ~new_n320_;
  assign new_n322_ = ~new_n317_ & ~new_n321_;
  assign new_n323_ = ng34 & ~new_n322_;
  assign g548 = new_n315_ | new_n323_;
  assign new_n325_ = ~g7 & new_n118_;
  assign new_n326_ = ~new_n316_ & ~new_n325_;
  assign new_n327_ = g9 & ~new_n326_;
  assign new_n328_ = ng34 & new_n327_;
  assign new_n329_ = g9 & new_n298_;
  assign new_n330_ = g10 & g9;
  assign new_n331_ = ~g10 & g11;
  assign new_n332_ = ~new_n330_ & ~new_n331_;
  assign new_n333_ = new_n216_ & ~new_n332_;
  assign new_n334_ = ~g8 & new_n100_1_;
  assign new_n335_ = new_n186_ & ~new_n216_;
  assign new_n336_ = ~new_n333_ & ~new_n334_;
  assign new_n337_ = ~new_n335_ & new_n336_;
  assign new_n338_ = g6 & ~new_n337_;
  assign new_n339_ = ~new_n329_ & ~new_n338_;
  assign new_n340_ = new_n314_ & ~new_n339_;
  assign g547 = new_n328_ | new_n340_;
  assign new_n342_ = ~new_n109_ & new_n154_;
  assign new_n343_ = ~g12 & new_n258_;
  assign new_n344_ = new_n260_ & new_n343_;
  assign new_n345_ = ~g12 & g13;
  assign new_n346_ = ~new_n221_ & new_n345_;
  assign new_n347_ = new_n192_ & new_n346_;
  assign new_n348_ = ~new_n342_ & ~new_n344_;
  assign g539 = new_n347_ | ~new_n348_;
  assign new_n350_ = g3 & g0;
  assign new_n351_ = new_n193_ & ~new_n350_;
  assign new_n352_ = new_n314_ & new_n351_;
  assign new_n353_ = g2 & new_n147_;
  assign new_n354_ = ~g3 & new_n99_;
  assign new_n355_ = ~new_n198_ & ~new_n354_;
  assign new_n356_ = g5 & ~new_n355_;
  assign new_n357_ = ~g6 & g5;
  assign new_n358_ = g6 & new_n197_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = ~new_n90_1_ & new_n359_;
  assign new_n361_ = ~g4 & ~new_n360_;
  assign new_n362_ = ~new_n353_ & ~new_n356_;
  assign new_n363_ = ~new_n361_ & new_n362_;
  assign new_n364_ = g1 & new_n221_;
  assign new_n365_ = new_n345_ & ~new_n363_;
  assign new_n366_ = new_n364_ & new_n365_;
  assign new_n367_ = g5 & g2;
  assign new_n368_ = g4 & g3;
  assign new_n369_ = ~g12 & new_n259_;
  assign new_n370_ = ~g13 & new_n369_;
  assign new_n371_ = new_n367_ & ~new_n368_;
  assign new_n372_ = new_n370_ & new_n371_;
  assign new_n373_ = g3 & ~g13;
  assign new_n374_ = ~ng33 & new_n373_;
  assign new_n375_ = ~new_n352_ & ~new_n366_;
  assign new_n376_ = ~new_n372_ & ~new_n374_;
  assign g549 = ~new_n375_ | ~new_n376_;
  assign new_n378_ = g2 & g0;
  assign new_n379_ = g1 & ~new_n378_;
  assign new_n380_ = g4 & new_n378_;
  assign new_n381_ = ~new_n379_ & ~new_n380_;
  assign new_n382_ = ~g3 & ~new_n381_;
  assign new_n383_ = ~new_n193_ & new_n350_;
  assign new_n384_ = ~g0 & new_n193_;
  assign new_n385_ = ~new_n382_ & ~new_n383_;
  assign new_n386_ = ~new_n384_ & new_n385_;
  assign new_n387_ = g5 & ~new_n386_;
  assign new_n388_ = new_n314_ & new_n387_;
  assign new_n389_ = g4 & ng39;
  assign new_n390_ = new_n370_ & new_n389_;
  assign new_n391_ = g4 & g2;
  assign new_n392_ = ~g1 & new_n391_;
  assign new_n393_ = new_n221_ & new_n392_;
  assign new_n394_ = new_n193_ & new_n221_;
  assign new_n395_ = new_n198_ & new_n394_;
  assign new_n396_ = ~new_n393_ & ~new_n395_;
  assign new_n397_ = g5 & ~new_n396_;
  assign new_n398_ = new_n147_ & ~new_n198_;
  assign new_n399_ = g6 & new_n198_;
  assign new_n400_ = ~g5 & new_n399_;
  assign new_n401_ = ~new_n398_ & ~new_n400_;
  assign new_n402_ = ~new_n354_ & new_n401_;
  assign new_n403_ = new_n364_ & ~new_n402_;
  assign new_n404_ = ~new_n397_ & ~new_n403_;
  assign new_n405_ = new_n345_ & ~new_n404_;
  assign new_n406_ = ~new_n388_ & ~new_n390_;
  assign g551 = new_n405_ | ~new_n406_;
  assign new_n408_ = g5 & ~g3;
  assign new_n409_ = ~g4 & ~new_n408_;
  assign new_n410_ = g1 & ~g0;
  assign new_n411_ = ~new_n409_ & new_n410_;
  assign new_n412_ = ~g4 & new_n90_1_;
  assign new_n413_ = ~g5 & new_n161_;
  assign new_n414_ = ~new_n412_ & ~new_n413_;
  assign new_n415_ = new_n139_ & new_n414_;
  assign new_n416_ = g0 & ~new_n415_;
  assign new_n417_ = ~new_n411_ & ~new_n416_;
  assign new_n418_ = g2 & ~new_n417_;
  assign new_n419_ = new_n314_ & new_n418_;
  assign new_n420_ = new_n255_ & new_n277_;
  assign g530 = new_n419_ | new_n420_;
  assign new_n422_ = ~ng40 & new_n314_;
  assign new_n423_ = g1 & ~new_n367_;
  assign new_n424_ = new_n99_ & new_n423_;
  assign new_n425_ = ~g4 & ~g3;
  assign new_n426_ = ~g1 & ~new_n147_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = g2 & ~new_n427_;
  assign new_n429_ = ~g4 & g1;
  assign new_n430_ = new_n90_1_ & new_n429_;
  assign new_n431_ = ~new_n428_ & ~new_n430_;
  assign new_n432_ = g6 & ~new_n431_;
  assign new_n433_ = ~new_n424_ & ~new_n432_;
  assign new_n434_ = new_n221_ & ~new_n433_;
  assign new_n435_ = new_n345_ & new_n434_;
  assign new_n436_ = ~new_n147_ & new_n399_;
  assign new_n437_ = g5 & ~g4;
  assign new_n438_ = ~new_n147_ & ~new_n437_;
  assign new_n439_ = g6 & ~new_n438_;
  assign new_n440_ = ~new_n354_ & ~new_n439_;
  assign new_n441_ = g2 & ~new_n440_;
  assign new_n442_ = ~new_n436_ & ~new_n441_;
  assign new_n443_ = new_n370_ & ~new_n442_;
  assign new_n444_ = ~new_n422_ & ~new_n435_;
  assign g552 = new_n443_ | ~new_n444_;
  assign new_n446_ = g7 & g9;
  assign new_n447_ = new_n118_ & ~new_n446_;
  assign new_n448_ = g7 & ~g8;
  assign new_n449_ = g11 & new_n448_;
  assign new_n450_ = g10 & ~g11;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = ~g9 & ~new_n451_;
  assign new_n453_ = ~new_n167_ & ~new_n447_;
  assign new_n454_ = ~new_n452_ & new_n453_;
  assign new_n455_ = g6 & new_n314_;
  assign new_n456_ = ~new_n454_ & new_n455_;
  assign new_n457_ = g9 & g8;
  assign new_n458_ = new_n102_ & ~new_n457_;
  assign new_n459_ = ng34 & new_n458_;
  assign new_n460_ = g8 & ng34;
  assign new_n461_ = ~new_n455_ & ~new_n460_;
  assign new_n462_ = new_n218_ & ~new_n461_;
  assign new_n463_ = ~new_n456_ & ~new_n459_;
  assign g542 = new_n462_ | ~new_n463_;
  assign new_n465_ = ~g2 & g1;
  assign new_n466_ = new_n408_ & new_n465_;
  assign new_n467_ = g2 & ~new_n161_;
  assign new_n468_ = ~g5 & ~g3;
  assign new_n469_ = ~g2 & new_n90_1_;
  assign new_n470_ = ~new_n467_ & ~new_n468_;
  assign new_n471_ = ~new_n469_ & new_n470_;
  assign new_n472_ = g4 & ~new_n471_;
  assign new_n473_ = ~new_n162_ & ~new_n466_;
  assign new_n474_ = ~new_n472_ & new_n473_;
  assign new_n475_ = g0 & ~new_n474_;
  assign new_n476_ = new_n314_ & new_n475_;
  assign new_n477_ = g11 & new_n264_;
  assign new_n478_ = g4 & new_n235_;
  assign new_n479_ = ~new_n477_ & ~new_n478_;
  assign new_n480_ = g2 & ~new_n479_;
  assign new_n481_ = ~new_n262_ & new_n480_;
  assign new_n482_ = new_n267_ & new_n481_;
  assign new_n483_ = g13 & new_n221_;
  assign new_n484_ = ~ng43 & new_n483_;
  assign new_n485_ = g3 & new_n224_;
  assign new_n486_ = new_n185_ & new_n485_;
  assign new_n487_ = new_n164_ & new_n276_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = new_n167_ & ~new_n488_;
  assign new_n490_ = new_n85_1_ & new_n489_;
  assign new_n491_ = g8 & new_n180_;
  assign new_n492_ = new_n251_ & new_n491_;
  assign new_n493_ = ng36 & new_n173_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = ~g3 & ~new_n494_;
  assign new_n496_ = new_n276_ & new_n495_;
  assign new_n497_ = ~new_n482_ & ~new_n484_;
  assign new_n498_ = ~new_n490_ & ~new_n496_;
  assign new_n499_ = new_n497_ & new_n498_;
  assign new_n500_ = ~g12 & ~new_n499_;
  assign g532 = new_n476_ | new_n500_;
  assign new_n502_ = g5 & ~new_n193_;
  assign new_n503_ = new_n221_ & new_n502_;
  assign new_n504_ = ~g5 & new_n394_;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = g2 & ~new_n505_;
  assign new_n507_ = new_n345_ & new_n506_;
  assign new_n508_ = g3 & new_n384_;
  assign new_n509_ = g0 & ~ng29;
  assign new_n510_ = ~new_n508_ & ~new_n509_;
  assign new_n511_ = new_n314_ & ~new_n510_;
  assign new_n512_ = new_n90_1_ & ~new_n391_;
  assign new_n513_ = new_n370_ & new_n512_;
  assign new_n514_ = ~new_n507_ & ~new_n511_;
  assign new_n515_ = ~new_n374_ & ~new_n513_;
  assign g550 = ~new_n514_ | ~new_n515_;
  assign n60 = new_n91_ & new_n96_;
  assign new_n518_ = g2 & ~new_n90_1_;
  assign n65 = new_n469_ | new_n518_;
  assign new_n520_ = ~g10 & new_n187_;
  assign new_n521_ = ~new_n103_ & ~new_n520_;
  assign n70 = ~g5 & ~new_n521_;
  assign new_n523_ = ~g6 & ~g8;
  assign new_n524_ = new_n179_ & new_n523_;
  assign new_n525_ = g6 & ~new_n244_;
  assign n75 = new_n524_ | new_n525_;
  assign new_n527_ = ~g6 & g9;
  assign n80 = new_n86_ | new_n527_;
  assign new_n529_ = g6 & ~new_n102_;
  assign new_n530_ = new_n100_1_ & new_n529_;
  assign new_n531_ = new_n110_1_ & ~new_n186_;
  assign new_n532_ = g6 & new_n118_;
  assign new_n533_ = ~new_n448_ & ~new_n532_;
  assign new_n534_ = ~g9 & ~new_n533_;
  assign new_n535_ = ~new_n531_ & ~new_n534_;
  assign new_n536_ = g11 & ~new_n535_;
  assign n85 = ~new_n530_ & ~new_n536_;
  assign new_n538_ = g6 & new_n147_;
  assign new_n539_ = ~g6 & new_n391_;
  assign new_n540_ = g5 & ~new_n99_;
  assign new_n541_ = ~new_n538_ & ~new_n539_;
  assign new_n542_ = ~new_n540_ & new_n541_;
  assign new_n543_ = new_n161_ & ~new_n542_;
  assign new_n544_ = g1 & new_n399_;
  assign new_n545_ = g3 & new_n212_;
  assign new_n546_ = ~new_n543_ & ~new_n544_;
  assign n90 = ~new_n545_ & new_n546_;
  assign new_n548_ = g6 & g9;
  assign new_n549_ = ~g11 & new_n548_;
  assign new_n550_ = ~g6 & ng30;
  assign new_n551_ = ~new_n549_ & ~new_n550_;
  assign new_n552_ = g7 & ~new_n551_;
  assign new_n553_ = g6 & ng31;
  assign new_n554_ = ~new_n552_ & ~new_n553_;
  assign new_n555_ = g8 & ~new_n554_;
  assign new_n556_ = g6 & new_n169_;
  assign n95 = ~new_n555_ & ~new_n556_;
  assign new_n558_ = ng34 & new_n447_;
  assign new_n559_ = new_n102_ & ~new_n548_;
  assign new_n560_ = new_n314_ & new_n559_;
  assign new_n561_ = ~new_n558_ & ~new_n560_;
  assign n100 = ~new_n462_ & new_n561_;
  assign new_n563_ = g11 & ~g9;
  assign n105 = g10 | new_n563_;
  assign new_n565_ = ~g5 & new_n174_;
  assign new_n566_ = g0 & ~new_n147_;
  assign new_n567_ = g1 & ~new_n566_;
  assign new_n568_ = g4 & ~new_n567_;
  assign new_n569_ = new_n90_1_ & new_n568_;
  assign new_n570_ = new_n135_1_ & ~new_n147_;
  assign new_n571_ = ~new_n565_ & ~new_n569_;
  assign new_n572_ = ~new_n570_ & new_n571_;
  assign new_n573_ = g2 & new_n139_;
  assign new_n574_ = ~new_n572_ & new_n573_;
  assign new_n575_ = ~g10 & new_n117_;
  assign new_n576_ = ~g7 & ~g6;
  assign new_n577_ = new_n141_ & ~new_n147_;
  assign new_n578_ = new_n198_ & ~new_n437_;
  assign new_n579_ = new_n147_ & new_n578_;
  assign new_n580_ = ~new_n577_ & ~new_n579_;
  assign new_n581_ = g0 & new_n580_;
  assign new_n582_ = ~g1 & ~new_n581_;
  assign new_n583_ = ~new_n574_ & ~new_n575_;
  assign new_n584_ = ~new_n576_ & ~new_n582_;
  assign n110 = new_n583_ & new_n584_;
  assign new_n586_ = ~new_n147_ & new_n198_;
  assign new_n587_ = ~new_n368_ & ~new_n437_;
  assign new_n588_ = new_n211_ & ~new_n587_;
  assign n115 = ~new_n586_ & ~new_n588_;
  assign new_n590_ = new_n103_ & new_n301_;
  assign new_n591_ = ~g6 & ~g5;
  assign new_n592_ = new_n113_ & new_n591_;
  assign new_n593_ = ~new_n304_ & ~new_n592_;
  assign new_n594_ = new_n125_1_ & ~new_n593_;
  assign n120 = ~new_n590_ & ~new_n594_;
  assign new_n596_ = ~g12 & new_n261_;
  assign new_n597_ = ~new_n192_ & new_n346_;
  assign new_n598_ = ~new_n155_ & ~new_n596_;
  assign n125 = new_n597_ | ~new_n598_;
  assign new_n600_ = g13 & ~new_n214_;
  assign new_n601_ = ~g13 & ng32;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = ~g12 & ~new_n602_;
  assign n130 = ~new_n220_ & new_n603_;
  assign new_n605_ = g0 & new_n429_;
  assign new_n606_ = new_n313_ & new_n605_;
  assign new_n607_ = new_n353_ & new_n369_;
  assign n135 = ~new_n606_ & ~new_n607_;
  assign new_n609_ = new_n198_ & ~new_n210_;
  assign new_n610_ = ~new_n164_ & new_n367_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign n140 = new_n353_ | ~new_n611_;
  assign new_n613_ = g10 & ~new_n100_1_;
  assign new_n614_ = ~g7 & g11;
  assign n145 = new_n613_ | new_n614_;
  assign g546 = ~ng41;
  assign g45 = ng45;
  always @ (posedge clock) begin
    ng38 <= n60;
    ng39 <= n65;
    ng36 <= n70;
    ng35 <= n75;
    ng37 <= n80;
    ng42 <= n85;
    ng43 <= n90;
    ng40 <= n95;
    ng41 <= n100;
    ng30 <= n105;
    ng46 <= n110;
    ng29 <= n115;
    ng44 <= n120;
    ng45 <= n125;
    ng34 <= n130;
    ng33 <= n135;
    ng32 <= n140;
    ng31 <= n145;
  end
endmodule

