// Benchmark "mem_ctrl" written by ABC on Thu Oct  8 22:04:11 2020

module mem_ctrl ( clock, 
    clk_i, rst_i, wb_we_i, wb_cyc_i, wb_stb_i, susp_req_i, resume_req_i,
    mc_clk_i, mc_br_pad_i, mc_ack_pad_i, mc_sts_pad_i, \wb_data_i[0] ,
    \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] , \wb_data_i[4] ,
    \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] , \wb_data_i[8] ,
    \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] , \wb_data_i[12] ,
    \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] , \wb_data_i[16] ,
    \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] , \wb_data_i[20] ,
    \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] , \wb_data_i[24] ,
    \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] , \wb_data_i[28] ,
    \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] , \wb_addr_i[0] ,
    \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] , \wb_addr_i[4] ,
    \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] , \wb_addr_i[8] ,
    \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] , \wb_addr_i[12] ,
    \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] , \wb_addr_i[16] ,
    \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] , \wb_addr_i[20] ,
    \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] , \wb_addr_i[24] ,
    \wb_addr_i[25] , \wb_addr_i[26] , \wb_addr_i[27] , \wb_addr_i[28] ,
    \wb_addr_i[29] , \wb_addr_i[30] , \wb_addr_i[31] , \mc_data_pad_i[0] ,
    \mc_data_pad_i[1] , \mc_data_pad_i[2] , \mc_data_pad_i[3] ,
    \mc_data_pad_i[4] , \mc_data_pad_i[5] , \mc_data_pad_i[6] ,
    \mc_data_pad_i[7] , \mc_data_pad_i[8] , \mc_data_pad_i[9] ,
    \mc_data_pad_i[10] , \mc_data_pad_i[11] , \mc_data_pad_i[12] ,
    \mc_data_pad_i[13] , \mc_data_pad_i[14] , \mc_data_pad_i[15] ,
    \mc_data_pad_i[16] , \mc_data_pad_i[17] , \mc_data_pad_i[18] ,
    \mc_data_pad_i[19] , \mc_data_pad_i[20] , \mc_data_pad_i[21] ,
    \mc_data_pad_i[22] , \mc_data_pad_i[23] , \mc_data_pad_i[24] ,
    \mc_data_pad_i[25] , \mc_data_pad_i[26] , \mc_data_pad_i[27] ,
    \mc_data_pad_i[28] , \mc_data_pad_i[29] , \mc_data_pad_i[30] ,
    \mc_data_pad_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] ,
    \wb_sel_i[3] , \mc_dp_pad_i[0] , \mc_dp_pad_i[1] , \mc_dp_pad_i[2] ,
    \mc_dp_pad_i[3] ,
    \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] ,
    \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] ,
    \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] ,
    \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] ,
    \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] ,
    \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] ,
    \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] ,
    \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] ,
    \poc_o[0] , \poc_o[1] , \poc_o[2] , \poc_o[3] , \poc_o[4] , \poc_o[5] ,
    \poc_o[6] , \poc_o[7] , \poc_o[8] , \poc_o[9] , \poc_o[10] ,
    \poc_o[11] , \poc_o[12] , \poc_o[13] , \poc_o[14] , \poc_o[15] ,
    \poc_o[16] , \poc_o[17] , \poc_o[18] , \poc_o[19] , \poc_o[20] ,
    \poc_o[21] , \poc_o[22] , \poc_o[23] , \poc_o[24] , \poc_o[25] ,
    \poc_o[26] , \poc_o[27] , \poc_o[28] , \poc_o[29] , \poc_o[30] ,
    \poc_o[31] , \mc_data_pad_o[0] , \mc_data_pad_o[1] ,
    \mc_data_pad_o[2] , \mc_data_pad_o[3] , \mc_data_pad_o[4] ,
    \mc_data_pad_o[5] , \mc_data_pad_o[6] , \mc_data_pad_o[7] ,
    \mc_data_pad_o[8] , \mc_data_pad_o[9] , \mc_data_pad_o[10] ,
    \mc_data_pad_o[11] , \mc_data_pad_o[12] , \mc_data_pad_o[13] ,
    \mc_data_pad_o[14] , \mc_data_pad_o[15] , \mc_data_pad_o[16] ,
    \mc_data_pad_o[17] , \mc_data_pad_o[18] , \mc_data_pad_o[19] ,
    \mc_data_pad_o[20] , \mc_data_pad_o[21] , \mc_data_pad_o[22] ,
    \mc_data_pad_o[23] , \mc_data_pad_o[24] , \mc_data_pad_o[25] ,
    \mc_data_pad_o[26] , \mc_data_pad_o[27] , \mc_data_pad_o[28] ,
    \mc_data_pad_o[29] , \mc_data_pad_o[30] , \mc_data_pad_o[31] ,
    wb_ack_o, wb_err_o, suspended_o, mc_bg_pad_o, mc_doe_pad_doe_o,
    mc_oe_pad_o_, mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_,
    mc_cke_pad_o_, mc_rp_pad_o_, mc_vpen_pad_o, mc_adsc_pad_o_,
    mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o, \mc_addr_pad_o[0] ,
    \mc_addr_pad_o[1] , \mc_addr_pad_o[2] , \mc_addr_pad_o[3] ,
    \mc_addr_pad_o[4] , \mc_addr_pad_o[5] , \mc_addr_pad_o[6] ,
    \mc_addr_pad_o[7] , \mc_addr_pad_o[8] , \mc_addr_pad_o[9] ,
    \mc_addr_pad_o[10] , \mc_addr_pad_o[11] , \mc_addr_pad_o[12] ,
    \mc_addr_pad_o[13] , \mc_addr_pad_o[14] , \mc_addr_pad_o[15] ,
    \mc_addr_pad_o[16] , \mc_addr_pad_o[17] , \mc_addr_pad_o[18] ,
    \mc_addr_pad_o[19] , \mc_addr_pad_o[20] , \mc_addr_pad_o[21] ,
    \mc_addr_pad_o[22] , \mc_addr_pad_o[23] , \mc_dp_pad_o[0] ,
    \mc_dp_pad_o[1] , \mc_dp_pad_o[2] , \mc_dp_pad_o[3] ,
    \mc_dqm_pad_o[0] , \mc_dqm_pad_o[1] , \mc_dqm_pad_o[2] ,
    \mc_dqm_pad_o[3] , \mc_cs_pad_o_[0] , \mc_cs_pad_o_[1] ,
    \mc_cs_pad_o_[2] , \mc_cs_pad_o_[3] , \mc_cs_pad_o_[4] ,
    \mc_cs_pad_o_[5] , \mc_cs_pad_o_[6] , \mc_cs_pad_o_[7]   );
  input  clock;
  input  clk_i, rst_i, wb_we_i, wb_cyc_i, wb_stb_i, susp_req_i,
    resume_req_i, mc_clk_i, mc_br_pad_i, mc_ack_pad_i, mc_sts_pad_i,
    \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] ,
    \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] ,
    \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] ,
    \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] ,
    \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] ,
    \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] ,
    \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] ,
    \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] ,
    \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] ,
    \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] ,
    \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] ,
    \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] ,
    \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] ,
    \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] ,
    \wb_addr_i[24] , \wb_addr_i[25] , \wb_addr_i[26] , \wb_addr_i[27] ,
    \wb_addr_i[28] , \wb_addr_i[29] , \wb_addr_i[30] , \wb_addr_i[31] ,
    \mc_data_pad_i[0] , \mc_data_pad_i[1] , \mc_data_pad_i[2] ,
    \mc_data_pad_i[3] , \mc_data_pad_i[4] , \mc_data_pad_i[5] ,
    \mc_data_pad_i[6] , \mc_data_pad_i[7] , \mc_data_pad_i[8] ,
    \mc_data_pad_i[9] , \mc_data_pad_i[10] , \mc_data_pad_i[11] ,
    \mc_data_pad_i[12] , \mc_data_pad_i[13] , \mc_data_pad_i[14] ,
    \mc_data_pad_i[15] , \mc_data_pad_i[16] , \mc_data_pad_i[17] ,
    \mc_data_pad_i[18] , \mc_data_pad_i[19] , \mc_data_pad_i[20] ,
    \mc_data_pad_i[21] , \mc_data_pad_i[22] , \mc_data_pad_i[23] ,
    \mc_data_pad_i[24] , \mc_data_pad_i[25] , \mc_data_pad_i[26] ,
    \mc_data_pad_i[27] , \mc_data_pad_i[28] , \mc_data_pad_i[29] ,
    \mc_data_pad_i[30] , \mc_data_pad_i[31] , \wb_sel_i[0] , \wb_sel_i[1] ,
    \wb_sel_i[2] , \wb_sel_i[3] , \mc_dp_pad_i[0] , \mc_dp_pad_i[1] ,
    \mc_dp_pad_i[2] , \mc_dp_pad_i[3] ;
  output \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] ,
    \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] ,
    \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] ,
    \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] ,
    \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] ,
    \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] ,
    \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] ,
    \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] ,
    \poc_o[0] , \poc_o[1] , \poc_o[2] , \poc_o[3] , \poc_o[4] , \poc_o[5] ,
    \poc_o[6] , \poc_o[7] , \poc_o[8] , \poc_o[9] , \poc_o[10] ,
    \poc_o[11] , \poc_o[12] , \poc_o[13] , \poc_o[14] , \poc_o[15] ,
    \poc_o[16] , \poc_o[17] , \poc_o[18] , \poc_o[19] , \poc_o[20] ,
    \poc_o[21] , \poc_o[22] , \poc_o[23] , \poc_o[24] , \poc_o[25] ,
    \poc_o[26] , \poc_o[27] , \poc_o[28] , \poc_o[29] , \poc_o[30] ,
    \poc_o[31] , \mc_data_pad_o[0] , \mc_data_pad_o[1] ,
    \mc_data_pad_o[2] , \mc_data_pad_o[3] , \mc_data_pad_o[4] ,
    \mc_data_pad_o[5] , \mc_data_pad_o[6] , \mc_data_pad_o[7] ,
    \mc_data_pad_o[8] , \mc_data_pad_o[9] , \mc_data_pad_o[10] ,
    \mc_data_pad_o[11] , \mc_data_pad_o[12] , \mc_data_pad_o[13] ,
    \mc_data_pad_o[14] , \mc_data_pad_o[15] , \mc_data_pad_o[16] ,
    \mc_data_pad_o[17] , \mc_data_pad_o[18] , \mc_data_pad_o[19] ,
    \mc_data_pad_o[20] , \mc_data_pad_o[21] , \mc_data_pad_o[22] ,
    \mc_data_pad_o[23] , \mc_data_pad_o[24] , \mc_data_pad_o[25] ,
    \mc_data_pad_o[26] , \mc_data_pad_o[27] , \mc_data_pad_o[28] ,
    \mc_data_pad_o[29] , \mc_data_pad_o[30] , \mc_data_pad_o[31] ,
    wb_ack_o, wb_err_o, suspended_o, mc_bg_pad_o, mc_doe_pad_doe_o,
    mc_oe_pad_o_, mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_,
    mc_cke_pad_o_, mc_rp_pad_o_, mc_vpen_pad_o, mc_adsc_pad_o_,
    mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o, \mc_addr_pad_o[0] ,
    \mc_addr_pad_o[1] , \mc_addr_pad_o[2] , \mc_addr_pad_o[3] ,
    \mc_addr_pad_o[4] , \mc_addr_pad_o[5] , \mc_addr_pad_o[6] ,
    \mc_addr_pad_o[7] , \mc_addr_pad_o[8] , \mc_addr_pad_o[9] ,
    \mc_addr_pad_o[10] , \mc_addr_pad_o[11] , \mc_addr_pad_o[12] ,
    \mc_addr_pad_o[13] , \mc_addr_pad_o[14] , \mc_addr_pad_o[15] ,
    \mc_addr_pad_o[16] , \mc_addr_pad_o[17] , \mc_addr_pad_o[18] ,
    \mc_addr_pad_o[19] , \mc_addr_pad_o[20] , \mc_addr_pad_o[21] ,
    \mc_addr_pad_o[22] , \mc_addr_pad_o[23] , \mc_dp_pad_o[0] ,
    \mc_dp_pad_o[1] , \mc_dp_pad_o[2] , \mc_dp_pad_o[3] ,
    \mc_dqm_pad_o[0] , \mc_dqm_pad_o[1] , \mc_dqm_pad_o[2] ,
    \mc_dqm_pad_o[3] , \mc_cs_pad_o_[0] , \mc_cs_pad_o_[1] ,
    \mc_cs_pad_o_[2] , \mc_cs_pad_o_[3] , \mc_cs_pad_o_[4] ,
    \mc_cs_pad_o_[5] , \mc_cs_pad_o_[6] , \mc_cs_pad_o_[7] ;
  reg \\u7_mc_addr_reg[10] , \\u7_mc_addr_reg[12] , \\u7_mc_addr_reg[11] ,
    \\u7_mc_addr_reg[9] , \\u7_mc_addr_reg[8] , \\u7_mc_addr_reg[7] ,
    \\u7_mc_addr_reg[6] , \\u7_mc_addr_reg[5] , \\u7_mc_addr_reg[4] ,
    \\u7_mc_addr_reg[3] , \\u7_mc_addr_reg[2] , \\u7_mc_addr_reg[1] ,
    \\u7_mc_addr_reg[0] , u7_mc_we__reg, \\u7_mc_cs__reg[1] ,
    \\u7_mc_cs__reg[0] , \\u7_mc_cs__reg[7] , \\u7_mc_cs__reg[6] ,
    \\u7_mc_cs__reg[5] , \\u7_mc_cs__reg[4] , \\u7_mc_cs__reg[3] ,
    \\u7_mc_cs__reg[2] , \\u5_cmd_del_reg[0] , \\u5_cmd_r_reg[0] ,
    u5_cmd_asserted_reg, u7_mc_cas__reg, \\u7_mc_dqm_reg[2] ,
    \\u7_mc_dqm_reg[1] , \\u7_mc_dqm_reg[0] , \\u7_mc_dqm_reg[3] ,
    \\u5_cmd_del_reg[3] , u6_wb_ack_o_reg, \\u5_state_reg[16] ,
    \\u5_timer_reg[0] , \\u5_timer_reg[1] , \\u5_state_reg[2] ,
    \\u5_state_reg[59] , \\u5_cmd_r_reg[3] , \\u5_state_reg[17] ,
    \\u5_state_reg[1] , \\u5_state_reg[35] , \\u5_burst_cnt_reg[2] ,
    \\u5_burst_cnt_reg[8] , \\u5_burst_cnt_reg[9] , \\u5_burst_cnt_reg[0] ,
    \\u5_state_reg[21] , \\u5_state_reg[29] , \\u5_state_reg[57] ,
    \\u5_state_reg[0] , \\u5_state_reg[10] , \\u5_state_reg[15] ,
    \\u5_state_reg[40] , \\u5_burst_cnt_reg[10] , \\u5_state_reg[18] ,
    \\u5_state_reg[20] , \\u5_state_reg[22] , \\u5_state_reg[23] ,
    \\u5_state_reg[24] , \\u5_state_reg[62] , \\u5_state_reg[26] ,
    \\u5_state_reg[27] , \\u5_state_reg[28] , \\u5_state_reg[25] ,
    \\u5_state_reg[30] , \\u5_state_reg[32] , \\u5_state_reg[33] ,
    \\u5_state_reg[38] , \\u5_state_reg[43] , \\u5_state_reg[36] ,
    \\u5_state_reg[46] , \\u5_state_reg[4] , \\u5_state_reg[45] ,
    \\u5_state_reg[52] , \\u5_state_reg[60] , \\u5_state_reg[9] ,
    \\u5_state_reg[13] , \\u5_state_reg[12] , \\u5_state_reg[48] ,
    u7_mc_data_oe_reg, \\u5_timer_reg[2] , u6_wb_err_reg,
    \\u5_state_reg[37] , \\u5_state_reg[39] , \\u5_state_reg[42] ,
    \\u5_state_reg[41] , \\u5_state_reg[44] , \\u5_state_reg[47] ,
    \\u5_state_reg[51] , \\u5_state_reg[56] , \\u5_state_reg[5] ,
    \\u5_state_reg[61] , \\u5_state_reg[58] , \\u5_state_reg[63] ,
    \\u5_state_reg[64] , \\u5_state_reg[11] , \\u5_state_reg[6] ,
    \\u5_state_reg[7] , \\u5_state_reg[8] , \\u5_state_reg[65] ,
    \\u5_burst_cnt_reg[3] , \\u5_state_reg[14] , \\u5_burst_cnt_reg[1] ,
    \\u5_state_reg[34] , \\u5_state_reg[50] , \\u5_state_reg[55] ,
    \\u5_cmd_del_reg[1] , \\u5_state_reg[19] , \\u5_state_reg[31] ,
    \\u5_state_reg[3] , \\u5_state_reg[49] , \\u5_state_reg[54] ,
    \\u5_state_reg[53] , u7_mc_oe__reg, \\u5_burst_cnt_reg[4] ,
    \\u5_burst_cnt_reg[7] , \\u5_burst_cnt_reg[6] , \\u5_burst_cnt_reg[5] ,
    \\u5_cmd_r_reg[1] , \\u5_timer_reg[3] , u5_data_oe_reg,
    u5_wb_stb_first_reg, \\u5_timer2_reg[2] , u5_mem_ack_r_reg,
    mem_ack_r_reg, u5_oe__reg, \\u5_timer2_reg[1] , \\u5_timer2_reg[3] ,
    u5_cke__reg, u5_data_oe_r2_reg, u5_cke_r_reg, \\u5_timer2_reg[5] ,
    u5_data_oe_r_reg, \\u5_timer2_reg[4] , \\u5_timer2_reg[0] ,
    \\u5_timer2_reg[8] , \\u5_timer2_reg[7] , \\u5_timer2_reg[6] ,
    u5_ap_en_reg, \\u5_timer_reg[5] , \\u5_timer_reg[4] ,
    \\u0_tms_reg[21] , \\u0_tms_reg[5] , \\u0_tms_reg[9] ,
    \\u0_tms_reg[27] , \\u0_tms_reg[1] , \\u0_tms_reg[16] ,
    \\u0_sp_tms_reg[9] , \\u0_sp_tms_reg[26] , \\u0_sp_tms_reg[5] ,
    \\u0_sp_tms_reg[20] , \\u0_sp_tms_reg[23] , \\u0_sp_tms_reg[11] ,
    \\u0_sp_tms_reg[0] , \\u0_sp_tms_reg[10] , \\u0_sp_tms_reg[12] ,
    \\u0_sp_tms_reg[13] , \\u0_sp_tms_reg[14] , \\u0_sp_tms_reg[15] ,
    \\u0_sp_tms_reg[17] , \\u0_sp_tms_reg[18] , \\u0_sp_tms_reg[19] ,
    \\u0_sp_tms_reg[1] , \\u0_sp_tms_reg[21] , \\u0_sp_tms_reg[22] ,
    \\u0_sp_tms_reg[24] , \\u0_sp_tms_reg[27] , \\u0_sp_tms_reg[2] ,
    \\u0_sp_tms_reg[25] , \\u0_sp_tms_reg[3] , \\u0_sp_tms_reg[4] ,
    \\u0_sp_tms_reg[6] , \\u0_sp_tms_reg[7] , \\u0_sp_tms_reg[8] ,
    \\u0_tms_reg[11] , \\u0_tms_reg[0] , \\u0_tms_reg[10] ,
    \\u0_tms_reg[12] , \\u0_tms_reg[13] , \\u0_tms_reg[15] ,
    \\u0_tms_reg[14] , \\u0_tms_reg[17] , \\u0_tms_reg[18] ,
    \\u0_tms_reg[19] , \\u0_tms_reg[20] , \\u0_tms_reg[22] ,
    \\u0_tms_reg[23] , \\u0_tms_reg[24] , \\u0_tms_reg[26] ,
    \\u0_tms_reg[25] , \\u0_tms_reg[2] , \\u0_tms_reg[3] ,
    \\u0_tms_reg[4] , \\u0_tms_reg[7] , \\u0_tms_reg[8] , \\u0_tms_reg[6] ,
    \\u5_timer_reg[7] , \\u5_timer_reg[6] , \\u0_sp_tms_reg[16] ,
    \\u0_csc_reg[10] , \\u0_csc_reg[5] , \\u0_csc_reg[4] ,
    u2_u0_bank0_open_reg, u2_u0_bank1_open_reg, u2_u0_bank3_open_reg,
    u2_u1_bank0_open_reg, u2_u1_bank1_open_reg, u2_u1_bank2_open_reg,
    \\u0_csc_reg[6] , \\u0_csc_reg[7] , \\u0_csc_reg[9] ,
    \\u0_sp_csc_reg[10] , \\u0_sp_csc_reg[4] , \\u0_sp_csc_reg[7] ,
    \\u0_sp_csc_reg[9] , \\u0_sp_csc_reg[6] , \\u0_sp_csc_reg[3] ,
    \\u0_sp_csc_reg[2] , \\u0_csc_reg[11] , u2_u1_bank3_open_reg,
    \\u0_sp_csc_reg[5] , u2_u0_bank2_open_reg, \\u0_sp_csc_reg[1] ,
    \\u0_csc_reg[1] , \\u0_csc_reg[3] , \\u0_csc_reg[2] , u5_cmd_a10_r_reg,
    u7_mc_ras__reg, u7_mc_adsc__reg, u5_wr_cycle_reg, u7_mc_c_oe_reg,
    u5_cs_le_reg, \\u5_cmd_del_reg[2] , u5_mc_c_oe_reg,
    \\u1_bank_adr_reg[0] , \\u1_row_adr_reg[10] , \\u1_row_adr_reg[11] ,
    \\u5_cmd_r_reg[2] , \\u1_bank_adr_reg[1] , \\u1_row_adr_reg[9] ,
    \\u1_row_adr_reg[12] , \\u1_row_adr_reg[3] , \\u1_row_adr_reg[7] ,
    \\u1_row_adr_reg[0] , \\u1_acs_addr_reg[23] , \\u1_row_adr_reg[1] ,
    \\u1_row_adr_reg[2] , \\u1_row_adr_reg[4] , \\u1_row_adr_reg[5] ,
    \\u1_row_adr_reg[6] , \\u1_row_adr_reg[8] , u5_cnt_reg,
    \\u3_byte1_reg[5] , u5_wb_cycle_reg, \\u1_acs_addr_reg[19] ,
    \\u1_acs_addr_reg[20] , \\u3_byte1_reg[0] , \\u3_byte1_reg[1] ,
    \\u3_byte1_reg[2] , \\u3_byte1_reg[3] , \\u3_byte1_reg[4] ,
    \\u3_byte1_reg[7] , \\u3_byte1_reg[6] , \\u1_col_adr_reg[8] ,
    \\u1_acs_addr_reg[22] , \\u1_acs_addr_reg[9] , \\u1_acs_addr_reg[10] ,
    \\u1_acs_addr_reg[2] , \\u1_acs_addr_reg[21] , \\u1_acs_addr_reg[18] ,
    \\u1_acs_addr_reg[4] , \\u1_acs_addr_reg[7] , \\u1_acs_addr_reg[13] ,
    \\u1_acs_addr_reg[16] , \\u1_acs_addr_reg[14] , \\u1_acs_addr_reg[11] ,
    \\u1_acs_addr_reg[17] , \\u1_acs_addr_reg[12] , \\u1_acs_addr_reg[8] ,
    \\u1_acs_addr_reg[0] , \\u1_acs_addr_reg[1] , \\u1_acs_addr_reg[3] ,
    \\u1_acs_addr_reg[5] , \\u1_acs_addr_reg[6] , \\u1_acs_addr_reg[15] ,
    \\u1_col_adr_reg[9] , \\u5_ack_cnt_reg[3] , \\u5_ack_cnt_reg[1] ,
    u4_rfr_req_reg, \\u5_ack_cnt_reg[0] , \\u5_ack_cnt_reg[2] ,
    \\u3_byte0_reg[1] , \\u3_byte0_reg[0] , \\u3_byte0_reg[2] ,
    \\u3_byte0_reg[4] , \\u3_byte0_reg[3] , \\u3_byte0_reg[5] ,
    \\u3_byte0_reg[6] , \\u3_byte0_reg[7] , \\u3_byte2_reg[7] ,
    u5_lmr_ack_reg, \\u5_ir_cnt_reg[1] , \\u5_ir_cnt_reg[2] ,
    \\u7_mc_addr_reg[14] , \\u3_byte2_reg[0] , \\u3_byte2_reg[1] ,
    \\u3_byte2_reg[2] , \\u3_byte2_reg[4] , \\u3_byte2_reg[5] ,
    \\u3_byte2_reg[6] , \\u3_byte2_reg[3] , \\u7_mc_addr_reg[13] ,
    \\u5_ir_cnt_reg[3] , \\u5_ir_cnt_reg[0] , u5_mc_adv_r1_reg,
    u5_tmr2_done_reg, \\u3_u0_r0_reg[16] , \\u3_u0_r0_reg[22] ,
    \\u3_u0_r1_reg[26] , \\u3_u0_r2_reg[25] , \\u3_u0_r2_reg[3] ,
    \\u3_u0_r0_reg[1] , \\u3_u0_r0_reg[18] , \\u3_u0_r0_reg[19] ,
    \\u3_u0_r0_reg[10] , \\u3_u0_r2_reg[32] , \\u3_u0_r2_reg[27] ,
    \\u3_u0_r2_reg[29] , \\u3_u0_r0_reg[14] , \\u3_u0_r2_reg[18] ,
    \\u3_u0_r2_reg[21] , \\u3_u0_wr_adr_reg[1] , \\u3_u0_wr_adr_reg[3] ,
    u5_rfr_ack_r_reg, \\u3_u0_r2_reg[14] , \\u3_u0_r2_reg[10] ,
    \\u3_u0_r2_reg[12] , \\u3_u0_r1_reg[9] , \\u3_u0_r1_reg[7] ,
    \\u3_u0_r1_reg[3] , \\u3_u0_r1_reg[32] , \\u3_u0_wr_adr_reg[0] ,
    \\u3_u0_wr_adr_reg[2] , \\u3_u0_r0_reg[0] , \\u3_u0_r0_reg[11] ,
    \\u3_u0_r0_reg[12] , \\u3_u0_r0_reg[13] , \\u3_u0_r0_reg[15] ,
    \\u3_u0_r0_reg[17] , \\u3_u0_r0_reg[20] , \\u3_u0_r0_reg[21] ,
    \\u3_u0_r0_reg[23] , \\u3_u0_r0_reg[24] , \\u3_u0_r0_reg[26] ,
    \\u3_u0_r0_reg[27] , \\u3_u0_r0_reg[28] , \\u3_u0_r0_reg[2] ,
    \\u3_u0_r0_reg[30] , \\u3_u0_r0_reg[31] , \\u3_u0_r0_reg[33] ,
    \\u3_u0_r0_reg[34] , \\u3_u0_r0_reg[35] , \\u3_u0_r0_reg[4] ,
    \\u3_u0_r0_reg[9] , \\u3_u0_r1_reg[0] , \\u3_u0_r1_reg[11] ,
    \\u3_u0_r1_reg[10] , \\u3_u0_r1_reg[12] , \\u3_u0_r1_reg[13] ,
    \\u3_u0_r1_reg[15] , \\u3_u0_r1_reg[16] , \\u3_u0_r1_reg[17] ,
    \\u3_u0_r1_reg[19] , \\u3_u0_r1_reg[1] , \\u3_u0_r1_reg[20] ,
    \\u3_u0_r1_reg[23] , \\u3_u0_r1_reg[22] , \\u3_u0_r1_reg[24] ,
    \\u3_u0_r1_reg[25] , \\u3_u0_r1_reg[27] , \\u3_u0_r1_reg[28] ,
    \\u3_u0_r1_reg[2] , \\u3_u0_r1_reg[30] , \\u3_u0_r1_reg[31] ,
    \\u3_u0_r1_reg[33] , \\u3_u0_r1_reg[34] , \\u3_u0_r1_reg[35] ,
    \\u3_u0_r1_reg[4] , \\u3_u0_r1_reg[5] , \\u3_u0_r1_reg[6] ,
    \\u3_u0_r1_reg[8] , \\u3_u0_r2_reg[0] , \\u3_u0_r2_reg[11] ,
    \\u3_u0_r2_reg[13] , \\u3_u0_r2_reg[15] , \\u3_u0_r2_reg[16] ,
    \\u3_u0_r2_reg[17] , \\u3_u0_r2_reg[19] , \\u3_u0_r2_reg[1] ,
    \\u3_u0_r2_reg[20] , \\u3_u0_r2_reg[22] , \\u3_u0_r2_reg[23] ,
    \\u3_u0_r2_reg[24] , \\u3_u0_r2_reg[26] , \\u3_u0_r2_reg[28] ,
    \\u3_u0_r2_reg[2] , \\u3_u0_r2_reg[30] , \\u3_u0_r2_reg[31] ,
    \\u3_u0_r2_reg[33] , \\u3_u0_r2_reg[34] , \\u3_u0_r2_reg[35] ,
    \\u3_u0_r2_reg[4] , \\u3_u0_r2_reg[5] , \\u3_u0_r2_reg[6] ,
    \\u3_u0_r2_reg[8] , \\u3_u0_r3_reg[0] , \\u3_u0_r3_reg[11] ,
    \\u3_u0_r3_reg[12] , \\u3_u0_r3_reg[13] , \\u3_u0_r3_reg[15] ,
    \\u3_u0_r3_reg[16] , \\u3_u0_r3_reg[17] , \\u3_u0_r3_reg[19] ,
    \\u3_u0_r3_reg[1] , \\u3_u0_r3_reg[20] , \\u3_u0_r3_reg[22] ,
    \\u3_u0_r3_reg[23] , \\u3_u0_r3_reg[24] , \\u3_u0_r3_reg[26] ,
    \\u3_u0_r3_reg[28] , \\u3_u0_r3_reg[2] , \\u3_u0_r3_reg[31] ,
    \\u3_u0_r3_reg[33] , \\u3_u0_r3_reg[34] , \\u3_u0_r3_reg[35] ,
    \\u3_u0_r3_reg[4] , \\u3_u0_r3_reg[5] , \\u3_u0_r3_reg[6] ,
    \\u3_u0_r3_reg[9] , \\u3_u0_r3_reg[8] , \\u3_u0_r1_reg[29] ,
    \\u3_u0_r1_reg[21] , \\u3_u0_r0_reg[7] , \\u3_u0_r1_reg[18] ,
    \\u3_u0_r3_reg[7] , \\u3_u0_r3_reg[3] , \\u3_u0_r3_reg[30] ,
    \\u3_u0_r3_reg[32] , \\u3_u0_r1_reg[14] , \\u3_u0_r3_reg[25] ,
    \\u3_u0_r3_reg[29] , \\u3_u0_r0_reg[8] , \\u3_u0_r3_reg[27] ,
    \\u3_u0_r0_reg[5] , \\u3_u0_r3_reg[14] , \\u3_u0_r3_reg[21] ,
    \\u3_u0_r0_reg[6] , \\u3_u0_r2_reg[7] , u4_rfr_clr_reg,
    \\u3_u0_r0_reg[3] , \\u3_u0_r3_reg[18] , \\u3_u0_r0_reg[32] ,
    \\u3_u0_r0_reg[29] , \\u3_u0_r0_reg[25] , \\u3_u0_r2_reg[9] ,
    \\u3_u0_r3_reg[10] , \\u7_mc_addr_reg[23] , \\u7_mc_addr_reg[17] ,
    u7_mc_bg_reg, u5_susp_sel_r_reg, \\u7_mc_addr_reg[22] ,
    \\u7_mc_addr_reg[21] , \\u7_mc_addr_reg[19] , \\u7_mc_addr_reg[20] ,
    \\u7_mc_addr_reg[18] , \\u7_mc_addr_reg[16] , \\u7_mc_addr_reg[15] ,
    u5_pack_le0_reg, u7_mc_adv__reg, u5_pack_le2_reg, u5_wb_wait_r_reg,
    u5_dv_r_reg, \\u2_u0_b0_last_row_reg[6] , \\u2_u0_b3_last_row_reg[8] ,
    \\u2_u1_b2_last_row_reg[0] , \\u2_u1_b2_last_row_reg[8] ,
    \\u2_u1_b3_last_row_reg[10] , \\u2_u1_b3_last_row_reg[1] ,
    \\u2_u0_b0_last_row_reg[4] , \\u2_u0_b0_last_row_reg[12] ,
    \\u2_u1_b3_last_row_reg[0] , \\u2_u1_b2_last_row_reg[7] ,
    \\u2_u1_b2_last_row_reg[9] , \\u2_u1_b2_last_row_reg[3] ,
    \\u2_u1_b2_last_row_reg[1] , \\u2_u1_b2_last_row_reg[12] ,
    \\u2_u1_b2_last_row_reg[11] , \\u2_u1_b1_last_row_reg[8] ,
    \\u2_u1_b1_last_row_reg[12] , \\u2_u0_b3_last_row_reg[9] ,
    \\u2_u1_b1_last_row_reg[4] , \\u2_u1_b1_last_row_reg[7] ,
    \\u2_u1_b1_last_row_reg[6] , \\u2_u1_b1_last_row_reg[5] ,
    \\u2_u1_b1_last_row_reg[2] , \\u2_u1_b0_last_row_reg[0] ,
    \\u2_u1_b1_last_row_reg[10] , \\u2_u1_b0_last_row_reg[7] ,
    \\u2_u1_b0_last_row_reg[9] , \\u2_u1_b0_last_row_reg[5] ,
    \\u2_u1_b0_last_row_reg[2] , \\u2_u0_b0_last_row_reg[0] ,
    \\u2_u0_b0_last_row_reg[10] , \\u2_u0_b0_last_row_reg[11] ,
    \\u2_u0_b0_last_row_reg[1] , \\u2_u0_b0_last_row_reg[2] ,
    \\u2_u0_b0_last_row_reg[3] , \\u2_u0_b0_last_row_reg[5] ,
    \\u2_u0_b0_last_row_reg[9] , \\u2_u0_b1_last_row_reg[10] ,
    \\u2_u0_b1_last_row_reg[12] , \\u2_u0_b1_last_row_reg[4] ,
    \\u2_u0_b1_last_row_reg[6] , \\u2_u0_b1_last_row_reg[9] ,
    \\u2_u0_b2_last_row_reg[10] , \\u2_u0_b2_last_row_reg[12] ,
    \\u2_u0_b2_last_row_reg[2] , \\u2_u0_b2_last_row_reg[4] ,
    \\u2_u0_b2_last_row_reg[5] , \\u2_u0_b2_last_row_reg[8] ,
    \\u2_u0_b2_last_row_reg[9] , \\u2_u0_b2_last_row_reg[3] ,
    \\u2_u0_b3_last_row_reg[11] , \\u2_u0_b3_last_row_reg[5] ,
    \\u2_u1_b0_last_row_reg[11] , \\u2_u1_b0_last_row_reg[12] ,
    \\u2_u1_b0_last_row_reg[3] , \\u2_u1_b0_last_row_reg[4] ,
    \\u2_u1_b0_last_row_reg[6] , \\u2_u1_b0_last_row_reg[8] ,
    \\u2_u1_b1_last_row_reg[0] , \\u2_u1_b1_last_row_reg[11] ,
    \\u2_u1_b1_last_row_reg[1] , \\u2_u1_b1_last_row_reg[3] ,
    \\u2_u1_b1_last_row_reg[9] , \\u2_u1_b2_last_row_reg[10] ,
    \\u2_u1_b2_last_row_reg[2] , \\u2_u1_b2_last_row_reg[4] ,
    \\u2_u1_b2_last_row_reg[5] , \\u2_u1_b2_last_row_reg[6] ,
    \\u2_u1_b3_last_row_reg[11] , \\u2_u1_b3_last_row_reg[12] ,
    \\u2_u1_b3_last_row_reg[3] , \\u2_u1_b3_last_row_reg[5] ,
    \\u2_u1_b3_last_row_reg[7] , \\u2_u1_b3_last_row_reg[6] ,
    \\u2_u1_b3_last_row_reg[8] , \\u2_u0_b3_last_row_reg[0] ,
    \\u2_u1_b0_last_row_reg[10] , \\u2_u1_b0_last_row_reg[1] ,
    \\u2_u0_b0_last_row_reg[7] , \\u2_u0_b3_last_row_reg[3] ,
    \\u2_u0_b1_last_row_reg[5] , \\u2_u0_b3_last_row_reg[7] ,
    \\u2_u1_b3_last_row_reg[4] , \\u2_u0_b3_last_row_reg[4] ,
    \\u2_u0_b3_last_row_reg[6] , \\u2_u0_b3_last_row_reg[1] ,
    u0_wp_err_reg, \\u2_u0_b3_last_row_reg[2] ,
    \\u2_u0_b3_last_row_reg[12] , \\u2_u0_b3_last_row_reg[10] ,
    \\u2_u0_b2_last_row_reg[7] , \\u2_u0_b2_last_row_reg[1] ,
    \\u2_u0_b2_last_row_reg[0] , \\u2_u0_b1_last_row_reg[7] ,
    \\u2_u0_b2_last_row_reg[11] , \\u2_u0_b2_last_row_reg[6] ,
    \\u2_u1_b3_last_row_reg[9] , \\u2_u0_b1_last_row_reg[8] ,
    \\u2_u0_b0_last_row_reg[8] , \\u2_u1_b3_last_row_reg[2] ,
    \\u2_u0_b1_last_row_reg[11] , \\u2_u0_b1_last_row_reg[3] ,
    u5_wb_wait_r2_reg, \\u2_u0_b1_last_row_reg[2] ,
    \\u2_u0_b1_last_row_reg[1] , \\u2_u0_b1_last_row_reg[0] ,
    \\u0_cs_reg[0] , \\u3_u0_rd_adr_reg[3] , u2_bank_open_reg,
    \\u3_u0_rd_adr_reg[0] , \\u3_u0_rd_adr_reg[2] , \\u3_u0_rd_adr_reg[1] ,
    u2_row_same_reg, \\u4_rfr_cnt_reg[3] , \\u4_rfr_cnt_reg[5] ,
    \\u4_rfr_cnt_reg[6] , \\u4_rfr_cnt_reg[4] , u0_u0_init_req_reg,
    \\u4_rfr_cnt_reg[7] , \\u4_rfr_cnt_reg[2] , \\u4_rfr_cnt_reg[1] ,
    \\u0_cs_reg[1] , \\u0_u0_csc_reg[0] , u0_u1_lmr_req_reg,
    \\u4_rfr_cnt_reg[0] , \\u0_u0_csc_reg[4] , \\u0_u0_csc_reg[7] ,
    \\u0_u0_csc_reg[16] , \\u0_u0_csc_reg[18] , \\u0_u0_csc_reg[13] ,
    \\u0_u0_csc_reg[14] , \\u0_u0_csc_reg[11] , \\u0_u0_csc_reg[15] ,
    \\u0_u0_csc_reg[2] , u0_u1_init_req_reg, \\u0_u0_csc_reg[1] ,
    \\u0_u0_csc_reg[5] , \\u0_u0_csc_reg[17] , \\u0_u0_csc_reg[22] ,
    \\u0_u0_csc_reg[12] , \\u0_u0_csc_reg[8] , \\u0_u0_csc_reg[9] ,
    \\u0_u0_csc_reg[6] , u0_u0_lmr_req_reg, \\u0_u1_csc_reg[16] ,
    \\u0_u0_csc_reg[21] , \\u0_u1_csc_reg[17] , \\u0_u1_csc_reg[19] ,
    \\u0_u0_csc_reg[19] , \\u0_u0_csc_reg[20] , \\u0_u1_csc_reg[13] ,
    \\u0_u1_csc_reg[15] , \\u0_u0_csc_reg[10] , \\u0_u1_csc_reg[10] ,
    \\u0_u1_csc_reg[12] , \\u0_u0_csc_reg[27] , \\u0_u1_csc_reg[5] ,
    \\u0_u1_csc_reg[7] , \\u0_u1_csc_reg[9] , \\u0_u0_csc_reg[28] ,
    \\u0_u1_csc_reg[21] , \\u0_u0_csc_reg[3] , \\u0_u1_csc_reg[4] ,
    \\u0_u0_csc_reg[23] , \\u0_u0_csc_reg[25] , \\u0_u1_csc_reg[14] ,
    \\u0_u1_csc_reg[20] , \\u0_u1_csc_reg[22] , \\u0_u1_csc_reg[26] ,
    \\u0_u1_csc_reg[27] , \\u0_u0_csc_reg[30] , \\u0_u0_csc_reg[31] ,
    \\u0_u0_csc_reg[29] , \\u0_u1_csc_reg[30] , \\u0_u1_csc_reg[24] ,
    \\u0_u0_csc_reg[26] , \\u0_u1_csc_reg[31] , \\u0_u0_csc_reg[24] ,
    \\u1_u0_out_r_reg[11] , \\u0_u1_csc_reg[18] , \\u0_u1_csc_reg[1] ,
    \\u0_u1_csc_reg[2] , \\u6_wb_data_o_reg[10] , \\u6_wb_data_o_reg[2] ,
    \\u0_u1_csc_reg[8] , \\u6_wb_data_o_reg[7] , \\u6_wb_data_o_reg[3] ,
    \\u6_wb_data_o_reg[0] , \\u0_u1_csc_reg[25] , \\u6_wb_data_o_reg[11] ,
    \\u6_wb_data_o_reg[14] , \\u6_wb_data_o_reg[1] ,
    \\u6_wb_data_o_reg[5] , \\u6_wb_data_o_reg[9] , \\u6_wb_data_o_reg[6] ,
    \\u6_wb_data_o_reg[4] , \\u6_wb_data_o_reg[12] ,
    \\u6_wb_data_o_reg[15] , \\u6_wb_data_o_reg[8] , \\u0_u1_csc_reg[0] ,
    \\u0_u1_csc_reg[3] , \\u6_wb_data_o_reg[13] , u5_wb_write_go_r_reg,
    \\u0_u1_tms_reg[30] , \\u6_wb_data_o_reg[31] , \\u0_u1_tms_reg[13] ,
    \\u0_u1_tms_reg[27] , \\u0_u1_tms_reg[15] , \\u6_wb_data_o_reg[24] ,
    \\u0_u1_tms_reg[8] , \\u0_u1_tms_reg[7] , \\u6_wb_data_o_reg[26] ,
    \\u0_u1_csc_reg[29] , \\u0_u1_tms_reg[28] , \\u0_u1_csc_reg[11] ,
    \\u0_u1_tms_reg[0] , \\u0_u1_tms_reg[29] , \\u0_u1_tms_reg[16] ,
    \\u0_u1_tms_reg[3] , \\u0_u1_tms_reg[10] , \\u0_u1_tms_reg[23] ,
    \\u0_u1_tms_reg[17] , \\u0_u1_tms_reg[24] , \\u0_u1_tms_reg[12] ,
    \\u0_u1_tms_reg[25] , \\u0_u1_tms_reg[5] , \\u6_wb_data_o_reg[17] ,
    \\u6_wb_data_o_reg[18] , \\u0_u1_tms_reg[18] , \\u0_u1_csc_reg[6] ,
    \\u6_wb_data_o_reg[20] , \\u6_wb_data_o_reg[23] ,
    \\u6_wb_data_o_reg[19] , \\u6_wb_data_o_reg[29] , \\u0_u1_csc_reg[23] ,
    \\u6_wb_data_o_reg[21] , \\u6_wb_data_o_reg[25] ,
    \\u6_wb_data_o_reg[16] , \\u6_wb_data_o_reg[27] ,
    \\u6_wb_data_o_reg[30] , \\u4_ps_cnt_reg[7] , \\u6_wb_data_o_reg[28] ,
    \\u0_u1_tms_reg[11] , \\u0_u1_tms_reg[14] , \\u0_u1_tms_reg[20] ,
    \\u0_u1_tms_reg[26] , \\u0_u1_tms_reg[2] , \\u0_u1_tms_reg[31] ,
    \\u0_u1_tms_reg[4] , \\u0_u1_tms_reg[6] , \\u4_ps_cnt_reg[4] ,
    \\u0_u1_csc_reg[28] , \\u6_wb_data_o_reg[22] , \\u0_u1_tms_reg[19] ,
    \\u0_u1_tms_reg[9] , \\u0_u1_tms_reg[1] , \\u0_u1_tms_reg[22] ,
    \\u0_u1_tms_reg[21] , \\u0_u0_tms_reg[8] , u0_u0_init_req_we_reg,
    \\u0_u0_tms_reg[14] , \\u0_u0_tms_reg[12] , \\u0_u0_tms_reg[9] ,
    \\u0_u0_tms_reg[31] , \\u0_u0_tms_reg[11] , \\u0_u0_tms_reg[4] ,
    \\u4_ps_cnt_reg[3] , \\u0_u0_tms_reg[6] , \\u0_u0_tms_reg[5] ,
    \\u0_u0_tms_reg[30] , \\u0_u0_tms_reg[23] , \\u0_u0_tms_reg[24] ,
    \\u0_u0_tms_reg[17] , \\u0_u0_tms_reg[18] , \\u0_u0_tms_reg[20] ,
    \\u0_u0_tms_reg[19] , \\u0_u0_tms_reg[13] , \\u0_u0_tms_reg[1] ,
    \\u0_u0_tms_reg[0] , \\u0_u0_tms_reg[15] , \\u0_u0_tms_reg[21] ,
    \\u0_u0_tms_reg[29] , \\u0_u0_tms_reg[3] , \\u0_u0_tms_reg[7] ,
    \\u4_ps_cnt_reg[0] , \\u0_u0_tms_reg[10] , \\u0_u0_tms_reg[16] ,
    \\u0_u0_tms_reg[25] , \\u4_ps_cnt_reg[6] , \\u0_u0_tms_reg[26] ,
    \\u4_ps_cnt_reg[1] , \\u0_u0_tms_reg[2] , \\u4_ps_cnt_reg[2] ,
    \\u0_u0_tms_reg[27] , \\u4_ps_cnt_reg[5] , \\u0_u0_tms_reg[28] ,
    \\u0_u0_tms_reg[22] , \\u0_csc_mask_r_reg[0] , u0_u1_inited_reg,
    u0_u0_inited_reg, \\u0_csc_mask_r_reg[1] , u0_sreq_cs_le_reg,
    \\u0_csc_mask_r_reg[9] , \\u0_csc_mask_r_reg[10] ,
    \\u0_csc_mask_r_reg[2] , u5_cmd_asserted2_reg, \\u0_csc_mask_r_reg[4] ,
    \\u0_csc_mask_r_reg[5] , \\u0_csc_mask_r_reg[6] ,
    \\u0_csc_mask_r_reg[7] , \\u0_csc_mask_r_reg[8] ,
    \\u0_csc_mask_r_reg[3] , u5_no_wb_cycle_reg, \\u0_csr_r2_reg[6] ,
    \\u0_csr_r2_reg[4] , \\u1_u0_out_r_reg[9] , u0_u1_init_req_we_reg,
    \\u0_csr_r2_reg[0] , \\u0_csr_r_reg[7] , \\u0_csr_r2_reg[1] ,
    \\u0_csr_r2_reg[2] , \\u1_u0_out_r_reg[12] , \\u0_csr_r_reg[6] ,
    \\u0_csr_r_reg[9] , \\u1_u0_out_r_reg[7] , u4_rfr_ce_reg,
    \\u0_csr_r2_reg[3] , \\u0_csr_r_reg[1] , \\u0_csr_r_reg[3] ,
    \\u0_csr_r_reg[8] , \\u0_csr_r_reg[2] , \\u0_csr_r_reg[4] ,
    \\u0_csr_r2_reg[7] , \\u0_csr_r_reg[5] , \\u0_csr_r_reg[10] ,
    \\u0_csr_r2_reg[5] , \\u1_u0_out_r_reg[4] , u6_wb_first_r_reg,
    \\u1_u0_out_r_reg[10] , \\u1_u0_out_r_reg[8] , u4_rfr_early_reg,
    u7_mc_rp_reg, u0_u1_lmr_req_we_reg, u6_read_go_r1_reg,
    \\u3_mc_dp_o_reg[3] , \\u3_mc_dp_o_reg[2] , \\u3_mc_dp_o_reg[0] ,
    \\u3_mc_dp_o_reg[1] , u6_write_go_r1_reg, \\u1_u0_out_r_reg[5] ,
    u0_u0_lmr_req_we_reg, u0_rf_we_reg, u6_wr_hold_reg, u7_mc_zz_o_reg,
    u5_lookup_ready2_reg, \\u1_u0_out_r_reg[6] , \\u0_poc_reg[0] ,
    \\u0_poc_reg[22] , \\u0_poc_reg[25] , \\u7_mc_dqm_r_reg[0] ,
    u5_tmr_done_reg, \\u0_poc_reg[23] , \\u0_poc_reg[24] ,
    \\u0_poc_reg[26] , \\u0_poc_reg[21] , \\u1_col_adr_reg[0] ,
    \\u0_poc_reg[17] , \\u0_poc_reg[13] , \\u7_mc_dqm_r_reg[2] ,
    \\u0_poc_reg[1] , \\u0_poc_reg[28] , \\u0_poc_reg[11] ,
    \\u0_poc_reg[16] , \\u0_poc_reg[19] , \\u0_poc_reg[10] ,
    \\u0_poc_reg[15] , \\u0_poc_reg[18] , \\u0_poc_reg[20] ,
    \\u0_poc_reg[9] , \\u0_poc_reg[31] , \\u1_col_adr_reg[7] ,
    \\u1_col_adr_reg[5] , \\u7_mc_dqm_r_reg[3] , \\u7_mc_dqm_r_reg[1] ,
    \\u0_poc_reg[14] , \\u0_poc_reg[5] , \\u0_poc_reg[29] ,
    \\u0_poc_reg[27] , \\u1_col_adr_reg[6] , \\u0_poc_reg[12] ,
    \\u0_poc_reg[3] , \\u0_poc_reg[2] , \\u0_poc_reg[7] , \\u0_poc_reg[8] ,
    \\u1_col_adr_reg[2] , \\u0_poc_reg[6] , \\u1_col_adr_reg[4] ,
    \\u1_col_adr_reg[3] , \\u1_col_adr_reg[1] , \\u0_poc_reg[30] ,
    \\u0_poc_reg[4] , u0_init_ack_r_reg, \\u3_mc_data_o_reg[7] ,
    \\u3_mc_data_o_reg[24] , \\u3_mc_data_o_reg[25] ,
    \\u3_mc_data_o_reg[9] , \\u3_mc_data_o_reg[0] ,
    \\u3_mc_data_o_reg[20] , \\u3_mc_data_o_reg[3] ,
    \\u3_mc_data_o_reg[26] , \\u3_mc_data_o_reg[16] ,
    \\u3_mc_data_o_reg[1] , u5_suspended_reg, \\u3_mc_data_o_reg[19] ,
    \\u3_mc_data_o_reg[13] , \\u3_mc_data_o_reg[18] , u5_pack_le1_reg,
    \\u3_mc_data_o_reg[29] , \\u3_mc_data_o_reg[15] ,
    \\u3_mc_data_o_reg[10] , u5_burst_act_rd_reg, \\u3_mc_data_o_reg[11] ,
    \\u3_mc_data_o_reg[21] , \\u3_mc_data_o_reg[27] ,
    \\u3_mc_data_o_reg[31] , \\u3_mc_data_o_reg[28] ,
    \\u0_spec_req_cs_reg[1] , \\u3_mc_data_o_reg[22] ,
    \\u3_mc_data_o_reg[5] , \\u3_mc_data_o_reg[17] ,
    \\u3_mc_data_o_reg[30] , \\u3_mc_data_o_reg[14] ,
    \\u3_mc_data_o_reg[6] , \\u1_u0_out_r_reg[3] , \\u3_mc_data_o_reg[8] ,
    \\u3_mc_data_o_reg[23] , \\u3_mc_data_o_reg[12] ,
    \\u3_mc_data_o_reg[4] , \\u3_mc_data_o_reg[2] , \\u1_sram_addr_reg[5] ,
    \\u1_sram_addr_reg[6] , \\u1_sram_addr_reg[18] ,
    \\u1_sram_addr_reg[20] , u5_ir_cnt_done_reg, \\u1_sram_addr_reg[21] ,
    \\u1_sram_addr_reg[23] , \\u1_sram_addr_reg[11] ,
    \\u1_sram_addr_reg[2] , \\u1_sram_addr_reg[10] ,
    \\u1_sram_addr_reg[0] , \\u1_sram_addr_reg[16] ,
    \\u1_sram_addr_reg[8] , \\u1_sram_addr_reg[3] ,
    \\u1_sram_addr_reg[13] , \\u1_sram_addr_reg[7] ,
    \\u1_sram_addr_reg[15] , \\u1_sram_addr_reg[14] ,
    \\u1_sram_addr_reg[1] , \\u1_sram_addr_reg[12] ,
    \\u1_sram_addr_reg[4] , \\u1_sram_addr_reg[19] ,
    \\u1_sram_addr_reg[22] , \\u1_sram_addr_reg[17] ,
    \\u1_sram_addr_reg[9] , u4_rfr_en_reg, u5_lookup_ready1_reg,
    \\u0_spec_req_cs_reg[0] , \\u1_u0_out_r_reg[2] , u5_mc_adv_r_reg,
    u6_rmw_r_reg, u6_write_go_r_reg, \\u0_u0_addr_r_reg[2] ,
    \\u0_u1_addr_r_reg[2] , u5_mc_le_reg, u0_rst_r3_reg,
    \\u0_wb_addr_r_reg[2] , u6_rmw_en_reg, \\u1_u0_out_r_reg[1] ,
    u5_cke_o_del_reg, \\u0_spec_req_cs_reg[5] , \\u0_cs_reg[6] ,
    u0_u1_rst_r2_reg, \\u0_spec_req_cs_reg[4] , u5_rsts_reg, u0_rst_r2_reg,
    u0_u0_rst_r2_reg, \\u0_cs_reg[7] , \\u0_wb_addr_r_reg[3] ,
    \\u0_cs_reg[4] , \\u0_spec_req_cs_reg[7] , \\u0_cs_reg[3] ,
    \\u0_spec_req_cs_reg[6] , \\u0_u1_addr_r_reg[3] , \\u0_cs_reg[2] ,
    \\u0_spec_req_cs_reg[3] , \\u1_u0_out_r_reg[0] , \\u0_cs_reg[5] ,
    \\u0_spec_req_cs_reg[2] , u0_init_req_reg, \\u0_u0_addr_r_reg[3] ,
    \\u0_csr_r_reg[0] , u6_read_go_r_reg, u0_lmr_ack_r_reg, u0_lmr_req_reg,
    u5_cke_o_r2_reg, u5_cs_le_r_reg, \\u7_mc_data_o_reg[8] ,
    \\u7_mc_dp_o_reg[3] , \\u7_mc_dp_o_reg[2] , \\u7_mc_data_o_reg[6] ,
    \\u7_mc_data_o_reg[19] , \\u7_mc_data_o_reg[31] , u5_resume_req_r_reg,
    \\u7_mc_data_o_reg[26] , u5_susp_req_r_reg, \\u7_mc_data_o_reg[28] ,
    \\u7_mc_data_o_reg[18] , u0_rst_r1_reg, \\u7_mc_data_o_reg[5] ,
    \\u7_mc_data_o_reg[30] , u0_u0_rst_r1_reg, \\u7_mc_data_o_reg[22] ,
    \\u7_mc_data_o_reg[16] , \\u7_mc_data_o_reg[11] ,
    \\u7_mc_data_o_reg[21] , \\u7_mc_data_o_reg[7] ,
    \\u7_mc_data_o_reg[20] , u0_u1_rst_r1_reg, \\u7_mc_data_o_reg[2] ,
    \\u7_mc_data_o_reg[9] , \\u7_mc_data_o_reg[14] ,
    \\u7_mc_data_o_reg[13] , \\u7_mc_data_o_reg[23] ,
    \\u7_mc_data_o_reg[3] , \\u7_mc_data_o_reg[10] ,
    \\u7_mc_data_o_reg[25] , \\u7_mc_data_o_reg[27] ,
    \\u7_mc_data_o_reg[15] , \\u7_mc_data_o_reg[4] ,
    \\u7_mc_data_o_reg[29] , \\u7_mc_data_o_reg[12] , \\u7_mc_dp_o_reg[0] ,
    u5_rsts1_reg, \\u7_mc_data_o_reg[0] , \\u7_mc_data_o_reg[24] ,
    \\u7_mc_data_o_reg[17] , \\u7_mc_dp_o_reg[1] , \\u7_mc_data_o_reg[1] ,
    \\u7_mc_data_ir_reg[23] , \\u7_mc_data_ir_reg[8] ,
    \\u7_mc_data_ir_reg[6] , \\u0_u0_addr_r_reg[6] ,
    \\u7_mc_data_ir_reg[13] , \\u7_mc_data_ir_reg[14] ,
    \\u7_mc_dqm_r2_reg[3] , \\u7_mc_data_ir_reg[35] ,
    \\u7_mc_data_ir_reg[21] , \\u7_mc_data_ir_reg[7] ,
    \\u7_mc_data_ir_reg[28] , \\u0_wb_addr_r_reg[5] ,
    \\u7_mc_data_ir_reg[22] , \\u7_mc_data_ir_reg[1] ,
    \\u7_mc_data_ir_reg[0] , u7_mc_ack_r_reg, \\u7_mc_data_ir_reg[19] ,
    u5_cs_le_r1_reg, \\u7_mc_data_ir_reg[5] , \\u0_u1_addr_r_reg[4] ,
    \\u7_mc_data_ir_reg[17] , \\u7_mc_dqm_r2_reg[2] ,
    \\u7_mc_data_ir_reg[29] , \\u7_mc_data_ir_reg[18] ,
    \\u7_mc_data_ir_reg[4] , \\u0_u0_addr_r_reg[5] ,
    \\u0_u0_addr_r_reg[4] , \\u7_mc_data_ir_reg[11] ,
    \\u7_mc_data_ir_reg[27] , u7_mc_sts_ir_reg, \\u7_mc_data_ir_reg[10] ,
    \\u0_u1_addr_r_reg[5] , \\u7_mc_data_ir_reg[15] ,
    \\u7_mc_data_ir_reg[34] , \\u7_mc_data_ir_reg[12] ,
    \\u7_mc_data_ir_reg[9] , \\u7_mc_data_ir_reg[33] ,
    \\u7_mc_data_ir_reg[3] , \\u7_mc_dqm_r2_reg[0] ,
    \\u7_mc_data_ir_reg[25] , u5_cke_o_r1_reg, \\u7_mc_data_ir_reg[31] ,
    \\u7_mc_dqm_r2_reg[1] , \\u7_mc_data_ir_reg[26] ,
    \\u7_mc_data_ir_reg[24] , \\u7_mc_data_ir_reg[16] ,
    \\u7_mc_data_ir_reg[30] , u7_mc_br_r_reg, \\u0_wb_addr_r_reg[6] ,
    \\u7_mc_data_ir_reg[2] , \\u0_wb_addr_r_reg[4] ,
    \\u7_mc_data_ir_reg[32] , \\u7_mc_data_ir_reg[20] ,
    \\u0_u1_addr_r_reg[6] ;
  wire new_u5_rsts1_reg_in_, \new_[1379]_ , \new_[1380]_ , \new_[1381]_ ,
    \new_[1382]_ , \new_[1383]_ , \new_[1384]_ , \new_[1385]_ ,
    \new_[1394]_ , \new_[1395]_ , \new_[1396]_ , \new_[1397]_ ,
    \new_[1398]_ , \new_[1399]_ , \new_[1400]_ , \new_[1410]_ ,
    \new_[1411]_ , \new_[1412]_ , \new_[1413]_ , \new_[1414]_ ,
    \new_[1415]_ , \new_[1416]_ , \new_[1417]_ , \new_[1418]_ ,
    \new_[1419]_ , \new_[1420]_ , \new_[1421]_ , \new_[1422]_ ,
    \new_[1423]_ , \new_[1424]_ , \new_[1425]_ , \new_[1426]_ ,
    \new_[1427]_ , \new_[1429]_ , \new_[1430]_ , \new_[1431]_ ,
    \new_[1432]_ , \new_[1433]_ , \new_[1434]_ , \new_[1442]_ ,
    \new_[1443]_ , \new_[1444]_ , \new_[1445]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1458]_ , \new_[1459]_ , \new_[1460]_ , \new_[1461]_ ,
    \new_[1462]_ , \new_[1463]_ , \new_[1464]_ , \new_[1465]_ ,
    \new_[1466]_ , \new_[1467]_ , \new_[1468]_ , \new_[1469]_ ,
    \new_[1470]_ , \new_[1471]_ , \new_[1472]_ , \new_[1473]_ ,
    \new_[1474]_ , \new_[1480]_ , \new_[1481]_ , \new_[1482]_ ,
    \new_[1483]_ , \new_[1484]_ , \new_[1485]_ , \new_[1486]_ ,
    \new_[1487]_ , \new_[1488]_ , \new_[1489]_ , \new_[1490]_ ,
    \new_[1491]_ , \new_[1492]_ , \new_[1493]_ , \new_[1494]_ ,
    \new_[1495]_ , \new_[1496]_ , \new_[1497]_ , \new_[1498]_ ,
    \new_[1499]_ , \new_[1500]_ , \new_[1501]_ , \new_[1502]_ ,
    \new_[1503]_ , \new_[1504]_ , \new_[1505]_ , \new_[1506]_ ,
    \new_[1507]_ , \new_[1519]_ , \new_[1521]_ , \new_[1522]_ ,
    \new_[1523]_ , \new_[1524]_ , \new_[1525]_ , \new_[1526]_ ,
    \new_[1527]_ , \new_[1528]_ , \new_[1529]_ , \new_[1530]_ ,
    \new_[1531]_ , \new_[1532]_ , \new_[1533]_ , \new_[1534]_ ,
    \new_[1535]_ , \new_[1536]_ , \new_[1537]_ , \new_[1538]_ ,
    \new_[1539]_ , \new_[1540]_ , \new_[1541]_ , \new_[1542]_ ,
    \new_[1543]_ , \new_[1544]_ , \new_[1545]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1552]_ , \new_[1554]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1564]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1579]_ , \new_[1580]_ , \new_[1581]_ ,
    \new_[1582]_ , \new_[1593]_ , \new_[1599]_ , \new_[1601]_ ,
    \new_[1602]_ , \new_[1603]_ , \new_[1604]_ , \new_[1605]_ ,
    \new_[1606]_ , \new_[1607]_ , \new_[1609]_ , \new_[1610]_ ,
    \new_[1611]_ , \new_[1612]_ , \new_[1622]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1641]_ ,
    \new_[1642]_ , \new_[1643]_ , \new_[1644]_ , \new_[1645]_ ,
    \new_[1646]_ , \new_[1647]_ , \new_[1648]_ , \new_[1649]_ ,
    \new_[1650]_ , \new_[1651]_ , \new_[1652]_ , \new_[1653]_ ,
    \new_[1655]_ , \new_[1656]_ , \new_[1657]_ , \new_[1658]_ ,
    \new_[1659]_ , \new_[1660]_ , \new_[1661]_ , \new_[1662]_ ,
    \new_[1663]_ , \new_[1664]_ , \new_[1665]_ , \new_[1666]_ ,
    \new_[1667]_ , \new_[1668]_ , \new_[1669]_ , \new_[1670]_ ,
    \new_[1672]_ , \new_[1673]_ , \new_[1674]_ , \new_[1675]_ ,
    \new_[1676]_ , \new_[1677]_ , \new_[1678]_ , \new_[1679]_ ,
    \new_[1680]_ , \new_[1681]_ , \new_[1682]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1690]_ , \new_[1691]_ , \new_[1692]_ , \new_[1693]_ ,
    \new_[1694]_ , \new_[1695]_ , \new_[1696]_ , \new_[1697]_ ,
    \new_[1698]_ , \new_[1699]_ , \new_[1700]_ , \new_[1701]_ ,
    \new_[1702]_ , \new_[1703]_ , \new_[1704]_ , \new_[1705]_ ,
    \new_[1706]_ , \new_[1707]_ , \new_[1708]_ , \new_[1709]_ ,
    \new_[1710]_ , \new_[1711]_ , \new_[1712]_ , \new_[1713]_ ,
    \new_[1714]_ , \new_[1715]_ , \new_[1716]_ , \new_[1717]_ ,
    \new_[1718]_ , \new_[1719]_ , \new_[1720]_ , \new_[1721]_ ,
    \new_[1722]_ , \new_[1723]_ , \new_[1724]_ , \new_[1725]_ ,
    \new_[1728]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1793]_ ,
    \new_[1796]_ , \new_[1797]_ , \new_[1798]_ , \new_[1799]_ ,
    \new_[1800]_ , \new_[1801]_ , \new_[1802]_ , \new_[1803]_ ,
    \new_[1804]_ , \new_[1805]_ , \new_[1806]_ , \new_[1807]_ ,
    \new_[1808]_ , \new_[1809]_ , \new_[1810]_ , \new_[1811]_ ,
    \new_[1812]_ , \new_[1813]_ , \new_[1814]_ , \new_[1815]_ ,
    \new_[1816]_ , \new_[1817]_ , \new_[1818]_ , \new_[1819]_ ,
    \new_[1820]_ , \new_[1821]_ , \new_[1822]_ , \new_[1823]_ ,
    \new_[1824]_ , \new_[1825]_ , \new_[1826]_ , \new_[1827]_ ,
    \new_[1828]_ , \new_[1829]_ , \new_[1830]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1837]_ ,
    \new_[1838]_ , \new_[1839]_ , \new_[1840]_ , \new_[1841]_ ,
    \new_[1842]_ , \new_[1843]_ , \new_[1844]_ , \new_[1845]_ ,
    \new_[1846]_ , \new_[1847]_ , \new_[1848]_ , \new_[1849]_ ,
    \new_[1850]_ , \new_[1851]_ , \new_[1852]_ , \new_[1853]_ ,
    \new_[1854]_ , \new_[1855]_ , \new_[1856]_ , \new_[1857]_ ,
    \new_[1858]_ , \new_[1859]_ , \new_[1860]_ , \new_[1861]_ ,
    \new_[1862]_ , \new_[1863]_ , \new_[1864]_ , \new_[1865]_ ,
    \new_[1866]_ , \new_[1867]_ , \new_[1868]_ , \new_[1869]_ ,
    \new_[1870]_ , \new_[1871]_ , \new_[1872]_ , \new_[1873]_ ,
    \new_[1874]_ , \new_[1875]_ , \new_[1876]_ , \new_[1877]_ ,
    \new_[1878]_ , \new_[1879]_ , \new_[1880]_ , \new_[1881]_ ,
    \new_[1882]_ , \new_[1883]_ , \new_[1884]_ , \new_[1885]_ ,
    \new_[1886]_ , \new_[1887]_ , \new_[1888]_ , \new_[1889]_ ,
    \new_[1890]_ , \new_[1891]_ , \new_[1892]_ , \new_[1893]_ ,
    \new_[1894]_ , \new_[1895]_ , \new_[1896]_ , \new_[1897]_ ,
    \new_[1898]_ , \new_[1899]_ , \new_[1900]_ , \new_[1901]_ ,
    \new_[1902]_ , \new_[1903]_ , \new_[1904]_ , \new_[1905]_ ,
    \new_[1906]_ , \new_[1907]_ , \new_[1908]_ , \new_[1909]_ ,
    \new_[1910]_ , \new_[1911]_ , \new_[1912]_ , \new_[1913]_ ,
    \new_[1914]_ , \new_[1915]_ , \new_[1916]_ , \new_[1917]_ ,
    \new_[1918]_ , \new_[1919]_ , \new_[1920]_ , \new_[1921]_ ,
    \new_[1922]_ , \new_[1923]_ , \new_[1924]_ , \new_[1925]_ ,
    \new_[1926]_ , \new_[1927]_ , \new_[1928]_ , \new_[1929]_ ,
    \new_[1930]_ , \new_[1931]_ , \new_[1932]_ , \new_[1933]_ ,
    \new_[1934]_ , \new_[1935]_ , \new_[1936]_ , \new_[1937]_ ,
    \new_[1938]_ , \new_[1939]_ , \new_[1940]_ , \new_[1941]_ ,
    \new_[1942]_ , \new_[1943]_ , \new_[1944]_ , \new_[1945]_ ,
    \new_[1946]_ , \new_[1947]_ , \new_[1948]_ , \new_[1949]_ ,
    \new_[1950]_ , \new_[1951]_ , \new_[1954]_ , \new_[1955]_ ,
    \new_[1956]_ , \new_[1957]_ , \new_[1958]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2021]_ ,
    \new_[2022]_ , \new_[2023]_ , \new_[2024]_ , \new_[2025]_ ,
    \new_[2026]_ , \new_[2027]_ , \new_[2028]_ , \new_[2029]_ ,
    \new_[2030]_ , \new_[2031]_ , \new_[2032]_ , \new_[2033]_ ,
    \new_[2034]_ , \new_[2035]_ , \new_[2036]_ , \new_[2037]_ ,
    \new_[2038]_ , \new_[2039]_ , \new_[2040]_ , \new_[2041]_ ,
    \new_[2042]_ , \new_[2043]_ , \new_[2044]_ , \new_[2045]_ ,
    \new_[2046]_ , \new_[2047]_ , \new_[2048]_ , \new_[2049]_ ,
    \new_[2050]_ , \new_[2051]_ , \new_[2052]_ , \new_[2053]_ ,
    \new_[2054]_ , \new_[2055]_ , \new_[2056]_ , \new_[2057]_ ,
    \new_[2058]_ , \new_[2059]_ , \new_[2060]_ , \new_[2061]_ ,
    \new_[2062]_ , \new_[2063]_ , \new_[2064]_ , \new_[2065]_ ,
    \new_[2066]_ , \new_[2067]_ , \new_[2068]_ , \new_[2069]_ ,
    \new_[2070]_ , \new_[2071]_ , \new_[2072]_ , \new_[2073]_ ,
    \new_[2074]_ , \new_[2075]_ , \new_[2076]_ , \new_[2077]_ ,
    \new_[2078]_ , \new_[2079]_ , \new_[2081]_ , \new_[2082]_ ,
    \new_[2083]_ , \new_[2084]_ , \new_[2085]_ , \new_[2087]_ ,
    \new_[2088]_ , \new_[2089]_ , \new_[2090]_ , \new_[2091]_ ,
    \new_[2092]_ , \new_[2093]_ , \new_[2094]_ , \new_[2095]_ ,
    \new_[2096]_ , \new_[2097]_ , \new_[2098]_ , \new_[2099]_ ,
    \new_[2100]_ , \new_[2101]_ , \new_[2102]_ , \new_[2103]_ ,
    \new_[2104]_ , \new_[2105]_ , \new_[2106]_ , \new_[2107]_ ,
    \new_[2108]_ , \new_[2109]_ , \new_[2110]_ , \new_[2111]_ ,
    \new_[2112]_ , \new_[2113]_ , \new_[2114]_ , \new_[2115]_ ,
    \new_[2116]_ , \new_[2117]_ , \new_[2118]_ , \new_[2119]_ ,
    \new_[2120]_ , \new_[2121]_ , \new_[2122]_ , \new_[2123]_ ,
    \new_[2124]_ , \new_[2125]_ , \new_[2126]_ , \new_[2127]_ ,
    \new_[2128]_ , \new_[2129]_ , \new_[2130]_ , \new_[2131]_ ,
    \new_[2132]_ , \new_[2133]_ , \new_[2134]_ , \new_[2135]_ ,
    \new_[2136]_ , \new_[2137]_ , \new_[2138]_ , \new_[2139]_ ,
    \new_[2140]_ , \new_[2141]_ , \new_[2142]_ , \new_[2143]_ ,
    \new_[2144]_ , \new_[2145]_ , \new_[2146]_ , \new_[2147]_ ,
    \new_[2148]_ , \new_[2149]_ , \new_[2150]_ , \new_[2151]_ ,
    \new_[2152]_ , \new_[2153]_ , \new_[2154]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2226]_ ,
    \new_[2227]_ , \new_[2228]_ , \new_[2229]_ , \new_[2230]_ ,
    \new_[2231]_ , \new_[2232]_ , \new_[2233]_ , \new_[2234]_ ,
    \new_[2235]_ , \new_[2236]_ , \new_[2237]_ , \new_[2238]_ ,
    \new_[2239]_ , \new_[2240]_ , \new_[2241]_ , \new_[2242]_ ,
    \new_[2243]_ , \new_[2244]_ , \new_[2245]_ , \new_[2246]_ ,
    \new_[2247]_ , \new_[2248]_ , \new_[2249]_ , \new_[2250]_ ,
    \new_[2251]_ , \new_[2252]_ , \new_[2253]_ , \new_[2254]_ ,
    \new_[2255]_ , \new_[2256]_ , \new_[2257]_ , \new_[2258]_ ,
    \new_[2259]_ , \new_[2260]_ , \new_[2261]_ , \new_[2262]_ ,
    \new_[2263]_ , \new_[2264]_ , \new_[2265]_ , \new_[2266]_ ,
    \new_[2267]_ , \new_[2268]_ , \new_[2269]_ , \new_[2270]_ ,
    \new_[2271]_ , \new_[2272]_ , \new_[2273]_ , \new_[2274]_ ,
    \new_[2275]_ , \new_[2276]_ , \new_[2277]_ , \new_[2278]_ ,
    \new_[2279]_ , \new_[2280]_ , \new_[2281]_ , \new_[2282]_ ,
    \new_[2283]_ , \new_[2284]_ , \new_[2285]_ , \new_[2286]_ ,
    \new_[2287]_ , \new_[2288]_ , \new_[2289]_ , \new_[2290]_ ,
    \new_[2291]_ , \new_[2292]_ , \new_[2293]_ , \new_[2294]_ ,
    \new_[2295]_ , \new_[2296]_ , \new_[2297]_ , \new_[2298]_ ,
    \new_[2299]_ , \new_[2300]_ , \new_[2301]_ , \new_[2302]_ ,
    \new_[2303]_ , \new_[2304]_ , \new_[2305]_ , \new_[2306]_ ,
    \new_[2307]_ , \new_[2308]_ , \new_[2309]_ , \new_[2310]_ ,
    \new_[2311]_ , \new_[2312]_ , \new_[2313]_ , \new_[2314]_ ,
    \new_[2315]_ , \new_[2316]_ , \new_[2317]_ , \new_[2318]_ ,
    \new_[2319]_ , \new_[2320]_ , \new_[2321]_ , \new_[2322]_ ,
    \new_[2323]_ , \new_[2324]_ , \new_[2325]_ , \new_[2326]_ ,
    \new_[2327]_ , \new_[2328]_ , \new_[2329]_ , \new_[2330]_ ,
    \new_[2331]_ , \new_[2332]_ , \new_[2333]_ , \new_[2334]_ ,
    \new_[2335]_ , \new_[2336]_ , \new_[2337]_ , \new_[2338]_ ,
    \new_[2339]_ , \new_[2340]_ , \new_[2341]_ , \new_[2342]_ ,
    \new_[2343]_ , \new_[2344]_ , \new_[2345]_ , \new_[2346]_ ,
    \new_[2347]_ , \new_[2348]_ , \new_[2349]_ , \new_[2350]_ ,
    \new_[2351]_ , \new_[2352]_ , \new_[2353]_ , \new_[2354]_ ,
    \new_[2355]_ , \new_[2356]_ , \new_[2357]_ , \new_[2358]_ ,
    \new_[2359]_ , \new_[2360]_ , \new_[2361]_ , \new_[2362]_ ,
    \new_[2363]_ , \new_[2364]_ , \new_[2365]_ , \new_[2366]_ ,
    \new_[2367]_ , \new_[2368]_ , \new_[2369]_ , \new_[2370]_ ,
    \new_[2371]_ , \new_[2372]_ , \new_[2373]_ , \new_[2374]_ ,
    \new_[2375]_ , \new_[2376]_ , \new_[2377]_ , \new_[2378]_ ,
    \new_[2379]_ , \new_[2380]_ , \new_[2381]_ , \new_[2382]_ ,
    \new_[2383]_ , \new_[2384]_ , \new_[2385]_ , \new_[2386]_ ,
    \new_[2387]_ , \new_[2388]_ , \new_[2389]_ , \new_[2390]_ ,
    \new_[2391]_ , \new_[2395]_ , \new_[2396]_ , \new_[2397]_ ,
    \new_[2398]_ , \new_[2399]_ , \new_[2400]_ , \new_[2401]_ ,
    \new_[2402]_ , \new_[2403]_ , \new_[2404]_ , \new_[2405]_ ,
    \new_[2406]_ , \new_[2407]_ , \new_[2408]_ , \new_[2409]_ ,
    \new_[2410]_ , \new_[2411]_ , \new_[2412]_ , \new_[2413]_ ,
    \new_[2414]_ , \new_[2415]_ , \new_[2416]_ , \new_[2417]_ ,
    \new_[2418]_ , \new_[2419]_ , \new_[2420]_ , \new_[2421]_ ,
    \new_[2422]_ , \new_[2423]_ , \new_[2424]_ , \new_[2425]_ ,
    \new_[2426]_ , \new_[2427]_ , \new_[2428]_ , \new_[2429]_ ,
    \new_[2430]_ , \new_[2431]_ , \new_[2432]_ , \new_[2433]_ ,
    \new_[2434]_ , \new_[2435]_ , \new_[2436]_ , \new_[2437]_ ,
    \new_[2438]_ , \new_[2451]_ , \new_[2452]_ , \new_[2453]_ ,
    \new_[2454]_ , \new_[2455]_ , \new_[2456]_ , \new_[2457]_ ,
    \new_[2458]_ , \new_[2459]_ , \new_[2460]_ , \new_[2461]_ ,
    \new_[2462]_ , \new_[2463]_ , \new_[2464]_ , \new_[2465]_ ,
    \new_[2466]_ , \new_[2467]_ , \new_[2468]_ , \new_[2469]_ ,
    \new_[2470]_ , \new_[2471]_ , \new_[2472]_ , \new_[2473]_ ,
    \new_[2474]_ , \new_[2475]_ , \new_[2476]_ , \new_[2477]_ ,
    \new_[2478]_ , \new_[2479]_ , \new_[2481]_ , \new_[2482]_ ,
    \new_[2483]_ , \new_[2484]_ , \new_[2485]_ , \new_[2486]_ ,
    \new_[2487]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2512]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2518]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2525]_ , \new_[2526]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2552]_ ,
    \new_[2553]_ , \new_[2554]_ , \new_[2555]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2559]_ , \new_[2560]_ ,
    \new_[2561]_ , \new_[2562]_ , \new_[2563]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2567]_ , \new_[2568]_ ,
    \new_[2569]_ , \new_[2573]_ , \new_[2574]_ , \new_[2575]_ ,
    \new_[2576]_ , \new_[2577]_ , \new_[2578]_ , \new_[2579]_ ,
    \new_[2580]_ , \new_[2581]_ , \new_[2582]_ , \new_[2583]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2587]_ , \new_[2588]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2599]_ , \new_[2600]_ ,
    \new_[2601]_ , \new_[2604]_ , \new_[2605]_ , \new_[2606]_ ,
    \new_[2607]_ , \new_[2608]_ , \new_[2609]_ , \new_[2610]_ ,
    \new_[2611]_ , \new_[2612]_ , \new_[2613]_ , \new_[2614]_ ,
    \new_[2615]_ , \new_[2616]_ , \new_[2617]_ , \new_[2618]_ ,
    \new_[2620]_ , \new_[2621]_ , \new_[2622]_ , \new_[2623]_ ,
    \new_[2625]_ , \new_[2626]_ , \new_[2627]_ , \new_[2628]_ ,
    \new_[2629]_ , \new_[2631]_ , \new_[2632]_ , \new_[2633]_ ,
    \new_[2634]_ , \new_[2635]_ , \new_[2636]_ , \new_[2639]_ ,
    \new_[2640]_ , \new_[2641]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2644]_ , \new_[2645]_ , \new_[2646]_ , \new_[2647]_ ,
    \new_[2648]_ , \new_[2649]_ , \new_[2650]_ , \new_[2651]_ ,
    \new_[2652]_ , \new_[2653]_ , \new_[2654]_ , \new_[2655]_ ,
    \new_[2656]_ , \new_[2657]_ , \new_[2658]_ , \new_[2659]_ ,
    \new_[2660]_ , \new_[2661]_ , \new_[2662]_ , \new_[2663]_ ,
    \new_[2664]_ , \new_[2665]_ , \new_[2666]_ , \new_[2667]_ ,
    \new_[2668]_ , \new_[2669]_ , \new_[2670]_ , \new_[2671]_ ,
    \new_[2672]_ , \new_[2673]_ , \new_[2674]_ , \new_[2675]_ ,
    \new_[2676]_ , \new_[2677]_ , \new_[2678]_ , \new_[2679]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2725]_ ,
    \new_[2726]_ , \new_[2727]_ , \new_[2728]_ , \new_[2729]_ ,
    \new_[2730]_ , \new_[2731]_ , \new_[2732]_ , \new_[2733]_ ,
    \new_[2734]_ , \new_[2735]_ , \new_[2736]_ , \new_[2737]_ ,
    \new_[2738]_ , \new_[2739]_ , \new_[2740]_ , \new_[2741]_ ,
    \new_[2742]_ , \new_[2743]_ , \new_[2744]_ , \new_[2745]_ ,
    \new_[2746]_ , \new_[2747]_ , \new_[2748]_ , \new_[2749]_ ,
    \new_[2750]_ , \new_[2751]_ , \new_[2752]_ , \new_[2753]_ ,
    \new_[2754]_ , \new_[2755]_ , \new_[2756]_ , \new_[2757]_ ,
    \new_[2758]_ , \new_[2759]_ , \new_[2760]_ , \new_[2761]_ ,
    \new_[2762]_ , \new_[2763]_ , \new_[2764]_ , \new_[2765]_ ,
    \new_[2766]_ , \new_[2767]_ , \new_[2768]_ , \new_[2769]_ ,
    \new_[2770]_ , \new_[2771]_ , \new_[2772]_ , \new_[2773]_ ,
    \new_[2774]_ , \new_[2775]_ , \new_[2776]_ , \new_[2777]_ ,
    \new_[2778]_ , \new_[2779]_ , \new_[2780]_ , \new_[2781]_ ,
    \new_[2782]_ , \new_[2783]_ , \new_[2784]_ , \new_[2785]_ ,
    \new_[2786]_ , \new_[2787]_ , \new_[2788]_ , \new_[2789]_ ,
    \new_[2790]_ , \new_[2791]_ , \new_[2792]_ , \new_[2793]_ ,
    \new_[2794]_ , \new_[2795]_ , \new_[2796]_ , \new_[2797]_ ,
    \new_[2798]_ , \new_[2799]_ , \new_[2800]_ , \new_[2802]_ ,
    \new_[2803]_ , \new_[2804]_ , \new_[2805]_ , \new_[2806]_ ,
    \new_[2807]_ , \new_[2808]_ , \new_[2809]_ , \new_[2810]_ ,
    \new_[2811]_ , \new_[2812]_ , \new_[2813]_ , \new_[2814]_ ,
    \new_[2815]_ , \new_[2816]_ , \new_[2817]_ , \new_[2818]_ ,
    \new_[2819]_ , \new_[2820]_ , \new_[2824]_ , \new_[2825]_ ,
    \new_[2826]_ , \new_[2827]_ , \new_[2828]_ , \new_[2829]_ ,
    \new_[2830]_ , \new_[2831]_ , \new_[2832]_ , \new_[2833]_ ,
    \new_[2834]_ , \new_[2835]_ , \new_[2836]_ , \new_[2837]_ ,
    \new_[2838]_ , \new_[2839]_ , \new_[2840]_ , \new_[2841]_ ,
    \new_[2842]_ , \new_[2843]_ , \new_[2844]_ , \new_[2845]_ ,
    \new_[2846]_ , \new_[2847]_ , \new_[2848]_ , \new_[2849]_ ,
    \new_[2850]_ , \new_[2851]_ , \new_[2852]_ , \new_[2853]_ ,
    \new_[2854]_ , \new_[2855]_ , \new_[2856]_ , \new_[2857]_ ,
    \new_[2858]_ , \new_[2859]_ , \new_[2860]_ , \new_[2861]_ ,
    \new_[2862]_ , \new_[2863]_ , \new_[2864]_ , \new_[2865]_ ,
    \new_[2866]_ , \new_[2868]_ , \new_[2869]_ , \new_[2870]_ ,
    \new_[2871]_ , \new_[2872]_ , \new_[2873]_ , \new_[2874]_ ,
    \new_[2875]_ , \new_[2876]_ , \new_[2877]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2880]_ , \new_[2881]_ , \new_[2882]_ ,
    \new_[2883]_ , \new_[2884]_ , \new_[2887]_ , \new_[2888]_ ,
    \new_[2889]_ , \new_[2890]_ , \new_[2891]_ , \new_[2892]_ ,
    \new_[2893]_ , \new_[2894]_ , \new_[2895]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2898]_ , \new_[2899]_ , \new_[2900]_ ,
    \new_[2901]_ , \new_[2902]_ , \new_[2903]_ , \new_[2904]_ ,
    \new_[2905]_ , \new_[2906]_ , \new_[2907]_ , \new_[2908]_ ,
    \new_[2909]_ , \new_[2910]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2915]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2934]_ , \new_[2935]_ , \new_[2936]_ ,
    \new_[2937]_ , \new_[2938]_ , \new_[2939]_ , \new_[2940]_ ,
    \new_[2941]_ , \new_[2942]_ , \new_[2943]_ , \new_[2944]_ ,
    \new_[2945]_ , \new_[2946]_ , \new_[2947]_ , \new_[2948]_ ,
    \new_[2950]_ , \new_[2951]_ , \new_[2952]_ , \new_[2953]_ ,
    \new_[2954]_ , \new_[2955]_ , \new_[2956]_ , \new_[2957]_ ,
    \new_[2958]_ , \new_[2959]_ , \new_[2960]_ , \new_[2961]_ ,
    \new_[2962]_ , \new_[2963]_ , \new_[2964]_ , \new_[2965]_ ,
    \new_[2966]_ , \new_[2967]_ , \new_[2968]_ , \new_[2969]_ ,
    \new_[2970]_ , \new_[2971]_ , \new_[2972]_ , \new_[2982]_ ,
    \new_[2983]_ , \new_[2984]_ , \new_[2985]_ , \new_[2986]_ ,
    \new_[2987]_ , \new_[2988]_ , \new_[2989]_ , \new_[2990]_ ,
    \new_[2991]_ , \new_[2992]_ , \new_[2993]_ , \new_[2994]_ ,
    \new_[2995]_ , \new_[2996]_ , \new_[2997]_ , \new_[2998]_ ,
    \new_[2999]_ , \new_[3000]_ , \new_[3001]_ , \new_[3002]_ ,
    \new_[3003]_ , \new_[3004]_ , \new_[3005]_ , \new_[3006]_ ,
    \new_[3007]_ , \new_[3008]_ , \new_[3009]_ , \new_[3010]_ ,
    \new_[3011]_ , \new_[3012]_ , \new_[3013]_ , \new_[3014]_ ,
    \new_[3015]_ , \new_[3016]_ , \new_[3017]_ , \new_[3018]_ ,
    \new_[3019]_ , \new_[3020]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3023]_ , \new_[3024]_ , \new_[3025]_ , \new_[3026]_ ,
    \new_[3027]_ , \new_[3028]_ , \new_[3029]_ , \new_[3030]_ ,
    \new_[3031]_ , \new_[3032]_ , \new_[3033]_ , \new_[3034]_ ,
    \new_[3035]_ , \new_[3036]_ , \new_[3037]_ , \new_[3038]_ ,
    \new_[3039]_ , \new_[3040]_ , \new_[3041]_ , \new_[3042]_ ,
    \new_[3043]_ , \new_[3044]_ , \new_[3045]_ , \new_[3046]_ ,
    \new_[3047]_ , \new_[3048]_ , \new_[3049]_ , \new_[3050]_ ,
    \new_[3051]_ , \new_[3052]_ , \new_[3053]_ , \new_[3054]_ ,
    \new_[3055]_ , \new_[3056]_ , \new_[3057]_ , \new_[3058]_ ,
    \new_[3059]_ , \new_[3060]_ , \new_[3061]_ , \new_[3062]_ ,
    \new_[3063]_ , \new_[3064]_ , \new_[3065]_ , \new_[3066]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3069]_ , \new_[3070]_ ,
    \new_[3071]_ , \new_[3072]_ , \new_[3073]_ , \new_[3074]_ ,
    \new_[3075]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3082]_ , \new_[3083]_ ,
    \new_[3084]_ , \new_[3085]_ , \new_[3086]_ , \new_[3087]_ ,
    \new_[3088]_ , \new_[3089]_ , \new_[3090]_ , \new_[3091]_ ,
    \new_[3092]_ , \new_[3093]_ , \new_[3094]_ , \new_[3095]_ ,
    \new_[3096]_ , \new_[3097]_ , \new_[3098]_ , \new_[3099]_ ,
    \new_[3100]_ , \new_[3101]_ , \new_[3102]_ , \new_[3103]_ ,
    \new_[3104]_ , \new_[3105]_ , \new_[3106]_ , \new_[3107]_ ,
    \new_[3108]_ , \new_[3109]_ , \new_[3110]_ , \new_[3111]_ ,
    \new_[3112]_ , \new_[3113]_ , \new_[3114]_ , \new_[3115]_ ,
    \new_[3116]_ , \new_[3117]_ , \new_[3118]_ , \new_[3119]_ ,
    \new_[3120]_ , \new_[3121]_ , \new_[3122]_ , \new_[3123]_ ,
    \new_[3124]_ , \new_[3125]_ , \new_[3126]_ , \new_[3127]_ ,
    \new_[3128]_ , \new_[3129]_ , \new_[3130]_ , \new_[3131]_ ,
    \new_[3132]_ , \new_[3133]_ , \new_[3134]_ , \new_[3135]_ ,
    \new_[3136]_ , \new_[3137]_ , \new_[3138]_ , \new_[3139]_ ,
    \new_[3140]_ , \new_[3141]_ , \new_[3142]_ , \new_[3143]_ ,
    \new_[3144]_ , \new_[3145]_ , \new_[3146]_ , \new_[3147]_ ,
    \new_[3148]_ , \new_[3149]_ , \new_[3150]_ , \new_[3151]_ ,
    \new_[3152]_ , \new_[3153]_ , \new_[3154]_ , \new_[3155]_ ,
    \new_[3156]_ , \new_[3157]_ , \new_[3158]_ , \new_[3159]_ ,
    \new_[3160]_ , \new_[3161]_ , \new_[3162]_ , \new_[3163]_ ,
    \new_[3164]_ , \new_[3165]_ , \new_[3166]_ , \new_[3167]_ ,
    \new_[3168]_ , \new_[3169]_ , \new_[3170]_ , \new_[3171]_ ,
    \new_[3172]_ , \new_[3173]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3177]_ , \new_[3178]_ , \new_[3179]_ ,
    \new_[3180]_ , \new_[3181]_ , \new_[3182]_ , \new_[3183]_ ,
    \new_[3184]_ , \new_[3185]_ , \new_[3186]_ , \new_[3187]_ ,
    \new_[3188]_ , \new_[3189]_ , \new_[3190]_ , \new_[3191]_ ,
    \new_[3192]_ , \new_[3193]_ , \new_[3194]_ , \new_[3195]_ ,
    \new_[3196]_ , \new_[3197]_ , \new_[3198]_ , \new_[3199]_ ,
    \new_[3200]_ , \new_[3201]_ , \new_[3202]_ , \new_[3203]_ ,
    \new_[3204]_ , \new_[3205]_ , \new_[3206]_ , \new_[3207]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3222]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3226]_ , \new_[3227]_ , \new_[3228]_ ,
    \new_[3229]_ , \new_[3230]_ , \new_[3231]_ , \new_[3232]_ ,
    \new_[3233]_ , \new_[3234]_ , \new_[3235]_ , \new_[3236]_ ,
    \new_[3237]_ , \new_[3238]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3246]_ , \new_[3247]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3251]_ , \new_[3252]_ ,
    \new_[3253]_ , \new_[3254]_ , \new_[3255]_ , \new_[3256]_ ,
    \new_[3257]_ , \new_[3258]_ , \new_[3259]_ , \new_[3260]_ ,
    \new_[3261]_ , \new_[3262]_ , \new_[3263]_ , \new_[3264]_ ,
    \new_[3265]_ , \new_[3266]_ , \new_[3267]_ , \new_[3268]_ ,
    \new_[3269]_ , \new_[3270]_ , \new_[3271]_ , \new_[3272]_ ,
    \new_[3273]_ , \new_[3274]_ , \new_[3275]_ , \new_[3276]_ ,
    \new_[3277]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3281]_ , \new_[3282]_ , \new_[3283]_ , \new_[3284]_ ,
    \new_[3285]_ , \new_[3286]_ , \new_[3287]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3294]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3299]_ , \new_[3301]_ ,
    \new_[3302]_ , \new_[3303]_ , \new_[3305]_ , \new_[3307]_ ,
    \new_[3308]_ , \new_[3317]_ , \new_[3318]_ , \new_[3319]_ ,
    \new_[3320]_ , \new_[3321]_ , \new_[3322]_ , \new_[3323]_ ,
    \new_[3326]_ , \new_[3327]_ , \new_[3328]_ , \new_[3329]_ ,
    \new_[3330]_ , \new_[3331]_ , \new_[3332]_ , \new_[3333]_ ,
    \new_[3335]_ , \new_[3336]_ , \new_[3337]_ , \new_[3338]_ ,
    \new_[3339]_ , \new_[3340]_ , \new_[3341]_ , \new_[3342]_ ,
    \new_[3343]_ , \new_[3344]_ , \new_[3345]_ , \new_[3346]_ ,
    \new_[3347]_ , \new_[3348]_ , \new_[3349]_ , \new_[3350]_ ,
    \new_[3351]_ , \new_[3352]_ , \new_[3353]_ , \new_[3354]_ ,
    \new_[3355]_ , \new_[3356]_ , \new_[3357]_ , \new_[3358]_ ,
    \new_[3359]_ , \new_[3360]_ , \new_[3361]_ , \new_[3362]_ ,
    \new_[3364]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3371]_ , \new_[3372]_ , \new_[3373]_ ,
    \new_[3374]_ , \new_[3375]_ , \new_[3376]_ , \new_[3377]_ ,
    \new_[3378]_ , \new_[3379]_ , \new_[3380]_ , \new_[3381]_ ,
    \new_[3382]_ , \new_[3383]_ , \new_[3384]_ , \new_[3385]_ ,
    \new_[3386]_ , \new_[3387]_ , \new_[3388]_ , \new_[3389]_ ,
    \new_[3390]_ , \new_[3391]_ , \new_[3392]_ , \new_[3393]_ ,
    \new_[3394]_ , \new_[3395]_ , \new_[3396]_ , \new_[3397]_ ,
    \new_[3398]_ , \new_[3399]_ , \new_[3400]_ , \new_[3401]_ ,
    \new_[3402]_ , \new_[3403]_ , \new_[3404]_ , \new_[3405]_ ,
    \new_[3406]_ , \new_[3407]_ , \new_[3408]_ , \new_[3409]_ ,
    \new_[3410]_ , \new_[3411]_ , \new_[3412]_ , \new_[3413]_ ,
    \new_[3414]_ , \new_[3415]_ , \new_[3416]_ , \new_[3417]_ ,
    \new_[3418]_ , \new_[3419]_ , \new_[3420]_ , \new_[3421]_ ,
    \new_[3422]_ , \new_[3423]_ , \new_[3424]_ , \new_[3425]_ ,
    \new_[3426]_ , \new_[3427]_ , \new_[3428]_ , \new_[3429]_ ,
    \new_[3430]_ , \new_[3431]_ , \new_[3432]_ , \new_[3433]_ ,
    \new_[3434]_ , \new_[3435]_ , \new_[3436]_ , \new_[3437]_ ,
    \new_[3438]_ , \new_[3439]_ , \new_[3440]_ , \new_[3441]_ ,
    \new_[3442]_ , \new_[3443]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3470]_ , \new_[3471]_ , \new_[3472]_ , \new_[3473]_ ,
    \new_[3474]_ , \new_[3475]_ , \new_[3476]_ , \new_[3477]_ ,
    \new_[3478]_ , \new_[3479]_ , \new_[3480]_ , \new_[3481]_ ,
    \new_[3482]_ , \new_[3483]_ , \new_[3484]_ , \new_[3485]_ ,
    \new_[3486]_ , \new_[3487]_ , \new_[3488]_ , \new_[3489]_ ,
    \new_[3490]_ , \new_[3491]_ , \new_[3492]_ , \new_[3493]_ ,
    \new_[3494]_ , \new_[3495]_ , \new_[3496]_ , \new_[3497]_ ,
    \new_[3498]_ , \new_[3499]_ , \new_[3500]_ , \new_[3501]_ ,
    \new_[3502]_ , \new_[3503]_ , \new_[3504]_ , \new_[3505]_ ,
    \new_[3506]_ , \new_[3507]_ , \new_[3508]_ , \new_[3509]_ ,
    \new_[3510]_ , \new_[3512]_ , \new_[3513]_ , \new_[3514]_ ,
    \new_[3515]_ , \new_[3516]_ , \new_[3517]_ , \new_[3518]_ ,
    \new_[3519]_ , \new_[3520]_ , \new_[3521]_ , \new_[3522]_ ,
    \new_[3523]_ , \new_[3524]_ , \new_[3525]_ , \new_[3526]_ ,
    \new_[3527]_ , \new_[3528]_ , \new_[3529]_ , \new_[3530]_ ,
    \new_[3531]_ , \new_[3532]_ , \new_[3533]_ , \new_[3534]_ ,
    \new_[3535]_ , \new_[3536]_ , \new_[3537]_ , \new_[3538]_ ,
    \new_[3539]_ , \new_[3540]_ , \new_[3541]_ , \new_[3542]_ ,
    \new_[3543]_ , \new_[3544]_ , \new_[3545]_ , \new_[3546]_ ,
    \new_[3547]_ , \new_[3548]_ , \new_[3549]_ , \new_[3550]_ ,
    \new_[3551]_ , \new_[3552]_ , \new_[3553]_ , \new_[3554]_ ,
    \new_[3555]_ , \new_[3556]_ , \new_[3557]_ , \new_[3558]_ ,
    \new_[3559]_ , \new_[3560]_ , \new_[3561]_ , \new_[3562]_ ,
    \new_[3563]_ , \new_[3564]_ , \new_[3565]_ , \new_[3566]_ ,
    \new_[3567]_ , \new_[3568]_ , \new_[3569]_ , \new_[3570]_ ,
    \new_[3571]_ , \new_[3572]_ , \new_[3573]_ , \new_[3574]_ ,
    \new_[3575]_ , \new_[3576]_ , \new_[3577]_ , \new_[3578]_ ,
    \new_[3579]_ , \new_[3580]_ , \new_[3581]_ , \new_[3582]_ ,
    \new_[3583]_ , \new_[3584]_ , \new_[3585]_ , \new_[3586]_ ,
    \new_[3587]_ , \new_[3588]_ , \new_[3589]_ , \new_[3590]_ ,
    \new_[3591]_ , \new_[3592]_ , \new_[3593]_ , \new_[3594]_ ,
    \new_[3595]_ , \new_[3596]_ , \new_[3597]_ , \new_[3598]_ ,
    \new_[3599]_ , \new_[3600]_ , \new_[3601]_ , \new_[3602]_ ,
    \new_[3603]_ , \new_[3604]_ , \new_[3605]_ , \new_[3606]_ ,
    \new_[3607]_ , \new_[3608]_ , \new_[3609]_ , \new_[3610]_ ,
    \new_[3611]_ , \new_[3612]_ , \new_[3613]_ , \new_[3614]_ ,
    \new_[3615]_ , \new_[3616]_ , \new_[3617]_ , \new_[3618]_ ,
    \new_[3619]_ , \new_[3620]_ , \new_[3621]_ , \new_[3622]_ ,
    \new_[3623]_ , \new_[3624]_ , \new_[3625]_ , \new_[3626]_ ,
    \new_[3631]_ , \new_[3632]_ , \new_[3633]_ , \new_[3634]_ ,
    \new_[3635]_ , \new_[3636]_ , \new_[3637]_ , \new_[3638]_ ,
    \new_[3639]_ , \new_[3640]_ , \new_[3641]_ , \new_[3642]_ ,
    \new_[3643]_ , \new_[3644]_ , \new_[3645]_ , \new_[3646]_ ,
    \new_[3647]_ , \new_[3648]_ , \new_[3649]_ , \new_[3650]_ ,
    \new_[3651]_ , \new_[3652]_ , \new_[3653]_ , \new_[3654]_ ,
    \new_[3655]_ , \new_[3656]_ , \new_[3657]_ , \new_[3658]_ ,
    \new_[3659]_ , \new_[3660]_ , \new_[3661]_ , \new_[3662]_ ,
    \new_[3663]_ , \new_[3664]_ , \new_[3665]_ , \new_[3666]_ ,
    \new_[3667]_ , \new_[3668]_ , \new_[3669]_ , \new_[3670]_ ,
    \new_[3671]_ , \new_[3672]_ , \new_[3673]_ , \new_[3674]_ ,
    \new_[3675]_ , \new_[3676]_ , \new_[3677]_ , \new_[3678]_ ,
    \new_[3679]_ , \new_[3680]_ , \new_[3681]_ , \new_[3682]_ ,
    \new_[3683]_ , \new_[3684]_ , \new_[3685]_ , \new_[3686]_ ,
    \new_[3687]_ , \new_[3688]_ , \new_[3689]_ , \new_[3690]_ ,
    \new_[3691]_ , \new_[3692]_ , \new_[3693]_ , \new_[3694]_ ,
    \new_[3695]_ , \new_[3696]_ , \new_[3697]_ , \new_[3698]_ ,
    \new_[3699]_ , \new_[3700]_ , \new_[3701]_ , \new_[3702]_ ,
    \new_[3703]_ , \new_[3704]_ , \new_[3705]_ , \new_[3706]_ ,
    \new_[3707]_ , \new_[3708]_ , \new_[3709]_ , \new_[3710]_ ,
    \new_[3711]_ , \new_[3712]_ , \new_[3713]_ , \new_[3714]_ ,
    \new_[3715]_ , \new_[3716]_ , \new_[3717]_ , \new_[3718]_ ,
    \new_[3719]_ , \new_[3720]_ , \new_[3721]_ , \new_[3722]_ ,
    \new_[3723]_ , \new_[3725]_ , \new_[3726]_ , \new_[3727]_ ,
    \new_[3728]_ , \new_[3729]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3732]_ , \new_[3733]_ , \new_[3734]_ , \new_[3735]_ ,
    \new_[3736]_ , \new_[3737]_ , \new_[3738]_ , \new_[3739]_ ,
    \new_[3740]_ , \new_[3741]_ , \new_[3742]_ , \new_[3743]_ ,
    \new_[3744]_ , \new_[3745]_ , \new_[3746]_ , \new_[3747]_ ,
    \new_[3748]_ , \new_[3749]_ , \new_[3750]_ , \new_[3751]_ ,
    \new_[3752]_ , \new_[3753]_ , \new_[3754]_ , \new_[3755]_ ,
    \new_[3756]_ , \new_[3757]_ , \new_[3758]_ , \new_[3759]_ ,
    \new_[3760]_ , \new_[3761]_ , \new_[3762]_ , \new_[3763]_ ,
    \new_[3764]_ , \new_[3765]_ , \new_[3766]_ , \new_[3767]_ ,
    \new_[3768]_ , \new_[3769]_ , \new_[3770]_ , \new_[3771]_ ,
    \new_[3772]_ , \new_[3773]_ , \new_[3774]_ , \new_[3775]_ ,
    \new_[3776]_ , \new_[3777]_ , \new_[3778]_ , \new_[3779]_ ,
    \new_[3780]_ , \new_[3781]_ , \new_[3782]_ , \new_[3783]_ ,
    \new_[3784]_ , \new_[3785]_ , \new_[3786]_ , \new_[3787]_ ,
    \new_[3788]_ , \new_[3789]_ , \new_[3790]_ , \new_[3791]_ ,
    \new_[3792]_ , \new_[3793]_ , \new_[3794]_ , \new_[3795]_ ,
    \new_[3796]_ , \new_[3797]_ , \new_[3798]_ , \new_[3799]_ ,
    \new_[3800]_ , \new_[3801]_ , \new_[3802]_ , \new_[3803]_ ,
    \new_[3804]_ , \new_[3805]_ , \new_[3806]_ , \new_[3807]_ ,
    \new_[3808]_ , \new_[3809]_ , \new_[3810]_ , \new_[3811]_ ,
    \new_[3812]_ , \new_[3813]_ , \new_[3814]_ , \new_[3815]_ ,
    \new_[3816]_ , \new_[3817]_ , \new_[3818]_ , \new_[3819]_ ,
    \new_[3820]_ , \new_[3821]_ , \new_[3822]_ , \new_[3823]_ ,
    \new_[3824]_ , \new_[3825]_ , \new_[3826]_ , \new_[3827]_ ,
    \new_[3828]_ , \new_[3829]_ , \new_[3830]_ , \new_[3831]_ ,
    \new_[3832]_ , \new_[3833]_ , \new_[3834]_ , \new_[3835]_ ,
    \new_[3836]_ , \new_[3837]_ , \new_[3838]_ , \new_[3839]_ ,
    \new_[3840]_ , \new_[3841]_ , \new_[3842]_ , \new_[3843]_ ,
    \new_[3844]_ , \new_[3845]_ , \new_[3846]_ , \new_[3847]_ ,
    \new_[3848]_ , \new_[3849]_ , \new_[3850]_ , \new_[3851]_ ,
    \new_[3852]_ , \new_[3853]_ , \new_[3854]_ , \new_[3855]_ ,
    \new_[3856]_ , \new_[3857]_ , \new_[3858]_ , \new_[3859]_ ,
    \new_[3860]_ , \new_[3861]_ , \new_[3862]_ , \new_[3863]_ ,
    \new_[3864]_ , \new_[3865]_ , \new_[3866]_ , \new_[3867]_ ,
    \new_[3868]_ , \new_[3869]_ , \new_[3870]_ , \new_[3871]_ ,
    \new_[3872]_ , \new_[3873]_ , \new_[3874]_ , \new_[3875]_ ,
    \new_[3876]_ , \new_[3877]_ , \new_[3878]_ , \new_[3879]_ ,
    \new_[3881]_ , \new_[3882]_ , \new_[3884]_ , \new_[3885]_ ,
    \new_[3886]_ , \new_[3887]_ , \new_[3888]_ , \new_[3889]_ ,
    \new_[3890]_ , \new_[3891]_ , \new_[3892]_ , \new_[3893]_ ,
    \new_[3894]_ , \new_[3895]_ , \new_[3896]_ , \new_[3897]_ ,
    \new_[3898]_ , \new_[3899]_ , \new_[3900]_ , \new_[3901]_ ,
    \new_[3902]_ , \new_[3903]_ , \new_[3904]_ , \new_[3905]_ ,
    \new_[3906]_ , \new_[3907]_ , \new_[3908]_ , \new_[3909]_ ,
    \new_[3910]_ , \new_[3911]_ , \new_[3912]_ , \new_[3913]_ ,
    \new_[3914]_ , \new_[3915]_ , \new_[3916]_ , \new_[3917]_ ,
    \new_[3918]_ , \new_[3919]_ , \new_[3920]_ , \new_[3921]_ ,
    \new_[3922]_ , \new_[3923]_ , \new_[3924]_ , \new_[3925]_ ,
    \new_[3926]_ , \new_[3927]_ , \new_[3928]_ , \new_[3929]_ ,
    \new_[3930]_ , \new_[3931]_ , \new_[3932]_ , \new_[3933]_ ,
    \new_[3934]_ , \new_[3935]_ , \new_[3937]_ , \new_[3938]_ ,
    \new_[3939]_ , \new_[3940]_ , \new_[3941]_ , \new_[3942]_ ,
    \new_[3943]_ , \new_[3944]_ , \new_[3945]_ , \new_[3946]_ ,
    \new_[3947]_ , \new_[3948]_ , \new_[3949]_ , \new_[3950]_ ,
    \new_[3951]_ , \new_[3952]_ , \new_[3953]_ , \new_[3954]_ ,
    \new_[3955]_ , \new_[3956]_ , \new_[3957]_ , \new_[3958]_ ,
    \new_[3959]_ , \new_[3960]_ , \new_[3961]_ , \new_[3962]_ ,
    \new_[3963]_ , \new_[3964]_ , \new_[3965]_ , \new_[3966]_ ,
    \new_[3967]_ , \new_[3968]_ , \new_[3969]_ , \new_[3970]_ ,
    \new_[3971]_ , \new_[3972]_ , \new_[3973]_ , \new_[3974]_ ,
    \new_[3975]_ , \new_[3976]_ , \new_[3977]_ , \new_[3978]_ ,
    \new_[3979]_ , \new_[3980]_ , \new_[3981]_ , \new_[3982]_ ,
    \new_[3983]_ , \new_[3984]_ , \new_[3985]_ , \new_[3986]_ ,
    \new_[3987]_ , \new_[3988]_ , \new_[3989]_ , \new_[3990]_ ,
    \new_[3991]_ , \new_[3992]_ , \new_[3993]_ , \new_[3994]_ ,
    \new_[3995]_ , \new_[3996]_ , \new_[3997]_ , \new_[3998]_ ,
    \new_[3999]_ , \new_[4000]_ , \new_[4001]_ , \new_[4002]_ ,
    \new_[4003]_ , \new_[4004]_ , \new_[4005]_ , \new_[4006]_ ,
    \new_[4007]_ , \new_[4008]_ , \new_[4009]_ , \new_[4010]_ ,
    \new_[4011]_ , \new_[4012]_ , \new_[4013]_ , \new_[4014]_ ,
    \new_[4015]_ , \new_[4016]_ , \new_[4017]_ , \new_[4018]_ ,
    \new_[4019]_ , \new_[4020]_ , \new_[4021]_ , \new_[4022]_ ,
    \new_[4023]_ , \new_[4024]_ , \new_[4025]_ , \new_[4026]_ ,
    \new_[4027]_ , \new_[4028]_ , \new_[4029]_ , \new_[4030]_ ,
    \new_[4031]_ , \new_[4032]_ , \new_[4033]_ , \new_[4034]_ ,
    \new_[4035]_ , \new_[4036]_ , \new_[4037]_ , \new_[4038]_ ,
    \new_[4039]_ , \new_[4040]_ , \new_[4041]_ , \new_[4042]_ ,
    \new_[4043]_ , \new_[4044]_ , \new_[4045]_ , \new_[4046]_ ,
    \new_[4047]_ , \new_[4048]_ , \new_[4049]_ , \new_[4050]_ ,
    \new_[4051]_ , \new_[4052]_ , \new_[4053]_ , \new_[4054]_ ,
    \new_[4055]_ , \new_[4056]_ , \new_[4057]_ , \new_[4058]_ ,
    \new_[4059]_ , \new_[4060]_ , \new_[4061]_ , \new_[4062]_ ,
    \new_[4063]_ , \new_[4064]_ , \new_[4065]_ , \new_[4066]_ ,
    \new_[4067]_ , \new_[4068]_ , \new_[4070]_ , \new_[4078]_ ,
    \new_[4079]_ , \new_[4080]_ , \new_[4081]_ , \new_[4082]_ ,
    \new_[4083]_ , \new_[4084]_ , \new_[4085]_ , \new_[4086]_ ,
    \new_[4087]_ , \new_[4088]_ , \new_[4089]_ , \new_[4090]_ ,
    \new_[4091]_ , \new_[4092]_ , \new_[4093]_ , \new_[4094]_ ,
    \new_[4095]_ , \new_[4096]_ , \new_[4097]_ , \new_[4098]_ ,
    \new_[4099]_ , \new_[4100]_ , \new_[4101]_ , \new_[4102]_ ,
    \new_[4103]_ , \new_[4104]_ , \new_[4105]_ , \new_[4106]_ ,
    \new_[4107]_ , \new_[4108]_ , \new_[4109]_ , \new_[4110]_ ,
    \new_[4111]_ , \new_[4112]_ , \new_[4113]_ , \new_[4114]_ ,
    \new_[4115]_ , \new_[4116]_ , \new_[4117]_ , \new_[4118]_ ,
    \new_[4119]_ , \new_[4120]_ , \new_[4121]_ , \new_[4122]_ ,
    \new_[4123]_ , \new_[4124]_ , \new_[4125]_ , \new_[4126]_ ,
    \new_[4127]_ , \new_[4128]_ , \new_[4129]_ , \new_[4130]_ ,
    \new_[4131]_ , \new_[4132]_ , \new_[4133]_ , \new_[4134]_ ,
    \new_[4135]_ , \new_[4136]_ , \new_[4137]_ , \new_[4138]_ ,
    \new_[4139]_ , \new_[4140]_ , \new_[4141]_ , \new_[4142]_ ,
    \new_[4143]_ , \new_[4144]_ , \new_[4145]_ , \new_[4146]_ ,
    \new_[4147]_ , \new_[4148]_ , \new_[4149]_ , \new_[4150]_ ,
    \new_[4151]_ , \new_[4152]_ , \new_[4153]_ , \new_[4154]_ ,
    \new_[4155]_ , \new_[4156]_ , \new_[4157]_ , \new_[4158]_ ,
    \new_[4159]_ , \new_[4160]_ , \new_[4161]_ , \new_[4162]_ ,
    \new_[4163]_ , \new_[4164]_ , \new_[4165]_ , \new_[4166]_ ,
    \new_[4167]_ , \new_[4168]_ , \new_[4169]_ , \new_[4170]_ ,
    \new_[4171]_ , \new_[4172]_ , \new_[4173]_ , \new_[4174]_ ,
    \new_[4175]_ , \new_[4176]_ , \new_[4177]_ , \new_[4178]_ ,
    \new_[4179]_ , \new_[4180]_ , \new_[4181]_ , \new_[4182]_ ,
    \new_[4183]_ , \new_[4185]_ , \new_[4186]_ , \new_[4187]_ ,
    \new_[4188]_ , \new_[4189]_ , \new_[4190]_ , \new_[4191]_ ,
    \new_[4193]_ , \new_[4194]_ , \new_[4195]_ , \new_[4196]_ ,
    \new_[4197]_ , \new_[4198]_ , \new_[4199]_ , \new_[4200]_ ,
    \new_[4201]_ , \new_[4202]_ , \new_[4203]_ , \new_[4204]_ ,
    \new_[4205]_ , \new_[4206]_ , \new_[4207]_ , \new_[4208]_ ,
    \new_[4209]_ , \new_[4210]_ , \new_[4211]_ , \new_[4212]_ ,
    \new_[4213]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4218]_ , \new_[4219]_ , \new_[4220]_ ,
    \new_[4221]_ , \new_[4222]_ , \new_[4223]_ , \new_[4224]_ ,
    \new_[4225]_ , \new_[4226]_ , \new_[4227]_ , \new_[4228]_ ,
    \new_[4229]_ , \new_[4230]_ , \new_[4231]_ , \new_[4232]_ ,
    \new_[4233]_ , \new_[4234]_ , \new_[4235]_ , \new_[4236]_ ,
    \new_[4237]_ , \new_[4238]_ , \new_[4239]_ , \new_[4240]_ ,
    \new_[4241]_ , \new_[4242]_ , \new_[4243]_ , \new_[4244]_ ,
    \new_[4245]_ , \new_[4248]_ , \new_[4249]_ , \new_[4250]_ ,
    \new_[4251]_ , \new_[4252]_ , \new_[4253]_ , \new_[4254]_ ,
    \new_[4255]_ , \new_[4256]_ , \new_[4257]_ , \new_[4258]_ ,
    \new_[4259]_ , \new_[4260]_ , \new_[4261]_ , \new_[4262]_ ,
    \new_[4263]_ , \new_[4264]_ , \new_[4265]_ , \new_[4266]_ ,
    \new_[4267]_ , \new_[4268]_ , \new_[4269]_ , \new_[4270]_ ,
    \new_[4271]_ , \new_[4272]_ , \new_[4273]_ , \new_[4274]_ ,
    \new_[4275]_ , \new_[4276]_ , \new_[4277]_ , \new_[4278]_ ,
    \new_[4279]_ , \new_[4280]_ , \new_[4281]_ , \new_[4282]_ ,
    \new_[4283]_ , \new_[4284]_ , \new_[4285]_ , \new_[4286]_ ,
    \new_[4287]_ , \new_[4288]_ , \new_[4289]_ , \new_[4290]_ ,
    \new_[4291]_ , \new_[4292]_ , \new_[4293]_ , \new_[4294]_ ,
    \new_[4295]_ , \new_[4296]_ , \new_[4297]_ , \new_[4298]_ ,
    \new_[4299]_ , \new_[4300]_ , \new_[4301]_ , \new_[4302]_ ,
    \new_[4303]_ , \new_[4304]_ , \new_[4305]_ , \new_[4306]_ ,
    \new_[4307]_ , \new_[4308]_ , \new_[4309]_ , \new_[4310]_ ,
    \new_[4311]_ , \new_[4312]_ , \new_[4313]_ , \new_[4314]_ ,
    \new_[4315]_ , \new_[4316]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4319]_ , \new_[4320]_ , \new_[4321]_ , \new_[4322]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4325]_ , \new_[4326]_ ,
    \new_[4327]_ , \new_[4328]_ , \new_[4329]_ , \new_[4330]_ ,
    \new_[4331]_ , \new_[4332]_ , \new_[4333]_ , \new_[4334]_ ,
    \new_[4335]_ , \new_[4336]_ , \new_[4337]_ , \new_[4338]_ ,
    \new_[4339]_ , \new_[4340]_ , \new_[4341]_ , \new_[4342]_ ,
    \new_[4343]_ , \new_[4344]_ , \new_[4345]_ , \new_[4346]_ ,
    \new_[4347]_ , \new_[4348]_ , \new_[4349]_ , \new_[4350]_ ,
    \new_[4351]_ , \new_[4352]_ , \new_[4353]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4356]_ , \new_[4357]_ , \new_[4358]_ ,
    \new_[4359]_ , \new_[4360]_ , \new_[4361]_ , \new_[4362]_ ,
    \new_[4363]_ , \new_[4364]_ , \new_[4365]_ , \new_[4366]_ ,
    \new_[4367]_ , \new_[4368]_ , \new_[4369]_ , \new_[4370]_ ,
    \new_[4371]_ , \new_[4372]_ , \new_[4373]_ , \new_[4374]_ ,
    \new_[4375]_ , \new_[4376]_ , \new_[4377]_ , \new_[4378]_ ,
    \new_[4379]_ , \new_[4380]_ , \new_[4381]_ , \new_[4382]_ ,
    \new_[4383]_ , \new_[4384]_ , \new_[4385]_ , \new_[4386]_ ,
    \new_[4387]_ , \new_[4388]_ , \new_[4389]_ , \new_[4390]_ ,
    \new_[4391]_ , \new_[4392]_ , \new_[4393]_ , \new_[4394]_ ,
    \new_[4395]_ , \new_[4396]_ , \new_[4397]_ , \new_[4398]_ ,
    \new_[4399]_ , \new_[4400]_ , \new_[4401]_ , \new_[4402]_ ,
    \new_[4403]_ , \new_[4404]_ , \new_[4405]_ , \new_[4406]_ ,
    \new_[4407]_ , \new_[4408]_ , \new_[4409]_ , \new_[4410]_ ,
    \new_[4411]_ , \new_[4412]_ , \new_[4413]_ , \new_[4414]_ ,
    \new_[4415]_ , \new_[4416]_ , \new_[4417]_ , \new_[4418]_ ,
    \new_[4419]_ , \new_[4420]_ , \new_[4421]_ , \new_[4422]_ ,
    \new_[4423]_ , \new_[4424]_ , \new_[4425]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4429]_ , \new_[4430]_ ,
    \new_[4431]_ , \new_[4432]_ , \new_[4433]_ , \new_[4434]_ ,
    \new_[4435]_ , \new_[4436]_ , \new_[4437]_ , \new_[4438]_ ,
    \new_[4439]_ , \new_[4440]_ , \new_[4441]_ , \new_[4442]_ ,
    \new_[4443]_ , \new_[4444]_ , \new_[4445]_ , \new_[4446]_ ,
    \new_[4447]_ , \new_[4448]_ , \new_[4449]_ , \new_[4450]_ ,
    \new_[4451]_ , \new_[4452]_ , \new_[4453]_ , \new_[4454]_ ,
    \new_[4455]_ , \new_[4456]_ , \new_[4457]_ , \new_[4458]_ ,
    \new_[4459]_ , \new_[4460]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4463]_ , \new_[4464]_ , \new_[4465]_ , \new_[4466]_ ,
    \new_[4467]_ , \new_[4468]_ , \new_[4469]_ , \new_[4470]_ ,
    \new_[4471]_ , \new_[4473]_ , \new_[4474]_ , \new_[4475]_ ,
    \new_[4476]_ , \new_[4477]_ , \new_[4478]_ , \new_[4479]_ ,
    \new_[4480]_ , \new_[4481]_ , \new_[4482]_ , \new_[4483]_ ,
    \new_[4484]_ , \new_[4485]_ , \new_[4486]_ , \new_[4487]_ ,
    \new_[4488]_ , \new_[4489]_ , \new_[4490]_ , \new_[4491]_ ,
    \new_[4492]_ , \new_[4493]_ , \new_[4494]_ , \new_[4495]_ ,
    \new_[4504]_ , \new_[4505]_ , \new_[4506]_ , \new_[4507]_ ,
    \new_[4508]_ , \new_[4509]_ , \new_[4510]_ , \new_[4511]_ ,
    \new_[4512]_ , \new_[4513]_ , \new_[4514]_ , \new_[4515]_ ,
    \new_[4516]_ , \new_[4517]_ , \new_[4518]_ , \new_[4519]_ ,
    \new_[4520]_ , \new_[4521]_ , \new_[4522]_ , \new_[4523]_ ,
    \new_[4524]_ , \new_[4525]_ , \new_[4526]_ , \new_[4527]_ ,
    \new_[4528]_ , \new_[4529]_ , \new_[4530]_ , \new_[4531]_ ,
    \new_[4532]_ , \new_[4533]_ , \new_[4534]_ , \new_[4535]_ ,
    \new_[4536]_ , \new_[4537]_ , \new_[4538]_ , \new_[4539]_ ,
    \new_[4540]_ , \new_[4541]_ , \new_[4542]_ , \new_[4543]_ ,
    \new_[4544]_ , \new_[4545]_ , \new_[4547]_ , \new_[4549]_ ,
    \new_[4551]_ , \new_[4553]_ , \new_[4555]_ , \new_[4556]_ ,
    \new_[4557]_ , \new_[4559]_ , \new_[4560]_ , \new_[4561]_ ,
    \new_[4562]_ , \new_[4563]_ , \new_[4564]_ , \new_[4565]_ ,
    \new_[4566]_ , \new_[4567]_ , \new_[4568]_ , \new_[4569]_ ,
    \new_[4570]_ , \new_[4571]_ , \new_[4572]_ , \new_[4573]_ ,
    \new_[4574]_ , \new_[4575]_ , \new_[4576]_ , \new_[4577]_ ,
    \new_[4578]_ , \new_[4579]_ , \new_[4580]_ , \new_[4581]_ ,
    \new_[4582]_ , \new_[4583]_ , \new_[4584]_ , \new_[4585]_ ,
    \new_[4586]_ , \new_[4587]_ , \new_[4588]_ , \new_[4589]_ ,
    \new_[4590]_ , \new_[4591]_ , \new_[4592]_ , \new_[4593]_ ,
    \new_[4594]_ , \new_[4595]_ , \new_[4596]_ , \new_[4597]_ ,
    \new_[4598]_ , \new_[4599]_ , \new_[4600]_ , \new_[4601]_ ,
    \new_[4602]_ , \new_[4603]_ , \new_[4604]_ , \new_[4605]_ ,
    \new_[4606]_ , \new_[4607]_ , \new_[4608]_ , \new_[4609]_ ,
    \new_[4610]_ , \new_[4611]_ , \new_[4612]_ , \new_[4613]_ ,
    \new_[4614]_ , \new_[4615]_ , \new_[4616]_ , \new_[4617]_ ,
    \new_[4618]_ , \new_[4619]_ , \new_[4620]_ , \new_[4621]_ ,
    \new_[4622]_ , \new_[4623]_ , \new_[4624]_ , \new_[4625]_ ,
    \new_[4626]_ , \new_[4627]_ , \new_[4628]_ , \new_[4629]_ ,
    \new_[4630]_ , \new_[4631]_ , \new_[4632]_ , \new_[4633]_ ,
    \new_[4634]_ , \new_[4635]_ , \new_[4636]_ , \new_[4637]_ ,
    \new_[4638]_ , \new_[4639]_ , \new_[4640]_ , \new_[4641]_ ,
    \new_[4642]_ , \new_[4643]_ , \new_[4644]_ , \new_[4645]_ ,
    \new_[4646]_ , \new_[4647]_ , \new_[4648]_ , \new_[4649]_ ,
    \new_[4650]_ , \new_[4651]_ , \new_[4652]_ , \new_[4653]_ ,
    \new_[4654]_ , \new_[4655]_ , \new_[4656]_ , \new_[4657]_ ,
    \new_[4658]_ , \new_[4659]_ , \new_[4660]_ , \new_[4661]_ ,
    \new_[4662]_ , \new_[4663]_ , \new_[4664]_ , \new_[4665]_ ,
    \new_[4666]_ , \new_[4667]_ , \new_[4668]_ , \new_[4669]_ ,
    \new_[4670]_ , \new_[4671]_ , \new_[4672]_ , \new_[4673]_ ,
    \new_[4674]_ , \new_[4675]_ , \new_[4676]_ , \new_[4677]_ ,
    \new_[4678]_ , \new_[4679]_ , \new_[4680]_ , \new_[4681]_ ,
    \new_[4682]_ , \new_[4683]_ , \new_[4684]_ , \new_[4685]_ ,
    \new_[4686]_ , \new_[4687]_ , \new_[4688]_ , \new_[4689]_ ,
    \new_[4691]_ , \new_[4692]_ , \new_[4700]_ , \new_[4701]_ ,
    \new_[4702]_ , \new_[4703]_ , \new_[4704]_ , \new_[4705]_ ,
    \new_[4706]_ , \new_[4707]_ , \new_[4708]_ , \new_[4709]_ ,
    \new_[4710]_ , \new_[4711]_ , \new_[4712]_ , \new_[4713]_ ,
    \new_[4714]_ , \new_[4715]_ , \new_[4716]_ , \new_[4717]_ ,
    \new_[4718]_ , \new_[4719]_ , \new_[4720]_ , \new_[4721]_ ,
    \new_[4722]_ , \new_[4723]_ , \new_[4724]_ , \new_[4725]_ ,
    \new_[4726]_ , \new_[4727]_ , \new_[4728]_ , \new_[4729]_ ,
    \new_[4730]_ , \new_[4731]_ , \new_[4732]_ , \new_[4733]_ ,
    \new_[4734]_ , \new_[4735]_ , \new_[4736]_ , \new_[4737]_ ,
    \new_[4738]_ , \new_[4739]_ , \new_[4740]_ , \new_[4741]_ ,
    \new_[4742]_ , \new_[4743]_ , \new_[4744]_ , \new_[4745]_ ,
    \new_[4746]_ , \new_[4747]_ , \new_[4748]_ , \new_[4749]_ ,
    \new_[4750]_ , \new_[4751]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4757]_ ,
    \new_[4758]_ , \new_[4759]_ , \new_[4760]_ , \new_[4761]_ ,
    \new_[4762]_ , \new_[4763]_ , \new_[4764]_ , \new_[4765]_ ,
    \new_[4766]_ , \new_[4767]_ , \new_[4768]_ , \new_[4769]_ ,
    \new_[4770]_ , \new_[4771]_ , \new_[4772]_ , \new_[4773]_ ,
    \new_[4774]_ , \new_[4775]_ , \new_[4776]_ , \new_[4777]_ ,
    \new_[4778]_ , \new_[4779]_ , \new_[4780]_ , \new_[4781]_ ,
    \new_[4782]_ , \new_[4783]_ , \new_[4784]_ , \new_[4785]_ ,
    \new_[4786]_ , \new_[4787]_ , \new_[4788]_ , \new_[4789]_ ,
    \new_[4790]_ , \new_[4791]_ , \new_[4792]_ , \new_[4793]_ ,
    \new_[4794]_ , \new_[4795]_ , \new_[4796]_ , \new_[4797]_ ,
    \new_[4798]_ , \new_[4799]_ , \new_[4800]_ , \new_[4801]_ ,
    \new_[4802]_ , \new_[4803]_ , \new_[4804]_ , \new_[4805]_ ,
    \new_[4806]_ , \new_[4807]_ , \new_[4808]_ , \new_[4809]_ ,
    \new_[4810]_ , \new_[4811]_ , \new_[4812]_ , \new_[4813]_ ,
    \new_[4814]_ , \new_[4815]_ , \new_[4816]_ , \new_[4817]_ ,
    \new_[4818]_ , \new_[4819]_ , \new_[4820]_ , \new_[4821]_ ,
    \new_[4822]_ , \new_[4823]_ , \new_[4824]_ , \new_[4825]_ ,
    \new_[4826]_ , \new_[4827]_ , \new_[4828]_ , \new_[4829]_ ,
    \new_[4830]_ , \new_[4831]_ , \new_[4832]_ , \new_[4833]_ ,
    \new_[4834]_ , \new_[4835]_ , \new_[4836]_ , \new_[4837]_ ,
    \new_[4838]_ , \new_[4839]_ , \new_[4840]_ , \new_[4841]_ ,
    \new_[4842]_ , \new_[4843]_ , \new_[4844]_ , \new_[4845]_ ,
    \new_[4846]_ , \new_[4847]_ , \new_[4848]_ , \new_[4849]_ ,
    \new_[4850]_ , \new_[4851]_ , \new_[4852]_ , \new_[4853]_ ,
    \new_[4854]_ , \new_[4855]_ , \new_[4856]_ , \new_[4857]_ ,
    \new_[4858]_ , \new_[4859]_ , \new_[4860]_ , \new_[4861]_ ,
    \new_[4862]_ , \new_[4863]_ , \new_[4864]_ , \new_[4865]_ ,
    \new_[4866]_ , \new_[4867]_ , \new_[4868]_ , \new_[4869]_ ,
    \new_[4870]_ , \new_[4871]_ , \new_[4872]_ , \new_[4873]_ ,
    \new_[4874]_ , \new_[4875]_ , \new_[4876]_ , \new_[4877]_ ,
    \new_[4878]_ , \new_[4879]_ , \new_[4880]_ , \new_[4881]_ ,
    \new_[4882]_ , \new_[4883]_ , \new_[4884]_ , \new_[4885]_ ,
    \new_[4886]_ , \new_[4887]_ , \new_[4888]_ , \new_[4889]_ ,
    \new_[4890]_ , \new_[4891]_ , \new_[4892]_ , \new_[4893]_ ,
    \new_[4894]_ , \new_[4895]_ , \new_[4896]_ , \new_[4897]_ ,
    \new_[4898]_ , \new_[4899]_ , \new_[4900]_ , \new_[4901]_ ,
    \new_[4902]_ , \new_[4903]_ , \new_[4904]_ , \new_[4905]_ ,
    \new_[4906]_ , \new_[4907]_ , \new_[4908]_ , \new_[4909]_ ,
    \new_[4910]_ , \new_[4911]_ , \new_[4912]_ , \new_[4913]_ ,
    \new_[4914]_ , \new_[4915]_ , \new_[4916]_ , \new_[4917]_ ,
    \new_[4918]_ , \new_[4919]_ , \new_[4920]_ , \new_[4921]_ ,
    \new_[4922]_ , \new_[4923]_ , \new_[4924]_ , \new_[4925]_ ,
    \new_[4926]_ , \new_[4927]_ , \new_[4928]_ , \new_[4929]_ ,
    \new_[4930]_ , \new_[4931]_ , \new_[4932]_ , \new_[4933]_ ,
    \new_[4934]_ , \new_[4935]_ , \new_[4936]_ , \new_[4937]_ ,
    \new_[4938]_ , \new_[4939]_ , \new_[4940]_ , \new_[4941]_ ,
    \new_[4942]_ , \new_[4943]_ , \new_[4944]_ , \new_[4945]_ ,
    \new_[4946]_ , \new_[4947]_ , \new_[4948]_ , \new_[4949]_ ,
    \new_[4950]_ , \new_[4951]_ , \new_[4952]_ , \new_[4953]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4956]_ , \new_[4957]_ ,
    \new_[4958]_ , \new_[4959]_ , \new_[4960]_ , \new_[4962]_ ,
    \new_[4963]_ , \new_[4964]_ , \new_[4965]_ , \new_[4966]_ ,
    \new_[4967]_ , \new_[4968]_ , \new_[4970]_ , \new_[4971]_ ,
    \new_[4972]_ , \new_[4973]_ , \new_[4974]_ , \new_[4975]_ ,
    \new_[4976]_ , \new_[4977]_ , \new_[4978]_ , \new_[4979]_ ,
    \new_[4981]_ , \new_[4982]_ , \new_[4983]_ , \new_[4984]_ ,
    \new_[4985]_ , \new_[4988]_ , \new_[4989]_ , \new_[4990]_ ,
    \new_[4991]_ , \new_[4992]_ , \new_[4993]_ , \new_[4994]_ ,
    \new_[4995]_ , \new_[4996]_ , \new_[4997]_ , \new_[4998]_ ,
    \new_[4999]_ , \new_[5000]_ , \new_[5001]_ , \new_[5002]_ ,
    \new_[5003]_ , \new_[5004]_ , \new_[5005]_ , \new_[5006]_ ,
    \new_[5007]_ , \new_[5008]_ , \new_[5009]_ , \new_[5010]_ ,
    \new_[5011]_ , \new_[5012]_ , \new_[5013]_ , \new_[5014]_ ,
    \new_[5015]_ , \new_[5016]_ , \new_[5017]_ , \new_[5018]_ ,
    \new_[5019]_ , \new_[5020]_ , \new_[5021]_ , \new_[5022]_ ,
    \new_[5023]_ , \new_[5024]_ , \new_[5025]_ , \new_[5026]_ ,
    \new_[5027]_ , \new_[5028]_ , \new_[5029]_ , \new_[5030]_ ,
    \new_[5031]_ , \new_[5032]_ , \new_[5033]_ , \new_[5034]_ ,
    \new_[5035]_ , \new_[5036]_ , \new_[5037]_ , \new_[5038]_ ,
    \new_[5039]_ , \new_[5040]_ , \new_[5041]_ , \new_[5042]_ ,
    \new_[5043]_ , \new_[5044]_ , \new_[5045]_ , \new_[5046]_ ,
    \new_[5047]_ , \new_[5048]_ , \new_[5049]_ , \new_[5050]_ ,
    \new_[5051]_ , \new_[5052]_ , \new_[5053]_ , \new_[5054]_ ,
    \new_[5055]_ , \new_[5056]_ , \new_[5057]_ , \new_[5058]_ ,
    \new_[5059]_ , \new_[5060]_ , \new_[5061]_ , \new_[5062]_ ,
    \new_[5063]_ , \new_[5064]_ , \new_[5065]_ , \new_[5066]_ ,
    \new_[5067]_ , \new_[5068]_ , \new_[5069]_ , \new_[5070]_ ,
    \new_[5071]_ , \new_[5072]_ , \new_[5073]_ , \new_[5074]_ ,
    \new_[5075]_ , \new_[5076]_ , \new_[5077]_ , \new_[5078]_ ,
    \new_[5079]_ , \new_[5080]_ , \new_[5081]_ , \new_[5082]_ ,
    \new_[5083]_ , \new_[5084]_ , \new_[5085]_ , \new_[5086]_ ,
    \new_[5087]_ , \new_[5088]_ , \new_[5093]_ , \new_[5096]_ ,
    \new_[5119]_ , \new_[5121]_ , \new_[5124]_ , \new_[5181]_ ,
    \new_[5239]_ , \new_[5240]_ , \new_[5241]_ , \new_[5242]_ ,
    \new_[5243]_ , \new_[5244]_ , \new_[5245]_ , \new_[5246]_ ,
    \new_[5247]_ , \new_[5248]_ , \new_[5249]_ , \new_[5250]_ ,
    \new_[5251]_ , \new_[5252]_ , \new_[5253]_ , \new_[5254]_ ,
    \new_[5255]_ , \new_[5256]_ , \new_[5257]_ , \new_[5258]_ ,
    \new_[5259]_ , \new_[5260]_ , \new_[5261]_ , \new_[5262]_ ,
    \new_[5263]_ , \new_[5264]_ , \new_[5265]_ , \new_[5266]_ ,
    \new_[5267]_ , \new_[5268]_ , \new_[5269]_ , \new_[5270]_ ,
    \new_[5271]_ , \new_[5272]_ , \new_[5273]_ , \new_[5274]_ ,
    \new_[5275]_ , \new_[5276]_ , \new_[5277]_ , \new_[5278]_ ,
    \new_[5279]_ , \new_[5280]_ , \new_[5281]_ , \new_[5282]_ ,
    \new_[5283]_ , \new_[5284]_ , \new_[5285]_ , \new_[5286]_ ,
    \new_[5287]_ , \new_[5288]_ , \new_[5289]_ , \new_[5290]_ ,
    \new_[5291]_ , \new_[5292]_ , \new_[5293]_ , \new_[5294]_ ,
    \new_[5295]_ , \new_[5296]_ , \new_[5297]_ , \new_[5298]_ ,
    \new_[5299]_ , \new_[5301]_ , \new_[5302]_ , \new_[5303]_ ,
    \new_[5304]_ , \new_[5305]_ , \new_[5306]_ , \new_[5307]_ ,
    \new_[5308]_ , \new_[5309]_ , \new_[5310]_ , \new_[5311]_ ,
    \new_[5312]_ , \new_[5313]_ , \new_[5314]_ , \new_[5315]_ ,
    \new_[5316]_ , \new_[5317]_ , \new_[5318]_ , \new_[5319]_ ,
    \new_[5320]_ , \new_[5321]_ , \new_[5322]_ , \new_[5323]_ ,
    \new_[5324]_ , \new_[5325]_ , \new_[5326]_ , \new_[5327]_ ,
    \new_[5328]_ , \new_[5329]_ , \new_[5330]_ , \new_[5331]_ ,
    \new_[5332]_ , \new_[5333]_ , \new_[5334]_ , \new_[5335]_ ,
    \new_[5336]_ , \new_[5337]_ , \new_[5338]_ , \new_[5339]_ ,
    \new_[5340]_ , \new_[5341]_ , \new_[5342]_ , \new_[5343]_ ,
    \new_[5344]_ , \new_[5345]_ , \new_[5346]_ , \new_[5347]_ ,
    \new_[5348]_ , \new_[5349]_ , \new_[5350]_ , \new_[5351]_ ,
    \new_[5352]_ , \new_[5353]_ , \new_[5354]_ , \new_[5355]_ ,
    \new_[5356]_ , \new_[5357]_ , \new_[5358]_ , \new_[5359]_ ,
    \new_[5360]_ , \new_[5361]_ , \new_[5362]_ , \new_[5363]_ ,
    \new_[5365]_ , \new_[5366]_ , \new_[5367]_ , \new_[5368]_ ,
    \new_[5369]_ , \new_[5370]_ , \new_[5371]_ , \new_[5372]_ ,
    \new_[5373]_ , \new_[5374]_ , \new_[5375]_ , \new_[5376]_ ,
    \new_[5377]_ , \new_[5378]_ , \new_[5379]_ , \new_[5380]_ ,
    \new_[5381]_ , \new_[5382]_ , \new_[5383]_ , \new_[5384]_ ,
    \new_[5385]_ , \new_[5386]_ , \new_[5387]_ , \new_[5388]_ ,
    \new_[5389]_ , \new_[5390]_ , \new_[5391]_ , \new_[5392]_ ,
    \new_[5393]_ , \new_[5394]_ , \new_[5395]_ , \new_[5396]_ ,
    \new_[5397]_ , \new_[5398]_ , \new_[5399]_ , \new_[5400]_ ,
    \new_[5401]_ , \new_[5402]_ , \new_[5403]_ , \new_[5404]_ ,
    \new_[5405]_ , \new_[5406]_ , \new_[5407]_ , \new_[5408]_ ,
    \new_[5409]_ , \new_[5410]_ , \new_[5411]_ , \new_[5412]_ ,
    \new_[5413]_ , \new_[5414]_ , \new_[5415]_ , \new_[5416]_ ,
    \new_[5417]_ , \new_[5418]_ , \new_[5419]_ , \new_[5420]_ ,
    \new_[5430]_ , \new_[5431]_ , \new_[5432]_ , \new_[5433]_ ,
    \new_[5434]_ , \new_[5435]_ , \new_[5436]_ , \new_[5437]_ ,
    \new_[5438]_ , \new_[5439]_ , \new_[5440]_ , \new_[5441]_ ,
    \new_[5442]_ , \new_[5443]_ , \new_[5444]_ , \new_[5445]_ ,
    \new_[5446]_ , \new_[5447]_ , \new_[5448]_ , \new_[5449]_ ,
    \new_[5450]_ , \new_[5451]_ , \new_[5452]_ , \new_[5453]_ ,
    \new_[5454]_ , \new_[5455]_ , \new_[5456]_ , \new_[5457]_ ,
    \new_[5458]_ , \new_[5459]_ , \new_[5460]_ , \new_[5461]_ ,
    \new_[5462]_ , \new_[5463]_ , \new_[5464]_ , \new_[5465]_ ,
    \new_[5466]_ , \new_[5467]_ , \new_[5468]_ , \new_[5469]_ ,
    \new_[5470]_ , \new_[5471]_ , \new_[5472]_ , \new_[5473]_ ,
    \new_[5474]_ , \new_[5475]_ , \new_[5476]_ , \new_[5477]_ ,
    \new_[5478]_ , \new_[5479]_ , \new_[5480]_ , \new_[5481]_ ,
    \new_[5482]_ , \new_[5483]_ , \new_[5484]_ , \new_[5485]_ ,
    \new_[5486]_ , \new_[5487]_ , \new_[5488]_ , \new_[5489]_ ,
    \new_[5490]_ , \new_[5491]_ , \new_[5492]_ , \new_[5493]_ ,
    \new_[5494]_ , \new_[5495]_ , \new_[5496]_ , \new_[5497]_ ,
    \new_[5498]_ , \new_[5499]_ , \new_[5500]_ , \new_[5501]_ ,
    \new_[5502]_ , \new_[5503]_ , \new_[5504]_ , \new_[5505]_ ,
    \new_[5506]_ , \new_[5507]_ , \new_[5508]_ , \new_[5509]_ ,
    \new_[5510]_ , \new_[5511]_ , \new_[5512]_ , \new_[5513]_ ,
    \new_[5514]_ , \new_[5515]_ , \new_[5516]_ , \new_[5517]_ ,
    \new_[5518]_ , \new_[5519]_ , \new_[5520]_ , \new_[5521]_ ,
    \new_[5522]_ , \new_[5523]_ , \new_[5524]_ , \new_[5525]_ ,
    \new_[5526]_ , \new_[5527]_ , \new_[5528]_ , \new_[5529]_ ,
    \new_[5530]_ , \new_[5531]_ , \new_[5532]_ , \new_[5533]_ ,
    \new_[5534]_ , \new_[5535]_ , \new_[5536]_ , \new_[5537]_ ,
    \new_[5538]_ , \new_[5539]_ , \new_[5540]_ , \new_[5541]_ ,
    \new_[5542]_ , \new_[5543]_ , \new_[5544]_ , \new_[5545]_ ,
    \new_[5546]_ , \new_[5547]_ , \new_[5548]_ , \new_[5549]_ ,
    \new_[5550]_ , \new_[5551]_ , \new_[5552]_ , \new_[5553]_ ,
    \new_[5554]_ , \new_[5555]_ , \new_[5556]_ , \new_[5557]_ ,
    \new_[5558]_ , \new_[5559]_ , \new_[5560]_ , \new_[5561]_ ,
    \new_[5562]_ , \new_[5563]_ , \new_[5564]_ , \new_[5565]_ ,
    \new_[5566]_ , \new_[5567]_ , \new_[5568]_ , \new_[5569]_ ,
    \new_[5570]_ , \new_[5571]_ , \new_[5572]_ , \new_[5573]_ ,
    \new_[5574]_ , \new_[5575]_ , \new_[5576]_ , \new_[5577]_ ,
    \new_[5578]_ , \new_[5579]_ , \new_[5580]_ , \new_[5581]_ ,
    \new_[5582]_ , \new_[5583]_ , \new_[5584]_ , \new_[5585]_ ,
    \new_[5586]_ , \new_[5587]_ , \new_[5588]_ , \new_[5589]_ ,
    \new_[5590]_ , \new_[5591]_ , \new_[5592]_ , \new_[5593]_ ,
    \new_[5594]_ , \new_[5595]_ , \new_[5596]_ , \new_[5597]_ ,
    \new_[5598]_ , \new_[5599]_ , \new_[5600]_ , \new_[5601]_ ,
    \new_[5602]_ , \new_[5603]_ , \new_[5604]_ , \new_[5605]_ ,
    \new_[5606]_ , \new_[5607]_ , \new_[5608]_ , \new_[5609]_ ,
    \new_[5610]_ , \new_[5611]_ , \new_[5612]_ , \new_[5613]_ ,
    \new_[5614]_ , \new_[5615]_ , \new_[5616]_ , \new_[5617]_ ,
    \new_[5618]_ , \new_[5619]_ , \new_[5620]_ , \new_[5621]_ ,
    \new_[5622]_ , \new_[5623]_ , \new_[5624]_ , \new_[5625]_ ,
    \new_[5626]_ , \new_[5627]_ , \new_[5628]_ , \new_[5629]_ ,
    \new_[5630]_ , \new_[5631]_ , \new_[5632]_ , \new_[5633]_ ,
    \new_[5634]_ , \new_[5635]_ , \new_[5637]_ , \new_[5638]_ ,
    \new_[5639]_ , \new_[5640]_ , \new_[5641]_ , \new_[5642]_ ,
    \new_[5643]_ , \new_[5644]_ , \new_[5645]_ , \new_[5646]_ ,
    \new_[5647]_ , \new_[5648]_ , \new_[5649]_ , \new_[5650]_ ,
    \new_[5651]_ , \new_[5652]_ , \new_[5653]_ , \new_[5654]_ ,
    \new_[5655]_ , \new_[5656]_ , \new_[5657]_ , \new_[5658]_ ,
    \new_[5659]_ , \new_[5660]_ , \new_[5661]_ , \new_[5662]_ ,
    \new_[5663]_ , \new_[5664]_ , \new_[5665]_ , \new_[5666]_ ,
    \new_[5667]_ , \new_[5668]_ , \new_[5669]_ , \new_[5670]_ ,
    \new_[5671]_ , \new_[5672]_ , \new_[5673]_ , \new_[5674]_ ,
    \new_[5675]_ , \new_[5676]_ , \new_[5677]_ , \new_[5678]_ ,
    \new_[5679]_ , \new_[5680]_ , \new_[5681]_ , \new_[5682]_ ,
    \new_[5683]_ , \new_[5684]_ , \new_[5685]_ , \new_[5686]_ ,
    \new_[5687]_ , \new_[5688]_ , \new_[5689]_ , \new_[5690]_ ,
    \new_[5691]_ , \new_[5692]_ , \new_[5693]_ , \new_[5694]_ ,
    \new_[5695]_ , \new_[5696]_ , \new_[5697]_ , \new_[5698]_ ,
    \new_[5699]_ , \new_[5700]_ , \new_[5701]_ , \new_[5702]_ ,
    \new_[5703]_ , \new_[5704]_ , \new_[5705]_ , \new_[5706]_ ,
    \new_[5707]_ , \new_[5708]_ , \new_[5709]_ , \new_[5710]_ ,
    \new_[5711]_ , \new_[5712]_ , \new_[5713]_ , \new_[5714]_ ,
    \new_[5715]_ , \new_[5716]_ , \new_[5717]_ , \new_[5718]_ ,
    \new_[5719]_ , \new_[5720]_ , \new_[5721]_ , \new_[5722]_ ,
    \new_[5723]_ , \new_[5724]_ , \new_[5725]_ , \new_[5726]_ ,
    \new_[5727]_ , \new_[5728]_ , \new_[5729]_ , \new_[5730]_ ,
    \new_[5731]_ , \new_[5732]_ , \new_[5733]_ , \new_[5734]_ ,
    \new_[5735]_ , \new_[5736]_ , \new_[5737]_ , \new_[5738]_ ,
    \new_[5739]_ , \new_[5740]_ , \new_[5741]_ , \new_[5742]_ ,
    \new_[5743]_ , \new_[5744]_ , \new_[5745]_ , \new_[5746]_ ,
    \new_[5747]_ , \new_[5748]_ , \new_[5749]_ , \new_[5750]_ ,
    \new_[5751]_ , \new_[5752]_ , \new_[5753]_ , \new_[5754]_ ,
    \new_[5755]_ , \new_[5756]_ , \new_[5757]_ , \new_[5758]_ ,
    \new_[5759]_ , \new_[5760]_ , \new_[5761]_ , \new_[5762]_ ,
    \new_[5763]_ , \new_[5764]_ , \new_[5765]_ , \new_[5766]_ ,
    \new_[5767]_ , \new_[5768]_ , \new_[5769]_ , \new_[5770]_ ,
    \new_[5771]_ , \new_[5772]_ , \new_[5773]_ , \new_[5774]_ ,
    \new_[5775]_ , \new_[5776]_ , \new_[5777]_ , \new_[5778]_ ,
    \new_[5779]_ , \new_[5780]_ , \new_[5781]_ , \new_[5782]_ ,
    \new_[5783]_ , \new_[5784]_ , \new_[5785]_ , \new_[5786]_ ,
    \new_[5787]_ , \new_[5788]_ , \new_[5789]_ , \new_[5790]_ ,
    \new_[5791]_ , \new_[5792]_ , \new_[5793]_ , \new_[5794]_ ,
    \new_[5795]_ , \new_[5796]_ , \new_[5797]_ , \new_[5798]_ ,
    \new_[5799]_ , \new_[5800]_ , \new_[5801]_ , \new_[5802]_ ,
    \new_[5803]_ , \new_[5804]_ , \new_[5806]_ , \new_[5807]_ ,
    \new_[5808]_ , \new_[5809]_ , \new_[5810]_ , \new_[5811]_ ,
    \new_[5812]_ , \new_[5813]_ , \new_[5814]_ , \new_[5815]_ ,
    \new_[5816]_ , \new_[5817]_ , \new_[5818]_ , \new_[5819]_ ,
    \new_[5820]_ , \new_[5821]_ , \new_[5822]_ , \new_[5823]_ ,
    \new_[5824]_ , \new_[5825]_ , \new_[5826]_ , \new_[5827]_ ,
    \new_[5828]_ , \new_[5829]_ , \new_[5830]_ , \new_[5831]_ ,
    \new_[5832]_ , \new_[5833]_ , \new_[5834]_ , \new_[5835]_ ,
    \new_[5836]_ , \new_[5837]_ , \new_[5838]_ , \new_[5839]_ ,
    \new_[5840]_ , \new_[5841]_ , \new_[5842]_ , \new_[5843]_ ,
    \new_[5844]_ , \new_[5845]_ , \new_[5846]_ , \new_[5847]_ ,
    \new_[5848]_ , \new_[5849]_ , \new_[5850]_ , \new_[5851]_ ,
    \new_[5852]_ , \new_[5853]_ , \new_[5854]_ , \new_[5855]_ ,
    \new_[5856]_ , \new_[5857]_ , \new_[5858]_ , \new_[5859]_ ,
    \new_[5860]_ , \new_[5861]_ , \new_[5862]_ , \new_[5863]_ ,
    \new_[5864]_ , \new_[5865]_ , \new_[5866]_ , \new_[5867]_ ,
    \new_[5868]_ , \new_[5869]_ , \new_[5870]_ , \new_[5871]_ ,
    \new_[5872]_ , \new_[5873]_ , \new_[5874]_ , \new_[5875]_ ,
    \new_[5876]_ , \new_[5877]_ , \new_[5878]_ , \new_[5879]_ ,
    \new_[5880]_ , \new_[5881]_ , \new_[5882]_ , \new_[5883]_ ,
    \new_[5884]_ , \new_[5885]_ , \new_[5886]_ , \new_[5887]_ ,
    \new_[5888]_ , \new_[5889]_ , \new_[5890]_ , \new_[5891]_ ,
    \new_[5892]_ , \new_[5893]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5896]_ , \new_[5897]_ , \new_[5898]_ , \new_[5899]_ ,
    \new_[5900]_ , \new_[5901]_ , \new_[5902]_ , \new_[5903]_ ,
    \new_[5904]_ , \new_[5905]_ , \new_[5906]_ , \new_[5907]_ ,
    \new_[5908]_ , \new_[5909]_ , \new_[5910]_ , \new_[5911]_ ,
    \new_[5912]_ , \new_[5913]_ , \new_[5914]_ , \new_[5915]_ ,
    \new_[5916]_ , \new_[5917]_ , \new_[5918]_ , \new_[5919]_ ,
    \new_[5920]_ , \new_[5921]_ , \new_[5922]_ , \new_[5923]_ ,
    \new_[5924]_ , \new_[5925]_ , \new_[5926]_ , \new_[5927]_ ,
    \new_[5928]_ , \new_[5929]_ , \new_[5930]_ , \new_[5931]_ ,
    \new_[5932]_ , \new_[5933]_ , \new_[5934]_ , \new_[5935]_ ,
    \new_[5936]_ , \new_[5937]_ , \new_[5938]_ , \new_[5939]_ ,
    \new_[5940]_ , \new_[5941]_ , \new_[5942]_ , \new_[5943]_ ,
    \new_[5944]_ , \new_[5945]_ , \new_[5946]_ , \new_[5947]_ ,
    \new_[5948]_ , \new_[5949]_ , \new_[5950]_ , \new_[5951]_ ,
    \new_[5952]_ , \new_[5953]_ , \new_[5954]_ , \new_[5955]_ ,
    \new_[5956]_ , \new_[5957]_ , \new_[5958]_ , \new_[5959]_ ,
    \new_[5960]_ , \new_[5961]_ , \new_[5962]_ , \new_[5963]_ ,
    \new_[5964]_ , \new_[5965]_ , \new_[5966]_ , \new_[5967]_ ,
    \new_[5968]_ , \new_[5969]_ , \new_[5970]_ , \new_[5971]_ ,
    \new_[5972]_ , \new_[5973]_ , \new_[5974]_ , \new_[5975]_ ,
    \new_[5976]_ , \new_[5977]_ , \new_[5978]_ , \new_[5979]_ ,
    \new_[5980]_ , \new_[5981]_ , \new_[5982]_ , \new_[5983]_ ,
    \new_[5984]_ , \new_[5985]_ , \new_[5986]_ , \new_[5987]_ ,
    \new_[5988]_ , \new_[5989]_ , \new_[5990]_ , \new_[5991]_ ,
    \new_[5992]_ , \new_[5993]_ , \new_[5994]_ , \new_[5995]_ ,
    \new_[5996]_ , \new_[5997]_ , \new_[5998]_ , \new_[5999]_ ,
    \new_[6000]_ , \new_[6001]_ , \new_[6002]_ , \new_[6003]_ ,
    \new_[6004]_ , \new_[6005]_ , \new_[6006]_ , \new_[6007]_ ,
    \new_[6008]_ , \new_[6009]_ , \new_[6010]_ , \new_[6011]_ ,
    \new_[6012]_ , \new_[6013]_ , \new_[6014]_ , \new_[6015]_ ,
    \new_[6016]_ , \new_[6017]_ , \new_[6018]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6021]_ , \new_[6022]_ , \new_[6023]_ ,
    \new_[6024]_ , \new_[6025]_ , \new_[6026]_ , \new_[6027]_ ,
    \new_[6029]_ , \new_[6030]_ , \new_[6031]_ , \new_[6032]_ ,
    \new_[6033]_ , \new_[6034]_ , \new_[6035]_ , \new_[6036]_ ,
    \new_[6037]_ , \new_[6038]_ , \new_[6039]_ , \new_[6040]_ ,
    \new_[6041]_ , \new_[6042]_ , \new_[6043]_ , \new_[6044]_ ,
    \new_[6045]_ , \new_[6046]_ , \new_[6047]_ , \new_[6048]_ ,
    \new_[6049]_ , \new_[6050]_ , \new_[6051]_ , \new_[6052]_ ,
    \new_[6053]_ , \new_[6054]_ , \new_[6055]_ , \new_[6056]_ ,
    \new_[6057]_ , \new_[6058]_ , \new_[6059]_ , \new_[6060]_ ,
    \new_[6062]_ , \new_[6063]_ , \new_[6064]_ , \new_[6065]_ ,
    \new_[6066]_ , \new_[6067]_ , \new_[6068]_ , \new_[6069]_ ,
    \new_[6070]_ , \new_[6071]_ , \new_[6072]_ , \new_[6073]_ ,
    \new_[6074]_ , \new_[6075]_ , \new_[6076]_ , \new_[6077]_ ,
    \new_[6078]_ , \new_[6079]_ , \new_[6080]_ , \new_[6081]_ ,
    \new_[6082]_ , \new_[6083]_ , \new_[6084]_ , \new_[6085]_ ,
    \new_[6086]_ , \new_[6087]_ , \new_[6088]_ , \new_[6089]_ ,
    \new_[6090]_ , \new_[6091]_ , \new_[6092]_ , \new_[6093]_ ,
    \new_[6094]_ , \new_[6095]_ , \new_[6096]_ , \new_[6097]_ ,
    \new_[6098]_ , \new_[6099]_ , \new_[6100]_ , \new_[6101]_ ,
    \new_[6102]_ , \new_[6103]_ , \new_[6104]_ , \new_[6105]_ ,
    \new_[6106]_ , \new_[6107]_ , \new_[6108]_ , \new_[6109]_ ,
    \new_[6110]_ , \new_[6111]_ , \new_[6112]_ , \new_[6113]_ ,
    \new_[6114]_ , \new_[6115]_ , \new_[6116]_ , \new_[6117]_ ,
    \new_[6118]_ , \new_[6119]_ , \new_[6120]_ , \new_[6121]_ ,
    \new_[6122]_ , \new_[6123]_ , \new_[6124]_ , \new_[6125]_ ,
    \new_[6126]_ , \new_[6127]_ , \new_[6128]_ , \new_[6129]_ ,
    \new_[6130]_ , \new_[6131]_ , \new_[6132]_ , \new_[6133]_ ,
    \new_[6134]_ , \new_[6135]_ , \new_[6136]_ , \new_[6137]_ ,
    \new_[6138]_ , \new_[6139]_ , \new_[6140]_ , \new_[6141]_ ,
    \new_[6142]_ , \new_[6143]_ , \new_[6144]_ , \new_[6145]_ ,
    \new_[6146]_ , \new_[6147]_ , \new_[6148]_ , \new_[6149]_ ,
    \new_[6150]_ , \new_[6151]_ , \new_[6152]_ , \new_[6153]_ ,
    \new_[6154]_ , \new_[6155]_ , \new_[6156]_ , \new_[6157]_ ,
    \new_[6158]_ , \new_[6159]_ , \new_[6160]_ , \new_[6161]_ ,
    \new_[6162]_ , \new_[6163]_ , \new_[6164]_ , \new_[6165]_ ,
    \new_[6166]_ , \new_[6167]_ , \new_[6168]_ , \new_[6169]_ ,
    \new_[6170]_ , \new_[6171]_ , \new_[6172]_ , \new_[6173]_ ,
    \new_[6174]_ , \new_[6175]_ , \new_[6176]_ , \new_[6177]_ ,
    \new_[6178]_ , \new_[6179]_ , \new_[6180]_ , \new_[6181]_ ,
    \new_[6182]_ , \new_[6183]_ , \new_[6184]_ , \new_[6185]_ ,
    \new_[6186]_ , \new_[6187]_ , \new_[6188]_ , \new_[6189]_ ,
    \new_[6190]_ , \new_[6191]_ , \new_[6192]_ , \new_[6193]_ ,
    \new_[6194]_ , \new_[6195]_ , \new_[6196]_ , \new_[6197]_ ,
    \new_[6198]_ , \new_[6199]_ , \new_[6200]_ , \new_[6201]_ ,
    \new_[6202]_ , \new_[6203]_ , \new_[6204]_ , \new_[6205]_ ,
    \new_[6206]_ , \new_[6207]_ , \new_[6208]_ , \new_[6209]_ ,
    \new_[6210]_ , \new_[6211]_ , \new_[6212]_ , \new_[6213]_ ,
    \new_[6214]_ , \new_[6215]_ , \new_[6216]_ , \new_[6217]_ ,
    \new_[6218]_ , \new_[6219]_ , \new_[6220]_ , \new_[6221]_ ,
    \new_[6222]_ , \new_[6223]_ , \new_[6224]_ , \new_[6225]_ ,
    \new_[6226]_ , \new_[6227]_ , \new_[6228]_ , \new_[6229]_ ,
    \new_[6230]_ , \new_[6231]_ , \new_[6232]_ , \new_[6233]_ ,
    \new_[6234]_ , \new_[6235]_ , \new_[6236]_ , \new_[6237]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6240]_ , \new_[6241]_ ,
    \new_[6242]_ , \new_[6243]_ , \new_[6244]_ , \new_[6245]_ ,
    \new_[6246]_ , \new_[6247]_ , \new_[6248]_ , \new_[6249]_ ,
    \new_[6250]_ , \new_[6251]_ , \new_[6252]_ , \new_[6253]_ ,
    \new_[6254]_ , \new_[6255]_ , \new_[6256]_ , \new_[6257]_ ,
    \new_[6258]_ , \new_[6259]_ , \new_[6260]_ , \new_[6261]_ ,
    \new_[6262]_ , \new_[6263]_ , \new_[6264]_ , \new_[6265]_ ,
    \new_[6266]_ , \new_[6267]_ , \new_[6268]_ , \new_[6269]_ ,
    \new_[6270]_ , \new_[6271]_ , \new_[6272]_ , \new_[6273]_ ,
    \new_[6274]_ , \new_[6275]_ , \new_[6276]_ , \new_[6277]_ ,
    \new_[6278]_ , \new_[6279]_ , \new_[6280]_ , \new_[6281]_ ,
    \new_[6282]_ , \new_[6283]_ , \new_[6284]_ , \new_[6285]_ ,
    \new_[6286]_ , \new_[6287]_ , \new_[6288]_ , \new_[6289]_ ,
    \new_[6290]_ , \new_[6291]_ , \new_[6292]_ , \new_[6293]_ ,
    \new_[6294]_ , \new_[6295]_ , \new_[6296]_ , \new_[6297]_ ,
    \new_[6298]_ , \new_[6299]_ , \new_[6300]_ , \new_[6301]_ ,
    \new_[6302]_ , \new_[6303]_ , \new_[6304]_ , \new_[6305]_ ,
    \new_[6306]_ , \new_[6307]_ , \new_[6308]_ , \new_[6309]_ ,
    \new_[6310]_ , \new_[6311]_ , \new_[6312]_ , \new_[6313]_ ,
    \new_[6314]_ , \new_[6315]_ , \new_[6316]_ , \new_[6317]_ ,
    \new_[6318]_ , \new_[6319]_ , \new_[6320]_ , \new_[6321]_ ,
    \new_[6322]_ , \new_[6323]_ , \new_[6324]_ , \new_[6325]_ ,
    \new_[6326]_ , \new_[6327]_ , \new_[6328]_ , \new_[6329]_ ,
    \new_[6330]_ , \new_[6331]_ , \new_[6332]_ , \new_[6333]_ ,
    \new_[6334]_ , \new_[6335]_ , \new_[6336]_ , \new_[6337]_ ,
    \new_[6338]_ , \new_[6339]_ , \new_[6340]_ , \new_[6341]_ ,
    \new_[6342]_ , \new_[6343]_ , \new_[6344]_ , \new_[6345]_ ,
    \new_[6346]_ , \new_[6347]_ , \new_[6348]_ , \new_[6349]_ ,
    \new_[6350]_ , \new_[6351]_ , \new_[6352]_ , \new_[6353]_ ,
    \new_[6354]_ , \new_[6355]_ , \new_[6356]_ , \new_[6357]_ ,
    \new_[6358]_ , \new_[6359]_ , \new_[6360]_ , \new_[6361]_ ,
    \new_[6362]_ , \new_[6363]_ , \new_[6364]_ , \new_[6365]_ ,
    \new_[6366]_ , \new_[6367]_ , \new_[6368]_ , \new_[6369]_ ,
    \new_[6370]_ , \new_[6371]_ , \new_[6372]_ , \new_[6373]_ ,
    \new_[6374]_ , \new_[6375]_ , \new_[6376]_ , \new_[6377]_ ,
    \new_[6378]_ , \new_[6379]_ , \new_[6380]_ , \new_[6381]_ ,
    \new_[6382]_ , \new_[6383]_ , \new_[6384]_ , \new_[6385]_ ,
    \new_[6386]_ , \new_[6387]_ , \new_[6388]_ , \new_[6389]_ ,
    \new_[6390]_ , \new_[6391]_ , \new_[6392]_ , \new_[6393]_ ,
    \new_[6394]_ , \new_[6395]_ , \new_[6396]_ , \new_[6397]_ ,
    \new_[6398]_ , \new_[6399]_ , \new_[6400]_ , \new_[6401]_ ,
    \new_[6402]_ , \new_[6403]_ , \new_[6404]_ , \new_[6405]_ ,
    \new_[6406]_ , \new_[6407]_ , \new_[6408]_ , \new_[6409]_ ,
    \new_[6410]_ , \new_[6411]_ , \new_[6412]_ , \new_[6413]_ ,
    \new_[6414]_ , \new_[6415]_ , \new_[6416]_ , \new_[6417]_ ,
    \new_[6418]_ , \new_[6419]_ , \new_[6420]_ , \new_[6421]_ ,
    \new_[6422]_ , \new_[6423]_ , \new_[6424]_ , \new_[6425]_ ,
    \new_[6426]_ , \new_[6427]_ , \new_[6428]_ , \new_[6429]_ ,
    \new_[6430]_ , \new_[6431]_ , \new_[6432]_ , \new_[6433]_ ,
    \new_[6434]_ , \new_[6435]_ , \new_[6436]_ , \new_[6437]_ ,
    \new_[6438]_ , \new_[6439]_ , \new_[6440]_ , \new_[6441]_ ,
    \new_[6442]_ , \new_[6443]_ , \new_[6444]_ , \new_[6445]_ ,
    \new_[6446]_ , \new_[6447]_ , \new_[6448]_ , \new_[6449]_ ,
    \new_[6450]_ , \new_[6451]_ , \new_[6452]_ , \new_[6453]_ ,
    \new_[6454]_ , \new_[6455]_ , \new_[6456]_ , \new_[6457]_ ,
    \new_[6458]_ , \new_[6459]_ , \new_[6460]_ , \new_[6461]_ ,
    \new_[6462]_ , \new_[6463]_ , \new_[6464]_ , \new_[6465]_ ,
    \new_[6466]_ , \new_[6467]_ , \new_[6468]_ , \new_[6469]_ ,
    \new_[6470]_ , \new_[6471]_ , \new_[6472]_ , \new_[6473]_ ,
    \new_[6474]_ , \new_[6475]_ , \new_[6476]_ , \new_[6477]_ ,
    \new_[6478]_ , \new_[6479]_ , \new_[6480]_ , \new_[6481]_ ,
    \new_[6482]_ , \new_[6483]_ , \new_[6484]_ , \new_[6485]_ ,
    \new_[6486]_ , \new_[6487]_ , \new_[6488]_ , \new_[6489]_ ,
    \new_[6490]_ , \new_[6491]_ , \new_[6492]_ , \new_[6493]_ ,
    \new_[6494]_ , \new_[6495]_ , \new_[6496]_ , \new_[6497]_ ,
    \new_[6498]_ , \new_[6499]_ , \new_[6500]_ , \new_[6501]_ ,
    \new_[6502]_ , \new_[6503]_ , \new_[6504]_ , \new_[6505]_ ,
    \new_[6506]_ , \new_[6507]_ , \new_[6508]_ , \new_[6509]_ ,
    \new_[6510]_ , \new_[6511]_ , \new_[6512]_ , \new_[6513]_ ,
    \new_[6514]_ , \new_[6515]_ , \new_[6516]_ , \new_[6517]_ ,
    \new_[6518]_ , \new_[6519]_ , \new_[6520]_ , \new_[6521]_ ,
    \new_[6522]_ , \new_[6523]_ , \new_[6524]_ , \new_[6525]_ ,
    \new_[6526]_ , \new_[6527]_ , \new_[6528]_ , \new_[6529]_ ,
    \new_[6530]_ , \new_[6531]_ , \new_[6532]_ , \new_[6533]_ ,
    \new_[6534]_ , \new_[6535]_ , \new_[6536]_ , \new_[6537]_ ,
    \new_[6538]_ , \new_[6539]_ , \new_[6540]_ , \new_[6541]_ ,
    \new_[6542]_ , \new_[6543]_ , \new_[6544]_ , \new_[6545]_ ,
    \new_[6546]_ , \new_[6547]_ , \new_[6548]_ , \new_[6549]_ ,
    \new_[6550]_ , \new_[6551]_ , \new_[6552]_ , \new_[6553]_ ,
    \new_[6554]_ , \new_[6555]_ , \new_[6556]_ , \new_[6557]_ ,
    \new_[6558]_ , \new_[6559]_ , \new_[6560]_ , \new_[6561]_ ,
    \new_[6562]_ , \new_[6563]_ , \new_[6564]_ , \new_[6565]_ ,
    \new_[6566]_ , \new_[6567]_ , \new_[6568]_ , \new_[6569]_ ,
    \new_[6570]_ , \new_[6571]_ , \new_[6572]_ , \new_[6573]_ ,
    \new_[6574]_ , \new_[6575]_ , \new_[6576]_ , \new_[6577]_ ,
    \new_[6578]_ , \new_[6579]_ , \new_[6580]_ , \new_[6581]_ ,
    \new_[6582]_ , \new_[6583]_ , \new_[6584]_ , \new_[6585]_ ,
    \new_[6586]_ , \new_[6587]_ , \new_[6588]_ , \new_[6589]_ ,
    \new_[6590]_ , \new_[6591]_ , \new_[6592]_ , \new_[6593]_ ,
    \new_[6594]_ , \new_[6595]_ , \new_[6596]_ , \new_[6597]_ ,
    \new_[6598]_ , \new_[6599]_ , \new_[6600]_ , \new_[6601]_ ,
    \new_[6602]_ , \new_[6603]_ , \new_[6604]_ , \new_[6605]_ ,
    \new_[6606]_ , \new_[6607]_ , \new_[6608]_ , \new_[6609]_ ,
    \new_[6610]_ , \new_[6611]_ , \new_[6612]_ , \new_[6613]_ ,
    \new_[6614]_ , \new_[6615]_ , \new_[6616]_ , \new_[6617]_ ,
    \new_[6618]_ , \new_[6619]_ , \new_[6620]_ , \new_[6621]_ ,
    \new_[6622]_ , \new_[6623]_ , \new_[6624]_ , \new_[6625]_ ,
    \new_[6626]_ , \new_[6627]_ , \new_[6628]_ , \new_[6629]_ ,
    \new_[6630]_ , \new_[6631]_ , \new_[6632]_ , \new_[6633]_ ,
    \new_[6634]_ , \new_[6635]_ , \new_[6636]_ , \new_[6637]_ ,
    \new_[6638]_ , \new_[6639]_ , \new_[6640]_ , \new_[6641]_ ,
    \new_[6642]_ , \new_[6643]_ , \new_[6644]_ , \new_[6645]_ ,
    \new_[6647]_ , \new_[6648]_ , \new_[6649]_ , \new_[6650]_ ,
    \new_[6651]_ , \new_[6652]_ , \new_[6653]_ , \new_[6654]_ ,
    \new_[6655]_ , \new_[6656]_ , \new_[6657]_ , \new_[6658]_ ,
    \new_[6659]_ , \new_[6660]_ , \new_[6661]_ , \new_[6662]_ ,
    \new_[6663]_ , \new_[6664]_ , \new_[6665]_ , \new_[6666]_ ,
    \new_[6667]_ , \new_[6668]_ , \new_[6669]_ , \new_[6670]_ ,
    \new_[6671]_ , \new_[6672]_ , \new_[6673]_ , \new_[6674]_ ,
    \new_[6675]_ , \new_[6676]_ , \new_[6677]_ , \new_[6678]_ ,
    \new_[6679]_ , \new_[6680]_ , \new_[6681]_ , \new_[6682]_ ,
    \new_[6683]_ , \new_[6684]_ , \new_[6685]_ , \new_[6686]_ ,
    \new_[6687]_ , \new_[6688]_ , \new_[6689]_ , \new_[6690]_ ,
    \new_[6691]_ , \new_[6692]_ , \new_[6693]_ , \new_[6694]_ ,
    \new_[6695]_ , \new_[6696]_ , \new_[6697]_ , \new_[6698]_ ,
    \new_[6699]_ , \new_[6700]_ , \new_[6701]_ , \new_[6702]_ ,
    \new_[6703]_ , \new_[6704]_ , \new_[6705]_ , \new_[6706]_ ,
    \new_[6707]_ , \new_[6708]_ , \new_[6709]_ , \new_[6710]_ ,
    \new_[6711]_ , \new_[6712]_ , \new_[6713]_ , \new_[6714]_ ,
    \new_[6715]_ , \new_[6716]_ , \new_[6717]_ , \new_[6718]_ ,
    \new_[6719]_ , \new_[6720]_ , \new_[6721]_ , \new_[6722]_ ,
    \new_[6723]_ , \new_[6724]_ , \new_[6725]_ , \new_[6726]_ ,
    \new_[6727]_ , \new_[6728]_ , \new_[6729]_ , \new_[6730]_ ,
    \new_[6731]_ , \new_[6732]_ , \new_[6733]_ , \new_[6734]_ ,
    \new_[6735]_ , \new_[6736]_ , \new_[6737]_ , \new_[6738]_ ,
    \new_[6739]_ , \new_[6740]_ , \new_[6741]_ , \new_[6742]_ ,
    \new_[6743]_ , \new_[6744]_ , \new_[6745]_ , \new_[6746]_ ,
    \new_[6747]_ , \new_[6748]_ , \new_[6749]_ , \new_[6750]_ ,
    \new_[6751]_ , \new_[6752]_ , \new_[6753]_ , \new_[6754]_ ,
    \new_[6755]_ , \new_[6756]_ , \new_[6757]_ , \new_[6758]_ ,
    \new_[6759]_ , \new_[6760]_ , \new_[6761]_ , \new_[6762]_ ,
    \new_[6763]_ , \new_[6764]_ , \new_[6765]_ , \new_[6766]_ ,
    \new_[6767]_ , \new_[6768]_ , \new_[6769]_ , \new_[6770]_ ,
    \new_[6771]_ , \new_[6772]_ , \new_[6773]_ , \new_[6774]_ ,
    \new_[6775]_ , \new_[6776]_ , \new_[6777]_ , \new_[6778]_ ,
    \new_[6779]_ , \new_[6780]_ , \new_[6781]_ , \new_[6782]_ ,
    \new_[6783]_ , \new_[6784]_ , \new_[6785]_ , \new_[6786]_ ,
    \new_[6787]_ , \new_[6788]_ , \new_[6789]_ , \new_[6790]_ ,
    \new_[6791]_ , \new_[6792]_ , \new_[6793]_ , \new_[6794]_ ,
    \new_[6795]_ , \new_[6796]_ , \new_[6797]_ , \new_[6798]_ ,
    \new_[6799]_ , \new_[6800]_ , \new_[6801]_ , \new_[6802]_ ,
    \new_[6803]_ , \new_[6804]_ , \new_[6805]_ , \new_[6806]_ ,
    \new_[6807]_ , \new_[6808]_ , \new_[6809]_ , \new_[6810]_ ,
    \new_[6811]_ , \new_[6812]_ , \new_[6813]_ , \new_[6814]_ ,
    \new_[6815]_ , \new_[6816]_ , \new_[6817]_ , \new_[6818]_ ,
    \new_[6819]_ , \new_[6820]_ , \new_[6821]_ , \new_[6822]_ ,
    \new_[6823]_ , \new_[6824]_ , \new_[6825]_ , \new_[6826]_ ,
    \new_[6827]_ , \new_[6828]_ , \new_[6829]_ , \new_[6830]_ ,
    \new_[6831]_ , \new_[6832]_ , \new_[6833]_ , \new_[6834]_ ,
    \new_[6835]_ , \new_[6836]_ , \new_[6837]_ , \new_[6838]_ ,
    \new_[6839]_ , \new_[6840]_ , \new_[6841]_ , \new_[6866]_ ,
    \new_[6894]_ , \new_[6948]_ , \new_[6949]_ , \new_[6950]_ ,
    \new_[6951]_ , \new_[6952]_ , \new_[6953]_ , \new_[6954]_ ,
    \new_[6955]_ , \new_[6956]_ , \new_[6957]_ , \new_[6958]_ ,
    \new_[6959]_ , \new_[6960]_ , \new_[6961]_ , \new_[6962]_ ,
    \new_[6963]_ , \new_[6964]_ , \new_[6965]_ , \new_[6966]_ ,
    \new_[6967]_ , \new_[6968]_ , \new_[6969]_ , \new_[6970]_ ,
    \new_[6971]_ , \new_[6972]_ , \new_[6973]_ , \new_[6974]_ ,
    \new_[6975]_ , \new_[6976]_ , \new_[6977]_ , \new_[6978]_ ,
    \new_[6979]_ , \new_[6980]_ , \new_[6981]_ , \new_[6982]_ ,
    \new_[6983]_ , \new_[6984]_ , \new_[6985]_ , \new_[6986]_ ,
    \new_[6987]_ , \new_[6988]_ , \new_[6989]_ , \new_[6990]_ ,
    \new_[6991]_ , \new_[6992]_ , \new_[6993]_ , \new_[6994]_ ,
    \new_[6995]_ , \new_[6996]_ , \new_[6997]_ , \new_[6998]_ ,
    \new_[6999]_ , \new_[7000]_ , \new_[7001]_ , \new_[7002]_ ,
    \new_[7003]_ , \new_[7004]_ , \new_[7005]_ , \new_[7006]_ ,
    \new_[7007]_ , \new_[7008]_ , \new_[7009]_ , \new_[7010]_ ,
    \new_[7011]_ , \new_[7012]_ , \new_[7013]_ , \new_[7014]_ ,
    \new_[7015]_ , \new_[7016]_ , \new_[7017]_ , \new_[7018]_ ,
    \new_[7019]_ , \new_[7020]_ , \new_[7021]_ , \new_[7022]_ ,
    \new_[7023]_ , \new_[7024]_ , \new_[7025]_ , \new_[7026]_ ,
    \new_[7027]_ , \new_[7028]_ , \new_[7029]_ , \new_[7030]_ ,
    \new_[7031]_ , \new_[7032]_ , \new_[7033]_ , \new_[7034]_ ,
    \new_[7035]_ , \new_[7036]_ , \new_[7037]_ , \new_[7038]_ ,
    \new_[7039]_ , \new_[7040]_ , \new_[7041]_ , \new_[7042]_ ,
    \new_[7043]_ , \new_[7044]_ , \new_[7045]_ , \new_[7046]_ ,
    \new_[7047]_ , \new_[7048]_ , \new_[7049]_ , \new_[7050]_ ,
    \new_[7051]_ , \new_[7052]_ , \new_[7053]_ , \new_[7054]_ ,
    \new_[7055]_ , \new_[7056]_ , \new_[7057]_ , \new_[7058]_ ,
    \new_[7059]_ , \new_[7060]_ , \new_[7061]_ , \new_[7063]_ ,
    \new_[7064]_ , \new_[7065]_ , \new_[7066]_ , \new_[7067]_ ,
    \new_[7068]_ , \new_[7069]_ , \new_[7070]_ , \new_[7071]_ ,
    \new_[7072]_ , \new_[7073]_ , \new_[7074]_ , \new_[7075]_ ,
    \new_[7076]_ , \new_[7077]_ , \new_[7078]_ , \new_[7079]_ ,
    \new_[7080]_ , \new_[7081]_ , \new_[7082]_ , \new_[7083]_ ,
    \new_[7084]_ , \new_[7085]_ , \new_[7086]_ , \new_[7087]_ ,
    \new_[7088]_ , \new_[7089]_ , \new_[7090]_ , \new_[7091]_ ,
    \new_[7092]_ , \new_[7093]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7096]_ , \new_[7097]_ , \new_[7098]_ , \new_[7099]_ ,
    \new_[7100]_ , \new_[7101]_ , \new_[7102]_ , \new_[7103]_ ,
    \new_[7104]_ , \new_[7105]_ , \new_[7106]_ , \new_[7107]_ ,
    \new_[7108]_ , \new_[7109]_ , \new_[7110]_ , \new_[7111]_ ,
    \new_[7112]_ , \new_[7113]_ , \new_[7114]_ , \new_[7115]_ ,
    \new_[7116]_ , \new_[7117]_ , \new_[7118]_ , \new_[7119]_ ,
    \new_[7120]_ , \new_[7121]_ , \new_[7122]_ , \new_[7123]_ ,
    \new_[7124]_ , \new_[7125]_ , \new_[7126]_ , \new_[7127]_ ,
    \new_[7128]_ , \new_[7129]_ , \new_[7130]_ , \new_[7131]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7134]_ , \new_[7135]_ ,
    \new_[7136]_ , \new_[7137]_ , \new_[7138]_ , \new_[7139]_ ,
    \new_[7140]_ , \new_[7141]_ , \new_[7142]_ , \new_[7143]_ ,
    \new_[7144]_ , \new_[7145]_ , \new_[7146]_ , \new_[7147]_ ,
    \new_[7148]_ , \new_[7149]_ , \new_[7150]_ , \new_[7151]_ ,
    \new_[7152]_ , \new_[7153]_ , \new_[7154]_ , \new_[7155]_ ,
    \new_[7156]_ , \new_[7157]_ , \new_[7158]_ , \new_[7159]_ ,
    \new_[7160]_ , \new_[7161]_ , \new_[7162]_ , \new_[7163]_ ,
    \new_[7164]_ , \new_[7165]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7168]_ , \new_[7169]_ , \new_[7170]_ , \new_[7171]_ ,
    \new_[7172]_ , \new_[7173]_ , \new_[7174]_ , \new_[7175]_ ,
    \new_[7176]_ , \new_[7177]_ , \new_[7178]_ , \new_[7179]_ ,
    \new_[7180]_ , \new_[7181]_ , \new_[7182]_ , \new_[7183]_ ,
    \new_[7184]_ , \new_[7185]_ , \new_[7186]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7189]_ , \new_[7190]_ , \new_[7191]_ ,
    \new_[7192]_ , \new_[7193]_ , \new_[7194]_ , \new_[7195]_ ,
    \new_[7196]_ , \new_[7197]_ , \new_[7198]_ , \new_[7199]_ ,
    \new_[7200]_ , \new_[7201]_ , \new_[7202]_ , \new_[7203]_ ,
    \new_[7204]_ , \new_[7205]_ , \new_[7206]_ , \new_[7207]_ ,
    \new_[7208]_ , \new_[7209]_ , \new_[7210]_ , \new_[7211]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7214]_ , \new_[7215]_ ,
    \new_[7216]_ , \new_[7217]_ , \new_[7218]_ , \new_[7219]_ ,
    \new_[7220]_ , \new_[7221]_ , \new_[7222]_ , \new_[7223]_ ,
    \new_[7224]_ , \new_[7225]_ , \new_[7226]_ , \new_[7227]_ ,
    \new_[7228]_ , \new_[7229]_ , \new_[7230]_ , \new_[7231]_ ,
    \new_[7232]_ , \new_[7233]_ , \new_[7234]_ , \new_[7235]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7241]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7244]_ , \new_[7245]_ , \new_[7246]_ , \new_[7247]_ ,
    \new_[7248]_ , \new_[7249]_ , \new_[7250]_ , \new_[7251]_ ,
    \new_[7252]_ , \new_[7253]_ , \new_[7254]_ , \new_[7255]_ ,
    \new_[7256]_ , \new_[7257]_ , \new_[7258]_ , \new_[7259]_ ,
    \new_[7260]_ , \new_[7261]_ , \new_[7262]_ , \new_[7263]_ ,
    \new_[7264]_ , \new_[7265]_ , \new_[7266]_ , \new_[7267]_ ,
    \new_[7268]_ , \new_[7269]_ , \new_[7270]_ , \new_[7271]_ ,
    \new_[7272]_ , \new_[7273]_ , \new_[7274]_ , \new_[7275]_ ,
    \new_[7277]_ , \new_[7278]_ , \new_[7279]_ , \new_[7280]_ ,
    \new_[7281]_ , \new_[7282]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7285]_ , \new_[7286]_ , \new_[7287]_ , \new_[7288]_ ,
    \new_[7289]_ , \new_[7290]_ , \new_[7291]_ , \new_[7292]_ ,
    \new_[7293]_ , \new_[7294]_ , \new_[7295]_ , \new_[7296]_ ,
    \new_[7297]_ , \new_[7298]_ , \new_[7299]_ , \new_[7300]_ ,
    \new_[7301]_ , \new_[7302]_ , \new_[7303]_ , \new_[7304]_ ,
    \new_[7305]_ , \new_[7306]_ , \new_[7307]_ , \new_[7308]_ ,
    \new_[7309]_ , \new_[7310]_ , \new_[7311]_ , \new_[7312]_ ,
    \new_[7313]_ , \new_[7314]_ , \new_[7315]_ , \new_[7316]_ ,
    \new_[7317]_ , \new_[7318]_ , \new_[7319]_ , \new_[7320]_ ,
    \new_[7321]_ , \new_[7322]_ , \new_[7323]_ , \new_[7324]_ ,
    \new_[7325]_ , \new_[7326]_ , \new_[7327]_ , \new_[7328]_ ,
    \new_[7329]_ , \new_[7330]_ , \new_[7331]_ , \new_[7332]_ ,
    \new_[7333]_ , \new_[7334]_ , \new_[7335]_ , \new_[7336]_ ,
    \new_[7337]_ , \new_[7338]_ , \new_[7339]_ , \new_[7340]_ ,
    \new_[7341]_ , \new_[7342]_ , \new_[7343]_ , \new_[7344]_ ,
    \new_[7345]_ , \new_[7346]_ , \new_[7347]_ , \new_[7348]_ ,
    \new_[7349]_ , \new_[7350]_ , \new_[7351]_ , \new_[7352]_ ,
    \new_[7353]_ , \new_[7354]_ , \new_[7355]_ , \new_[7356]_ ,
    \new_[7357]_ , \new_[7358]_ , \new_[7359]_ , \new_[7360]_ ,
    \new_[7361]_ , \new_[7362]_ , \new_[7363]_ , \new_[7364]_ ,
    \new_[7365]_ , \new_[7366]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7369]_ , \new_[7370]_ , \new_[7372]_ , \new_[7373]_ ,
    \new_[7374]_ , \new_[7375]_ , \new_[7376]_ , \new_[7377]_ ,
    \new_[7378]_ , \new_[7379]_ , \new_[7380]_ , \new_[7381]_ ,
    \new_[7382]_ , \new_[7383]_ , \new_[7384]_ , \new_[7385]_ ,
    \new_[7386]_ , \new_[7387]_ , \new_[7388]_ , \new_[7389]_ ,
    \new_[7390]_ , \new_[7391]_ , \new_[7392]_ , \new_[7393]_ ,
    \new_[7394]_ , \new_[7395]_ , \new_[7396]_ , \new_[7397]_ ,
    \new_[7398]_ , \new_[7399]_ , \new_[7400]_ , \new_[7401]_ ,
    \new_[7402]_ , \new_[7403]_ , \new_[7404]_ , \new_[7405]_ ,
    \new_[7406]_ , \new_[7407]_ , \new_[7408]_ , \new_[7409]_ ,
    \new_[7410]_ , \new_[7411]_ , \new_[7412]_ , \new_[7413]_ ,
    \new_[7414]_ , \new_[7415]_ , \new_[7416]_ , \new_[7417]_ ,
    \new_[7418]_ , \new_[7419]_ , \new_[7420]_ , \new_[7421]_ ,
    \new_[7422]_ , \new_[7423]_ , \new_[7424]_ , \new_[7425]_ ,
    \new_[7426]_ , \new_[7427]_ , \new_[7428]_ , \new_[7429]_ ,
    \new_[7430]_ , \new_[7431]_ , \new_[7432]_ , \new_[7433]_ ,
    \new_[7438]_ , \new_[7439]_ , \new_[7440]_ , \new_[7442]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7445]_ , \new_[7446]_ ,
    \new_[7447]_ , \new_[7448]_ , \new_[7449]_ , \new_[7450]_ ,
    \new_[7451]_ , \new_[7452]_ , \new_[7453]_ , \new_[7454]_ ,
    \new_[7455]_ , \new_[7456]_ , \new_[7457]_ , \new_[7458]_ ,
    \new_[7459]_ , \new_[7460]_ , \new_[7461]_ , \new_[7462]_ ,
    \new_[7463]_ , \new_[7464]_ , \new_[7465]_ , \new_[7466]_ ,
    \new_[7467]_ , \new_[7468]_ , \new_[7469]_ , \new_[7470]_ ,
    \new_[7471]_ , \new_[7472]_ , \new_[7473]_ , \new_[7474]_ ,
    \new_[7475]_ , \new_[7476]_ , \new_[7477]_ , \new_[7478]_ ,
    \new_[7479]_ , \new_[7480]_ , \new_[7481]_ , \new_[7482]_ ,
    \new_[7483]_ , \new_[7484]_ , \new_[7485]_ , \new_[7486]_ ,
    \new_[7487]_ , \new_[7488]_ , \new_[7489]_ , \new_[7490]_ ,
    \new_[7491]_ , \new_[7492]_ , \new_[7493]_ , \new_[7494]_ ,
    \new_[7495]_ , \new_[7496]_ , \new_[7497]_ , \new_[7498]_ ,
    \new_[7499]_ , \new_[7500]_ , \new_[7501]_ , \new_[7502]_ ,
    \new_[7503]_ , \new_[7504]_ , \new_[7505]_ , \new_[7506]_ ,
    \new_[7507]_ , \new_[7508]_ , \new_[7509]_ , \new_[7510]_ ,
    \new_[7511]_ , \new_[7512]_ , \new_[7513]_ , \new_[7514]_ ,
    \new_[7515]_ , \new_[7516]_ , \new_[7517]_ , \new_[7518]_ ,
    \new_[7519]_ , \new_[7520]_ , \new_[7521]_ , \new_[7522]_ ,
    \new_[7523]_ , \new_[7524]_ , \new_[7525]_ , \new_[7526]_ ,
    \new_[7527]_ , \new_[7528]_ , \new_[7529]_ , \new_[7530]_ ,
    \new_[7531]_ , \new_[7532]_ , \new_[7533]_ , \new_[7534]_ ,
    \new_[7535]_ , \new_[7536]_ , \new_[7537]_ , \new_[7538]_ ,
    \new_[7539]_ , \new_[7540]_ , \new_[7541]_ , \new_[7542]_ ,
    \new_[7543]_ , \new_[7544]_ , \new_[7545]_ , \new_[7546]_ ,
    \new_[7547]_ , \new_[7548]_ , \new_[7549]_ , \new_[7550]_ ,
    \new_[7551]_ , \new_[7552]_ , \new_[7553]_ , \new_[7554]_ ,
    \new_[7555]_ , \new_[7556]_ , \new_[7557]_ , \new_[7558]_ ,
    \new_[7559]_ , \new_[7560]_ , \new_[7561]_ , \new_[7562]_ ,
    \new_[7563]_ , \new_[7564]_ , \new_[7565]_ , \new_[7566]_ ,
    \new_[7567]_ , \new_[7568]_ , \new_[7569]_ , \new_[7570]_ ,
    \new_[7571]_ , \new_[7572]_ , \new_[7573]_ , \new_[7574]_ ,
    \new_[7575]_ , \new_[7576]_ , \new_[7577]_ , \new_[7578]_ ,
    \new_[7579]_ , \new_[7580]_ , \new_[7581]_ , \new_[7582]_ ,
    \new_[7583]_ , \new_[7584]_ , \new_[7585]_ , \new_[7586]_ ,
    \new_[7587]_ , \new_[7588]_ , \new_[7589]_ , \new_[7590]_ ,
    \new_[7591]_ , \new_[7592]_ , \new_[7593]_ , \new_[7594]_ ,
    \new_[7595]_ , \new_[7596]_ , \new_[7597]_ , \new_[7598]_ ,
    \new_[7599]_ , \new_[7600]_ , \new_[7601]_ , \new_[7602]_ ,
    \new_[7603]_ , \new_[7604]_ , \new_[7605]_ , \new_[7606]_ ,
    \new_[7607]_ , \new_[7608]_ , \new_[7610]_ , \new_[7612]_ ,
    \new_[7613]_ , \new_[7614]_ , \new_[7615]_ , \new_[7616]_ ,
    \new_[7617]_ , \new_[7618]_ , \new_[7619]_ , \new_[7620]_ ,
    \new_[7621]_ , \new_[7622]_ , \new_[7623]_ , \new_[7624]_ ,
    \new_[7625]_ , \new_[7626]_ , \new_[7627]_ , \new_[7628]_ ,
    \new_[7629]_ , \new_[7630]_ , \new_[7631]_ , \new_[7632]_ ,
    \new_[7633]_ , \new_[7634]_ , \new_[7635]_ , \new_[7636]_ ,
    \new_[7637]_ , \new_[7639]_ , \new_[7640]_ , \new_[7641]_ ,
    \new_[7642]_ , \new_[7647]_ , \new_[7648]_ , \new_[7649]_ ,
    \new_[7650]_ , \new_[7651]_ , \new_[7652]_ , \new_[7653]_ ,
    \new_[7654]_ , \new_[7655]_ , \new_[7656]_ , \new_[7657]_ ,
    \new_[7658]_ , \new_[7659]_ , \new_[7660]_ , \new_[7661]_ ,
    \new_[7662]_ , \new_[7663]_ , \new_[7664]_ , \new_[7665]_ ,
    \new_[7666]_ , \new_[7668]_ , \new_[7669]_ , \new_[7670]_ ,
    \new_[7671]_ , \new_[7672]_ , \new_[7673]_ , \new_[7674]_ ,
    \new_[7675]_ , \new_[7676]_ , \new_[7677]_ , \new_[7678]_ ,
    \new_[7679]_ , \new_[7680]_ , \new_[7681]_ , \new_[7682]_ ,
    \new_[7683]_ , \new_[7684]_ , \new_[7685]_ , \new_[7686]_ ,
    \new_[7687]_ , \new_[7688]_ , \new_[7689]_ , \new_[7690]_ ,
    \new_[7691]_ , \new_[7692]_ , \new_[7693]_ , \new_[7694]_ ,
    \new_[7695]_ , \new_[7696]_ , \new_[7697]_ , \new_[7698]_ ,
    \new_[7699]_ , \new_[7700]_ , \new_[7701]_ , \new_[7702]_ ,
    \new_[7703]_ , \new_[7704]_ , \new_[7705]_ , \new_[7706]_ ,
    \new_[7707]_ , \new_[7708]_ , \new_[7709]_ , \new_[7710]_ ,
    \new_[7711]_ , \new_[7712]_ , \new_[7713]_ , \new_[7714]_ ,
    \new_[7715]_ , \new_[7716]_ , \new_[7717]_ , \new_[7718]_ ,
    \new_[7720]_ , \new_[7721]_ , \new_[7722]_ , \new_[7723]_ ,
    \new_[7724]_ , \new_[7725]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7731]_ , \new_[7732]_ ,
    \new_[7733]_ , \new_[7734]_ , \new_[7735]_ , \new_[7736]_ ,
    \new_[7737]_ , \new_[7738]_ , \new_[7739]_ , \new_[7740]_ ,
    \new_[7741]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7745]_ , \new_[7746]_ , \new_[7747]_ , \new_[7748]_ ,
    \new_[7749]_ , \new_[7750]_ , \new_[7751]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7754]_ , \new_[7755]_ , \new_[7756]_ ,
    \new_[7757]_ , \new_[7758]_ , \new_[7759]_ , \new_[7760]_ ,
    \new_[7761]_ , \new_[7763]_ , \new_[7765]_ , \new_[7766]_ ,
    \new_[7767]_ , \new_[7768]_ , \new_[7769]_ , \new_[7770]_ ,
    \new_[7771]_ , \new_[7772]_ , \new_[7773]_ , \new_[7774]_ ,
    \new_[7775]_ , \new_[7776]_ , \new_[7777]_ , \new_[7778]_ ,
    \new_[7779]_ , \new_[7780]_ , \new_[7781]_ , \new_[7782]_ ,
    \new_[7783]_ , \new_[7784]_ , \new_[7785]_ , \new_[7786]_ ,
    \new_[7787]_ , \new_[7788]_ , \new_[7789]_ , \new_[7798]_ ,
    \new_[7804]_ , \new_[7805]_ , \new_[7806]_ , \new_[7807]_ ,
    \new_[7808]_ , \new_[7809]_ , \new_[7810]_ , \new_[7811]_ ,
    \new_[7812]_ , \new_[7813]_ , \new_[7814]_ , \new_[7816]_ ,
    \new_[7817]_ , \new_[7818]_ , \new_[7819]_ , \new_[7820]_ ,
    \new_[7821]_ , \new_[7822]_ , \new_[7823]_ , \new_[7824]_ ,
    \new_[7825]_ , \new_[7826]_ , \new_[7827]_ , \new_[7828]_ ,
    \new_[7830]_ , \new_[7833]_ , \new_[7837]_ , \new_[7838]_ ,
    \new_[7839]_ , \new_[7850]_ , \new_[7851]_ , \new_[7852]_ ,
    \new_[7854]_ , \new_[7855]_ , \new_[7856]_ , \new_[7857]_ ,
    \new_[7858]_ , \new_[7859]_ , \new_[7861]_ , \new_[7862]_ ,
    \new_[7863]_ , \new_[7864]_ , \new_[7865]_ , \new_[7866]_ ,
    \new_[7871]_ , \new_[7872]_ , \new_[7873]_ , \new_[7874]_ ,
    \new_[7875]_ , \new_[7885]_ , \new_[7886]_ , \new_[7907]_ ,
    \new_[7908]_ , \new_[7909]_ , \new_[7910]_ , \new_[7911]_ ,
    \new_[7912]_ , \new_[7913]_ , \new_[7914]_ , \new_[7915]_ ,
    \new_[7917]_ , \new_[7918]_ , \new_[7919]_ , \new_[7920]_ ,
    \new_[7921]_ , \new_[7922]_ , \new_[7924]_ , \new_[7925]_ ,
    \new_[7926]_ , \new_[7927]_ , \new_[7929]_ , \new_[7930]_ ,
    \new_[7931]_ , \new_[7932]_ , \new_[7933]_ , \new_[7934]_ ,
    \new_[7935]_ , \new_[7936]_ , \new_[7937]_ , \new_[7938]_ ,
    \new_[7939]_ , \new_[7941]_ , \new_[7942]_ , \new_[7943]_ ,
    \new_[7944]_ , \new_[7945]_ , \new_[7950]_ , \new_[7951]_ ,
    \new_[7956]_ , \new_[7957]_ , \new_[7960]_ , \new_[7966]_ ,
    \new_[7968]_ , \new_[7969]_ , \new_[7970]_ , \new_[7971]_ ,
    \new_[7972]_ , \new_[7973]_ , \new_[7974]_ , \new_[7975]_ ,
    \new_[7976]_ , \new_[7977]_ , \new_[7978]_ , \new_[7979]_ ,
    \new_[7981]_ , \new_[7982]_ , \new_[7983]_ , \new_[7984]_ ,
    \new_[7985]_ , \new_[7986]_ , \new_[7987]_ , \new_[7988]_ ,
    \new_[7989]_ , \new_[7990]_ , \new_[7991]_ , \new_[7992]_ ,
    \new_[7993]_ , \new_[7994]_ , \new_[7995]_ , \new_[7996]_ ,
    \new_[7997]_ , \new_[7998]_ , \new_[7999]_ , \new_[8000]_ ,
    \new_[8001]_ , \new_[8002]_ , \new_[8003]_ , \new_[8004]_ ,
    \new_[8005]_ , \new_[8013]_ , \new_[8014]_ , \new_[8015]_ ,
    \new_[8016]_ , \new_[8017]_ , \new_[8018]_ , \new_[8019]_ ,
    \new_[8020]_ , \new_[8021]_ , \new_[8022]_ , \new_[8023]_ ,
    \new_[8024]_ , \new_[8025]_ , \new_[8026]_ , \new_[8027]_ ,
    \new_[8028]_ , \new_[8029]_ , \new_[8030]_ , \new_[8031]_ ,
    \new_[8032]_ , \new_[8034]_ , \new_[8035]_ , \new_[8036]_ ,
    \new_[8037]_ , \new_[8038]_ , \new_[8039]_ , \new_[8040]_ ,
    \new_[8041]_ , \new_[8042]_ , \new_[8043]_ , \new_[8044]_ ,
    \new_[8045]_ , \new_[8046]_ , \new_[8047]_ , \new_[8048]_ ,
    \new_[8049]_ , \new_[8050]_ , \new_[8051]_ , \new_[8052]_ ,
    \new_[8053]_ , \new_[8054]_ , \new_[8055]_ , \new_[8056]_ ,
    \new_[8057]_ , \new_[8058]_ , \new_[8059]_ , \new_[8060]_ ,
    \new_[8061]_ , \new_[8063]_ , \new_[8064]_ , \new_[8065]_ ,
    \new_[8066]_ , \new_[8067]_ , \new_[8068]_ , \new_[8070]_ ,
    \new_[8071]_ , \new_[8072]_ , \new_[8073]_ , \new_[8074]_ ,
    \new_[8075]_ , \new_[8076]_ , \new_[8077]_ , \new_[8078]_ ,
    \new_[8079]_ , \new_[8080]_ , \new_[8081]_ , \new_[8082]_ ,
    \new_[8083]_ , \new_[8084]_ , \new_[8085]_ , \new_[8092]_ ,
    \new_[8093]_ , \new_[8094]_ , \new_[8102]_ , \new_[8104]_ ,
    \new_[8105]_ , \new_[8106]_ , \new_[8107]_ , \new_[8108]_ ,
    \new_[8109]_ , \new_[8110]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8143]_ , \new_[8144]_ , \new_[8145]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8148]_ , \new_[8149]_ , \new_[8150]_ ,
    \new_[8151]_ , \new_[8152]_ , \new_[8153]_ , \new_[8154]_ ,
    \new_[8155]_ , \new_[8156]_ , \new_[8157]_ , \new_[8158]_ ,
    \new_[8159]_ , \new_[8160]_ , \new_[8161]_ , \new_[8162]_ ,
    \new_[8163]_ , \new_[8164]_ , \new_[8165]_ , \new_[8166]_ ,
    \new_[8167]_ , \new_[8168]_ , \new_[8169]_ , \new_[8170]_ ,
    \new_[8171]_ , \new_[8172]_ , \new_[8173]_ , \new_[8174]_ ,
    \new_[8175]_ , \new_[8177]_ , \new_[8179]_ , \new_[8185]_ ,
    \new_[8186]_ , \new_[8187]_ , \new_[8188]_ , \new_[8189]_ ,
    \new_[8190]_ , \new_[8191]_ , \new_[8192]_ , \new_[8194]_ ,
    \new_[8195]_ , \new_[8196]_ , \new_[8197]_ , \new_[8198]_ ,
    \new_[8199]_ , \new_[8200]_ , \new_[8201]_ , \new_[8202]_ ,
    \new_[8203]_ , \new_[8204]_ , \new_[8205]_ , \new_[8215]_ ,
    \new_[8216]_ , \new_[8217]_ , \new_[8218]_ , \new_[8219]_ ,
    \new_[8220]_ , \new_[8229]_ , \new_[8230]_ , \new_[8231]_ ,
    \new_[8232]_ , \new_[8258]_ , \new_[8259]_ , \new_[8260]_ ,
    \new_[8261]_ , \new_[8262]_ , \new_[8263]_ , \new_[8264]_ ,
    \new_[8265]_ , \new_[8266]_ , \new_[8267]_ , \new_[8268]_ ,
    \new_[8269]_ , \new_[8270]_ , \new_[8271]_ , \new_[8272]_ ,
    \new_[8273]_ , \new_[8274]_ , \new_[8275]_ , \new_[8276]_ ,
    \new_[8277]_ , \new_[8278]_ , \new_[8279]_ , \new_[8280]_ ,
    \new_[8281]_ , \new_[8282]_ , \new_[8283]_ , \new_[8284]_ ,
    \new_[8285]_ , \new_[8286]_ , \new_[8287]_ , \new_[8288]_ ,
    \new_[8289]_ , \new_[8290]_ , \new_[8291]_ , \new_[8292]_ ,
    \new_[8293]_ , \new_[8294]_ , \new_[8295]_ , \new_[8296]_ ,
    \new_[8297]_ , \new_[8298]_ , \new_[8299]_ , \new_[8300]_ ,
    \new_[8301]_ , \new_[8302]_ , \new_[8303]_ , \new_[8304]_ ,
    \new_[8305]_ , \new_[8306]_ , \new_[8307]_ , \new_[8308]_ ,
    \new_[8309]_ , \new_[8310]_ , \new_[8311]_ , \new_[8312]_ ,
    \new_[8313]_ , \new_[8314]_ , \new_[8315]_ , \new_[8316]_ ,
    \new_[8317]_ , \new_[8318]_ , \new_[8319]_ , \new_[8320]_ ,
    \new_[8321]_ , \new_[8322]_ , \new_[8323]_ , \new_[8324]_ ,
    \new_[8325]_ , \new_[8326]_ , \new_[8327]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8330]_ , \new_[8331]_ , \new_[8332]_ ,
    \new_[8333]_ , \new_[8334]_ , \new_[8335]_ , \new_[8336]_ ,
    \new_[8337]_ , \new_[8338]_ , \new_[8339]_ , \new_[8340]_ ,
    \new_[8341]_ , \new_[8342]_ , \new_[8343]_ , \new_[8344]_ ,
    \new_[8345]_ , \new_[8346]_ , \new_[8347]_ , \new_[8348]_ ,
    \new_[8349]_ , \new_[8350]_ , \new_[8351]_ , \new_[8352]_ ,
    \new_[8353]_ , \new_[8354]_ , \new_[8355]_ , \new_[8356]_ ,
    \new_[8357]_ , \new_[8358]_ , \new_[8359]_ , \new_[8360]_ ,
    \new_[8361]_ , \new_[8362]_ , \new_[8364]_ , \new_[8365]_ ,
    \new_[8366]_ , \new_[8367]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8378]_ , \new_[8380]_ , \new_[8382]_ , \new_[8385]_ ,
    \new_[8387]_ , \new_[8388]_ , \new_[8389]_ , \new_[8390]_ ,
    \new_[8391]_ , \new_[8392]_ , \new_[8393]_ , \new_[8394]_ ,
    \new_[8395]_ , \new_[8396]_ , \new_[8397]_ , \new_[8398]_ ,
    \new_[8399]_ , \new_[8400]_ , \new_[8401]_ , \new_[8402]_ ,
    \new_[8403]_ , \new_[8404]_ , \new_[8405]_ , \new_[8406]_ ,
    \new_[8407]_ , \new_[8408]_ , \new_[8409]_ , \new_[8410]_ ,
    \new_[8413]_ , \new_[8414]_ , \new_[8415]_ , \new_[8416]_ ,
    \new_[8417]_ , \new_[8418]_ , \new_[8419]_ , \new_[8420]_ ,
    \new_[8421]_ , \new_[8423]_ , \new_[8424]_ , \new_[8425]_ ,
    \new_[8426]_ , \new_[8427]_ , \new_[8428]_ , \new_[8429]_ ,
    \new_[8430]_ , \new_[8431]_ , \new_[8432]_ , \new_[8433]_ ,
    \new_[8434]_ , \new_[8435]_ , \new_[8436]_ , \new_[8437]_ ,
    \new_[8438]_ , \new_[8439]_ , \new_[8440]_ , \new_[8441]_ ,
    \new_[8442]_ , \new_[8443]_ , \new_[8444]_ , \new_[8445]_ ,
    \new_[8446]_ , \new_[8447]_ , \new_[8448]_ , \new_[8449]_ ,
    \new_[8450]_ , \new_[8451]_ , \new_[8452]_ , \new_[8453]_ ,
    \new_[8454]_ , \new_[8455]_ , \new_[8456]_ , \new_[8457]_ ,
    \new_[8469]_ , \new_[8470]_ , \new_[8471]_ , \new_[8472]_ ,
    \new_[8473]_ , \new_[8474]_ , \new_[8475]_ , \new_[8476]_ ,
    \new_[8477]_ , \new_[8479]_ , \new_[8480]_ , \new_[8481]_ ,
    \new_[8482]_ , \new_[8483]_ , \new_[8484]_ , \new_[8485]_ ,
    \new_[8486]_ , \new_[8487]_ , \new_[8488]_ , \new_[8489]_ ,
    \new_[8490]_ , \new_[8491]_ , \new_[8492]_ , \new_[8493]_ ,
    \new_[8495]_ , \new_[8496]_ , \new_[8497]_ , \new_[8498]_ ,
    \new_[8499]_ , \new_[8500]_ , \new_[8501]_ , \new_[8502]_ ,
    \new_[8503]_ , \new_[8504]_ , \new_[8505]_ , \new_[8506]_ ,
    \new_[8507]_ , \new_[8508]_ , \new_[8509]_ , \new_[8510]_ ,
    \new_[8511]_ , \new_[8512]_ , \new_[8513]_ , \new_[8514]_ ,
    \new_[8515]_ , \new_[8516]_ , \new_[8517]_ , \new_[8518]_ ,
    \new_[8519]_ , \new_[8520]_ , \new_[8521]_ , \new_[8522]_ ,
    \new_[8524]_ , \new_[8525]_ , \new_[8526]_ , \new_[8527]_ ,
    \new_[8528]_ , \new_[8529]_ , \new_[8530]_ , \new_[8531]_ ,
    \new_[8532]_ , \new_[8533]_ , \new_[8534]_ , \new_[8535]_ ,
    \new_[8536]_ , \new_[8537]_ , \new_[8538]_ , \new_[8539]_ ,
    \new_[8540]_ , \new_[8541]_ , \new_[8542]_ , \new_[8543]_ ,
    \new_[8544]_ , \new_[8545]_ , \new_[8546]_ , \new_[8547]_ ,
    \new_[8548]_ , \new_[8549]_ , \new_[8550]_ , \new_[8551]_ ,
    \new_[8552]_ , \new_[8553]_ , \new_[8554]_ , \new_[8555]_ ,
    \new_[8556]_ , \new_[8557]_ , \new_[8558]_ , \new_[8559]_ ,
    \new_[8560]_ , \new_[8561]_ , \new_[8562]_ , \new_[8563]_ ,
    \new_[8564]_ , \new_[8565]_ , \new_[8566]_ , \new_[8567]_ ,
    \new_[8568]_ , \new_[8569]_ , \new_[8570]_ , \new_[8571]_ ,
    \new_[8572]_ , \new_[8573]_ , \new_[8574]_ , \new_[8575]_ ,
    \new_[8576]_ , \new_[8577]_ , \new_[8578]_ , \new_[8579]_ ,
    \new_[8580]_ , \new_[8581]_ , \new_[8582]_ , \new_[8583]_ ,
    \new_[8584]_ , \new_[8585]_ , \new_[8586]_ , \new_[8587]_ ,
    \new_[8588]_ , \new_[8589]_ , \new_[8590]_ , \new_[8591]_ ,
    \new_[8592]_ , \new_[8593]_ , \new_[8594]_ , \new_[8595]_ ,
    \new_[8596]_ , \new_[8597]_ , \new_[8598]_ , \new_[8599]_ ,
    \new_[8600]_ , \new_[8601]_ , \new_[8602]_ , \new_[8603]_ ,
    \new_[8604]_ , \new_[8605]_ , \new_[8606]_ , \new_[8607]_ ,
    \new_[8608]_ , \new_[8609]_ , \new_[8610]_ , \new_[8611]_ ,
    \new_[8612]_ , \new_[8613]_ , \new_[8614]_ , \new_[8615]_ ,
    \new_[8616]_ , \new_[8617]_ , \new_[8618]_ , \new_[8619]_ ,
    \new_[8620]_ , \new_[8621]_ , \new_[8622]_ , \new_[8623]_ ,
    \new_[8624]_ , \new_[8625]_ , \new_[8626]_ , \new_[8627]_ ,
    \new_[8628]_ , \new_[8629]_ , \new_[8630]_ , \new_[8631]_ ,
    \new_[8632]_ , \new_[8633]_ , \new_[8635]_ , \new_[8636]_ ,
    \new_[8637]_ , \new_[8638]_ , \new_[8639]_ , \new_[8640]_ ,
    \new_[8641]_ , \new_[8642]_ , \new_[8643]_ , \new_[8644]_ ,
    \new_[8645]_ , \new_[8646]_ , \new_[8647]_ , \new_[8648]_ ,
    \new_[8649]_ , \new_[8650]_ , \new_[8651]_ , \new_[8652]_ ,
    \new_[8653]_ , \new_[8654]_ , \new_[8655]_ , \new_[8656]_ ,
    \new_[8657]_ , \new_[8658]_ , \new_[8659]_ , \new_[8660]_ ,
    \new_[8661]_ , \new_[8662]_ , \new_[8663]_ , \new_[8664]_ ,
    \new_[8665]_ , \new_[8666]_ , \new_[8667]_ , \new_[8668]_ ,
    \new_[8669]_ , \new_[8670]_ , \new_[8671]_ , \new_[8672]_ ,
    \new_[8673]_ , \new_[8674]_ , \new_[8675]_ , \new_[8676]_ ,
    \new_[8688]_ , \new_[8694]_ , \new_[8695]_ , \new_[8696]_ ,
    \new_[8697]_ , \new_[8698]_ , \new_[8699]_ , \new_[8700]_ ,
    \new_[8701]_ , \new_[8702]_ , \new_[8703]_ , \new_[8704]_ ,
    \new_[8705]_ , \new_[8706]_ , \new_[8707]_ , \new_[8708]_ ,
    \new_[8709]_ , \new_[8710]_ , \new_[8711]_ , \new_[8712]_ ,
    \new_[8713]_ , \new_[8714]_ , \new_[8717]_ , \new_[8718]_ ,
    \new_[8720]_ , \new_[8721]_ , \new_[8723]_ , \new_[8724]_ ,
    \new_[8725]_ , \new_[8726]_ , \new_[8727]_ , \new_[8728]_ ,
    \new_[8730]_ , \new_[8731]_ , \new_[8732]_ , \new_[8733]_ ,
    \new_[8734]_ , \new_[8735]_ , \new_[8737]_ , \new_[8738]_ ,
    \new_[8739]_ , \new_[8740]_ , \new_[8741]_ , \new_[8742]_ ,
    \new_[8743]_ , \new_[8744]_ , \new_[8745]_ , \new_[8746]_ ,
    \new_[8747]_ , \new_[8748]_ , \new_[8749]_ , \new_[8750]_ ,
    \new_[8751]_ , \new_[8752]_ , \new_[8753]_ , \new_[8754]_ ,
    \new_[8755]_ , \new_[8756]_ , \new_[8757]_ , \new_[8758]_ ,
    \new_[8759]_ , \new_[8760]_ , \new_[8761]_ , \new_[8762]_ ,
    \new_[8763]_ , \new_[8764]_ , \new_[8765]_ , \new_[8766]_ ,
    \new_[8767]_ , \new_[8768]_ , \new_[8769]_ , \new_[8770]_ ,
    \new_[8771]_ , \new_[8772]_ , \new_[8773]_ , \new_[8774]_ ,
    \new_[8775]_ , \new_[8776]_ , \new_[8777]_ , \new_[8778]_ ,
    \new_[8779]_ , \new_[8780]_ , \new_[8781]_ , \new_[8782]_ ,
    \new_[8783]_ , \new_[8784]_ , \new_[8785]_ , \new_[8786]_ ,
    \new_[8789]_ , \new_[8790]_ , \new_[8791]_ , \new_[8792]_ ,
    \new_[8794]_ , \new_[8795]_ , \new_[8796]_ , \new_[8797]_ ,
    \new_[8798]_ , \new_[8799]_ , \new_[8800]_ , \new_[8801]_ ,
    \new_[8802]_ , \new_[8803]_ , \new_[8804]_ , \new_[8805]_ ,
    \new_[8806]_ , \new_[8807]_ , \new_[8809]_ , \new_[8810]_ ,
    \new_[8812]_ , \new_[8813]_ , \new_[8816]_ , \new_[8817]_ ,
    \new_[8818]_ , \new_[8820]_ , \new_[8821]_ , \new_[8822]_ ,
    \new_[8824]_ , \new_[8828]_ , \new_[8829]_ , \new_[8830]_ ,
    \new_[8831]_ , \new_[8832]_ , \new_[8833]_ , \new_[8834]_ ,
    \new_[8835]_ , \new_[8836]_ , \new_[8837]_ , \new_[8838]_ ,
    \new_[8840]_ , \new_[8841]_ , \new_[8842]_ , \new_[8843]_ ,
    \new_[8844]_ , \new_[8845]_ , \new_[8847]_ , \new_[8848]_ ,
    \new_[8850]_ , \new_[8851]_ , \new_[8853]_ , \new_[8854]_ ,
    \new_[8855]_ , \new_[8856]_ , \new_[8857]_ , \new_[8858]_ ,
    \new_[8861]_ , \new_[8862]_ , \new_[8863]_ , \new_[8864]_ ,
    \new_[8866]_ , \new_[8867]_ , \new_[8868]_ , \new_[8869]_ ,
    \new_[8870]_ , \new_[8871]_ , \new_[8872]_ , \new_[8873]_ ,
    \new_[8874]_ , \new_[8875]_ , \new_[8876]_ , \new_[8877]_ ,
    \new_[8880]_ , \new_[8881]_ , \new_[8882]_ , \new_[8883]_ ,
    \new_[8884]_ , \new_[8885]_ , \new_[8887]_ , \new_[8888]_ ,
    \new_[8889]_ , \new_[8890]_ , \new_[8891]_ , \new_[8892]_ ,
    \new_[8893]_ , \new_[8894]_ , \new_[8895]_ , \new_[8896]_ ,
    \new_[8897]_ , \new_[8898]_ , \new_[8899]_ , \new_[8900]_ ,
    \new_[8901]_ , \new_[8902]_ , \new_[8903]_ , \new_[8904]_ ,
    \new_[8905]_ , \new_[8906]_ , \new_[8907]_ , \new_[8908]_ ,
    \new_[8909]_ , \new_[8910]_ , \new_[8912]_ , \new_[8913]_ ,
    \new_[8914]_ , \new_[8917]_ , \new_[8918]_ , \new_[8919]_ ,
    \new_[8920]_ , \new_[8921]_ , \new_[8922]_ , \new_[8923]_ ,
    \new_[8926]_ , \new_[8929]_ , \new_[8930]_ , \new_[8931]_ ,
    \new_[8939]_ , \new_[8940]_ , \new_[8943]_ , \new_[8945]_ ,
    \new_[8947]_ , \new_[8950]_ , \new_[8951]_ , \new_[8953]_ ,
    \new_[8955]_ , \new_[8956]_ , \new_[8957]_ , \new_[8958]_ ,
    \new_[8959]_ , \new_[8961]_ , \new_[8966]_ , \new_[8967]_ ,
    \new_[8969]_ , \new_[8970]_ , \new_[8971]_ , \new_[8972]_ ,
    \new_[8973]_ , \new_[8976]_ , \new_[8977]_ , \new_[8978]_ ,
    \new_[8979]_ , \new_[8980]_ , \new_[8981]_ , \new_[8982]_ ,
    \new_[8983]_ , \new_[8984]_ , \new_[8985]_ , \new_[8986]_ ,
    \new_[8987]_ , \new_[8988]_ , \new_[8989]_ , \new_[8990]_ ,
    \new_[8991]_ , \new_[8992]_ , \new_[8993]_ , \new_[8994]_ ,
    \new_[8995]_ , \new_[8996]_ , \new_[8997]_ , \new_[8998]_ ,
    \new_[8999]_ , \new_[9000]_ , \new_[9001]_ , \new_[9002]_ ,
    \new_[9003]_ , \new_[9004]_ , \new_[9005]_ , \new_[9007]_ ,
    \new_[9008]_ , \new_[9009]_ , \new_[9010]_ , \new_[9011]_ ,
    \new_[9012]_ , \new_[9013]_ , \new_[9014]_ , \new_[9015]_ ,
    \new_[9016]_ , \new_[9017]_ , \new_[9018]_ , \new_[9019]_ ,
    \new_[9020]_ , \new_[9021]_ , \new_[9022]_ , \new_[9023]_ ,
    \new_[9024]_ , \new_[9025]_ , \new_[9026]_ , \new_[9027]_ ,
    \new_[9028]_ , \new_[9029]_ , \new_[9030]_ , \new_[9031]_ ,
    \new_[9032]_ , \new_[9034]_ , \new_[9035]_ , \new_[9036]_ ,
    \new_[9037]_ , \new_[9040]_ , \new_[9041]_ , \new_[9042]_ ,
    \new_[9043]_ , \new_[9044]_ , \new_[9045]_ , \new_[9046]_ ,
    \new_[9047]_ , \new_[9048]_ , \new_[9049]_ , \new_[9050]_ ,
    \new_[9051]_ , \new_[9052]_ , \new_[9054]_ , \new_[9055]_ ,
    \new_[9056]_ , \new_[9057]_ , \new_[9058]_ , \new_[9059]_ ,
    \new_[9060]_ , \new_[9061]_ , \new_[9062]_ , \new_[9063]_ ,
    \new_[9064]_ , \new_[9065]_ , \new_[9066]_ , \new_[9067]_ ,
    \new_[9068]_ , \new_[9069]_ , \new_[9070]_ , \new_[9071]_ ,
    \new_[9072]_ , \new_[9073]_ , \new_[9074]_ , \new_[9075]_ ,
    \new_[9076]_ , \new_[9077]_ , \new_[9078]_ , \new_[9079]_ ,
    \new_[9080]_ , \new_[9081]_ , \new_[9082]_ , \new_[9083]_ ,
    \new_[9084]_ , \new_[9085]_ , \new_[9086]_ , \new_[9087]_ ,
    \new_[9088]_ , \new_[9089]_ , \new_[9090]_ , \new_[9091]_ ,
    \new_[9092]_ , \new_[9093]_ , \new_[9094]_ , \new_[9095]_ ,
    \new_[9096]_ , \new_[9097]_ , \new_[9098]_ , \new_[9099]_ ,
    \new_[9100]_ , \new_[9101]_ , \new_[9102]_ , \new_[9103]_ ,
    \new_[9104]_ , \new_[9106]_ , \new_[9107]_ , \new_[9108]_ ,
    \new_[9109]_ , \new_[9110]_ , \new_[9111]_ , \new_[9112]_ ,
    \new_[9113]_ , \new_[9114]_ , \new_[9115]_ , \new_[9116]_ ,
    \new_[9117]_ , \new_[9118]_ , \new_[9119]_ , \new_[9120]_ ,
    \new_[9121]_ , \new_[9122]_ , \new_[9123]_ , \new_[9124]_ ,
    \new_[9125]_ , \new_[9126]_ , \new_[9127]_ , \new_[9128]_ ,
    \new_[9129]_ , \new_[9130]_ , \new_[9131]_ , \new_[9132]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9137]_ , \new_[9138]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9143]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9146]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9150]_ , \new_[9151]_ , \new_[9152]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9163]_ , \new_[9164]_ ,
    \new_[9165]_ , \new_[9166]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9170]_ , \new_[9171]_ , \new_[9173]_ ,
    \new_[9175]_ , \new_[9176]_ , \new_[9177]_ , \new_[9178]_ ,
    \new_[9179]_ , \new_[9184]_ , \new_[9186]_ , \new_[9187]_ ,
    \new_[9188]_ , \new_[9190]_ , \new_[9191]_ , \new_[9192]_ ,
    \new_[9193]_ , \new_[9194]_ , \new_[9195]_ , \new_[9196]_ ,
    \new_[9198]_ , \new_[9199]_ , \new_[9201]_ , \new_[9202]_ ,
    \new_[9204]_ , \new_[9205]_ , \new_[9206]_ , \new_[9207]_ ,
    \new_[9208]_ , \new_[9209]_ , \new_[9210]_ , \new_[9211]_ ,
    \new_[9212]_ , \new_[9213]_ , \new_[9214]_ , \new_[9215]_ ,
    \new_[9216]_ , \new_[9217]_ , \new_[9218]_ , \new_[9219]_ ,
    \new_[9227]_ , \new_[9235]_ , \new_[9236]_ , \new_[9237]_ ,
    \new_[9238]_ , \new_[9239]_ , \new_[9240]_ , \new_[9241]_ ,
    \new_[9242]_ , \new_[9243]_ , \new_[9244]_ , \new_[9245]_ ,
    \new_[9246]_ , \new_[9247]_ , \new_[9248]_ , \new_[9249]_ ,
    \new_[9255]_ , \new_[9257]_ , \new_[9260]_ , \new_[9261]_ ,
    \new_[9262]_ , \new_[9263]_ , \new_[9265]_ , \new_[9266]_ ,
    \new_[9267]_ , \new_[9268]_ , \new_[9269]_ , \new_[9270]_ ,
    \new_[9272]_ , \new_[9273]_ , \new_[9274]_ , \new_[9275]_ ,
    \new_[9276]_ , \new_[9277]_ , \new_[9278]_ , \new_[9279]_ ,
    \new_[9280]_ , \new_[9281]_ , \new_[9282]_ , \new_[9284]_ ,
    \new_[9285]_ , \new_[9286]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9290]_ , \new_[9291]_ , \new_[9292]_ ,
    \new_[9293]_ , \new_[9294]_ , \new_[9295]_ , \new_[9296]_ ,
    \new_[9297]_ , \new_[9298]_ , \new_[9299]_ , \new_[9300]_ ,
    \new_[9302]_ , \new_[9303]_ , \new_[9304]_ , \new_[9305]_ ,
    \new_[9306]_ , \new_[9307]_ , \new_[9308]_ , \new_[9309]_ ,
    \new_[9311]_ , \new_[9312]_ , \new_[9314]_ , \new_[9315]_ ,
    \new_[9316]_ , \new_[9317]_ , \new_[9318]_ , \new_[9319]_ ,
    \new_[9320]_ , \new_[9321]_ , \new_[9322]_ , \new_[9323]_ ,
    \new_[9324]_ , \new_[9325]_ , \new_[9326]_ , \new_[9327]_ ,
    \new_[9328]_ , \new_[9329]_ , \new_[9330]_ , \new_[9331]_ ,
    \new_[9332]_ , \new_[9333]_ , \new_[9334]_ , \new_[9335]_ ,
    \new_[9336]_ , \new_[9337]_ , \new_[9338]_ , \new_[9339]_ ,
    \new_[9340]_ , \new_[9341]_ , \new_[9342]_ , \new_[9343]_ ,
    \new_[9344]_ , \new_[9345]_ , \new_[9346]_ , \new_[9347]_ ,
    \new_[9348]_ , \new_[9349]_ , \new_[9350]_ , \new_[9351]_ ,
    \new_[9353]_ , \new_[9354]_ , \new_[9355]_ , \new_[9357]_ ,
    \new_[9358]_ , \new_[9361]_ , \new_[9362]_ , \new_[9363]_ ,
    \new_[9364]_ , \new_[9365]_ , \new_[9366]_ , \new_[9367]_ ,
    \new_[9369]_ , \new_[9370]_ , \new_[9371]_ , \new_[9372]_ ,
    \new_[9373]_ , \new_[9374]_ , \new_[9375]_ , \new_[9376]_ ,
    \new_[9378]_ , \new_[9379]_ , \new_[9380]_ , \new_[9382]_ ,
    \new_[9383]_ , \new_[9384]_ , \new_[9385]_ , \new_[9387]_ ,
    \new_[9388]_ , \new_[9389]_ , \new_[9390]_ , \new_[9391]_ ,
    \new_[9392]_ , \new_[9393]_ , \new_[9394]_ , \new_[9396]_ ,
    \new_[9397]_ , \new_[9398]_ , \new_[9399]_ , \new_[9400]_ ,
    \new_[9401]_ , \new_[9402]_ , \new_[9403]_ , \new_[9404]_ ,
    \new_[9405]_ , \new_[9406]_ , \new_[9407]_ , \new_[9408]_ ,
    \new_[9409]_ , \new_[9410]_ , \new_[9411]_ , \new_[9412]_ ,
    \new_[9413]_ , \new_[9414]_ , \new_[9415]_ , \new_[9416]_ ,
    \new_[9417]_ , \new_[9418]_ , \new_[9419]_ , \new_[9421]_ ,
    \new_[9422]_ , \new_[9423]_ , \new_[9424]_ , \new_[9425]_ ,
    \new_[9426]_ , \new_[9427]_ , \new_[9428]_ , \new_[9429]_ ,
    \new_[9430]_ , \new_[9431]_ , \new_[9432]_ , \new_[9433]_ ,
    \new_[9434]_ , \new_[9435]_ , \new_[9436]_ , \new_[9437]_ ,
    \new_[9438]_ , \new_[9439]_ , \new_[9440]_ , \new_[9441]_ ,
    \new_[9442]_ , \new_[9443]_ , \new_[9444]_ , \new_[9445]_ ,
    \new_[9446]_ , \new_[9447]_ , \new_[9448]_ , \new_[9449]_ ,
    \new_[9450]_ , \new_[9451]_ , \new_[9452]_ , \new_[9453]_ ,
    \new_[9454]_ , \new_[9455]_ , \new_[9456]_ , \new_[9457]_ ,
    \new_[9458]_ , \new_[9459]_ , \new_[9460]_ , \new_[9461]_ ,
    \new_[9462]_ , \new_[9463]_ , \new_[9464]_ , \new_[9465]_ ,
    \new_[9466]_ , \new_[9467]_ , \new_[9468]_ , \new_[9469]_ ,
    \new_[9470]_ , \new_[9471]_ , \new_[9472]_ , \new_[9473]_ ,
    \new_[9474]_ , \new_[9475]_ , \new_[9479]_ , \new_[9489]_ ,
    \new_[9493]_ , \new_[9494]_ , \new_[9495]_ , \new_[9496]_ ,
    \new_[9497]_ , \new_[9498]_ , \new_[9499]_ , \new_[9500]_ ,
    \new_[9501]_ , \new_[9502]_ , \new_[9503]_ , \new_[9504]_ ,
    \new_[9505]_ , \new_[9506]_ , \new_[9507]_ , \new_[9508]_ ,
    \new_[9509]_ , \new_[9510]_ , \new_[9511]_ , \new_[9512]_ ,
    \new_[9513]_ , \new_[9514]_ , \new_[9515]_ , \new_[9516]_ ,
    \new_[9517]_ , \new_[9518]_ , \new_[9519]_ , \new_[9520]_ ,
    \new_[9521]_ , \new_[9522]_ , \new_[9523]_ , \new_[9524]_ ,
    \new_[9525]_ , \new_[9526]_ , \new_[9527]_ , \new_[9528]_ ,
    \new_[9529]_ , \new_[9530]_ , \new_[9531]_ , \new_[9532]_ ,
    \new_[9533]_ , \new_[9534]_ , \new_[9535]_ , \new_[9536]_ ,
    \new_[9537]_ , \new_[9538]_ , \new_[9539]_ , \new_[9540]_ ,
    \new_[9541]_ , \new_[9542]_ , \new_[9543]_ , \new_[9544]_ ,
    \new_[9545]_ , \new_[9546]_ , \new_[9547]_ , \new_[9548]_ ,
    \new_[9549]_ , \new_[9550]_ , \new_[9551]_ , \new_[9552]_ ,
    \new_[9553]_ , \new_[9554]_ , \new_[9555]_ , \new_[9556]_ ,
    \new_[9557]_ , \new_[9559]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9562]_ , \new_[9563]_ , \new_[9564]_ , \new_[9565]_ ,
    \new_[9566]_ , \new_[9567]_ , \new_[9568]_ , \new_[9569]_ ,
    \new_[9570]_ , \new_[9571]_ , \new_[9573]_ , \new_[9574]_ ,
    \new_[9575]_ , \new_[9576]_ , \new_[9577]_ , \new_[9578]_ ,
    \new_[9579]_ , \new_[9580]_ , \new_[9581]_ , \new_[9582]_ ,
    \new_[9583]_ , \new_[9584]_ , \new_[9585]_ , \new_[9586]_ ,
    \new_[9587]_ , \new_[9588]_ , \new_[9589]_ , \new_[9590]_ ,
    \new_[9591]_ , \new_[9592]_ , \new_[9593]_ , \new_[9594]_ ,
    \new_[9595]_ , \new_[9596]_ , \new_[9597]_ , \new_[9598]_ ,
    \new_[9599]_ , \new_[9600]_ , \new_[9601]_ , \new_[9602]_ ,
    \new_[9603]_ , \new_[9604]_ , \new_[9605]_ , \new_[9606]_ ,
    \new_[9607]_ , \new_[9608]_ , \new_[9609]_ , \new_[9610]_ ,
    \new_[9611]_ , \new_[9612]_ , \new_[9613]_ , \new_[9614]_ ,
    \new_[9615]_ , \new_[9616]_ , \new_[9617]_ , \new_[9618]_ ,
    \new_[9619]_ , \new_[9620]_ , \new_[9621]_ , \new_[9622]_ ,
    \new_[9623]_ , \new_[9624]_ , \new_[9625]_ , \new_[9626]_ ,
    \new_[9627]_ , \new_[9628]_ , \new_[9629]_ , \new_[9630]_ ,
    \new_[9631]_ , \new_[9632]_ , \new_[9633]_ , \new_[9634]_ ,
    \new_[9635]_ , \new_[9636]_ , \new_[9637]_ , \new_[9638]_ ,
    \new_[9639]_ , \new_[9640]_ , \new_[9641]_ , \new_[9642]_ ,
    \new_[9643]_ , \new_[9644]_ , \new_[9645]_ , \new_[9646]_ ,
    \new_[9647]_ , \new_[9648]_ , \new_[9649]_ , \new_[9650]_ ,
    \new_[9651]_ , \new_[9652]_ , \new_[9653]_ , \new_[9654]_ ,
    \new_[9655]_ , \new_[9656]_ , \new_[9657]_ , \new_[9658]_ ,
    \new_[9659]_ , \new_[9660]_ , \new_[9661]_ , \new_[9663]_ ,
    \new_[9664]_ , \new_[9665]_ , \new_[9666]_ , \new_[9667]_ ,
    \new_[9668]_ , \new_[9669]_ , \new_[9670]_ , \new_[9673]_ ,
    \new_[9674]_ , \new_[9675]_ , \new_[9677]_ , \new_[9678]_ ,
    \new_[9680]_ , \new_[9681]_ , \new_[9682]_ , \new_[9684]_ ,
    \new_[9685]_ , \new_[9687]_ , \new_[9688]_ , \new_[9690]_ ,
    \new_[9691]_ , \new_[9692]_ , \new_[9693]_ , \new_[9694]_ ,
    \new_[9695]_ , \new_[9698]_ , \new_[9701]_ , \new_[9706]_ ,
    \new_[9707]_ , \new_[9708]_ , \new_[9709]_ , \new_[9710]_ ,
    \new_[9711]_ , \new_[9712]_ , \new_[9713]_ , \new_[9714]_ ,
    \new_[9715]_ , \new_[9716]_ , \new_[9717]_ , \new_[9718]_ ,
    \new_[9720]_ , \new_[9721]_ , \new_[9722]_ , \new_[9723]_ ,
    \new_[9724]_ , \new_[9725]_ , \new_[9726]_ , \new_[9727]_ ,
    \new_[9728]_ , \new_[9730]_ , \new_[9732]_ , \new_[9733]_ ,
    \new_[9734]_ , \new_[9735]_ , \new_[9736]_ , \new_[9737]_ ,
    \new_[9738]_ , \new_[9739]_ , \new_[9741]_ , \new_[9742]_ ,
    \new_[9743]_ , \new_[9744]_ , \new_[9745]_ , \new_[9746]_ ,
    \new_[9747]_ , \new_[9748]_ , \new_[9749]_ , \new_[9750]_ ,
    \new_[9751]_ , \new_[9752]_ , \new_[9754]_ , \new_[9755]_ ,
    \new_[9756]_ , \new_[9757]_ , \new_[9758]_ , \new_[9759]_ ,
    \new_[9760]_ , \new_[9761]_ , \new_[9762]_ , \new_[9763]_ ,
    \new_[9764]_ , \new_[9765]_ , \new_[9766]_ , \new_[9767]_ ,
    \new_[9768]_ , \new_[9769]_ , \new_[9770]_ , \new_[9771]_ ,
    \new_[9772]_ , \new_[9773]_ , \new_[9774]_ , \new_[9775]_ ,
    \new_[9776]_ , \new_[9777]_ , \new_[9778]_ , \new_[9779]_ ,
    \new_[9780]_ , \new_[9781]_ , \new_[9782]_ , \new_[9783]_ ,
    \new_[9784]_ , \new_[9785]_ , \new_[9786]_ , \new_[9787]_ ,
    \new_[9788]_ , \new_[9789]_ , \new_[9790]_ , \new_[9791]_ ,
    \new_[9792]_ , \new_[9793]_ , \new_[9794]_ , \new_[9795]_ ,
    \new_[9796]_ , \new_[9797]_ , \new_[9798]_ , \new_[9799]_ ,
    \new_[9800]_ , \new_[9801]_ , \new_[9802]_ , \new_[9803]_ ,
    \new_[9804]_ , \new_[9805]_ , \new_[9806]_ , \new_[9807]_ ,
    \new_[9808]_ , \new_[9809]_ , \new_[9810]_ , \new_[9811]_ ,
    \new_[9812]_ , \new_[9813]_ , \new_[9814]_ , \new_[9815]_ ,
    \new_[9816]_ , \new_[9817]_ , \new_[9818]_ , \new_[9819]_ ,
    \new_[9820]_ , \new_[9821]_ , \new_[9822]_ , \new_[9823]_ ,
    \new_[9824]_ , \new_[9835]_ , \new_[9836]_ , \new_[9837]_ ,
    \new_[9838]_ , \new_[9839]_ , \new_[9840]_ , \new_[9841]_ ,
    \new_[9842]_ , \new_[9843]_ , \new_[9844]_ , \new_[9845]_ ,
    \new_[9846]_ , \new_[9847]_ , \new_[9848]_ , \new_[9849]_ ,
    \new_[9850]_ , \new_[9851]_ , \new_[9852]_ , \new_[9853]_ ,
    \new_[9854]_ , \new_[9855]_ , \new_[9856]_ , \new_[9857]_ ,
    \new_[9858]_ , \new_[9859]_ , \new_[9860]_ , \new_[9861]_ ,
    \new_[9862]_ , \new_[9863]_ , \new_[9864]_ , \new_[9865]_ ,
    \new_[9866]_ , \new_[9867]_ , \new_[9868]_ , \new_[9869]_ ,
    \new_[9870]_ , \new_[9871]_ , \new_[9872]_ , \new_[9873]_ ,
    \new_[9874]_ , \new_[9875]_ , \new_[9876]_ , \new_[9877]_ ,
    \new_[9878]_ , \new_[9879]_ , \new_[9880]_ , \new_[9881]_ ,
    \new_[9882]_ , \new_[9883]_ , \new_[9884]_ , \new_[9885]_ ,
    \new_[9886]_ , \new_[9887]_ , \new_[9889]_ , \new_[9890]_ ,
    \new_[9891]_ , \new_[9892]_ , \new_[9893]_ , \new_[9894]_ ,
    \new_[9895]_ , \new_[9896]_ , \new_[9898]_ , \new_[9899]_ ,
    \new_[9900]_ , \new_[9901]_ , \new_[9902]_ , \new_[9903]_ ,
    \new_[9904]_ , \new_[9905]_ , \new_[9906]_ , \new_[9907]_ ,
    \new_[9908]_ , \new_[9909]_ , \new_[9910]_ , \new_[9911]_ ,
    \new_[9912]_ , \new_[9913]_ , \new_[9914]_ , \new_[9915]_ ,
    \new_[9916]_ , \new_[9918]_ , \new_[9919]_ , \new_[9920]_ ,
    \new_[9921]_ , \new_[9922]_ , \new_[9924]_ , \new_[9925]_ ,
    \new_[9926]_ , \new_[9927]_ , \new_[9929]_ , \new_[9930]_ ,
    \new_[9932]_ , \new_[9933]_ , \new_[9934]_ , \new_[9935]_ ,
    \new_[9936]_ , \new_[9937]_ , \new_[9938]_ , \new_[9939]_ ,
    \new_[9940]_ , \new_[9941]_ , \new_[9942]_ , \new_[9943]_ ,
    \new_[9944]_ , \new_[9946]_ , \new_[9947]_ , \new_[9949]_ ,
    \new_[9950]_ , \new_[9951]_ , \new_[9953]_ , \new_[9954]_ ,
    \new_[9955]_ , \new_[9956]_ , \new_[9957]_ , \new_[9958]_ ,
    \new_[9959]_ , \new_[9960]_ , \new_[9961]_ , \new_[9962]_ ,
    \new_[9963]_ , \new_[9965]_ , \new_[9966]_ , \new_[9967]_ ,
    \new_[9968]_ , \new_[9969]_ , \new_[9970]_ , \new_[9971]_ ,
    \new_[9972]_ , \new_[9973]_ , \new_[9975]_ , \new_[9978]_ ,
    \new_[9979]_ , \new_[9980]_ , \new_[9981]_ , \new_[9982]_ ,
    \new_[9983]_ , \new_[9984]_ , \new_[9985]_ , \new_[9986]_ ,
    \new_[9987]_ , \new_[9988]_ , \new_[9989]_ , \new_[9990]_ ,
    \new_[9991]_ , \new_[9992]_ , \new_[9993]_ , \new_[9994]_ ,
    \new_[9995]_ , \new_[9996]_ , \new_[9997]_ , \new_[9998]_ ,
    \new_[9999]_ , \new_[10000]_ , \new_[10001]_ , \new_[10002]_ ,
    \new_[10003]_ , \new_[10004]_ , \new_[10005]_ , \new_[10006]_ ,
    \new_[10007]_ , \new_[10008]_ , \new_[10009]_ , \new_[10010]_ ,
    \new_[10011]_ , \new_[10012]_ , \new_[10013]_ , \new_[10014]_ ,
    \new_[10015]_ , \new_[10016]_ , \new_[10017]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10020]_ , \new_[10021]_ , \new_[10022]_ ,
    \new_[10023]_ , \new_[10024]_ , \new_[10025]_ , \new_[10026]_ ,
    \new_[10027]_ , \new_[10028]_ , \new_[10029]_ , \new_[10030]_ ,
    \new_[10031]_ , \new_[10032]_ , \new_[10033]_ , \new_[10034]_ ,
    \new_[10035]_ , \new_[10036]_ , \new_[10037]_ , \new_[10038]_ ,
    \new_[10039]_ , \new_[10040]_ , \new_[10041]_ , \new_[10042]_ ,
    \new_[10043]_ , \new_[10044]_ , \new_[10045]_ , \new_[10046]_ ,
    \new_[10047]_ , \new_[10048]_ , \new_[10049]_ , \new_[10050]_ ,
    \new_[10051]_ , \new_[10052]_ , \new_[10053]_ , \new_[10054]_ ,
    \new_[10055]_ , \new_[10056]_ , \new_[10057]_ , \new_[10058]_ ,
    \new_[10059]_ , \new_[10060]_ , \new_[10061]_ , \new_[10062]_ ,
    \new_[10063]_ , \new_[10064]_ , \new_[10065]_ , \new_[10066]_ ,
    \new_[10067]_ , \new_[10068]_ , \new_[10069]_ , \new_[10070]_ ,
    \new_[10071]_ , \new_[10072]_ , \new_[10073]_ , \new_[10074]_ ,
    \new_[10075]_ , \new_[10076]_ , \new_[10077]_ , \new_[10078]_ ,
    \new_[10079]_ , \new_[10080]_ , \new_[10081]_ , \new_[10082]_ ,
    \new_[10083]_ , \new_[10084]_ , \new_[10085]_ , \new_[10086]_ ,
    \new_[10087]_ , \new_[10088]_ , \new_[10089]_ , \new_[10090]_ ,
    \new_[10091]_ , \new_[10092]_ , \new_[10093]_ , \new_[10094]_ ,
    \new_[10095]_ , \new_[10096]_ , \new_[10097]_ , \new_[10098]_ ,
    \new_[10099]_ , \new_[10100]_ , \new_[10101]_ , \new_[10102]_ ,
    \new_[10103]_ , \new_[10104]_ , \new_[10105]_ , \new_[10106]_ ,
    \new_[10107]_ , \new_[10108]_ , \new_[10109]_ , \new_[10110]_ ,
    \new_[10111]_ , \new_[10112]_ , \new_[10113]_ , \new_[10114]_ ,
    \new_[10115]_ , \new_[10116]_ , \new_[10118]_ , \new_[10119]_ ,
    \new_[10120]_ , \new_[10121]_ , \new_[10122]_ , \new_[10123]_ ,
    \new_[10124]_ , \new_[10125]_ , \new_[10126]_ , \new_[10127]_ ,
    \new_[10128]_ , \new_[10129]_ , \new_[10130]_ , \new_[10131]_ ,
    \new_[10132]_ , \new_[10133]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10136]_ , \new_[10137]_ , \new_[10138]_ , \new_[10139]_ ,
    \new_[10140]_ , \new_[10141]_ , \new_[10142]_ , \new_[10143]_ ,
    \new_[10144]_ , \new_[10145]_ , \new_[10146]_ , \new_[10147]_ ,
    \new_[10148]_ , \new_[10149]_ , \new_[10150]_ , \new_[10151]_ ,
    \new_[10152]_ , \new_[10153]_ , \new_[10154]_ , \new_[10155]_ ,
    \new_[10156]_ , \new_[10157]_ , \new_[10158]_ , \new_[10159]_ ,
    \new_[10160]_ , \new_[10161]_ , \new_[10162]_ , \new_[10163]_ ,
    \new_[10164]_ , \new_[10165]_ , \new_[10166]_ , \new_[10167]_ ,
    \new_[10168]_ , \new_[10169]_ , \new_[10170]_ , \new_[10171]_ ,
    \new_[10172]_ , \new_[10173]_ , \new_[10174]_ , \new_[10175]_ ,
    \new_[10176]_ , \new_[10177]_ , \new_[10178]_ , \new_[10179]_ ,
    \new_[10180]_ , \new_[10181]_ , \new_[10182]_ , \new_[10183]_ ,
    \new_[10184]_ , \new_[10185]_ , \new_[10186]_ , \new_[10187]_ ,
    \new_[10188]_ , \new_[10189]_ , \new_[10190]_ , \new_[10191]_ ,
    \new_[10192]_ , \new_[10193]_ , \new_[10194]_ , \new_[10195]_ ,
    \new_[10196]_ , \new_[10197]_ , \new_[10198]_ , \new_[10199]_ ,
    \new_[10200]_ , \new_[10201]_ , \new_[10202]_ , \new_[10203]_ ,
    \new_[10204]_ , \new_[10205]_ , \new_[10206]_ , \new_[10207]_ ,
    \new_[10208]_ , \new_[10209]_ , \new_[10210]_ , \new_[10211]_ ,
    \new_[10212]_ , \new_[10213]_ , \new_[10214]_ , \new_[10215]_ ,
    \new_[10216]_ , \new_[10217]_ , \new_[10218]_ , \new_[10219]_ ,
    \new_[10221]_ , \new_[10222]_ , \new_[10223]_ , \new_[10224]_ ,
    \new_[10225]_ , \new_[10226]_ , \new_[10227]_ , \new_[10228]_ ,
    \new_[10229]_ , \new_[10230]_ , \new_[10231]_ , \new_[10232]_ ,
    \new_[10233]_ , \new_[10234]_ , \new_[10235]_ , \new_[10236]_ ,
    \new_[10237]_ , \new_[10238]_ , \new_[10239]_ , \new_[10240]_ ,
    \new_[10242]_ , \new_[10243]_ , \new_[10244]_ , \new_[10245]_ ,
    \new_[10246]_ , \new_[10247]_ , \new_[10248]_ , \new_[10249]_ ,
    \new_[10250]_ , \new_[10251]_ , \new_[10252]_ , \new_[10253]_ ,
    \new_[10254]_ , \new_[10255]_ , \new_[10256]_ , \new_[10257]_ ,
    \new_[10258]_ , \new_[10259]_ , \new_[10260]_ , \new_[10261]_ ,
    \new_[10262]_ , \new_[10263]_ , \new_[10264]_ , \new_[10265]_ ,
    \new_[10266]_ , \new_[10267]_ , \new_[10268]_ , \new_[10269]_ ,
    \new_[10270]_ , \new_[10271]_ , \new_[10272]_ , \new_[10273]_ ,
    \new_[10274]_ , \new_[10275]_ , \new_[10276]_ , \new_[10277]_ ,
    \new_[10278]_ , \new_[10279]_ , \new_[10280]_ , \new_[10281]_ ,
    \new_[10282]_ , \new_[10283]_ , \new_[10284]_ , \new_[10285]_ ,
    \new_[10286]_ , \new_[10287]_ , \new_[10288]_ , \new_[10289]_ ,
    \new_[10291]_ , \new_[10293]_ , \new_[10294]_ , \new_[10295]_ ,
    \new_[10296]_ , \new_[10297]_ , \new_[10298]_ , \new_[10299]_ ,
    \new_[10300]_ , \new_[10301]_ , \new_[10302]_ , \new_[10303]_ ,
    \new_[10304]_ , \new_[10305]_ , \new_[10306]_ , \new_[10307]_ ,
    \new_[10308]_ , \new_[10309]_ , \new_[10310]_ , \new_[10311]_ ,
    \new_[10313]_ , \new_[10314]_ , \new_[10315]_ , \new_[10316]_ ,
    \new_[10317]_ , \new_[10318]_ , \new_[10319]_ , \new_[10320]_ ,
    \new_[10321]_ , \new_[10322]_ , \new_[10323]_ , \new_[10324]_ ,
    \new_[10325]_ , \new_[10326]_ , \new_[10327]_ , \new_[10328]_ ,
    \new_[10329]_ , \new_[10330]_ , \new_[10331]_ , \new_[10332]_ ,
    \new_[10333]_ , \new_[10334]_ , \new_[10335]_ , \new_[10336]_ ,
    \new_[10337]_ , \new_[10338]_ , \new_[10339]_ , \new_[10340]_ ,
    \new_[10341]_ , \new_[10342]_ , \new_[10343]_ , \new_[10344]_ ,
    \new_[10345]_ , \new_[10346]_ , \new_[10347]_ , \new_[10348]_ ,
    \new_[10349]_ , \new_[10350]_ , \new_[10351]_ , \new_[10352]_ ,
    \new_[10353]_ , \new_[10354]_ , \new_[10355]_ , \new_[10356]_ ,
    \new_[10357]_ , \new_[10358]_ , \new_[10359]_ , \new_[10360]_ ,
    \new_[10361]_ , \new_[10362]_ , \new_[10363]_ , \new_[10364]_ ,
    \new_[10365]_ , \new_[10366]_ , \new_[10367]_ , \new_[10368]_ ,
    \new_[10369]_ , \new_[10370]_ , \new_[10371]_ , \new_[10372]_ ,
    \new_[10373]_ , \new_[10374]_ , \new_[10375]_ , \new_[10376]_ ,
    \new_[10377]_ , \new_[10378]_ , \new_[10379]_ , \new_[10380]_ ,
    \new_[10381]_ , \new_[10382]_ , \new_[10383]_ , \new_[10384]_ ,
    \new_[10385]_ , \new_[10386]_ , \new_[10387]_ , \new_[10388]_ ,
    \new_[10389]_ , \new_[10390]_ , \new_[10391]_ , \new_[10392]_ ,
    \new_[10393]_ , \new_[10394]_ , \new_[10395]_ , \new_[10396]_ ,
    \new_[10397]_ , \new_[10398]_ , \new_[10399]_ , \new_[10400]_ ,
    \new_[10401]_ , \new_[10402]_ , \new_[10403]_ , \new_[10404]_ ,
    \new_[10405]_ , \new_[10406]_ , \new_[10407]_ , \new_[10408]_ ,
    \new_[10409]_ , \new_[10410]_ , \new_[10411]_ , \new_[10412]_ ,
    \new_[10413]_ , \new_[10414]_ , \new_[10415]_ , \new_[10416]_ ,
    \new_[10417]_ , \new_[10418]_ , \new_[10419]_ , \new_[10420]_ ,
    \new_[10421]_ , \new_[10422]_ , \new_[10423]_ , \new_[10424]_ ,
    \new_[10425]_ , \new_[10426]_ , \new_[10427]_ , \new_[10428]_ ,
    \new_[10429]_ , \new_[10430]_ , \new_[10431]_ , \new_[10432]_ ,
    \new_[10433]_ , \new_[10434]_ , \new_[10435]_ , \new_[10436]_ ,
    \new_[10437]_ , \new_[10438]_ , \new_[10439]_ , \new_[10440]_ ,
    \new_[10441]_ , \new_[10442]_ , \new_[10443]_ , \new_[10444]_ ,
    \new_[10445]_ , \new_[10446]_ , \new_[10447]_ , \new_[10448]_ ,
    \new_[10449]_ , \new_[10450]_ , \new_[10451]_ , \new_[10452]_ ,
    \new_[10453]_ , \new_[10454]_ , \new_[10455]_ , \new_[10456]_ ,
    \new_[10457]_ , \new_[10458]_ , \new_[10459]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10462]_ , \new_[10463]_ , \new_[10464]_ ,
    \new_[10465]_ , \new_[10466]_ , \new_[10467]_ , \new_[10468]_ ,
    \new_[10469]_ , \new_[10470]_ , \new_[10471]_ , \new_[10472]_ ,
    \new_[10473]_ , \new_[10474]_ , \new_[10475]_ , \new_[10476]_ ,
    \new_[10477]_ , \new_[10478]_ , \new_[10479]_ , \new_[10480]_ ,
    \new_[10481]_ , \new_[10482]_ , \new_[10483]_ , \new_[10484]_ ,
    \new_[10485]_ , \new_[10486]_ , \new_[10487]_ , \new_[10488]_ ,
    \new_[10489]_ , \new_[10490]_ , \new_[10491]_ , \new_[10492]_ ,
    \new_[10493]_ , \new_[10494]_ , \new_[10495]_ , \new_[10496]_ ,
    \new_[10497]_ , \new_[10498]_ , \new_[10499]_ , \new_[10500]_ ,
    \new_[10501]_ , \new_[10502]_ , \new_[10503]_ , \new_[10504]_ ,
    \new_[10505]_ , \new_[10506]_ , \new_[10507]_ , \new_[10508]_ ,
    \new_[10509]_ , \new_[10510]_ , \new_[10511]_ , \new_[10512]_ ,
    \new_[10513]_ , \new_[10514]_ , \new_[10515]_ , \new_[10516]_ ,
    \new_[10517]_ , \new_[10518]_ , \new_[10519]_ , \new_[10520]_ ,
    \new_[10521]_ , \new_[10522]_ , \new_[10523]_ , \new_[10524]_ ,
    \new_[10525]_ , \new_[10526]_ , \new_[10528]_ , \new_[10529]_ ,
    \new_[10531]_ , \new_[10532]_ , \new_[10533]_ , \new_[10534]_ ,
    \new_[10535]_ , \new_[10536]_ , \new_[10537]_ , \new_[10538]_ ,
    \new_[10540]_ , \new_[10542]_ , \new_[10543]_ , \new_[10545]_ ,
    \new_[10549]_ , \new_[10550]_ , \new_[10551]_ , \new_[10552]_ ,
    \new_[10553]_ , \new_[10554]_ , \new_[10555]_ , \new_[10556]_ ,
    \new_[10558]_ , \new_[10559]_ , \new_[10560]_ , \new_[10561]_ ,
    \new_[10562]_ , \new_[10563]_ , \new_[10564]_ , \new_[10567]_ ,
    \new_[10568]_ , \new_[10570]_ , \new_[10571]_ , \new_[10572]_ ,
    \new_[10573]_ , \new_[10574]_ , \new_[10575]_ , \new_[10576]_ ,
    \new_[10577]_ , \new_[10578]_ , \new_[10579]_ , \new_[10582]_ ,
    \new_[10583]_ , \new_[10584]_ , \new_[10585]_ , \new_[10587]_ ,
    \new_[10588]_ , \new_[10590]_ , \new_[10591]_ , \new_[10592]_ ,
    \new_[10593]_ , \new_[10594]_ , \new_[10595]_ , \new_[10597]_ ,
    \new_[10598]_ , \new_[10599]_ , \new_[10600]_ , \new_[10601]_ ,
    \new_[10602]_ , \new_[10604]_ , \new_[10605]_ , \new_[10608]_ ,
    \new_[10610]_ , \new_[10611]_ , \new_[10612]_ , \new_[10613]_ ,
    \new_[10614]_ , \new_[10615]_ , \new_[10616]_ , \new_[10617]_ ,
    \new_[10618]_ , \new_[10619]_ , \new_[10620]_ , \new_[10621]_ ,
    \new_[10622]_ , \new_[10623]_ , \new_[10624]_ , \new_[10625]_ ,
    \new_[10626]_ , \new_[10628]_ , \new_[10629]_ , \new_[10631]_ ,
    \new_[10634]_ , \new_[10635]_ , \new_[10636]_ , \new_[10638]_ ,
    \new_[10639]_ , \new_[10640]_ , \new_[10641]_ , \new_[10642]_ ,
    \new_[10643]_ , \new_[10644]_ , \new_[10645]_ , \new_[10646]_ ,
    \new_[10647]_ , \new_[10648]_ , \new_[10649]_ , \new_[10650]_ ,
    \new_[10651]_ , \new_[10652]_ , \new_[10653]_ , \new_[10654]_ ,
    \new_[10655]_ , \new_[10656]_ , \new_[10657]_ , \new_[10658]_ ,
    \new_[10662]_ , \new_[10663]_ , \new_[10665]_ , \new_[10666]_ ,
    \new_[10667]_ , \new_[10669]_ , \new_[10670]_ , \new_[10671]_ ,
    \new_[10672]_ , \new_[10673]_ , \new_[10674]_ , \new_[10676]_ ,
    \new_[10677]_ , \new_[10678]_ , \new_[10679]_ , \new_[10680]_ ,
    \new_[10681]_ , \new_[10682]_ , \new_[10683]_ , \new_[10684]_ ,
    \new_[10685]_ , \new_[10686]_ , \new_[10687]_ , \new_[10689]_ ,
    \new_[10690]_ , \new_[10691]_ , \new_[10692]_ , \new_[10693]_ ,
    \new_[10694]_ , \new_[10695]_ , \new_[10696]_ , \new_[10697]_ ,
    \new_[10698]_ , \new_[10699]_ , \new_[10700]_ , \new_[10701]_ ,
    \new_[10703]_ , \new_[10704]_ , \new_[10705]_ , \new_[10708]_ ,
    \new_[10709]_ , \new_[10710]_ , \new_[10711]_ , \new_[10712]_ ,
    \new_[10713]_ , \new_[10714]_ , \new_[10715]_ , \new_[10719]_ ,
    \new_[10720]_ , \new_[10721]_ , \new_[10722]_ , \new_[10723]_ ,
    \new_[10724]_ , \new_[10725]_ , \new_[10727]_ , \new_[10728]_ ,
    \new_[10729]_ , \new_[10731]_ , \new_[10733]_ , \new_[10734]_ ,
    \new_[10735]_ , \new_[10736]_ , \new_[10737]_ , \new_[10738]_ ,
    \new_[10739]_ , \new_[10740]_ , \new_[10741]_ , \new_[10742]_ ,
    \new_[10743]_ , \new_[10745]_ , \new_[10746]_ , \new_[10747]_ ,
    \new_[10748]_ , \new_[10749]_ , \new_[10750]_ , \new_[10751]_ ,
    \new_[10752]_ , \new_[10753]_ , \new_[10754]_ , \new_[10757]_ ,
    \new_[10758]_ , \new_[10759]_ , \new_[10760]_ , \new_[10761]_ ,
    \new_[10762]_ , \new_[10763]_ , \new_[10764]_ , \new_[10767]_ ,
    \new_[10768]_ , \new_[10769]_ , \new_[10771]_ , \new_[10772]_ ,
    \new_[10773]_ , \new_[10775]_ , \new_[10776]_ , \new_[10779]_ ,
    \new_[10780]_ , \new_[10781]_ , \new_[10782]_ , \new_[10783]_ ,
    \new_[10784]_ , \new_[10785]_ , \new_[10786]_ , \new_[10787]_ ,
    \new_[10788]_ , \new_[10792]_ , \new_[10793]_ , \new_[10794]_ ,
    \new_[10795]_ , \new_[10796]_ , \new_[10797]_ , \new_[10799]_ ,
    \new_[10800]_ , \new_[10801]_ , \new_[10802]_ , \new_[10803]_ ,
    \new_[10804]_ , \new_[10805]_ , \new_[10806]_ , \new_[10807]_ ,
    \new_[10808]_ , \new_[10809]_ , \new_[10810]_ , \new_[10811]_ ,
    \new_[10813]_ , \new_[10814]_ , \new_[10815]_ , \new_[10816]_ ,
    \new_[10817]_ , \new_[10818]_ , \new_[10819]_ , \new_[10820]_ ,
    \new_[10821]_ , \new_[10822]_ , \new_[10823]_ , \new_[10824]_ ,
    \new_[10825]_ , \new_[10826]_ , \new_[10827]_ , \new_[10828]_ ,
    \new_[10829]_ , \new_[10830]_ , \new_[10831]_ , \new_[10832]_ ,
    \new_[10833]_ , \new_[10834]_ , \new_[10835]_ , \new_[10836]_ ,
    \new_[10837]_ , \new_[10838]_ , \new_[10839]_ , \new_[10840]_ ,
    \new_[10841]_ , \new_[10842]_ , \new_[10843]_ , \new_[10844]_ ,
    \new_[10845]_ , \new_[10846]_ , \new_[10847]_ , \new_[10848]_ ,
    \new_[10849]_ , \new_[10851]_ , \new_[10852]_ , \new_[10853]_ ,
    \new_[10854]_ , \new_[10855]_ , \new_[10856]_ , \new_[10857]_ ,
    \new_[10858]_ , \new_[10859]_ , \new_[10860]_ , \new_[10861]_ ,
    \new_[10862]_ , \new_[10863]_ , \new_[10864]_ , \new_[10865]_ ,
    \new_[10866]_ , \new_[10867]_ , \new_[10868]_ , \new_[10869]_ ,
    \new_[10870]_ , \new_[10871]_ , \new_[10872]_ , \new_[10873]_ ,
    \new_[10874]_ , \new_[10875]_ , \new_[10876]_ , \new_[10877]_ ,
    \new_[10878]_ , \new_[10879]_ , \new_[10880]_ , \new_[10881]_ ,
    \new_[10883]_ , \new_[10884]_ , \new_[10885]_ , \new_[10886]_ ,
    \new_[10887]_ , \new_[10888]_ , \new_[10889]_ , \new_[10890]_ ,
    \new_[10891]_ , \new_[10892]_ , \new_[10893]_ , \new_[10894]_ ,
    \new_[10895]_ , \new_[10896]_ , \new_[10897]_ , \new_[10898]_ ,
    \new_[10899]_ , \new_[10900]_ , \new_[10901]_ , \new_[10902]_ ,
    \new_[10903]_ , \new_[10904]_ , \new_[10905]_ , \new_[10906]_ ,
    \new_[10907]_ , \new_[10908]_ , \new_[10909]_ , \new_[10910]_ ,
    \new_[10911]_ , \new_[10912]_ , \new_[10913]_ , \new_[10914]_ ,
    \new_[10915]_ , \new_[10916]_ , \new_[10917]_ , \new_[10918]_ ,
    \new_[10919]_ , \new_[10920]_ , \new_[10921]_ , \new_[10922]_ ,
    \new_[10923]_ , \new_[10924]_ , \new_[10926]_ , \new_[10927]_ ,
    \new_[10928]_ , \new_[10929]_ , \new_[10930]_ , \new_[10931]_ ,
    \new_[10932]_ , \new_[10933]_ , \new_[10934]_ , \new_[10935]_ ,
    \new_[10936]_ , \new_[10937]_ , \new_[10938]_ , \new_[10939]_ ,
    \new_[10940]_ , \new_[10941]_ , \new_[10942]_ , \new_[10943]_ ,
    \new_[10944]_ , \new_[10945]_ , \new_[10946]_ , \new_[10947]_ ,
    \new_[10948]_ , \new_[10949]_ , \new_[10950]_ , \new_[10951]_ ,
    \new_[10952]_ , \new_[10953]_ , \new_[10954]_ , \new_[10955]_ ,
    \new_[10956]_ , \new_[10957]_ , \new_[10958]_ , \new_[10959]_ ,
    \new_[10960]_ , \new_[10961]_ , \new_[10962]_ , \new_[10963]_ ,
    \new_[10964]_ , \new_[10965]_ , \new_[10966]_ , \new_[10968]_ ,
    \new_[10969]_ , \new_[10970]_ , \new_[10971]_ , \new_[10972]_ ,
    \new_[10973]_ , \new_[10974]_ , \new_[10975]_ , \new_[10977]_ ,
    \new_[10978]_ , \new_[10979]_ , \new_[10980]_ , \new_[10981]_ ,
    \new_[10982]_ , \new_[10983]_ , \new_[10985]_ , \new_[10986]_ ,
    \new_[10988]_ , \new_[10989]_ , \new_[10990]_ , \new_[10991]_ ,
    \new_[10993]_ , \new_[10994]_ , \new_[10995]_ , \new_[10996]_ ,
    \new_[10999]_ , \new_[11000]_ , \new_[11001]_ , \new_[11002]_ ,
    \new_[11004]_ , \new_[11005]_ , \new_[11006]_ , \new_[11007]_ ,
    \new_[11008]_ , \new_[11010]_ , \new_[11011]_ , \new_[11012]_ ,
    \new_[11013]_ , \new_[11014]_ , \new_[11015]_ , \new_[11016]_ ,
    \new_[11018]_ , \new_[11019]_ , \new_[11020]_ , \new_[11022]_ ,
    \new_[11023]_ , \new_[11024]_ , \new_[11025]_ , \new_[11026]_ ,
    \new_[11027]_ , \new_[11028]_ , \new_[11029]_ , \new_[11030]_ ,
    \new_[11031]_ , \new_[11032]_ , \new_[11033]_ , \new_[11034]_ ,
    \new_[11035]_ , \new_[11036]_ , \new_[11037]_ , \new_[11038]_ ,
    \new_[11039]_ , \new_[11040]_ , \new_[11041]_ , \new_[11042]_ ,
    \new_[11043]_ , \new_[11044]_ , \new_[11045]_ , \new_[11046]_ ,
    \new_[11047]_ , \new_[11048]_ , \new_[11050]_ , \new_[11051]_ ,
    \new_[11052]_ , \new_[11053]_ , \new_[11054]_ , \new_[11055]_ ,
    \new_[11056]_ , \new_[11057]_ , \new_[11058]_ , \new_[11059]_ ,
    \new_[11060]_ , \new_[11061]_ , \new_[11062]_ , \new_[11063]_ ,
    \new_[11064]_ , \new_[11065]_ , \new_[11066]_ , \new_[11067]_ ,
    \new_[11068]_ , \new_[11070]_ , \new_[11071]_ , \new_[11072]_ ,
    \new_[11073]_ , \new_[11074]_ , \new_[11076]_ , \new_[11077]_ ,
    \new_[11078]_ , \new_[11079]_ , \new_[11080]_ , \new_[11081]_ ,
    \new_[11082]_ , \new_[11083]_ , \new_[11084]_ , \new_[11086]_ ,
    \new_[11088]_ , \new_[11089]_ , \new_[11090]_ , \new_[11091]_ ,
    \new_[11092]_ , \new_[11093]_ , \new_[11096]_ , \new_[11097]_ ,
    \new_[11098]_ , \new_[11099]_ , \new_[11100]_ , \new_[11101]_ ,
    \new_[11102]_ , \new_[11103]_ , \new_[11104]_ , \new_[11105]_ ,
    \new_[11106]_ , \new_[11107]_ , \new_[11108]_ , \new_[11109]_ ,
    \new_[11111]_ , \new_[11113]_ , \new_[11114]_ , \new_[11117]_ ,
    \new_[11118]_ , \new_[11119]_ , \new_[11120]_ , \new_[11121]_ ,
    \new_[11122]_ , \new_[11123]_ , \new_[11124]_ , \new_[11126]_ ,
    \new_[11127]_ , \new_[11128]_ , \new_[11129]_ , \new_[11130]_ ,
    \new_[11131]_ , \new_[11132]_ , \new_[11133]_ , \new_[11134]_ ,
    \new_[11135]_ , \new_[11136]_ , \new_[11137]_ , \new_[11139]_ ,
    \new_[11140]_ , \new_[11141]_ , \new_[11142]_ , \new_[11143]_ ,
    \new_[11145]_ , \new_[11146]_ , \new_[11147]_ , \new_[11148]_ ,
    \new_[11149]_ , \new_[11150]_ , \new_[11151]_ , \new_[11152]_ ,
    \new_[11153]_ , \new_[11154]_ , \new_[11155]_ , \new_[11156]_ ,
    \new_[11157]_ , \new_[11158]_ , \new_[11159]_ , \new_[11160]_ ,
    \new_[11161]_ , \new_[11162]_ , \new_[11163]_ , \new_[11164]_ ,
    \new_[11165]_ , \new_[11166]_ , \new_[11167]_ , \new_[11168]_ ,
    \new_[11169]_ , \new_[11170]_ , \new_[11171]_ , \new_[11172]_ ,
    \new_[11173]_ , \new_[11174]_ , \new_[11175]_ , \new_[11176]_ ,
    \new_[11177]_ , \new_[11178]_ , \new_[11179]_ , \new_[11180]_ ,
    \new_[11181]_ , \new_[11182]_ , \new_[11183]_ , \new_[11184]_ ,
    \new_[11185]_ , \new_[11186]_ , \new_[11188]_ , \new_[11189]_ ,
    \new_[11190]_ , \new_[11192]_ , \new_[11193]_ , \new_[11194]_ ,
    \new_[11195]_ , \new_[11197]_ , \new_[11198]_ , \new_[11199]_ ,
    \new_[11200]_ , \new_[11201]_ , \new_[11202]_ , \new_[11203]_ ,
    \new_[11205]_ , \new_[11206]_ , \new_[11207]_ , \new_[11209]_ ,
    \new_[11212]_ , \new_[11213]_ , \new_[11214]_ , \new_[11215]_ ,
    \new_[11216]_ , \new_[11217]_ , \new_[11218]_ , \new_[11219]_ ,
    \new_[11220]_ , \new_[11221]_ , \new_[11223]_ , \new_[11224]_ ,
    \new_[11225]_ , \new_[11226]_ , \new_[11227]_ , \new_[11231]_ ,
    \new_[11232]_ , \new_[11233]_ , \new_[11234]_ , \new_[11235]_ ,
    \new_[11238]_ , \new_[11240]_ , \new_[11241]_ , \new_[11243]_ ,
    \new_[11244]_ , \new_[11245]_ , \new_[11246]_ , \new_[11247]_ ,
    \new_[11248]_ , \new_[11249]_ , \new_[11250]_ , \new_[11251]_ ,
    \new_[11252]_ , \new_[11253]_ , \new_[11254]_ , \new_[11255]_ ,
    \new_[11256]_ , \new_[11257]_ , \new_[11258]_ , \new_[11259]_ ,
    \new_[11260]_ , \new_[11261]_ , \new_[11262]_ , \new_[11263]_ ,
    \new_[11264]_ , \new_[11266]_ , \new_[11267]_ , \new_[11268]_ ,
    \new_[11269]_ , \new_[11270]_ , \new_[11271]_ , \new_[11272]_ ,
    \new_[11273]_ , \new_[11274]_ , \new_[11275]_ , \new_[11276]_ ,
    \new_[11277]_ , \new_[11278]_ , \new_[11279]_ , \new_[11280]_ ,
    \new_[11281]_ , \new_[11282]_ , \new_[11283]_ , \new_[11284]_ ,
    \new_[11285]_ , \new_[11286]_ , \new_[11287]_ , \new_[11288]_ ,
    \new_[11289]_ , \new_[11290]_ , \new_[11291]_ , \new_[11292]_ ,
    \new_[11293]_ , \new_[11294]_ , \new_[11295]_ , \new_[11296]_ ,
    \new_[11297]_ , \new_[11298]_ , \new_[11299]_ , \new_[11300]_ ,
    \new_[11301]_ , \new_[11302]_ , \new_[11303]_ , \new_[11304]_ ,
    \new_[11305]_ , \new_[11306]_ , \new_[11307]_ , \new_[11308]_ ,
    \new_[11309]_ , \new_[11310]_ , \new_[11311]_ , \new_[11312]_ ,
    \new_[11313]_ , \new_[11314]_ , \new_[11315]_ , \new_[11316]_ ,
    \new_[11317]_ , \new_[11318]_ , \new_[11319]_ , \new_[11320]_ ,
    \new_[11321]_ , \new_[11322]_ , \new_[11323]_ , \new_[11324]_ ,
    \new_[11325]_ , \new_[11326]_ , \new_[11327]_ , \new_[11328]_ ,
    \new_[11329]_ , \new_[11330]_ , \new_[11331]_ , \new_[11332]_ ,
    \new_[11333]_ , \new_[11334]_ , \new_[11335]_ , \new_[11336]_ ,
    \new_[11337]_ , \new_[11338]_ , \new_[11339]_ , \new_[11340]_ ,
    \new_[11341]_ , \new_[11342]_ , \new_[11343]_ , \new_[11344]_ ,
    \new_[11345]_ , \new_[11346]_ , \new_[11347]_ , \new_[11348]_ ,
    \new_[11349]_ , \new_[11350]_ , \new_[11351]_ , \new_[11352]_ ,
    \new_[11353]_ , \new_[11354]_ , \new_[11355]_ , \new_[11356]_ ,
    \new_[11357]_ , \new_[11358]_ , \new_[11359]_ , \new_[11360]_ ,
    \new_[11361]_ , \new_[11362]_ , \new_[11363]_ , \new_[11364]_ ,
    \new_[11365]_ , \new_[11366]_ , \new_[11367]_ , \new_[11368]_ ,
    \new_[11369]_ , \new_[11370]_ , \new_[11371]_ , \new_[11372]_ ,
    \new_[11373]_ , \new_[11374]_ , \new_[11375]_ , \new_[11376]_ ,
    \new_[11377]_ , \new_[11378]_ , \new_[11379]_ , \new_[11380]_ ,
    \new_[11381]_ , \new_[11382]_ , \new_[11383]_ , \new_[11384]_ ,
    \new_[11385]_ , \new_[11386]_ , \new_[11387]_ , \new_[11388]_ ,
    \new_[11389]_ , \new_[11390]_ , \new_[11391]_ , \new_[11392]_ ,
    \new_[11393]_ , \new_[11394]_ , \new_[11395]_ , \new_[11396]_ ,
    \new_[11397]_ , \new_[11398]_ , \new_[11399]_ , \new_[11400]_ ,
    \new_[11401]_ , \new_[11402]_ , \new_[11403]_ , \new_[11404]_ ,
    \new_[11405]_ , \new_[11406]_ , \new_[11407]_ , \new_[11408]_ ,
    \new_[11409]_ , \new_[11410]_ , \new_[11411]_ , \new_[11412]_ ,
    \new_[11413]_ , \new_[11414]_ , \new_[11415]_ , \new_[11416]_ ,
    \new_[11417]_ , \new_[11418]_ , \new_[11419]_ , \new_[11420]_ ,
    \new_[11422]_ , \new_[11423]_ , \new_[11424]_ , \new_[11425]_ ,
    \new_[11426]_ , \new_[11427]_ , \new_[11428]_ , \new_[11429]_ ,
    \new_[11430]_ , \new_[11431]_ , \new_[11432]_ , \new_[11433]_ ,
    \new_[11434]_ , \new_[11435]_ , \new_[11436]_ , \new_[11437]_ ,
    \new_[11438]_ , \new_[11439]_ , \new_[11440]_ , \new_[11441]_ ,
    \new_[11442]_ , \new_[11443]_ , \new_[11445]_ , \new_[11446]_ ,
    \new_[11447]_ , \new_[11448]_ , \new_[11449]_ , \new_[11450]_ ,
    \new_[11451]_ , \new_[11452]_ , \new_[11453]_ , \new_[11454]_ ,
    \new_[11455]_ , \new_[11456]_ , \new_[11457]_ , \new_[11458]_ ,
    \new_[11459]_ , \new_[11460]_ , \new_[11461]_ , \new_[11462]_ ,
    \new_[11463]_ , \new_[11464]_ , \new_[11465]_ , \new_[11466]_ ,
    \new_[11467]_ , \new_[11468]_ , \new_[11469]_ , \new_[11470]_ ,
    \new_[11471]_ , \new_[11472]_ , \new_[11473]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11476]_ , \new_[11477]_ , \new_[11478]_ ,
    \new_[11479]_ , \new_[11480]_ , \new_[11481]_ , \new_[11482]_ ,
    \new_[11483]_ , \new_[11484]_ , \new_[11485]_ , \new_[11486]_ ,
    \new_[11487]_ , \new_[11488]_ , \new_[11489]_ , \new_[11490]_ ,
    \new_[11491]_ , \new_[11492]_ , \new_[11493]_ , \new_[11494]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11497]_ , \new_[11498]_ ,
    \new_[11499]_ , \new_[11500]_ , \new_[11501]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11504]_ , \new_[11505]_ , \new_[11506]_ ,
    \new_[11507]_ , \new_[11508]_ , \new_[11509]_ , \new_[11510]_ ,
    \new_[11511]_ , \new_[11512]_ , \new_[11513]_ , \new_[11514]_ ,
    \new_[11515]_ , \new_[11516]_ , \new_[11517]_ , \new_[11518]_ ,
    \new_[11519]_ , \new_[11520]_ , \new_[11521]_ , \new_[11522]_ ,
    \new_[11523]_ , \new_[11524]_ , \new_[11525]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11528]_ , \new_[11529]_ , \new_[11530]_ ,
    \new_[11532]_ , \new_[11533]_ , \new_[11534]_ , \new_[11535]_ ,
    \new_[11536]_ , \new_[11537]_ , \new_[11538]_ , \new_[11540]_ ,
    \new_[11541]_ , \new_[11542]_ , \new_[11543]_ , \new_[11544]_ ,
    \new_[11545]_ , \new_[11546]_ , \new_[11548]_ , \new_[11549]_ ,
    \new_[11550]_ , \new_[11551]_ , \new_[11552]_ , \new_[11553]_ ,
    \new_[11554]_ , \new_[11555]_ , \new_[11556]_ , \new_[11557]_ ,
    \new_[11558]_ , \new_[11559]_ , \new_[11560]_ , \new_[11562]_ ,
    \new_[11563]_ , \new_[11564]_ , \new_[11565]_ , \new_[11566]_ ,
    \new_[11567]_ , \new_[11568]_ , \new_[11569]_ , \new_[11570]_ ,
    \new_[11571]_ , \new_[11572]_ , \new_[11573]_ , \new_[11574]_ ,
    \new_[11575]_ , \new_[11576]_ , \new_[11577]_ , \new_[11578]_ ,
    \new_[11579]_ , \new_[11580]_ , \new_[11581]_ , \new_[11582]_ ,
    \new_[11583]_ , \new_[11584]_ , \new_[11585]_ , \new_[11586]_ ,
    \new_[11588]_ , \new_[11589]_ , \new_[11590]_ , \new_[11592]_ ,
    \new_[11593]_ , \new_[11594]_ , \new_[11595]_ , \new_[11596]_ ,
    \new_[11597]_ , \new_[11598]_ , \new_[11600]_ , \new_[11601]_ ,
    \new_[11602]_ , \new_[11603]_ , \new_[11604]_ , \new_[11605]_ ,
    \new_[11607]_ , \new_[11608]_ , \new_[11609]_ , \new_[11610]_ ,
    \new_[11611]_ , \new_[11612]_ , \new_[11613]_ , \new_[11615]_ ,
    \new_[11616]_ , \new_[11617]_ , \new_[11618]_ , \new_[11619]_ ,
    \new_[11620]_ , \new_[11621]_ , \new_[11623]_ , \new_[11624]_ ,
    \new_[11625]_ , \new_[11626]_ , \new_[11627]_ , \new_[11628]_ ,
    \new_[11629]_ , \new_[11630]_ , \new_[11632]_ , \new_[11633]_ ,
    \new_[11634]_ , \new_[11635]_ , \new_[11636]_ , \new_[11637]_ ,
    \new_[11638]_ , \new_[11640]_ , \new_[11641]_ , \new_[11642]_ ,
    \new_[11643]_ , \new_[11644]_ , \new_[11645]_ , \new_[11647]_ ,
    \new_[11648]_ , \new_[11649]_ , \new_[11650]_ , \new_[11651]_ ,
    \new_[11652]_ , \new_[11654]_ , \new_[11655]_ , \new_[11656]_ ,
    \new_[11657]_ , \new_[11658]_ , \new_[11659]_ , \new_[11660]_ ,
    \new_[11662]_ , \new_[11663]_ , \new_[11664]_ , \new_[11665]_ ,
    \new_[11666]_ , \new_[11667]_ , \new_[11668]_ , \new_[11669]_ ,
    \new_[11670]_ , \new_[11672]_ , \new_[11673]_ , \new_[11674]_ ,
    \new_[11675]_ , \new_[11676]_ , \new_[11677]_ , \new_[11678]_ ,
    \new_[11680]_ , \new_[11681]_ , \new_[11682]_ , \new_[11683]_ ,
    \new_[11684]_ , \new_[11685]_ , \new_[11686]_ , \new_[11687]_ ,
    \new_[11689]_ , \new_[11690]_ , \new_[11691]_ , \new_[11692]_ ,
    \new_[11693]_ , \new_[11694]_ , \new_[11696]_ , \new_[11697]_ ,
    \new_[11698]_ , \new_[11699]_ , \new_[11700]_ , \new_[11701]_ ,
    \new_[11702]_ , \new_[11703]_ , \new_[11704]_ , \new_[11705]_ ,
    \new_[11706]_ , \new_[11707]_ , \new_[11708]_ , \new_[11709]_ ,
    \new_[11710]_ , \new_[11711]_ , \new_[11712]_ , \new_[11713]_ ,
    \new_[11714]_ , \new_[11715]_ , \new_[11716]_ , \new_[11717]_ ,
    \new_[11718]_ , \new_[11719]_ , \new_[11720]_ , \new_[11721]_ ,
    \new_[11722]_ , \new_[11723]_ , \new_[11724]_ , \new_[11725]_ ,
    \new_[11726]_ , \new_[11727]_ , \new_[11728]_ , \new_[11729]_ ,
    \new_[11730]_ , \new_[11731]_ , \new_[11732]_ , \new_[11733]_ ,
    \new_[11734]_ , \new_[11735]_ , \new_[11736]_ , \new_[11737]_ ,
    \new_[11738]_ , \new_[11739]_ , \new_[11740]_ , \new_[11741]_ ,
    \new_[11742]_ , \new_[11743]_ , \new_[11744]_ , \new_[11745]_ ,
    \new_[11746]_ , \new_[11747]_ , \new_[11748]_ , \new_[11749]_ ,
    \new_[11750]_ , \new_[11751]_ , \new_[11752]_ , \new_[11753]_ ,
    \new_[11754]_ , \new_[11755]_ , \new_[11756]_ , \new_[11757]_ ,
    \new_[11758]_ , \new_[11759]_ , \new_[11760]_ , \new_[11761]_ ,
    \new_[11762]_ , \new_[11763]_ , \new_[11764]_ , \new_[11765]_ ,
    \new_[11766]_ , \new_[11767]_ , \new_[11768]_ , \new_[11769]_ ,
    \new_[11770]_ , \new_[11771]_ , \new_[11772]_ , \new_[11773]_ ,
    \new_[11774]_ , \new_[11775]_ , \new_[11776]_ , \new_[11777]_ ,
    \new_[11778]_ , \new_[11779]_ , \new_[11781]_ , \new_[11782]_ ,
    \new_[11783]_ , \new_[11784]_ , \new_[11785]_ , \new_[11786]_ ,
    \new_[11787]_ , \new_[11788]_ , \new_[11789]_ , \new_[11790]_ ,
    \new_[11791]_ , \new_[11792]_ , \new_[11793]_ , \new_[11794]_ ,
    \new_[11795]_ , \new_[11796]_ , \new_[11797]_ , \new_[11798]_ ,
    \new_[11799]_ , \new_[11800]_ , \new_[11801]_ , \new_[11802]_ ,
    \new_[11803]_ , \new_[11804]_ , \new_[11805]_ , \new_[11806]_ ,
    \new_[11807]_ , \new_[11808]_ , \new_[11809]_ , \new_[11810]_ ,
    \new_[11811]_ , \new_[11812]_ , \new_[11813]_ , \new_[11814]_ ,
    \new_[11815]_ , \new_[11816]_ , \new_[11817]_ , \new_[11818]_ ,
    \new_[11819]_ , \new_[11820]_ , \new_[11821]_ , \new_[11822]_ ,
    \new_[11823]_ , \new_[11824]_ , \new_[11825]_ , \new_[11826]_ ,
    \new_[11827]_ , \new_[11828]_ , \new_[11829]_ , \new_[11830]_ ,
    \new_[11831]_ , \new_[11832]_ , \new_[11833]_ , \new_[11834]_ ,
    \new_[11835]_ , \new_[11836]_ , \new_[11837]_ , \new_[11838]_ ,
    \new_[11839]_ , \new_[11840]_ , \new_[11841]_ , \new_[11842]_ ,
    \new_[11843]_ , \new_[11844]_ , \new_[11845]_ , \new_[11846]_ ,
    \new_[11847]_ , \new_[11848]_ , \new_[11849]_ , \new_[11850]_ ,
    \new_[11851]_ , \new_[11852]_ , \new_[11853]_ , \new_[11854]_ ,
    \new_[11855]_ , \new_[11856]_ , \new_[11857]_ , \new_[11858]_ ,
    \new_[11859]_ , \new_[11860]_ , \new_[11861]_ , \new_[11862]_ ,
    \new_[11863]_ , \new_[11864]_ , \new_[11865]_ , \new_[11866]_ ,
    \new_[11867]_ , \new_[11868]_ , \new_[11869]_ , \new_[11870]_ ,
    \new_[11871]_ , \new_[11872]_ , \new_[11873]_ , \new_[11874]_ ,
    \new_[11876]_ , \new_[11877]_ , \new_[11878]_ , \new_[11879]_ ,
    \new_[11880]_ , \new_[11881]_ , \new_[11882]_ , \new_[11883]_ ,
    \new_[11884]_ , \new_[11885]_ , \new_[11886]_ , \new_[11887]_ ,
    \new_[11888]_ , \new_[11889]_ , \new_[11890]_ , \new_[11891]_ ,
    \new_[11892]_ , \new_[11893]_ , \new_[11894]_ , \new_[11895]_ ,
    \new_[11896]_ , \new_[11897]_ , \new_[11898]_ , \new_[11899]_ ,
    \new_[11900]_ , \new_[11901]_ , \new_[11902]_ , \new_[11903]_ ,
    \new_[11904]_ , \new_[11905]_ , \new_[11906]_ , \new_[11907]_ ,
    \new_[11908]_ , \new_[11909]_ , \new_[11910]_ , \new_[11911]_ ,
    \new_[11912]_ , \new_[11913]_ , \new_[11914]_ , \new_[11915]_ ,
    \new_[11916]_ , \new_[11917]_ , \new_[11918]_ , \new_[11919]_ ,
    \new_[11920]_ , \new_[11921]_ , \new_[11922]_ , \new_[11923]_ ,
    \new_[11924]_ , \new_[11925]_ , \new_[11926]_ , \new_[11927]_ ,
    \new_[11928]_ , \new_[11929]_ , \new_[11930]_ , \new_[11931]_ ,
    \new_[11932]_ , \new_[11933]_ , \new_[11934]_ , \new_[11935]_ ,
    \new_[11936]_ , \new_[11937]_ , \new_[11938]_ , \new_[11939]_ ,
    \new_[11940]_ , \new_[11941]_ , \new_[11942]_ , \new_[11943]_ ,
    \new_[11944]_ , \new_[11946]_ , \new_[11947]_ , \new_[11948]_ ,
    \new_[11949]_ , \new_[11950]_ , \new_[11951]_ , \new_[11952]_ ,
    \new_[11953]_ , \new_[11954]_ , \new_[11955]_ , \new_[11956]_ ,
    \new_[11957]_ , \new_[11958]_ , \new_[11959]_ , \new_[11960]_ ,
    \new_[11961]_ , \new_[11962]_ , \new_[11963]_ , \new_[11964]_ ,
    \new_[11965]_ , \new_[11966]_ , \new_[11967]_ , \new_[11968]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11971]_ , \new_[11972]_ ,
    \new_[11973]_ , \new_[11974]_ , \new_[11975]_ , \new_[11976]_ ,
    \new_[11977]_ , \new_[11978]_ , \new_[11979]_ , \new_[11980]_ ,
    \new_[11981]_ , \new_[11982]_ , \new_[11983]_ , \new_[11984]_ ,
    \new_[11985]_ , \new_[11986]_ , \new_[11987]_ , \new_[11988]_ ,
    \new_[11989]_ , \new_[11990]_ , \new_[11991]_ , \new_[11992]_ ,
    \new_[11993]_ , \new_[11994]_ , \new_[11995]_ , \new_[11996]_ ,
    \new_[11997]_ , \new_[11998]_ , \new_[11999]_ , \new_[12000]_ ,
    \new_[12001]_ , \new_[12002]_ , \new_[12003]_ , \new_[12005]_ ,
    \new_[12006]_ , \new_[12007]_ , \new_[12008]_ , \new_[12009]_ ,
    \new_[12010]_ , \new_[12011]_ , \new_[12013]_ , \new_[12014]_ ,
    \new_[12015]_ , \new_[12016]_ , \new_[12017]_ , \new_[12018]_ ,
    \new_[12019]_ , \new_[12020]_ , \new_[12021]_ , \new_[12022]_ ,
    \new_[12023]_ , \new_[12024]_ , \new_[12025]_ , \new_[12026]_ ,
    \new_[12027]_ , \new_[12028]_ , \new_[12029]_ , \new_[12030]_ ,
    \new_[12031]_ , \new_[12032]_ , \new_[12033]_ , \new_[12034]_ ,
    \new_[12035]_ , \new_[12036]_ , \new_[12037]_ , \new_[12038]_ ,
    \new_[12039]_ , \new_[12040]_ , \new_[12041]_ , \new_[12042]_ ,
    \new_[12043]_ , \new_[12044]_ , \new_[12045]_ , \new_[12046]_ ,
    \new_[12047]_ , \new_[12048]_ , \new_[12049]_ , \new_[12050]_ ,
    \new_[12051]_ , \new_[12052]_ , \new_[12053]_ , \new_[12054]_ ,
    \new_[12055]_ , \new_[12056]_ , \new_[12057]_ , \new_[12058]_ ,
    \new_[12059]_ , \new_[12060]_ , \new_[12061]_ , \new_[12062]_ ,
    \new_[12063]_ , \new_[12064]_ , \new_[12066]_ , \new_[12067]_ ,
    \new_[12068]_ , \new_[12069]_ , \new_[12070]_ , \new_[12071]_ ,
    \new_[12072]_ , \new_[12073]_ , \new_[12074]_ , \new_[12075]_ ,
    \new_[12077]_ , \new_[12078]_ , \new_[12079]_ , \new_[12080]_ ,
    \new_[12081]_ , \new_[12082]_ , \new_[12083]_ , \new_[12084]_ ,
    \new_[12085]_ , \new_[12086]_ , \new_[12087]_ , \new_[12088]_ ,
    \new_[12089]_ , \new_[12090]_ , \new_[12091]_ , \new_[12092]_ ,
    \new_[12093]_ , \new_[12094]_ , \new_[12095]_ , \new_[12096]_ ,
    \new_[12097]_ , \new_[12098]_ , \new_[12099]_ , \new_[12100]_ ,
    \new_[12101]_ , \new_[12102]_ , \new_[12103]_ , \new_[12104]_ ,
    \new_[12105]_ , \new_[12106]_ , \new_[12107]_ , \new_[12108]_ ,
    \new_[12109]_ , \new_[12110]_ , \new_[12111]_ , \new_[12112]_ ,
    \new_[12113]_ , \new_[12114]_ , \new_[12115]_ , \new_[12116]_ ,
    \new_[12117]_ , \new_[12118]_ , \new_[12119]_ , \new_[12120]_ ,
    \new_[12121]_ , \new_[12122]_ , \new_[12123]_ , \new_[12124]_ ,
    \new_[12125]_ , \new_[12126]_ , \new_[12127]_ , \new_[12128]_ ,
    \new_[12129]_ , \new_[12130]_ , \new_[12131]_ , \new_[12132]_ ,
    \new_[12133]_ , \new_[12134]_ , \new_[12135]_ , \new_[12136]_ ,
    \new_[12137]_ , \new_[12138]_ , \new_[12139]_ , \new_[12140]_ ,
    \new_[12141]_ , \new_[12142]_ , \new_[12143]_ , \new_[12144]_ ,
    \new_[12145]_ , \new_[12146]_ , \new_[12147]_ , \new_[12148]_ ,
    \new_[12149]_ , \new_[12150]_ , \new_[12151]_ , \new_[12152]_ ,
    \new_[12153]_ , \new_[12154]_ , \new_[12155]_ , \new_[12156]_ ,
    \new_[12157]_ , \new_[12158]_ , \new_[12159]_ , \new_[12160]_ ,
    \new_[12161]_ , \new_[12162]_ , \new_[12163]_ , \new_[12164]_ ,
    \new_[12165]_ , \new_[12166]_ , \new_[12167]_ , \new_[12168]_ ,
    \new_[12169]_ , \new_[12170]_ , \new_[12171]_ , \new_[12172]_ ,
    \new_[12173]_ , \new_[12174]_ , \new_[12175]_ , \new_[12176]_ ,
    \new_[12177]_ , \new_[12178]_ , \new_[12179]_ , \new_[12180]_ ,
    \new_[12181]_ , \new_[12182]_ , \new_[12183]_ , \new_[12184]_ ,
    \new_[12185]_ , \new_[12186]_ , \new_[12187]_ , \new_[12188]_ ,
    \new_[12189]_ , \new_[12190]_ , \new_[12191]_ , \new_[12192]_ ,
    \new_[12193]_ , \new_[12194]_ , \new_[12195]_ , \new_[12197]_ ,
    \new_[12198]_ , \new_[12199]_ , \new_[12200]_ , \new_[12201]_ ,
    \new_[12202]_ , \new_[12204]_ , \new_[12205]_ , \new_[12206]_ ,
    \new_[12207]_ , \new_[12208]_ , \new_[12209]_ , \new_[12210]_ ,
    \new_[12211]_ , \new_[12212]_ , \new_[12213]_ , \new_[12214]_ ,
    \new_[12215]_ , \new_[12216]_ , \new_[12217]_ , \new_[12218]_ ,
    \new_[12219]_ , \new_[12220]_ , \new_[12221]_ , \new_[12222]_ ,
    \new_[12223]_ , \new_[12224]_ , \new_[12225]_ , \new_[12226]_ ,
    \new_[12227]_ , \new_[12228]_ , \new_[12229]_ , \new_[12230]_ ,
    \new_[12231]_ , \new_[12232]_ , \new_[12233]_ , \new_[12234]_ ,
    \new_[12235]_ , \new_[12236]_ , \new_[12237]_ , \new_[12238]_ ,
    \new_[12239]_ , \new_[12240]_ , \new_[12242]_ , \new_[12243]_ ,
    \new_[12244]_ , \new_[12245]_ , \new_[12246]_ , \new_[12247]_ ,
    \new_[12248]_ , \new_[12250]_ , \new_[12251]_ , \new_[12252]_ ,
    \new_[12253]_ , \new_[12254]_ , \new_[12255]_ , \new_[12256]_ ,
    \new_[12257]_ , \new_[12258]_ , \new_[12259]_ , \new_[12261]_ ,
    \new_[12262]_ , \new_[12263]_ , \new_[12264]_ , \new_[12265]_ ,
    \new_[12266]_ , \new_[12267]_ , \new_[12268]_ , \new_[12269]_ ,
    \new_[12270]_ , \new_[12271]_ , \new_[12272]_ , \new_[12273]_ ,
    \new_[12274]_ , \new_[12275]_ , \new_[12276]_ , \new_[12277]_ ,
    \new_[12278]_ , \new_[12279]_ , \new_[12280]_ , \new_[12281]_ ,
    \new_[12282]_ , \new_[12283]_ , \new_[12284]_ , \new_[12285]_ ,
    \new_[12286]_ , \new_[12287]_ , \new_[12288]_ , \new_[12289]_ ,
    \new_[12290]_ , \new_[12291]_ , \new_[12292]_ , \new_[12293]_ ,
    \new_[12294]_ , \new_[12295]_ , \new_[12296]_ , \new_[12297]_ ,
    \new_[12298]_ , \new_[12299]_ , \new_[12300]_ , \new_[12301]_ ,
    \new_[12302]_ , \new_[12303]_ , \new_[12304]_ , \new_[12305]_ ,
    \new_[12306]_ , \new_[12307]_ , \new_[12308]_ , \new_[12309]_ ,
    \new_[12310]_ , \new_[12311]_ , \new_[12312]_ , \new_[12313]_ ,
    \new_[12314]_ , \new_[12315]_ , \new_[12316]_ , \new_[12317]_ ,
    \new_[12318]_ , \new_[12319]_ , \new_[12320]_ , \new_[12321]_ ,
    \new_[12322]_ , \new_[12323]_ , \new_[12324]_ , \new_[12326]_ ,
    \new_[12327]_ , \new_[12328]_ , \new_[12329]_ , \new_[12330]_ ,
    \new_[12331]_ , \new_[12332]_ , \new_[12333]_ , \new_[12334]_ ,
    \new_[12335]_ , \new_[12336]_ , \new_[12337]_ , \new_[12338]_ ,
    \new_[12339]_ , \new_[12340]_ , \new_[12341]_ , \new_[12342]_ ,
    \new_[12343]_ , \new_[12344]_ , \new_[12345]_ , \new_[12346]_ ,
    \new_[12347]_ , \new_[12348]_ , \new_[12349]_ , \new_[12350]_ ,
    \new_[12351]_ , \new_[12352]_ , \new_[12353]_ , \new_[12354]_ ,
    \new_[12355]_ , \new_[12356]_ , \new_[12357]_ , \new_[12358]_ ,
    \new_[12359]_ , \new_[12360]_ , \new_[12361]_ , \new_[12362]_ ,
    \new_[12363]_ , \new_[12364]_ , \new_[12365]_ , \new_[12366]_ ,
    \new_[12367]_ , \new_[12368]_ , \new_[12369]_ , \new_[12370]_ ,
    \new_[12371]_ , \new_[12372]_ , \new_[12373]_ , \new_[12374]_ ,
    \new_[12375]_ , \new_[12376]_ , \new_[12377]_ , \new_[12378]_ ,
    \new_[12379]_ , \new_[12380]_ , \new_[12381]_ , \new_[12382]_ ,
    \new_[12383]_ , \new_[12384]_ , \new_[12385]_ , \new_[12386]_ ,
    \new_[12387]_ , \new_[12388]_ , \new_[12389]_ , \new_[12390]_ ,
    \new_[12391]_ , \new_[12392]_ , \new_[12393]_ , \new_[12394]_ ,
    \new_[12395]_ , \new_[12396]_ , \new_[12397]_ , \new_[12398]_ ,
    \new_[12399]_ , \new_[12400]_ , \new_[12401]_ , \new_[12402]_ ,
    \new_[12403]_ , \new_[12405]_ , \new_[12406]_ , \new_[12407]_ ,
    \new_[12408]_ , \new_[12409]_ , \new_[12410]_ , \new_[12411]_ ,
    \new_[12412]_ , \new_[12413]_ , \new_[12414]_ , \new_[12415]_ ,
    \new_[12416]_ , \new_[12417]_ , \new_[12418]_ , \new_[12419]_ ,
    \new_[12420]_ , \new_[12421]_ , \new_[12422]_ , \new_[12423]_ ,
    \new_[12424]_ , \new_[12425]_ , \new_[12426]_ , \new_[12427]_ ,
    \new_[12428]_ , \new_[12429]_ , \new_[12430]_ , \new_[12431]_ ,
    \new_[12432]_ , \new_[12433]_ , \new_[12434]_ , \new_[12435]_ ,
    \new_[12436]_ , \new_[12437]_ , \new_[12438]_ , \new_[12439]_ ,
    \new_[12440]_ , \new_[12441]_ , \new_[12442]_ , \new_[12443]_ ,
    \new_[12444]_ , \new_[12445]_ , \new_[12446]_ , \new_[12447]_ ,
    \new_[12448]_ , \new_[12449]_ , \new_[12450]_ , \new_[12451]_ ,
    \new_[12452]_ , \new_[12453]_ , \new_[12454]_ , \new_[12455]_ ,
    \new_[12456]_ , \new_[12457]_ , \new_[12458]_ , \new_[12459]_ ,
    \new_[12460]_ , \new_[12461]_ , \new_[12462]_ , \new_[12463]_ ,
    \new_[12464]_ , \new_[12465]_ , \new_[12466]_ , \new_[12467]_ ,
    \new_[12468]_ , \new_[12469]_ , \new_[12470]_ , \new_[12471]_ ,
    \new_[12472]_ , \new_[12473]_ , \new_[12474]_ , \new_[12475]_ ,
    \new_[12476]_ , \new_[12477]_ , \new_[12478]_ , \new_[12479]_ ,
    \new_[12480]_ , \new_[12481]_ , \new_[12482]_ , \new_[12483]_ ,
    \new_[12484]_ , \new_[12485]_ , \new_[12486]_ , \new_[12487]_ ,
    \new_[12488]_ , \new_[12489]_ , \new_[12490]_ , \new_[12491]_ ,
    \new_[12492]_ , \new_[12493]_ , \new_[12494]_ , \new_[12495]_ ,
    \new_[12496]_ , \new_[12497]_ , \new_[12498]_ , \new_[12499]_ ,
    \new_[12500]_ , \new_[12501]_ , \new_[12503]_ , \new_[12504]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12507]_ , \new_[12508]_ ,
    \new_[12509]_ , \new_[12510]_ , \new_[12511]_ , \new_[12512]_ ,
    \new_[12513]_ , \new_[12514]_ , \new_[12515]_ , \new_[12516]_ ,
    \new_[12517]_ , \new_[12518]_ , \new_[12519]_ , \new_[12520]_ ,
    \new_[12522]_ , \new_[12523]_ , \new_[12524]_ , \new_[12525]_ ,
    \new_[12526]_ , \new_[12527]_ , \new_[12528]_ , \new_[12529]_ ,
    \new_[12530]_ , \new_[12531]_ , \new_[12532]_ , \new_[12533]_ ,
    \new_[12534]_ , \new_[12535]_ , \new_[12536]_ , \new_[12537]_ ,
    \new_[12538]_ , \new_[12539]_ , \new_[12540]_ , \new_[12541]_ ,
    \new_[12542]_ , \new_[12543]_ , \new_[12544]_ , \new_[12545]_ ,
    \new_[12546]_ , \new_[12547]_ , \new_[12548]_ , \new_[12549]_ ,
    \new_[12550]_ , \new_[12551]_ , \new_[12552]_ , \new_[12553]_ ,
    \new_[12554]_ , \new_[12555]_ , \new_[12556]_ , \new_[12557]_ ,
    \new_[12558]_ , \new_[12559]_ , \new_[12560]_ , \new_[12561]_ ,
    \new_[12562]_ , \new_[12563]_ , \new_[12564]_ , \new_[12565]_ ,
    \new_[12566]_ , \new_[12567]_ , \new_[12568]_ , \new_[12569]_ ,
    \new_[12570]_ , \new_[12571]_ , \new_[12572]_ , \new_[12573]_ ,
    \new_[12574]_ , \new_[12575]_ , \new_[12576]_ , \new_[12577]_ ,
    \new_[12578]_ , \new_[12579]_ , \new_[12580]_ , \new_[12581]_ ,
    \new_[12582]_ , \new_[12583]_ , \new_[12584]_ , \new_[12585]_ ,
    \new_[12586]_ , \new_[12587]_ , \new_[12588]_ , \new_[12589]_ ,
    \new_[12590]_ , \new_[12591]_ , \new_[12592]_ , \new_[12593]_ ,
    \new_[12594]_ , \new_[12595]_ , \new_[12596]_ , \new_[12597]_ ,
    \new_[12598]_ , \new_[12599]_ , \new_[12600]_ , \new_[12601]_ ,
    \new_[12602]_ , \new_[12603]_ , \new_[12604]_ , \new_[12605]_ ,
    \new_[12606]_ , \new_[12607]_ , \new_[12608]_ , \new_[12609]_ ,
    \new_[12610]_ , \new_[12611]_ , \new_[12612]_ , \new_[12613]_ ,
    \new_[12614]_ , \new_[12615]_ , \new_[12616]_ , \new_[12617]_ ,
    \new_[12618]_ , \new_[12619]_ , \new_[12620]_ , \new_[12621]_ ,
    \new_[12622]_ , \new_[12623]_ , \new_[12624]_ , \new_[12625]_ ,
    \new_[12626]_ , \new_[12627]_ , \new_[12628]_ , \new_[12629]_ ,
    \new_[12630]_ , \new_[12631]_ , \new_[12632]_ , \new_[12633]_ ,
    \new_[12634]_ , \new_[12635]_ , \new_[12636]_ , \new_[12637]_ ,
    \new_[12638]_ , \new_[12639]_ , \new_[12640]_ , \new_[12641]_ ,
    \new_[12642]_ , \new_[12643]_ , \new_[12644]_ , \new_[12645]_ ,
    \new_[12646]_ , \new_[12647]_ , \new_[12648]_ , \new_[12649]_ ,
    \new_[12650]_ , \new_[12651]_ , \new_[12652]_ , \new_[12653]_ ,
    \new_[12654]_ , \new_[12655]_ , \new_[12656]_ , \new_[12657]_ ,
    \new_[12658]_ , \new_[12659]_ , \new_[12660]_ , \new_[12661]_ ,
    \new_[12662]_ , \new_[12663]_ , \new_[12664]_ , \new_[12665]_ ,
    \new_[12666]_ , \new_[12667]_ , \new_[12668]_ , \new_[12669]_ ,
    \new_[12670]_ , \new_[12671]_ , \new_[12672]_ , \new_[12673]_ ,
    \new_[12674]_ , \new_[12675]_ , \new_[12676]_ , \new_[12677]_ ,
    \new_[12678]_ , \new_[12679]_ , \new_[12680]_ , \new_[12681]_ ,
    \new_[12682]_ , \new_[12683]_ , \new_[12684]_ , \new_[12685]_ ,
    \new_[12686]_ , \new_[12687]_ , \new_[12688]_ , \new_[12689]_ ,
    \new_[12690]_ , \new_[12691]_ , \new_[12692]_ , \new_[12693]_ ,
    \new_[12694]_ , \new_[12695]_ , \new_[12696]_ , \new_[12697]_ ,
    \new_[12698]_ , \new_[12699]_ , \new_[12700]_ , \new_[12701]_ ,
    \new_[12702]_ , \new_[12703]_ , \new_[12704]_ , \new_[12705]_ ,
    \new_[12706]_ , \new_[12707]_ , \new_[12708]_ , \new_[12709]_ ,
    \new_[12710]_ , \new_[12711]_ , \new_[12712]_ , \new_[12713]_ ,
    \new_[12714]_ , \new_[12715]_ , \new_[12716]_ , \new_[12717]_ ,
    \new_[12718]_ , \new_[12719]_ , \new_[12720]_ , \new_[12721]_ ,
    \new_[12722]_ , \new_[12723]_ , \new_[12724]_ , \new_[12725]_ ,
    \new_[12726]_ , \new_[12727]_ , \new_[12728]_ , \new_[12729]_ ,
    \new_[12730]_ , \new_[12731]_ , \new_[12732]_ , \new_[12733]_ ,
    \new_[12734]_ , \new_[12735]_ , \new_[12736]_ , \new_[12737]_ ,
    \new_[12738]_ , \new_[12739]_ , \new_[12740]_ , \new_[12741]_ ,
    \new_[12742]_ , \new_[12743]_ , \new_[12744]_ , \new_[12745]_ ,
    \new_[12746]_ , \new_[12747]_ , \new_[12748]_ , \new_[12749]_ ,
    \new_[12750]_ , \new_[12751]_ , \new_[12752]_ , \new_[12753]_ ,
    \new_[12754]_ , \new_[12755]_ , \new_[12756]_ , \new_[12757]_ ,
    \new_[12758]_ , \new_[12759]_ , \new_[12760]_ , \new_[12761]_ ,
    \new_[12762]_ , \new_[12763]_ , \new_[12764]_ , \new_[12765]_ ,
    \new_[12766]_ , \new_[12767]_ , \new_[12768]_ , \new_[12769]_ ,
    \new_[12770]_ , \new_[12771]_ , \new_[12772]_ , \new_[12773]_ ,
    \new_[12774]_ , \new_[12775]_ , \new_[12776]_ , \new_[12777]_ ,
    \new_[12778]_ , \new_[12779]_ , \new_[12780]_ , \new_[12781]_ ,
    \new_[12782]_ , \new_[12783]_ , \new_[12784]_ , \new_[12785]_ ,
    \new_[12786]_ , \new_[12787]_ , \new_[12788]_ , \new_[12789]_ ,
    \new_[12790]_ , \new_[12791]_ , \new_[12792]_ , \new_[12793]_ ,
    \new_[12794]_ , n536, n541, n546, n551, n556, n561, n566, n571, n576,
    n581, n586, n591, n596, n601, n606, n611, n616, n621, n626, n631, n636,
    n641, n646, n651, n656, n661, n666, n671, n676, n681, n686, n691, n696,
    n701, n706, n711, n716, n721, n726, n731, n736, n741, n746, n751, n756,
    n761, n766, n771, n776, n781, n786, n791, n796, n801, n806, n811, n816,
    n821, n826, n831, n836, n841, n846, n851, n856, n861, n866, n871, n876,
    n881, n886, n891, n896, n901, n906, n911, n916, n921, n926, n931, n936,
    n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996,
    n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046,
    n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096,
    n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146,
    n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196,
    n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246,
    n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296,
    n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346,
    n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396,
    n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446,
    n1451, n1456, n1461, n1466, n1471, n1476, n1481, n1486, n1491, n1496,
    n1501, n1506, n1511, n1516, n1521, n1526, n1531, n1536, n1541, n1546,
    n1551, n1556, n1561, n1566, n1571, n1576, n1581, n1586, n1591, n1596,
    n1601, n1606, n1611, n1616, n1621, n1626, n1631, n1636, n1641, n1646,
    n1651, n1656, n1661, n1666, n1671, n1676, n1681, n1686, n1691, n1696,
    n1701, n1706, n1711, n1716, n1721, n1726, n1731, n1736, n1741, n1746,
    n1751, n1756, n1761, n1766, n1771, n1776, n1781, n1786, n1791, n1796,
    n1801, n1806, n1811, n1816, n1821, n1826, n1831, n1836, n1841, n1846,
    n1851, n1856, n1861, n1866, n1871, n1876, n1881, n1886, n1891, n1896,
    n1901, n1906, n1911, n1916, n1921, n1926, n1931, n1936, n1941, n1946,
    n1951, n1956, n1961, n1966, n1971, n1976, n1981, n1986, n1991, n1996,
    n2001, n2006, n2011, n2016, n2021, n2026, n2031, n2036, n2041, n2046,
    n2051, n2056, n2061, n2066, n2071, n2076, n2081, n2086, n2091, n2096,
    n2101, n2106, n2111, n2116, n2121, n2126, n2131, n2136, n2141, n2146,
    n2151, n2156, n2161, n2166, n2171, n2176, n2181, n2186, n2191, n2196,
    n2201, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246,
    n2251, n2256, n2261, n2266, n2271, n2276, n2281, n2286, n2291, n2296,
    n2301, n2306, n2311, n2316, n2321, n2326, n2331, n2336, n2341, n2346,
    n2351, n2356, n2361, n2366, n2371, n2376, n2381, n2386, n2391, n2396,
    n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436, n2441, n2446,
    n2451, n2456, n2461, n2466, n2471, n2476, n2481, n2486, n2491, n2496,
    n2501, n2506, n2511, n2516, n2521, n2526, n2531, n2536, n2541, n2546,
    n2551, n2556, n2561, n2566, n2571, n2576, n2581, n2586, n2591, n2596,
    n2601, n2606, n2611, n2616, n2621, n2626, n2631, n2636, n2641, n2646,
    n2651, n2656, n2661, n2666, n2671, n2676, n2681, n2686, n2691, n2696,
    n2701, n2706, n2711, n2716, n2721, n2726, n2731, n2736, n2741, n2746,
    n2751, n2756, n2761, n2766, n2771, n2776, n2781, n2786, n2791, n2796,
    n2801, n2806, n2811, n2816, n2821, n2826, n2831, n2836, n2841, n2846,
    n2851, n2856, n2861, n2866, n2871, n2876, n2881, n2886, n2891, n2896,
    n2901, n2906, n2911, n2916, n2921, n2926, n2931, n2936, n2941, n2946,
    n2951, n2956, n2961, n2966, n2971, n2976, n2981, n2986, n2991, n2996,
    n3001, n3006, n3011, n3016, n3021, n3026, n3031, n3036, n3041, n3046,
    n3051, n3056, n3061, n3066, n3071, n3076, n3081, n3086, n3091, n3096,
    n3101, n3106, n3111, n3116, n3121, n3126, n3131, n3136, n3141, n3146,
    n3151, n3156, n3161, n3166, n3171, n3176, n3181, n3186, n3191, n3196,
    n3201, n3206, n3211, n3216, n3221, n3226, n3231, n3236, n3241, n3246,
    n3251, n3256, n3261, n3266, n3271, n3276, n3281, n3286, n3291, n3296,
    n3301, n3306, n3311, n3316, n3321, n3326, n3331, n3336, n3341, n3346,
    n3351, n3356, n3361, n3366, n3371, n3376, n3381, n3386, n3391, n3396,
    n3401, n3406, n3411, n3416, n3421, n3426, n3431, n3436, n3441, n3446,
    n3451, n3456, n3461, n3466, n3471, n3476, n3481, n3486, n3491, n3496,
    n3501, n3506, n3511, n3516, n3521, n3526, n3531, n3536, n3541, n3546,
    n3551, n3556, n3561, n3566, n3571, n3576, n3581, n3586, n3591, n3596,
    n3601, n3606, n3611, n3616, n3621, n3626, n3631, n3636, n3641, n3646,
    n3651, n3656, n3661, n3666, n3671, n3676, n3681, n3686, n3691, n3696,
    n3701, n3706, n3711, n3716, n3721, n3726, n3731, n3736, n3741, n3746,
    n3751, n3756, n3761, n3766, n3771, n3776, n3781, n3786, n3791, n3796,
    n3801, n3806, n3811, n3816, n3821, n3826, n3831, n3836, n3841, n3846,
    n3851, n3856, n3861, n3866, n3871, n3876, n3881, n3886, n3891, n3896,
    n3901, n3906, n3911, n3916, n3921, n3926, n3931, n3936, n3941, n3946,
    n3951, n3956, n3961, n3966, n3971, n3976, n3981, n3986, n3991, n3996,
    n4001, n4006, n4011, n4016, n4021, n4026, n4031, n4036, n4041, n4046,
    n4051, n4056, n4061, n4066, n4071, n4076, n4081, n4086, n4091, n4096,
    n4101, n4106, n4111, n4116, n4121, n4126, n4131, n4136, n4141, n4146,
    n4151, n4156, n4161, n4166, n4171, n4176, n4181, n4186, n4191, n4196,
    n4201, n4206, n4211, n4216, n4221, n4226, n4231, n4236, n4241, n4246,
    n4251, n4256, n4261, n4266, n4271, n4276, n4281, n4286, n4291, n4296,
    n4301, n4306, n4311, n4316, n4321, n4326, n4331, n4336, n4341, n4346,
    n4351, n4356, n4361, n4366, n4371, n4376, n4381, n4386, n4391, n4396,
    n4401, n4406, n4411, n4416, n4421, n4426, n4431, n4436, n4441, n4446,
    n4451, n4456, n4461, n4466, n4471, n4476, n4481, n4486, n4491, n4496,
    n4501, n4506, n4511, n4516, n4521, n4526, n4531, n4536, n4541, n4546,
    n4551, n4556, n4561, n4566, n4571, n4576, n4581, n4586, n4591, n4596,
    n4601, n4606, n4611, n4616, n4621, n4626, n4631, n4636, n4641, n4646,
    n4651, n4656, n4661, n4666, n4671, n4676, n4681, n4686, n4691, n4696,
    n4701, n4706, n4711, n4716, n4721, n4726, n4731, n4736, n4741, n4746,
    n4751, n4756, n4761, n4766, n4771, n4776, n4781, n4786, n4791, n4796,
    n4801, n4806, n4811, n4816, n4821, n4826, n4831, n4836, n4841, n4846,
    n4851, n4856, n4861, n4866, n4871, n4876, n4881, n4886, n4891, n4896,
    n4901, n4906, n4911, n4916, n4921, n4926, n4931, n4936, n4941, n4946,
    n4951, n4956, n4961, n4966, n4971, n4976, n4981, n4986, n4991, n4996,
    n5001, n5006, n5011, n5016, n5021, n5026, n5031, n5036, n5041, n5046,
    n5051, n5056, n5061, n5066, n5071, n5076, n5081, n5086, n5091, n5096,
    n5101, n5106, n5111, n5116, n5121, n5126, n5131, n5136, n5141, n5146,
    n5151, n5156, n5161, n5166, n5171, n5176, n5181, n5186, n5191, n5196,
    n5201, n5206, n5211, n5216, n5221, n5226, n5231, n5236, n5241, n5246,
    n5251, n5256, n5261, n5266, n5271, n5276, n5281, n5286, n5291, n5296,
    n5301, n5306, n5311, n5316, n5321, n5326, n5331, n5336, n5341, n5346,
    n5351, n5356, n5361, n5366, n5371, n5376, n5381, n5386, n5391, n5396,
    n5401, n5406, n5411, n5416, n5421, n5426, n5431, n5436, n5441, n5446,
    n5451, n5456, n5461, n5466, n5471, n5476, n5481, n5486, n5491, n5496,
    n5501, n5506, n5511, n5516, n5521, n5526, n5531, n5536, n5541, n5546,
    n5551, n5556, n5561, n5566, n5571, n5576, n5581, n5586, n5591, n5596,
    n5601, n5606, n5611, n5616, n5621, n5626, n5631, n5636, n5641, n5646,
    n5651, n5656, n5661, n5666, n5671, n5676, n5681, n5686, n5691, n5696,
    n5701, n5706, n5711, n5716, n5721, n5726, n5731, n5736, n5741, n5746,
    n5751, n5756, n5761, n5766, n5771, n5776, n5781, n5786, n5791, n5796,
    n5801, n5806, n5811, n5816, n5821, n5826, n5831, n5836, n5841, n5846,
    n5851, n5856, n5861, n5866, n5871, n5876, n5881, n5886, n5891, n5896,
    n5901, n5906, n5911, n5916, n5921, n5926, n5931, n5936, n5941, n5946;
  assign new_u5_rsts1_reg_in_ = 1'b0;
  assign \mc_addr_pad_o[10]  = \\u7_mc_addr_reg[10] ;
  assign \mc_addr_pad_o[12]  = \\u7_mc_addr_reg[12] ;
  assign \mc_addr_pad_o[11]  = \\u7_mc_addr_reg[11] ;
  assign n536 = ~\new_[6650]_  | ~\new_[10805]_  | ~\new_[1382]_  | ~\new_[6473]_ ;
  assign \mc_addr_pad_o[9]  = \\u7_mc_addr_reg[9] ;
  assign \mc_addr_pad_o[8]  = \\u7_mc_addr_reg[8] ;
  assign \mc_addr_pad_o[7]  = \\u7_mc_addr_reg[7] ;
  assign \mc_addr_pad_o[6]  = \\u7_mc_addr_reg[6] ;
  assign \mc_addr_pad_o[5]  = \\u7_mc_addr_reg[5] ;
  assign \mc_addr_pad_o[4]  = \\u7_mc_addr_reg[4] ;
  assign \mc_addr_pad_o[3]  = \\u7_mc_addr_reg[3] ;
  assign \mc_addr_pad_o[2]  = \\u7_mc_addr_reg[2] ;
  assign \mc_addr_pad_o[1]  = \\u7_mc_addr_reg[1] ;
  assign \mc_addr_pad_o[0]  = \\u7_mc_addr_reg[0] ;
  assign n541 = ~\new_[6474]_  | ~\new_[1381]_  | ~\new_[6649]_ ;
  assign n546 = ~\new_[6489]_  | ~\new_[1379]_  | ~\new_[6648]_ ;
  assign n581 = ~\new_[1384]_  | ~\new_[6485]_ ;
  assign n596 = ~\new_[1398]_  | ~\new_[6472]_ ;
  assign n576 = ~\new_[1385]_  | ~\new_[6486]_ ;
  assign n571 = ~\new_[1394]_  | ~\new_[6487]_ ;
  assign n566 = ~\new_[1395]_  | ~\new_[6488]_ ;
  assign n561 = ~\new_[1396]_  | ~\new_[6494]_ ;
  assign n591 = ~\new_[1380]_  | ~\new_[6479]_ ;
  assign n556 = ~\new_[1397]_  | ~\new_[6493]_ ;
  assign n551 = ~\new_[1399]_  | ~\new_[6491]_ ;
  assign n586 = ~\new_[1383]_  | ~\new_[6484]_ ;
  assign mc_we_pad_o_ = u7_mc_we__reg;
  assign \new_[1379]_  = ~\new_[1425]_  | ~\new_[1420]_  | ~\new_[7286]_ ;
  assign \new_[1380]_  = (~\new_[1411]_  | ~\new_[7286]_ ) & (~\new_[3183]_  | ~\new_[6830]_ );
  assign \new_[1381]_  = ~\new_[1422]_  | ~\new_[1421]_  | ~\new_[7286]_ ;
  assign \new_[1382]_  = ~\new_[1400]_  | ~\new_[6064]_ ;
  assign \new_[1383]_  = (~\new_[1412]_  | ~\new_[7286]_ ) & (~\new_[3114]_  | ~\new_[6830]_ );
  assign \new_[1384]_  = (~\new_[1413]_  | ~\new_[7286]_ ) & (~\new_[10710]_  | ~\new_[7115]_ );
  assign \new_[1385]_  = (~\new_[1414]_  | ~\new_[7286]_ ) & (~\new_[10836]_  | ~\new_[7115]_ );
  assign \mc_cs_pad_o_[1]  = \\u7_mc_cs__reg[1] ;
  assign \mc_cs_pad_o_[0]  = \\u7_mc_cs__reg[0] ;
  assign \mc_cs_pad_o_[7]  = \\u7_mc_cs__reg[7] ;
  assign \mc_cs_pad_o_[6]  = \\u7_mc_cs__reg[6] ;
  assign \mc_cs_pad_o_[5]  = \\u7_mc_cs__reg[5] ;
  assign \mc_cs_pad_o_[4]  = \\u7_mc_cs__reg[4] ;
  assign \mc_cs_pad_o_[3]  = \\u7_mc_cs__reg[3] ;
  assign \mc_cs_pad_o_[2]  = \\u7_mc_cs__reg[2] ;
  assign \new_[1394]_  = (~\new_[1415]_  | ~\new_[7286]_ ) & (~\new_[11100]_  | ~\new_[6831]_ );
  assign \new_[1395]_  = (~\new_[1416]_  | ~\new_[7286]_ ) & (~\new_[10820]_  | ~\new_[6831]_ );
  assign \new_[1396]_  = (~\new_[1417]_  | ~\new_[7286]_ ) & (~\new_[11131]_  | ~\new_[6831]_ );
  assign \new_[1397]_  = (~\new_[1418]_  | ~\new_[7286]_ ) & (~\new_[11205]_  | ~\new_[6830]_ );
  assign \new_[1398]_  = (~\new_[1410]_  | ~\new_[7286]_ ) & (~\new_[3182]_  | ~\new_[6831]_ );
  assign \new_[1399]_  = (~\new_[1419]_  | ~\new_[7286]_ ) & (~\new_[11051]_  | ~\new_[6830]_ );
  assign \new_[1400]_  = ~\new_[1442]_  | ~\new_[1424]_ ;
  assign n611 = \new_[1423]_  | \new_[11404]_ ;
  assign n606 = \new_[1423]_  | \new_[11403]_ ;
  assign n641 = \new_[7912]_  | \new_[1423]_ ;
  assign n636 = \new_[7910]_  | \new_[1423]_ ;
  assign n631 = \new_[7699]_  | \new_[1423]_ ;
  assign n626 = \new_[7855]_  | \new_[1423]_ ;
  assign n621 = \new_[7808]_  | \new_[1423]_ ;
  assign n616 = \new_[7810]_  | \new_[1423]_ ;
  assign \new_[1410]_  = \new_[12467]_  ? \new_[1430]_  : \new_[3617]_ ;
  assign \new_[1411]_  = \new_[11406]_  ? \new_[1429]_  : \new_[3618]_ ;
  assign \new_[1412]_  = \new_[11409]_  ? \new_[1429]_  : \new_[3619]_ ;
  assign \new_[1413]_  = \new_[5701]_  ? \new_[1430]_  : \new_[3620]_ ;
  assign \new_[1414]_  = \new_[7376]_  ? \new_[1430]_  : \new_[3621]_ ;
  assign \new_[1415]_  = \new_[7375]_  ? \new_[1432]_  : \new_[3622]_ ;
  assign \new_[1416]_  = \new_[5695]_  ? \new_[1430]_  : \new_[3623]_ ;
  assign \new_[1417]_  = \new_[5703]_  ? \new_[1432]_  : \new_[3624]_ ;
  assign \new_[1418]_  = \new_[6337]_  ? \new_[1429]_  : \new_[3625]_ ;
  assign \new_[1419]_  = \new_[12499]_  ? \new_[1429]_  : \new_[3626]_ ;
  assign \new_[1420]_  = ~\new_[6076]_  | ~\new_[1426]_ ;
  assign \new_[1421]_  = ~\new_[4819]_  | ~\new_[1426]_ ;
  assign \new_[1422]_  = ~\new_[3825]_  | ~\new_[1432]_ ;
  assign \new_[1423]_  = \new_[1427]_ ;
  assign \new_[1424]_  = ~\new_[2495]_  | ~\new_[1431]_ ;
  assign \new_[1425]_  = ~\new_[3824]_  | ~\new_[1432]_ ;
  assign \new_[1426]_  = ~\new_[1432]_ ;
  assign \new_[1427]_  = (~\new_[1554]_  | ~\new_[10283]_ ) & (~\new_[1444]_  | ~\new_[10420]_ );
  assign n646 = \\u5_cmd_r_reg[0] ;
  assign \new_[1429]_  = ~\new_[1434]_ ;
  assign \new_[1430]_  = ~\new_[1434]_ ;
  assign \new_[1431]_  = ~\new_[1434]_ ;
  assign \new_[1432]_  = ~\new_[1434]_ ;
  assign \new_[1433]_  = ~u5_cmd_asserted_reg;
  assign \new_[1434]_  = ~\new_[1443]_ ;
  assign n651 = ~\new_[1445]_ ;
  assign n601 = ~\new_[1445]_ ;
  assign mc_cas_pad_o_ = u7_mc_cas__reg;
  assign \mc_dqm_pad_o[2]  = \\u7_mc_dqm_reg[2] ;
  assign \mc_dqm_pad_o[1]  = \\u7_mc_dqm_reg[1] ;
  assign \mc_dqm_pad_o[0]  = \\u7_mc_dqm_reg[0] ;
  assign \mc_dqm_pad_o[3]  = \\u7_mc_dqm_reg[3] ;
  assign \new_[1442]_  = ~\new_[12619]_  | ~\new_[6336]_  | ~\new_[11266]_ ;
  assign \new_[1443]_  = ~\new_[12224]_  | ~\new_[12619]_ ;
  assign \new_[1444]_  = \\u5_cmd_del_reg[3] ;
  assign \new_[1445]_  = ~\new_[1545]_  & ~\new_[5807]_  & ~\new_[2860]_  & ~\new_[3414]_ ;
  assign n656 = ~\new_[8480]_  | ~\new_[1458]_ ;
  assign n676 = ~\new_[1472]_  | ~\new_[11113]_ ;
  assign n671 = ~\new_[1471]_  | ~\new_[11113]_ ;
  assign n666 = ~\new_[1473]_  | ~\new_[11113]_ ;
  assign n681 = ~\new_[1474]_  | ~\new_[11113]_ ;
  assign wb_ack_o = u6_wb_ack_o_reg;
  assign \new_[1452]_  = \\u5_state_reg[16] ;
  assign \new_[1453]_  = \\u5_timer_reg[0] ;
  assign \new_[1454]_  = \\u5_timer_reg[1] ;
  assign \new_[1455]_  = \\u5_state_reg[2] ;
  assign \new_[1456]_  = \\u5_state_reg[59] ;
  assign n686 = \\u5_cmd_r_reg[3] ;
  assign \new_[1458]_  = ~n721 | ~n5306;
  assign \new_[1459]_  = \\u5_state_reg[17] ;
  assign \new_[1460]_  = \\u5_state_reg[1] ;
  assign \new_[1461]_  = \\u5_state_reg[35] ;
  assign \new_[1462]_  = \\u5_burst_cnt_reg[2] ;
  assign \new_[1463]_  = \\u5_burst_cnt_reg[8] ;
  assign \new_[1464]_  = \\u5_burst_cnt_reg[9] ;
  assign \new_[1465]_  = \\u5_burst_cnt_reg[0] ;
  assign \new_[1466]_  = \\u5_state_reg[21] ;
  assign \new_[1467]_  = \\u5_state_reg[29] ;
  assign \new_[1468]_  = \\u5_state_reg[57] ;
  assign \new_[1469]_  = \\u5_state_reg[0] ;
  assign \new_[1470]_  = \\u5_state_reg[10] ;
  assign \new_[1471]_  = ~\new_[1556]_  & (~\new_[10937]_  | ~\new_[1612]_ );
  assign \new_[1472]_  = ~\new_[1556]_  & (~\new_[10921]_  | ~\new_[1612]_ );
  assign \new_[1473]_  = ~\new_[1556]_  & (~\new_[10865]_  | ~\new_[1612]_ );
  assign \new_[1474]_  = ~\new_[1556]_  & (~\new_[10830]_  | ~\new_[1612]_ );
  assign n691 = ~\new_[1564]_  | ~\new_[9041]_ ;
  assign n711 = \new_[2620]_  | \new_[1549]_ ;
  assign n716 = ~\new_[5382]_  | ~\new_[2635]_  | ~\new_[1576]_ ;
  assign n701 = ~\new_[1548]_  | ~\new_[2256]_ ;
  assign n706 = ~\new_[11741]_  | ~\new_[2256]_ ;
  assign \new_[1480]_  = \\u5_state_reg[15] ;
  assign \new_[1481]_  = \\u5_state_reg[40] ;
  assign \new_[1482]_  = \\u5_burst_cnt_reg[10] ;
  assign \new_[1483]_  = \\u5_state_reg[18] ;
  assign \new_[1484]_  = \\u5_state_reg[20] ;
  assign \new_[1485]_  = \\u5_state_reg[22] ;
  assign \new_[1486]_  = \\u5_state_reg[23] ;
  assign \new_[1487]_  = \\u5_state_reg[24] ;
  assign \new_[1488]_  = \\u5_state_reg[62] ;
  assign \new_[1489]_  = \\u5_state_reg[26] ;
  assign \new_[1490]_  = \\u5_state_reg[27] ;
  assign \new_[1491]_  = \\u5_state_reg[28] ;
  assign \new_[1492]_  = \\u5_state_reg[25] ;
  assign \new_[1493]_  = \\u5_state_reg[30] ;
  assign \new_[1494]_  = \\u5_state_reg[32] ;
  assign \new_[1495]_  = \\u5_state_reg[33] ;
  assign \new_[1496]_  = \\u5_state_reg[38] ;
  assign \new_[1497]_  = \\u5_state_reg[43] ;
  assign \new_[1498]_  = \\u5_state_reg[36] ;
  assign \new_[1499]_  = \\u5_state_reg[46] ;
  assign \new_[1500]_  = \\u5_state_reg[4] ;
  assign \new_[1501]_  = \\u5_state_reg[45] ;
  assign \new_[1502]_  = \\u5_state_reg[52] ;
  assign \new_[1503]_  = \\u5_state_reg[60] ;
  assign \new_[1504]_  = \\u5_state_reg[9] ;
  assign \new_[1505]_  = \\u5_state_reg[13] ;
  assign \new_[1506]_  = \\u5_state_reg[12] ;
  assign \new_[1507]_  = \\u5_state_reg[48] ;
  assign mc_doe_pad_doe_o = u7_mc_data_oe_reg;
  assign n696 = \new_[12055]_  | \new_[1698]_  | \new_[2784]_  | \new_[2744]_ ;
  assign n746 = ~\new_[9674]_  & (~\new_[1602]_  | ~\new_[2237]_ );
  assign n756 = ~\new_[9674]_  & (~\new_[1601]_  | ~\new_[2235]_ );
  assign n726 = ~\new_[12345]_  | ~\new_[2618]_ ;
  assign n731 = ~\new_[1577]_  | ~\new_[1710]_ ;
  assign n741 = \new_[1599]_  | \new_[9674]_ ;
  assign n751 = ~\new_[9674]_  & (~\new_[2064]_  | ~\new_[1603]_ );
  assign n736 = ~\new_[12366]_  | ~\new_[2650]_ ;
  assign n721 = \new_[1554]_ ;
  assign n771 = ~\new_[5380]_  | ~\new_[2664]_  | ~\new_[1609]_ ;
  assign \new_[1519]_  = \\u5_timer_reg[2] ;
  assign wb_err_o = u6_wb_err_reg;
  assign \new_[1521]_  = \\u5_state_reg[37] ;
  assign \new_[1522]_  = \\u5_state_reg[39] ;
  assign \new_[1523]_  = \\u5_state_reg[42] ;
  assign \new_[1524]_  = \\u5_state_reg[41] ;
  assign \new_[1525]_  = \\u5_state_reg[44] ;
  assign \new_[1526]_  = \\u5_state_reg[47] ;
  assign \new_[1527]_  = \\u5_state_reg[51] ;
  assign \new_[1528]_  = \\u5_state_reg[56] ;
  assign \new_[1529]_  = \\u5_state_reg[5] ;
  assign \new_[1530]_  = \\u5_state_reg[61] ;
  assign \new_[1531]_  = \\u5_state_reg[58] ;
  assign \new_[1532]_  = \\u5_state_reg[63] ;
  assign \new_[1533]_  = \\u5_state_reg[64] ;
  assign \new_[1534]_  = \\u5_state_reg[11] ;
  assign \new_[1535]_  = \\u5_state_reg[6] ;
  assign \new_[1536]_  = \\u5_state_reg[7] ;
  assign \new_[1537]_  = \\u5_state_reg[8] ;
  assign \new_[1538]_  = \\u5_state_reg[65] ;
  assign \new_[1539]_  = \\u5_burst_cnt_reg[3] ;
  assign \new_[1540]_  = \\u5_state_reg[14] ;
  assign \new_[1541]_  = \\u5_burst_cnt_reg[1] ;
  assign \new_[1542]_  = \\u5_state_reg[34] ;
  assign \new_[1543]_  = \\u5_state_reg[50] ;
  assign \new_[1544]_  = \\u5_state_reg[55] ;
  assign \new_[1545]_  = ~\new_[7998]_  | ~\new_[12736]_  | ~\new_[1593]_  | ~\new_[6678]_ ;
  assign n796 = ~\new_[9674]_  & (~\new_[2223]_  | ~\new_[1638]_ );
  assign n786 = ~\new_[4209]_  | ~\new_[5023]_  | ~\new_[1629]_  | ~\new_[2674]_ ;
  assign \new_[1548]_  = ~\new_[3482]_  & ~\new_[1610]_ ;
  assign \new_[1549]_  = ~\new_[1977]_  | ~\new_[1653]_  | ~\new_[1634]_  | ~\new_[1859]_ ;
  assign n791 = ~\new_[12355]_  | ~\new_[2651]_ ;
  assign n921 = \new_[1651]_  | \new_[2711]_  | \new_[2863]_  | \new_[2728]_ ;
  assign \new_[1552]_  = \\u5_cmd_del_reg[1] ;
  assign n926 = \new_[2634]_  & \new_[1612]_ ;
  assign \new_[1554]_  = ~\new_[5481]_  | ~\new_[1625]_  | ~\new_[7222]_ ;
  assign n826 = \new_[12186]_  | \new_[2685]_ ;
  assign \new_[1556]_  = ~\new_[1612]_  & (~\new_[3036]_  | ~\new_[10804]_ );
  assign \new_[1557]_  = \\u5_state_reg[19] ;
  assign \new_[1558]_  = \\u5_state_reg[31] ;
  assign \new_[1559]_  = \\u5_state_reg[3] ;
  assign \new_[1560]_  = \\u5_state_reg[49] ;
  assign \new_[1561]_  = \\u5_state_reg[54] ;
  assign \new_[1562]_  = \\u5_state_reg[53] ;
  assign n821 = ~\new_[5379]_  | ~\new_[2682]_  | ~\new_[1633]_ ;
  assign \new_[1564]_  = ~\new_[9932]_  | ~n1151 | ~\new_[1632]_ ;
  assign n871 = \new_[1604]_  | \new_[2652]_ ;
  assign n891 = \new_[1605]_  | \new_[2645]_ ;
  assign n881 = \new_[11905]_  | \new_[2654]_ ;
  assign n896 = \new_[1606]_  | \new_[2656]_ ;
  assign n901 = \new_[1607]_  | \new_[2657]_ ;
  assign n906 = ~\new_[2684]_  | ~\new_[1636]_  | ~\new_[4179]_ ;
  assign n936 = ~\new_[9944]_  & ~\new_[1632]_ ;
  assign n1056 = \new_[1666]_  | \new_[2736]_  | \new_[2785]_  | \new_[2758]_ ;
  assign n931 = ~\new_[11935]_  | ~\new_[2256]_ ;
  assign n1036 = \new_[1667]_  | \new_[1696]_  | \new_[2786]_  | \new_[2742]_ ;
  assign n971 = ~\new_[2660]_  | ~\new_[4869]_  | ~\new_[1635]_  | ~\new_[6325]_ ;
  assign \new_[1576]_  = ~\new_[2813]_  & ~\new_[1637]_ ;
  assign \new_[1577]_  = ~\new_[2673]_  & ~\new_[1639]_ ;
  assign mc_oe_pad_o_ = u7_mc_oe__reg;
  assign \new_[1579]_  = \\u5_burst_cnt_reg[4] ;
  assign \new_[1580]_  = \\u5_burst_cnt_reg[7] ;
  assign \new_[1581]_  = \\u5_burst_cnt_reg[6] ;
  assign \new_[1582]_  = \\u5_burst_cnt_reg[5] ;
  assign n956 = \new_[12144]_  | \new_[2633]_ ;
  assign n961 = \new_[1624]_  | \new_[2653]_ ;
  assign n966 = \new_[12121]_  | \new_[2655]_ ;
  assign n991 = \new_[1626]_  | \new_[2646]_ ;
  assign n981 = \new_[12128]_  | \new_[2683]_ ;
  assign n986 = \new_[1627]_  | \new_[2661]_ ;
  assign n996 = \new_[12136]_  | \new_[2658]_ ;
  assign n1016 = \new_[1631]_  | \new_[2659]_ ;
  assign n1021 = \new_[1628]_  | \new_[2639]_ ;
  assign n951 = \new_[12114]_  | \new_[2626]_ ;
  assign \new_[1593]_  = ~\new_[4526]_  & ~\new_[1622]_ ;
  assign n1001 = \new_[1630]_  | \new_[2662]_ ;
  assign n1026 = \new_[12412]_  | \new_[2663]_ ;
  assign n1011 = \new_[2438]_  | \new_[12158]_ ;
  assign n1006 = \new_[12102]_  | \new_[12041]_  | \new_[2727]_  | \new_[4882]_ ;
  assign n1041 = (~\new_[1641]_  & ~\new_[8917]_ ) | (~\new_[2376]_  & ~\new_[2380]_ );
  assign \new_[1599]_  = ~\new_[2236]_  | (~\new_[1642]_  & ~\new_[9658]_ );
  assign n1031 = (~\new_[1647]_  & ~\new_[8917]_ ) | (~\new_[2380]_  & ~\new_[2377]_ );
  assign \new_[1601]_  = ~\new_[1650]_  | ~\new_[9902]_ ;
  assign \new_[1602]_  = ~\new_[1648]_  | ~\new_[9902]_ ;
  assign \new_[1603]_  = ~\new_[1649]_  | ~\new_[9902]_ ;
  assign \new_[1604]_  = ~\new_[1928]_  | ~\new_[1692]_  | ~\new_[4861]_  | ~\new_[2803]_ ;
  assign \new_[1605]_  = ~\new_[4865]_  | ~\new_[1693]_  | ~\new_[1866]_  | ~\new_[2804]_ ;
  assign \new_[1606]_  = ~\new_[1935]_  | ~\new_[1694]_  | ~\new_[4870]_  | ~\new_[2820]_ ;
  assign \new_[1607]_  = ~\new_[1941]_  | ~\new_[1695]_  | ~\new_[4876]_  | ~\new_[2814]_ ;
  assign n1061 = \\u5_cmd_r_reg[1] ;
  assign \new_[1609]_  = ~\new_[2808]_  & ~\new_[1652]_ ;
  assign \new_[1610]_  = ~\new_[11944]_  & (~\new_[1668]_  | ~\new_[11940]_ );
  assign \new_[1611]_  = \\u5_timer_reg[3] ;
  assign \new_[1612]_  = u5_data_oe_reg;
  assign n1066 = ~\new_[4210]_  | ~\new_[5027]_  | ~\new_[1658]_  | ~\new_[2675]_ ;
  assign n1071 = ~\new_[4212]_  | ~\new_[5051]_  | ~\new_[1660]_  | ~\new_[2676]_ ;
  assign n1081 = ~\new_[4213]_  | ~\new_[5087]_  | ~\new_[1661]_  | ~\new_[2677]_ ;
  assign n1091 = ~\new_[4214]_  | ~\new_[5093]_  | ~\new_[1662]_  | ~\new_[2678]_ ;
  assign n1086 = ~\new_[4215]_  | ~\new_[5096]_  | ~\new_[1663]_  | ~\new_[2679]_ ;
  assign n1116 = ~\new_[8917]_  & (~\new_[1677]_  | ~\new_[1678]_ );
  assign n1111 = ~\new_[8917]_  & (~\new_[1687]_  | ~\new_[1679]_ );
  assign n1096 = ~\new_[1655]_  | ~\new_[11113]_ ;
  assign n1106 = ~\new_[8917]_  & (~\new_[1688]_  | ~\new_[1680]_ );
  assign \new_[1622]_  = \new_[1728]_  | \new_[7577]_  | \new_[12479]_  | \new_[5765]_ ;
  assign n1101 = ~\new_[8917]_  & (~\new_[1686]_  | ~\new_[1676]_ );
  assign \new_[1624]_  = ~\new_[1929]_  | ~\new_[1716]_  | ~\new_[2811]_  | ~\new_[4863]_ ;
  assign \new_[1625]_  = ~\new_[1670]_  & ~\new_[3345]_  & ~\new_[2083]_ ;
  assign \new_[1626]_  = ~\new_[1939]_  | ~\new_[1720]_  | ~\new_[4874]_  | ~\new_[2812]_ ;
  assign \new_[1627]_  = ~\new_[1942]_  | ~\new_[1721]_  | ~\new_[4878]_  | ~\new_[2809]_ ;
  assign \new_[1628]_  = ~\new_[1946]_  | ~\new_[1724]_  | ~\new_[4884]_  | ~\new_[2817]_ ;
  assign \new_[1629]_  = ~\new_[11781]_  & ~\new_[1699]_ ;
  assign \new_[1630]_  = ~\new_[1944]_  | ~\new_[1722]_  | ~\new_[4880]_  | ~\new_[2815]_ ;
  assign \new_[1631]_  = ~\new_[1868]_  | ~\new_[1723]_  | ~\new_[4881]_  | ~\new_[2816]_ ;
  assign \new_[1632]_  = \new_[11866]_  & \new_[9134]_ ;
  assign \new_[1633]_  = ~\new_[2866]_  & ~\new_[1659]_ ;
  assign \new_[1634]_  = ~\new_[11764]_  & ~\new_[2810]_ ;
  assign \new_[1635]_  = ~\new_[2735]_  & ~\new_[1664]_ ;
  assign \new_[1636]_  = ~\new_[2636]_  & ~\new_[1665]_ ;
  assign \new_[1637]_  = ~\new_[1669]_  | ~\new_[1940]_  | ~\new_[1989]_ ;
  assign \new_[1638]_  = ~\new_[1685]_  | ~\new_[9902]_  | ~\new_[1684]_ ;
  assign \new_[1639]_  = ~\new_[1725]_  | ~\new_[3317]_  | ~\new_[6133]_  | ~\new_[4563]_ ;
  assign n1126 = ~\new_[2484]_  | (~\new_[1707]_  & ~\new_[11944]_ );
  assign \new_[1641]_  = ~\new_[1673]_  & (~\new_[11294]_  | ~\new_[1541]_ );
  assign \new_[1642]_  = ~\new_[1674]_  & (~\new_[11293]_  | ~\new_[1462]_ );
  assign \new_[1643]_  = u5_wb_stb_first_reg;
  assign \new_[1644]_  = \\u5_timer2_reg[2] ;
  assign \new_[1645]_  = u5_mem_ack_r_reg;
  assign \new_[1646]_  = ~mem_ack_r_reg;
  assign \new_[1647]_  = ~\new_[1675]_  & (~\new_[11294]_  | ~\new_[1539]_ );
  assign \new_[1648]_  = ~\new_[1681]_  | (~\new_[11294]_  & ~\new_[8861]_ );
  assign \new_[1649]_  = ~\new_[1682]_  | (~\new_[11293]_  & ~\new_[8982]_ );
  assign \new_[1650]_  = ~\new_[1672]_  | (~\new_[11294]_  & ~\new_[1465]_ );
  assign \new_[1651]_  = ~\new_[1703]_  | ~\new_[1835]_  | ~\new_[1930]_ ;
  assign \new_[1652]_  = ~\new_[1700]_  | ~\new_[1938]_  | ~\new_[1988]_ ;
  assign \new_[1653]_  = ~\new_[1697]_  & (~\new_[12064]_  | ~\new_[9848]_ );
  assign n1131 = \new_[1709]_  ? \new_[10283]_  : n1191;
  assign \new_[1655]_  = ~u5_oe__reg;
  assign \new_[1656]_  = \\u5_timer2_reg[1] ;
  assign \new_[1657]_  = \\u5_timer2_reg[3] ;
  assign \new_[1658]_  = ~\new_[1714]_  & ~\new_[1858]_ ;
  assign \new_[1659]_  = ~\new_[1971]_  | ~\new_[1713]_ ;
  assign \new_[1660]_  = ~\new_[1715]_  & ~\new_[1845]_ ;
  assign \new_[1661]_  = ~\new_[1717]_  & ~\new_[1839]_ ;
  assign \new_[1662]_  = ~\new_[1718]_  & ~\new_[11511]_ ;
  assign \new_[1663]_  = ~\new_[1719]_  & ~\new_[1833]_ ;
  assign \new_[1664]_  = ~\new_[1750]_  | ~\new_[1934]_  | ~\new_[2011]_ ;
  assign \new_[1665]_  = ~\new_[1755]_  | ~\new_[1948]_  | ~\new_[2016]_ ;
  assign \new_[1666]_  = ~\new_[2013]_  | ~\new_[1704]_  | ~\new_[1867]_ ;
  assign \new_[1667]_  = ~\new_[3152]_  | ~\new_[5616]_  | ~\new_[1708]_  | ~\new_[1950]_ ;
  assign \new_[1668]_  = ~\new_[5840]_  & (~\new_[1758]_  | ~\new_[6282]_ );
  assign \new_[1669]_  = ~\new_[1757]_  & (~\new_[12064]_  | ~\new_[9871]_ );
  assign \new_[1670]_  = \new_[12230]_  | \new_[6098]_  | \new_[4143]_  | \new_[7303]_ ;
  assign n5881 = u5_cke__reg;
  assign \new_[1672]_  = ~\new_[11293]_  | ~\new_[1465]_ ;
  assign \new_[1673]_  = ~\new_[10335]_  & ~\new_[11293]_ ;
  assign \new_[1674]_  = ~\new_[10005]_  & ~\new_[11293]_ ;
  assign \new_[1675]_  = ~\new_[9720]_  & ~\new_[11295]_ ;
  assign \new_[1676]_  = ~\new_[11295]_  | ~\new_[1579]_ ;
  assign \new_[1677]_  = \new_[11294]_  | \new_[9419]_ ;
  assign \new_[1678]_  = ~\new_[11295]_  | ~\new_[1582]_ ;
  assign \new_[1679]_  = ~\new_[11295]_  | ~\new_[1581]_ ;
  assign \new_[1680]_  = ~\new_[11295]_  | ~\new_[1580]_ ;
  assign \new_[1681]_  = ~\new_[11293]_  | ~\new_[1463]_ ;
  assign \new_[1682]_  = ~\new_[11293]_  | ~\new_[1464]_ ;
  assign n1136 = ~\new_[8258]_  & ~n1151;
  assign \new_[1684]_  = \new_[11293]_  | \new_[9164]_ ;
  assign \new_[1685]_  = ~\new_[11295]_  | ~\new_[11209]_ ;
  assign \new_[1686]_  = \new_[11294]_  | \new_[9363]_ ;
  assign \new_[1687]_  = \new_[11294]_  | \new_[9272]_ ;
  assign \new_[1688]_  = \new_[11294]_  | \new_[9385]_ ;
  assign n1141 = \new_[1763]_  ? \new_[7018]_  : \new_[12762]_ ;
  assign \new_[1690]_  = ~\new_[1741]_  | ~\new_[5882]_ ;
  assign \new_[1691]_  = ~\new_[1749]_  | ~\new_[5893]_ ;
  assign \new_[1692]_  = ~\new_[1745]_  & (~\new_[12628]_  | ~\new_[8507]_ );
  assign \new_[1693]_  = ~\new_[1746]_  & (~\new_[12628]_  | ~\new_[8509]_ );
  assign \new_[1694]_  = ~\new_[1751]_  & (~\new_[8511]_  | ~\new_[11267]_ );
  assign \new_[1695]_  = ~\new_[1752]_  & (~\new_[8516]_  | ~\new_[11267]_ );
  assign \new_[1696]_  = ~\new_[4972]_  | ~\new_[7467]_  | ~\new_[1991]_  | ~\new_[1790]_ ;
  assign \new_[1697]_  = ~\new_[4761]_  | ~\new_[1760]_ ;
  assign \new_[1698]_  = ~\new_[1829]_  | ~\new_[3238]_  | ~\new_[2004]_  | ~\new_[4047]_ ;
  assign \new_[1699]_  = ~\new_[4208]_  | ~\new_[1827]_  | ~\new_[1963]_  | ~\new_[3087]_ ;
  assign \new_[1700]_  = ~\new_[1789]_  & (~\new_[12064]_  | ~\new_[9967]_ );
  assign \new_[1701]_  = ~\new_[1782]_  & (~\new_[12064]_  | ~\new_[10065]_ );
  assign \new_[1702]_  = ~\new_[1783]_  & (~\new_[12064]_  | ~\new_[9849]_ );
  assign \new_[1703]_  = ~\new_[1784]_  & (~\new_[12064]_  | ~\new_[10153]_ );
  assign \new_[1704]_  = ~\new_[1785]_  & (~\new_[12064]_  | ~\new_[9847]_ );
  assign \new_[1705]_  = ~\new_[1786]_  & (~\new_[12064]_  | ~\new_[10050]_ );
  assign \new_[1706]_  = ~\new_[1787]_  & (~\new_[12064]_  | ~\new_[10140]_ );
  assign \new_[1707]_  = ~\new_[2160]_  & (~\new_[1797]_  | ~\new_[6736]_ );
  assign \new_[1708]_  = ~\new_[1788]_  & (~\new_[12064]_  | ~\new_[9953]_ );
  assign \new_[1709]_  = u5_data_oe_r2_reg;
  assign \new_[1710]_  = ~\new_[2666]_  & ~\new_[1793]_ ;
  assign \new_[1711]_  = u5_cke_r_reg;
  assign \new_[1712]_  = \\u5_timer2_reg[5] ;
  assign \new_[1713]_  = ~\new_[1762]_  & (~\new_[12628]_  | ~\new_[8502]_ );
  assign \new_[1714]_  = \new_[1765]_  | \new_[1861]_ ;
  assign \new_[1715]_  = \new_[1766]_  | \new_[2878]_ ;
  assign \new_[1716]_  = ~\new_[1769]_  & (~\new_[12628]_  | ~\new_[8508]_ );
  assign \new_[1717]_  = \new_[1771]_  | \new_[1862]_ ;
  assign \new_[1718]_  = \new_[1772]_  | \new_[1863]_ ;
  assign \new_[1719]_  = \new_[12480]_  | \new_[1864]_ ;
  assign \new_[1720]_  = ~\new_[1774]_  & (~\new_[8514]_  | ~\new_[11267]_ );
  assign \new_[1721]_  = ~\new_[1776]_  & (~\new_[8517]_  | ~\new_[11267]_ );
  assign \new_[1722]_  = ~\new_[1778]_  & (~\new_[8519]_  | ~\new_[12420]_ );
  assign \new_[1723]_  = ~\new_[1780]_  & (~\new_[8727]_  | ~\new_[12628]_ );
  assign \new_[1724]_  = ~\new_[1781]_  & (~\new_[8520]_  | ~\new_[11267]_ );
  assign \new_[1725]_  = ~\new_[1761]_  & (~\new_[7067]_  | ~\new_[9388]_ );
  assign n1161 = ~\new_[2227]_  | (~\new_[1821]_  & ~\new_[5748]_ );
  assign n1166 = \new_[1822]_  ? \new_[7018]_  : \new_[2383]_ ;
  assign \new_[1728]_  = ~\new_[1828]_  | ~\new_[4471]_  | ~\new_[6121]_  | ~\new_[8001]_ ;
  assign n1171 = \new_[1823]_  & \new_[1711]_ ;
  assign \new_[1730]_  = ~\new_[1798]_  & (~\new_[12064]_  | ~\new_[10054]_ );
  assign \new_[1731]_  = ~\new_[1799]_  & (~\new_[12064]_  | ~\new_[9912]_ );
  assign \new_[1732]_  = ~\new_[1800]_  & (~\new_[12064]_  | ~\new_[10053]_ );
  assign \new_[1733]_  = ~\new_[1801]_  & (~\new_[12064]_  | ~\new_[10046]_ );
  assign \new_[1734]_  = ~\new_[1802]_  & (~\new_[12064]_  | ~\new_[9737]_ );
  assign \new_[1735]_  = ~\new_[1803]_  & (~\new_[12064]_  | ~\new_[9854]_ );
  assign \new_[1736]_  = ~\new_[1804]_  & (~\new_[12064]_  | ~\new_[10078]_ );
  assign \new_[1737]_  = ~\new_[1805]_  & (~\new_[12064]_  | ~\new_[9880]_ );
  assign \new_[1738]_  = ~\new_[1806]_  & (~\new_[12064]_  | ~\new_[10081]_ );
  assign \new_[1739]_  = ~\new_[1807]_  & (~\new_[12064]_  | ~\new_[10130]_ );
  assign \new_[1740]_  = ~\new_[1808]_  & (~\new_[12064]_  | ~\new_[10082]_ );
  assign \new_[1741]_  = ~\new_[1809]_  & (~\new_[12064]_  | ~\new_[10061]_ );
  assign \new_[1742]_  = ~\new_[1810]_  & (~\new_[12064]_  | ~\new_[9807]_ );
  assign \new_[1743]_  = ~\new_[1812]_  & (~\new_[12064]_  | ~\new_[10071]_ );
  assign \new_[1744]_  = ~\new_[3989]_  | ~\new_[1846]_  | ~\new_[5754]_  | ~\new_[4763]_ ;
  assign \new_[1745]_  = ~\new_[3994]_  | ~\new_[1847]_  | ~\new_[5757]_  | ~\new_[5272]_ ;
  assign \new_[1746]_  = ~\new_[3996]_  | ~\new_[1848]_  | ~\new_[5759]_  | ~\new_[5274]_ ;
  assign \new_[1747]_  = ~\new_[3997]_  | ~\new_[1849]_  | ~\new_[5760]_  | ~\new_[5275]_ ;
  assign \new_[1748]_  = ~\new_[1814]_  & (~\new_[12064]_  | ~\new_[10118]_ );
  assign \new_[1749]_  = ~\new_[1815]_  & (~\new_[12064]_  | ~\new_[9904]_ );
  assign \new_[1750]_  = ~\new_[1816]_  & (~\new_[12064]_  | ~\new_[9839]_ );
  assign \new_[1751]_  = ~\new_[11883]_  | ~\new_[11839]_  | ~\new_[5762]_  | ~\new_[4765]_ ;
  assign \new_[1752]_  = ~\new_[3813]_  | ~\new_[1852]_  | ~\new_[5770]_  | ~\new_[5289]_ ;
  assign \new_[1753]_  = ~\new_[3815]_  | ~\new_[1853]_  | ~\new_[5772]_  | ~\new_[5291]_ ;
  assign \new_[1754]_  = ~\new_[1818]_  & (~\new_[12064]_  | ~\new_[10107]_ );
  assign \new_[1755]_  = ~\new_[1819]_  & (~\new_[12064]_  | ~\new_[9608]_ );
  assign \new_[1756]_  = ~\new_[1820]_  & (~\new_[12064]_  | ~\new_[10063]_ );
  assign \new_[1757]_  = ~\new_[3811]_  | ~\new_[7009]_  | ~\new_[1851]_  | ~\new_[5898]_ ;
  assign \new_[1758]_  = ~\new_[12024]_  | (~\new_[3703]_  & ~\new_[2552]_ );
  assign \new_[1759]_  = ~\new_[12334]_  | (~\new_[3879]_  & ~\new_[2553]_ );
  assign \new_[1760]_  = ~\new_[1791]_ ;
  assign \new_[1761]_  = ~\new_[3801]_  | ~\new_[4824]_  | ~\new_[1875]_  | ~\new_[5250]_ ;
  assign \new_[1762]_  = ~\new_[3975]_  | ~\new_[1878]_  | ~\new_[4818]_  | ~\new_[5240]_ ;
  assign \new_[1763]_  = ~\new_[4647]_  | ~\new_[1918]_  | ~\new_[5908]_  | ~\new_[2255]_ ;
  assign \new_[1764]_  = ~\new_[1825]_  & (~\new_[4646]_  | ~\new_[9998]_ );
  assign \new_[1765]_  = ~\new_[3970]_  | ~\new_[1874]_  | ~\new_[5750]_  | ~\new_[5253]_ ;
  assign \new_[1766]_  = ~\new_[3982]_  | ~\new_[1884]_  | ~\new_[5753]_  | ~\new_[5263]_ ;
  assign \new_[1767]_  = ~\new_[3992]_  | ~\new_[1893]_  | ~\new_[5755]_  | ~\new_[5270]_ ;
  assign \new_[1768]_  = ~\new_[3993]_  | ~\new_[5756]_  | ~\new_[1894]_  | ~\new_[5271]_ ;
  assign \new_[1769]_  = ~\new_[3995]_  | ~\new_[12279]_  | ~\new_[5758]_  | ~\new_[5273]_ ;
  assign \new_[1770]_  = ~\new_[3806]_  | ~\new_[1895]_  | ~\new_[5761]_  | ~\new_[5276]_ ;
  assign \new_[1771]_  = ~\new_[4000]_  | ~\new_[1896]_  | ~\new_[11448]_  | ~\new_[5278]_ ;
  assign \new_[1772]_  = ~\new_[4003]_  | ~\new_[1899]_  | ~\new_[5764]_  | ~\new_[5281]_ ;
  assign \new_[1773]_  = ~\new_[4005]_  | ~\new_[1900]_  | ~\new_[5767]_  | ~\new_[5284]_ ;
  assign \new_[1774]_  = ~\new_[4006]_  | ~\new_[1902]_  | ~\new_[5768]_  | ~\new_[5286]_ ;
  assign \new_[1775]_  = ~\new_[4008]_  | ~\new_[1903]_  | ~\new_[5769]_  | ~\new_[5288]_ ;
  assign \new_[1776]_  = ~\new_[4009]_  | ~\new_[1904]_  | ~\new_[5771]_  | ~\new_[5290]_ ;
  assign \new_[1777]_  = ~\new_[4011]_  | ~\new_[1905]_  | ~\new_[5774]_  | ~\new_[4767]_ ;
  assign \new_[1778]_  = ~\new_[4013]_  | ~\new_[1906]_  | ~\new_[5775]_  | ~\new_[4768]_ ;
  assign \new_[1779]_  = ~\new_[3817]_  | ~\new_[1908]_  | ~\new_[5777]_  | ~\new_[4769]_ ;
  assign \new_[1780]_  = ~\new_[3818]_  | ~\new_[1909]_  | ~\new_[5778]_  | ~\new_[5295]_ ;
  assign \new_[1781]_  = ~\new_[4016]_  | ~\new_[1911]_  | ~\new_[5779]_  | ~\new_[4770]_ ;
  assign \new_[1782]_  = ~\new_[1840]_  | ~\new_[5255]_  | ~\new_[3972]_ ;
  assign \new_[1783]_  = ~\new_[1844]_  | ~\new_[5262]_  | ~\new_[3980]_ ;
  assign \new_[1784]_  = ~\new_[12450]_  | ~\new_[5277]_  | ~\new_[3999]_ ;
  assign \new_[1785]_  = ~\new_[1850]_  | ~\new_[4766]_  | ~\new_[4004]_ ;
  assign \new_[1786]_  = ~\new_[1854]_  | ~\new_[5292]_  | ~\new_[4010]_ ;
  assign \new_[1787]_  = ~\new_[1855]_  | ~\new_[5294]_  | ~\new_[4015]_ ;
  assign \new_[1788]_  = ~\new_[1856]_  | ~\new_[4771]_  | ~\new_[4019]_ ;
  assign \new_[1789]_  = ~\new_[4174]_  | ~\new_[7015]_  | ~\new_[1901]_  | ~\new_[5808]_ ;
  assign \new_[1790]_  = ~\new_[1826]_  & (~\new_[11864]_  | ~\new_[10136]_ );
  assign \new_[1791]_  = ~\new_[5639]_  & (~\new_[1857]_  | ~\new_[3826]_ );
  assign n1176 = u5_data_oe_r_reg;
  assign \new_[1793]_  = ~\new_[2915]_  | ~\new_[4583]_  | ~\new_[1834]_  | ~\new_[1966]_ ;
  assign n1181 = ~\new_[1830]_  | ~\new_[2649]_ ;
  assign n1186 = ~\new_[2320]_  | ~\new_[1832]_ ;
  assign \new_[1796]_  = \\u5_timer2_reg[4] ;
  assign \new_[1797]_  = ~\new_[2030]_  | ~\new_[1962]_  | ~\new_[2382]_  | ~\new_[3496]_ ;
  assign \new_[1798]_  = ~\new_[1873]_  | ~\new_[5252]_  | ~\new_[3969]_ ;
  assign \new_[1799]_  = ~\new_[12183]_  | ~\new_[5254]_  | ~\new_[3971]_ ;
  assign \new_[1800]_  = ~\new_[1876]_  | ~\new_[5256]_  | ~\new_[3973]_ ;
  assign \new_[1801]_  = ~\new_[1877]_  | ~\new_[5257]_  | ~\new_[3974]_ ;
  assign \new_[1802]_  = ~\new_[1879]_  | ~\new_[5258]_  | ~\new_[3976]_ ;
  assign \new_[1803]_  = ~\new_[1880]_  | ~\new_[5259]_  | ~\new_[3977]_ ;
  assign \new_[1804]_  = ~\new_[1881]_  | ~\new_[5260]_  | ~\new_[3978]_ ;
  assign \new_[1805]_  = ~\new_[1882]_  | ~\new_[5261]_  | ~\new_[3979]_ ;
  assign \new_[1806]_  = ~\new_[1883]_  | ~\new_[5241]_  | ~\new_[3981]_ ;
  assign \new_[1807]_  = ~\new_[1885]_  | ~\new_[5264]_  | ~\new_[3983]_ ;
  assign \new_[1808]_  = ~\new_[1886]_  | ~\new_[5265]_  | ~\new_[3984]_ ;
  assign \new_[1809]_  = ~\new_[4762]_  | ~\new_[1887]_  | ~\new_[3985]_ ;
  assign \new_[1810]_  = ~\new_[1888]_  | ~\new_[5266]_  | ~\new_[3987]_ ;
  assign \new_[1811]_  = ~\new_[1889]_  | ~\new_[5267]_  | ~\new_[3803]_ ;
  assign \new_[1812]_  = ~\new_[1890]_  | ~\new_[5268]_  | ~\new_[3988]_ ;
  assign \new_[1813]_  = ~\new_[1891]_  | ~\new_[5269]_  | ~\new_[3804]_ ;
  assign \new_[1814]_  = ~\new_[1897]_  | ~\new_[5279]_  | ~\new_[4001]_ ;
  assign \new_[1815]_  = ~\new_[4764]_  | ~\new_[1898]_  | ~\new_[4002]_ ;
  assign \new_[1816]_  = ~\new_[12546]_  | ~\new_[5280]_  | ~\new_[3809]_ ;
  assign \new_[1817]_  = ~\new_[1910]_  | ~\new_[5296]_  | ~\new_[3819]_ ;
  assign \new_[1818]_  = ~\new_[1913]_  | ~\new_[5298]_  | ~\new_[4017]_ ;
  assign \new_[1819]_  = ~\new_[1912]_  | ~\new_[5297]_  | ~\new_[3821]_ ;
  assign \new_[1820]_  = ~\new_[1914]_  | ~\new_[5299]_  | ~\new_[4018]_ ;
  assign \new_[1821]_  = \new_[1838]_  & \new_[2255]_ ;
  assign \new_[1822]_  = ~\new_[2485]_  | (~\new_[1919]_  & ~\new_[6159]_ );
  assign \new_[1823]_  = \new_[1915]_  ? \new_[7072]_  : \new_[2726]_ ;
  assign \new_[1824]_  = ~\new_[1860]_  | ~\new_[6282]_ ;
  assign \new_[1825]_  = ~\new_[4646]_  & (~\new_[1957]_  | ~\new_[1954]_ );
  assign \new_[1826]_  = ~\new_[7330]_  | ~\new_[4288]_  | ~\new_[1870]_  | ~\new_[4544]_ ;
  assign \new_[1827]_  = ~\new_[1871]_  & ~\new_[3698]_ ;
  assign \new_[1828]_  = ~\new_[1872]_  | ~\new_[5242]_ ;
  assign \new_[1829]_  = ~\new_[1920]_  & (~\new_[7077]_  | ~\new_[9979]_ );
  assign \new_[1830]_  = ~\new_[1951]_  | ~\new_[6809]_  | ~\new_[5639]_ ;
  assign n1191 = ~\new_[7681]_  | ~\new_[4453]_  | ~\new_[1921]_  | ~\new_[6316]_ ;
  assign \new_[1832]_  = ~\new_[1994]_  | ~\new_[6738]_  | ~\new_[6123]_  | ~\new_[5908]_ ;
  assign \new_[1833]_  = ~\new_[7345]_  | ~\new_[1987]_  | ~\new_[2818]_  | ~\new_[6143]_ ;
  assign \new_[1834]_  = ~\new_[1922]_  & (~\new_[11997]_  | ~\new_[12306]_ );
  assign \new_[1835]_  = ~\new_[1923]_  & (~\new_[11997]_  | ~\new_[10084]_ );
  assign n1196 = ~\new_[2427]_  | (~\new_[4809]_  & ~\new_[1961]_ );
  assign \new_[1837]_  = ~\new_[11588]_ ;
  assign \new_[1838]_  = ~\new_[1956]_  & (~\new_[6642]_  | ~\new_[11750]_ );
  assign \new_[1839]_  = ~\new_[2028]_  | ~\new_[12384]_  | ~\new_[2882]_  | ~\new_[5891]_ ;
  assign \new_[1840]_  = ~\new_[12553]_  | ~\new_[11348]_  | ~\new_[11840]_  | ~\new_[11292]_ ;
  assign \new_[1841]_  = \\u5_timer2_reg[0] ;
  assign \new_[1842]_  = \\u5_timer2_reg[8] ;
  assign \new_[1843]_  = \\u5_timer2_reg[7] ;
  assign \new_[1844]_  = ~\new_[12553]_  | ~\new_[10808]_  | ~\new_[11840]_  | ~\new_[11292]_ ;
  assign \new_[1845]_  = ~\new_[6635]_  | ~\new_[2039]_  | ~\new_[1979]_  | ~\new_[3091]_ ;
  assign \new_[1846]_  = ~\new_[12695]_  | ~\new_[9785]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[1847]_  = ~\new_[12695]_  | ~n5021 | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1848]_  = ~\new_[12695]_  | ~\new_[10164]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1849]_  = ~\new_[12553]_  | ~\new_[11363]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1850]_  = ~\new_[12553]_  | ~\new_[12598]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1851]_  = ~\new_[12695]_  | ~\new_[11323]_  | ~\new_[12451]_  | ~\new_[11840]_ ;
  assign \new_[1852]_  = ~\new_[12553]_  | ~\new_[11328]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1853]_  = ~\new_[12695]_  | ~\new_[11356]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1854]_  = ~\new_[12553]_  | ~\new_[10419]_  | ~\new_[11840]_  | ~\new_[11292]_ ;
  assign \new_[1855]_  = ~\new_[12695]_  | ~\new_[11526]_  | ~\new_[11840]_  | ~\new_[11292]_ ;
  assign \new_[1856]_  = ~\new_[12553]_  | ~\new_[10634]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[1857]_  = ~\new_[4187]_  & (~\new_[2003]_  | ~\new_[2062]_ );
  assign \new_[1858]_  = ~\new_[6576]_  | ~\new_[2031]_  | ~\new_[2819]_  | ~\new_[5907]_ ;
  assign \new_[1859]_  = ~\new_[1960]_  & (~\new_[11997]_  | ~\new_[9975]_ );
  assign \new_[1860]_  = ~\new_[2428]_  & (~\new_[1986]_  | ~\new_[3879]_ );
  assign \new_[1861]_  = ~\new_[5950]_  | ~\new_[1965]_  | ~\new_[3382]_ ;
  assign \new_[1862]_  = ~\new_[5951]_  | ~\new_[1931]_  | ~\new_[3384]_ ;
  assign \new_[1863]_  = ~\new_[5957]_  | ~\new_[1936]_  | ~\new_[3386]_ ;
  assign \new_[1864]_  = ~\new_[5958]_  | ~\new_[1937]_  | ~\new_[3387]_ ;
  assign \new_[1865]_  = ~\new_[7440]_  | ~\new_[4471]_  | ~\new_[2027]_  | ~\new_[7564]_ ;
  assign \new_[1866]_  = ~\new_[10164]_  | ~\new_[12606]_  | ~\new_[12635]_ ;
  assign \new_[1867]_  = ~\new_[1993]_  | ~\new_[12602]_ ;
  assign \new_[1868]_  = ~\new_[9946]_  | ~\new_[12606]_  | ~\new_[12641]_ ;
  assign \new_[1869]_  = \new_[1995]_  & \new_[2072]_ ;
  assign \new_[1870]_  = ~\new_[1999]_  & (~\new_[9574]_  | ~\new_[12792]_ );
  assign \new_[1871]_  = ~\new_[1997]_  | (~\new_[7020]_  & ~\new_[12003]_ );
  assign \new_[1872]_  = ~\new_[1996]_  | ~\new_[12508]_ ;
  assign \new_[1873]_  = ~\new_[12553]_  | ~\new_[10827]_  | ~\new_[12660]_  | ~\new_[11292]_ ;
  assign \new_[1874]_  = ~\new_[12695]_  | ~\new_[10922]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1875]_  = ~\new_[12553]_  | ~\new_[10743]_  | ~\new_[12661]_  | ~\new_[12451]_ ;
  assign \new_[1876]_  = ~\new_[12553]_  | ~\new_[10928]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1877]_  = ~\new_[12553]_  | ~\new_[9997]_  | ~\new_[12660]_  | ~\new_[11292]_ ;
  assign \new_[1878]_  = ~\new_[12695]_  | ~\new_[11576]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[1879]_  = ~\new_[12553]_  | ~\new_[9379]_  | ~\new_[12660]_  | ~\new_[11292]_ ;
  assign \new_[1880]_  = ~\new_[12553]_  | ~\new_[11332]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1881]_  = ~\new_[12553]_  | ~\new_[10177]_  | ~\new_[12661]_  | ~\new_[12451]_ ;
  assign \new_[1882]_  = ~\new_[12695]_  | ~\new_[11343]_  | ~\new_[12661]_  | ~\new_[12451]_ ;
  assign \new_[1883]_  = ~\new_[12695]_  | ~\new_[11340]_  | ~\new_[12659]_  | ~\new_[11292]_ ;
  assign \new_[1884]_  = ~\new_[12695]_  | ~\new_[11492]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1885]_  = ~\new_[12553]_  | ~\new_[10243]_  | ~\new_[12659]_  | ~\new_[11292]_ ;
  assign \new_[1886]_  = ~\new_[12553]_  | ~\new_[11320]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1887]_  = ~\new_[12553]_  | ~\new_[10938]_  | ~\new_[12661]_  | ~\new_[12451]_ ;
  assign \new_[1888]_  = ~\new_[12553]_  | ~\new_[9913]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1889]_  = ~\new_[12695]_  | ~\new_[11298]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1890]_  = ~\new_[12553]_  | ~\new_[11316]_  | ~\new_[12659]_  | ~\new_[12451]_ ;
  assign \new_[1891]_  = ~\new_[12553]_  | ~\new_[12089]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1892]_  = ~\new_[12695]_  | ~\new_[10108]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[1893]_  = ~\new_[12695]_  | ~\new_[10802]_  | ~\new_[12660]_  | ~\new_[12451]_ ;
  assign \new_[1894]_  = ~\new_[12553]_  | ~\new_[12093]_  | ~\new_[12451]_  | ~\new_[12660]_ ;
  assign \new_[1895]_  = ~\new_[12553]_  | ~\new_[10411]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[1896]_  = ~\new_[12553]_  | ~\new_[10496]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[1897]_  = ~\new_[12553]_  | ~\new_[10902]_  | ~\new_[12659]_  | ~\new_[12451]_ ;
  assign \new_[1898]_  = ~\new_[12553]_  | ~\new_[9903]_  | ~\new_[12661]_  | ~\new_[12451]_ ;
  assign \new_[1899]_  = ~\new_[12553]_  | ~\new_[10250]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[1900]_  = ~\new_[12695]_  | ~\new_[12610]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[1901]_  = ~\new_[12695]_  | ~\new_[11337]_  | ~\new_[12451]_  | ~\new_[11840]_ ;
  assign \new_[1902]_  = ~\new_[12695]_  | ~\new_[11353]_  | ~\new_[12659]_  | ~\new_[12278]_ ;
  assign \new_[1903]_  = ~\new_[12553]_  | ~\new_[10955]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1904]_  = ~\new_[12695]_  | ~\new_[11366]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[1905]_  = ~\new_[12553]_  | ~\new_[11310]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[1906]_  = ~\new_[12695]_  | ~\new_[11313]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[1907]_  = ~\new_[12695]_  | ~\new_[11361]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[1908]_  = ~\new_[12553]_  | ~\new_[10933]_  | ~\new_[12660]_  | ~\new_[12451]_ ;
  assign \new_[1909]_  = ~\new_[12553]_  | ~\new_[9946]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[1910]_  = ~\new_[12695]_  | ~\new_[12044]_  | ~\new_[12660]_  | ~\new_[11292]_ ;
  assign \new_[1911]_  = ~\new_[12695]_  | ~\new_[10960]_  | ~\new_[12659]_  | ~\new_[12278]_ ;
  assign \new_[1912]_  = ~\new_[12695]_  | ~\new_[10509]_  | ~\new_[11292]_  | ~\new_[11840]_ ;
  assign \new_[1913]_  = ~\new_[12695]_  | ~\new_[10526]_  | ~\new_[12661]_  | ~\new_[12451]_ ;
  assign \new_[1914]_  = ~\new_[12553]_  | ~\new_[10919]_  | ~\new_[12660]_  | ~\new_[11292]_ ;
  assign \new_[1915]_  = \new_[7708]_  ? \new_[2012]_  : n5881;
  assign \new_[1916]_  = ~\new_[2000]_  & (~\new_[11997]_  | ~\new_[9621]_ );
  assign \new_[1917]_  = ~\new_[2001]_  & (~\new_[11997]_  | ~\new_[9586]_ );
  assign \new_[1918]_  = ~\new_[2244]_  & (~\new_[2018]_  | ~\new_[6738]_ );
  assign \new_[1919]_  = ~\new_[2246]_  & (~\new_[2019]_  | ~\new_[6738]_ );
  assign \new_[1920]_  = ~\new_[1958]_ ;
  assign \new_[1921]_  = ~\new_[7242]_  & ~\new_[1992]_ ;
  assign \new_[1922]_  = ~\new_[6287]_  | ~\new_[2006]_ ;
  assign \new_[1923]_  = ~\new_[1984]_  | (~\new_[6827]_  & ~\new_[10150]_ );
  assign \new_[1924]_  = ~\new_[10938]_  | ~\new_[12602]_  | ~\new_[12645]_ ;
  assign \new_[1925]_  = ~\new_[9913]_  | ~\new_[12606]_  | ~\new_[12638]_ ;
  assign \new_[1926]_  = ~\new_[11316]_  | ~\new_[12604]_  | ~\new_[12635]_ ;
  assign \new_[1927]_  = ~\new_[9785]_  | ~\new_[12604]_  | ~\new_[12643]_ ;
  assign \new_[1928]_  = ~n5021 | ~\new_[12606]_  | ~\new_[12641]_ ;
  assign \new_[1929]_  = ~\new_[12567]_  | ~\new_[12603]_  | ~\new_[12636]_ ;
  assign \new_[1930]_  = ~\new_[12453]_  | ~\new_[12604]_  | ~\new_[12645]_ ;
  assign \new_[1931]_  = ~\new_[10496]_  | ~\new_[12606]_  | ~\new_[12635]_ ;
  assign \new_[1932]_  = ~\new_[10902]_  | ~\new_[12606]_  | ~\new_[12639]_ ;
  assign \new_[1933]_  = ~\new_[9903]_  | ~\new_[12602]_  | ~\new_[12645]_ ;
  assign \new_[1934]_  = ~\new_[9648]_  | ~\new_[12603]_  | ~\new_[12638]_ ;
  assign \new_[1935]_  = ~\new_[9674]_  | ~\new_[12606]_  | ~\new_[12641]_ ;
  assign \new_[1936]_  = ~\new_[10250]_  | ~\new_[12606]_  | ~\new_[12636]_ ;
  assign \new_[1937]_  = ~\new_[12755]_  | ~\new_[12606]_  | ~\new_[12636]_ ;
  assign \new_[1938]_  = ~\new_[11337]_  | ~\new_[12606]_  | ~\new_[12636]_ ;
  assign \new_[1939]_  = ~\new_[11353]_  | ~\new_[12602]_  | ~\new_[12646]_ ;
  assign \new_[1940]_  = ~\new_[11323]_  | ~\new_[12603]_  | ~\new_[12636]_ ;
  assign \new_[1941]_  = ~\new_[11328]_  | ~\new_[12602]_  | ~\new_[12641]_ ;
  assign \new_[1942]_  = ~\new_[11367]_  | ~\new_[12602]_  | ~\new_[12646]_ ;
  assign \new_[1943]_  = ~\new_[10419]_  | ~\new_[12606]_  | ~\new_[12635]_ ;
  assign \new_[1944]_  = ~\new_[11313]_  | ~\new_[12602]_  | ~\new_[12646]_ ;
  assign \new_[1945]_  = ~\new_[11526]_  | ~\new_[12603]_  | ~\new_[12636]_ ;
  assign \new_[1946]_  = ~\new_[10960]_  | ~\new_[12606]_  | ~\new_[12646]_ ;
  assign \new_[1947]_  = ~\new_[10526]_  | ~\new_[12604]_  | ~\new_[12636]_ ;
  assign \new_[1948]_  = ~\new_[10509]_  | ~\new_[12602]_  | ~\new_[12641]_ ;
  assign \new_[1949]_  = ~\new_[10919]_  | ~\new_[12604]_  | ~\new_[12635]_ ;
  assign \new_[1950]_  = ~\new_[10634]_  | ~\new_[12602]_  | ~\new_[12641]_ ;
  assign \new_[1951]_  = \new_[1711]_  ? \new_[2051]_  : \new_[7708]_ ;
  assign n1211 = ~\new_[2025]_  | ~\new_[2250]_ ;
  assign n1206 = ~\new_[2026]_  | ~\new_[2322]_ ;
  assign \new_[1954]_  = ~\new_[12721]_  | ~\new_[9998]_  | ~\new_[2077]_  | ~\new_[11814]_ ;
  assign \new_[1955]_  = \\u5_timer2_reg[6] ;
  assign \new_[1956]_  = (~\new_[2047]_  & ~\new_[7186]_ ) | (~\new_[6685]_  & ~\new_[2486]_ );
  assign \new_[1957]_  = ~\new_[2029]_  | ~\new_[2217]_ ;
  assign \new_[1958]_  = ~\new_[11776]_  | ~\new_[10119]_  | ~\new_[2060]_  | ~\new_[2048]_ ;
  assign n1201 = ~\new_[1998]_ ;
  assign \new_[1960]_  = ~\new_[6288]_  | ~\new_[2037]_ ;
  assign \new_[1961]_  = ~\new_[2140]_  & (~\new_[2054]_  | ~\new_[7426]_ );
  assign \new_[1962]_  = ~\new_[9205]_  | ~\new_[2024]_  | ~\new_[3703]_ ;
  assign \new_[1963]_  = ~\new_[10291]_  | ~\new_[12603]_  | ~\new_[12638]_ ;
  assign \new_[1964]_  = ~\new_[10827]_  | ~\new_[12606]_  | ~\new_[12639]_ ;
  assign \new_[1965]_  = ~\new_[10922]_  | ~\new_[12606]_  | ~\new_[12647]_ ;
  assign \new_[1966]_  = ~\new_[9658]_  | ~\new_[12602]_  | ~\new_[12641]_ ;
  assign \new_[1967]_  = ~\new_[11355]_  | ~\new_[12606]_  | ~\new_[12647]_ ;
  assign \new_[1968]_  = ~\new_[11348]_  | ~\new_[12604]_  | ~\new_[12635]_ ;
  assign \new_[1969]_  = ~\new_[10928]_  | ~\new_[12602]_  | ~\new_[12647]_ ;
  assign \new_[1970]_  = ~\new_[9997]_  | ~\new_[12604]_  | ~\new_[12635]_ ;
  assign \new_[1971]_  = ~\new_[11576]_  | ~\new_[12604]_  | ~\new_[12644]_ ;
  assign \new_[1972]_  = ~\new_[9379]_  | ~\new_[12603]_  | ~\new_[12635]_ ;
  assign \new_[1973]_  = ~\new_[11332]_  | ~\new_[12606]_  | ~\new_[12635]_ ;
  assign \new_[1974]_  = ~\new_[10177]_  | ~\new_[12606]_  | ~\new_[12638]_ ;
  assign \new_[1975]_  = ~\new_[11343]_  | ~\new_[12603]_  | ~\new_[12647]_ ;
  assign \new_[1976]_  = ~\new_[10808]_  | ~\new_[12603]_  | ~\new_[12639]_ ;
  assign \new_[1977]_  = ~\new_[10818]_  | ~\new_[12604]_  | ~\new_[12644]_ ;
  assign \new_[1978]_  = ~\new_[11340]_  | ~\new_[12603]_  | ~\new_[12635]_ ;
  assign \new_[1979]_  = ~\new_[11492]_  | ~\new_[12606]_  | ~\new_[12638]_ ;
  assign \new_[1980]_  = ~\new_[10243]_  | ~\new_[12604]_  | ~\new_[12635]_ ;
  assign \new_[1981]_  = ~\new_[11320]_  | ~\new_[12606]_  | ~\new_[12638]_ ;
  assign \new_[1982]_  = ~\new_[9913]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[1983]_  = ~\new_[11316]_  | ~\new_[12629]_  | ~\new_[11777]_ ;
  assign \new_[1984]_  = ~\new_[12453]_  | ~\new_[12420]_  | ~\new_[11777]_ ;
  assign \new_[1985]_  = ~\new_[10902]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[1986]_  = \new_[2065]_  ? \new_[12338]_  : \new_[2071]_ ;
  assign \new_[1987]_  = ~\new_[12755]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[1988]_  = ~\new_[11337]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[1989]_  = ~\new_[11323]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[1990]_  = ~\new_[11777]_  | ~\new_[2050]_  | ~\new_[2218]_ ;
  assign \new_[1991]_  = ~\new_[10634]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[1992]_  = ~\new_[4976]_  | ~\new_[6620]_  | ~\new_[2053]_  | ~\new_[7421]_ ;
  assign \new_[1993]_  = ~\new_[12638]_  | ~\new_[12599]_ ;
  assign \new_[1994]_  = ~\new_[2052]_  & (~\new_[2386]_  | ~\new_[9648]_ );
  assign \new_[1995]_  = ~\new_[2057]_  & (~\new_[11885]_  | ~\new_[10291]_ );
  assign \new_[1996]_  = ~\new_[12512]_  | ~\new_[5652]_  | ~\new_[12722]_ ;
  assign \new_[1997]_  = ~\new_[2076]_  | ~\new_[8311]_  | ~\new_[2060]_  | ~\new_[11776]_ ;
  assign \new_[1998]_  = ~\new_[2046]_  & (~\new_[2429]_  | ~\new_[7018]_ );
  assign \new_[1999]_  = ~\new_[7078]_  & (~\new_[2061]_  | ~\new_[10167]_ );
  assign \new_[2000]_  = ~\new_[2042]_  | (~\new_[6829]_  & ~\new_[9924]_ );
  assign \new_[2001]_  = ~\new_[2045]_  | (~\new_[6829]_  & ~\new_[9742]_ );
  assign \new_[2002]_  = ~\new_[2048]_  | ~\new_[10200]_ ;
  assign \new_[2003]_  = ~\new_[2217]_  & ~\new_[12720]_ ;
  assign \new_[2004]_  = ~\new_[10838]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2005]_  = ~\new_[10827]_  | ~\new_[12629]_  | ~\new_[11777]_ ;
  assign \new_[2006]_  = ~\new_[9658]_  | ~\new_[12420]_  | ~\new_[11777]_ ;
  assign \new_[2007]_  = ~\new_[10928]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[2008]_  = ~\new_[9997]_  | ~\new_[12630]_  | ~\new_[11777]_ ;
  assign \new_[2009]_  = ~\new_[11332]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2010]_  = ~\new_[11343]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[2011]_  = ~\new_[9648]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2012]_  = ~\new_[2927]_  | ~\new_[2152]_  | ~\new_[2218]_ ;
  assign \new_[2013]_  = ~\new_[12598]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2014]_  = ~\new_[10419]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2015]_  = ~\new_[11526]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2016]_  = ~\new_[10509]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[2017]_  = ~\new_[10919]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2018]_  = \new_[2245]_  | \new_[2058]_ ;
  assign \new_[2019]_  = \new_[2247]_  | \new_[2059]_ ;
  assign n1216 = ~\new_[2248]_  | (~\new_[2079]_  & ~\new_[7444]_ );
  assign \new_[2021]_  = \new_[12640]_  & \new_[12273]_ ;
  assign \new_[2022]_  = \new_[12640]_  & \new_[11735]_ ;
  assign \new_[2023]_  = \new_[12636]_  & \new_[10108]_ ;
  assign \new_[2024]_  = \new_[12217]_  ^ \new_[2141]_ ;
  assign \new_[2025]_  = \new_[2068]_  | \new_[5748]_ ;
  assign \new_[2026]_  = \new_[2069]_  | \new_[5748]_ ;
  assign \new_[2027]_  = ~\new_[12233]_  | (~\new_[2142]_  & ~\new_[5348]_ );
  assign \new_[2028]_  = (~\new_[12628]_  | ~\new_[8515]_ ) & (~\new_[12385]_  | ~\new_[10496]_ );
  assign \new_[2029]_  = \new_[11814]_  & \new_[12721]_ ;
  assign \new_[2030]_  = ~\new_[2063]_  | ~\new_[3879]_ ;
  assign \new_[2031]_  = ~\new_[10922]_  | ~\new_[12629]_  | ~\new_[11777]_ ;
  assign \new_[2032]_  = ~\new_[11355]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[2033]_  = ~\new_[11348]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[2034]_  = ~\new_[9379]_  | ~\new_[12420]_  | ~\new_[11777]_ ;
  assign \new_[2035]_  = ~\new_[10177]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2036]_  = ~\new_[10808]_  | ~\new_[11268]_  | ~\new_[11777]_ ;
  assign \new_[2037]_  = ~\new_[10818]_  | ~\new_[12420]_  | ~\new_[11777]_ ;
  assign \new_[2038]_  = ~\new_[11340]_  | ~\new_[12420]_  | ~\new_[11777]_ ;
  assign \new_[2039]_  = ~\new_[11492]_  | ~\new_[12629]_  | ~\new_[11777]_ ;
  assign \new_[2040]_  = ~\new_[10243]_  | ~\new_[12630]_  | ~\new_[11777]_ ;
  assign \new_[2041]_  = ~\new_[11320]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2042]_  = ~\new_[10938]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2043]_  = ~\new_[11735]_  | ~\new_[12420]_  | ~\new_[11777]_ ;
  assign \new_[2044]_  = ~\new_[10108]_  | ~\new_[12630]_  | ~\new_[11777]_ ;
  assign \new_[2045]_  = ~\new_[9903]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[2046]_  = ~\new_[5748]_  & (~\new_[2150]_  | ~\new_[2255]_ );
  assign \new_[2047]_  = (~\new_[2148]_  | ~\new_[12384]_ ) & (~\new_[12674]_  | ~\new_[7443]_ );
  assign \new_[2048]_  = ~\new_[2076]_  & ~n3951;
  assign \new_[2049]_  = ~\new_[2146]_  & (~\new_[2152]_  | ~\new_[10291]_ );
  assign \new_[2050]_  = ~\new_[7564]_  & (~\new_[2152]_  | ~\new_[10715]_ );
  assign \new_[2051]_  = ~\new_[2084]_  & ~\new_[10640]_ ;
  assign \new_[2052]_  = ~\new_[2088]_  & ~\new_[9648]_ ;
  assign \new_[2053]_  = ~\new_[2083]_  & (~\new_[6975]_  | ~\new_[3940]_ );
  assign \new_[2054]_  = ~\new_[2226]_  | ~\new_[2087]_ ;
  assign \new_[2055]_  = u5_ap_en_reg;
  assign \new_[2056]_  = \\u5_timer_reg[5] ;
  assign \new_[2057]_  = ~\new_[2143]_  & ~\new_[6091]_ ;
  assign \new_[2058]_  = \new_[2149]_  & \new_[12384]_ ;
  assign \new_[2059]_  = \new_[2151]_  & \new_[12384]_ ;
  assign \new_[2060]_  = \new_[11773]_  & \new_[2147]_ ;
  assign \new_[2061]_  = ~n3951 | ~\new_[2147]_  | ~\new_[11776]_ ;
  assign \new_[2062]_  = ~\new_[4926]_  & (~\new_[7520]_  | ~\new_[2219]_ );
  assign \new_[2063]_  = (~\new_[12217]_  & ~\new_[11474]_  & ~\new_[12338]_ ) | (~\new_[12338]_  & ~\new_[3905]_  & ~\new_[2239]_ );
  assign \new_[2064]_  = ~\new_[2156]_  | ~\new_[9658]_ ;
  assign \new_[2065]_  = ~\new_[2159]_  | (~\new_[3905]_  & ~\new_[2234]_ );
  assign \new_[2066]_  = ~\new_[2153]_  & (~\new_[2385]_  | ~\new_[10964]_ );
  assign \new_[2067]_  = ~\new_[2154]_  & (~\new_[2434]_  | ~\new_[10964]_ );
  assign \new_[2068]_  = \new_[2157]_  | \new_[7444]_ ;
  assign \new_[2069]_  = \new_[2158]_  | \new_[7444]_ ;
  assign \new_[2070]_  = \\u5_timer_reg[4] ;
  assign \new_[2071]_  = \new_[11416]_  ^ \new_[11820]_ ;
  assign \new_[2072]_  = ~\new_[12549]_  | ~\new_[12723]_  | ~\new_[11814]_ ;
  assign \new_[2073]_  = ~\\u0_tms_reg[21] ;
  assign \new_[2074]_  = ~\\u0_tms_reg[5] ;
  assign \new_[2075]_  = \\u0_tms_reg[9] ;
  assign \new_[2076]_  = \new_[12520]_  & \new_[11418]_ ;
  assign \new_[2077]_  = \new_[2219]_  & \new_[12695]_ ;
  assign \new_[2078]_  = ~\\u0_tms_reg[27] ;
  assign \new_[2079]_  = ~\new_[5908]_  | ~\new_[6738]_  | ~\new_[6733]_  | ~\new_[2242]_ ;
  assign n1221 = (~\new_[2235]_  & ~\new_[11510]_ ) | (~\new_[10119]_  & ~\new_[9658]_ );
  assign \new_[2081]_  = \\u0_tms_reg[1] ;
  assign \new_[2082]_  = ~\\u0_tms_reg[16] ;
  assign \new_[2083]_  = ~\new_[8002]_  & (~\new_[2318]_  | ~\new_[2243]_ );
  assign \new_[2084]_  = ~\new_[2152]_ ;
  assign \new_[2085]_  = \\u0_sp_tms_reg[9] ;
  assign n1226 = ~\new_[3481]_  & (~\new_[2254]_  | ~\new_[3241]_ );
  assign \new_[2087]_  = ~\new_[2220]_  & (~\new_[8391]_  | ~\new_[9566]_ );
  assign \new_[2088]_  = ~\new_[2221]_  | (~\new_[8385]_  & ~\new_[10108]_ );
  assign \new_[2089]_  = ~\\u0_sp_tms_reg[26] ;
  assign \new_[2090]_  = ~\\u0_sp_tms_reg[5] ;
  assign \new_[2091]_  = ~\\u0_sp_tms_reg[20] ;
  assign \new_[2092]_  = ~\\u0_sp_tms_reg[23] ;
  assign \new_[2093]_  = ~\\u0_sp_tms_reg[11] ;
  assign \new_[2094]_  = \\u0_sp_tms_reg[0] ;
  assign \new_[2095]_  = ~\\u0_sp_tms_reg[10] ;
  assign \new_[2096]_  = ~\\u0_sp_tms_reg[12] ;
  assign \new_[2097]_  = ~\\u0_sp_tms_reg[13] ;
  assign \new_[2098]_  = ~\\u0_sp_tms_reg[14] ;
  assign \new_[2099]_  = ~\\u0_sp_tms_reg[15] ;
  assign \new_[2100]_  = ~\\u0_sp_tms_reg[17] ;
  assign \new_[2101]_  = ~\\u0_sp_tms_reg[18] ;
  assign \new_[2102]_  = ~\\u0_sp_tms_reg[19] ;
  assign \new_[2103]_  = \\u0_sp_tms_reg[1] ;
  assign \new_[2104]_  = ~\\u0_sp_tms_reg[21] ;
  assign \new_[2105]_  = ~\\u0_sp_tms_reg[22] ;
  assign \new_[2106]_  = ~\\u0_sp_tms_reg[24] ;
  assign \new_[2107]_  = ~\\u0_sp_tms_reg[27] ;
  assign \new_[2108]_  = \\u0_sp_tms_reg[2] ;
  assign \new_[2109]_  = ~\\u0_sp_tms_reg[25] ;
  assign \new_[2110]_  = ~\\u0_sp_tms_reg[3] ;
  assign \new_[2111]_  = ~\\u0_sp_tms_reg[4] ;
  assign \new_[2112]_  = ~\\u0_sp_tms_reg[6] ;
  assign \new_[2113]_  = ~\\u0_sp_tms_reg[7] ;
  assign \new_[2114]_  = ~\\u0_sp_tms_reg[8] ;
  assign \new_[2115]_  = ~\\u0_tms_reg[11] ;
  assign \new_[2116]_  = \\u0_tms_reg[0] ;
  assign \new_[2117]_  = ~\\u0_tms_reg[10] ;
  assign \new_[2118]_  = ~\\u0_tms_reg[12] ;
  assign \new_[2119]_  = ~\\u0_tms_reg[13] ;
  assign \new_[2120]_  = ~\\u0_tms_reg[15] ;
  assign \new_[2121]_  = ~\\u0_tms_reg[14] ;
  assign \new_[2122]_  = ~\\u0_tms_reg[17] ;
  assign \new_[2123]_  = ~\\u0_tms_reg[18] ;
  assign \new_[2124]_  = ~\\u0_tms_reg[19] ;
  assign \new_[2125]_  = ~\\u0_tms_reg[20] ;
  assign \new_[2126]_  = ~\\u0_tms_reg[22] ;
  assign \new_[2127]_  = ~\\u0_tms_reg[23] ;
  assign \new_[2128]_  = ~\\u0_tms_reg[24] ;
  assign \new_[2129]_  = ~\\u0_tms_reg[26] ;
  assign \new_[2130]_  = ~\\u0_tms_reg[25] ;
  assign \new_[2131]_  = \\u0_tms_reg[2] ;
  assign \new_[2132]_  = ~\\u0_tms_reg[3] ;
  assign \new_[2133]_  = ~\\u0_tms_reg[4] ;
  assign \new_[2134]_  = ~\\u0_tms_reg[7] ;
  assign \new_[2135]_  = ~\\u0_tms_reg[8] ;
  assign \new_[2136]_  = ~\\u0_tms_reg[6] ;
  assign \new_[2137]_  = \\u5_timer_reg[7] ;
  assign \new_[2138]_  = \\u5_timer_reg[6] ;
  assign \new_[2139]_  = ~\\u0_sp_tms_reg[16] ;
  assign \new_[2140]_  = \new_[2228]_  | \new_[2319]_ ;
  assign \new_[2141]_  = \new_[11416]_  | \new_[11820]_ ;
  assign \new_[2142]_  = ~\new_[6072]_  & (~\new_[12551]_  | ~\new_[7003]_ );
  assign \new_[2143]_  = ~\new_[11736]_  | ~\new_[2219]_  | ~\new_[12549]_ ;
  assign \new_[2144]_  = ~\new_[12520]_  | ~\new_[7921]_  | ~\new_[7993]_  | ~\new_[11773]_ ;
  assign \new_[2145]_  = ~\new_[12520]_  | ~\new_[7547]_  | ~\new_[12233]_ ;
  assign \new_[2146]_  = ~\new_[2218]_ ;
  assign \new_[2147]_  = ~\new_[12519]_  | ~\new_[3036]_ ;
  assign \new_[2148]_  = ~\new_[2232]_  | (~\new_[2325]_  & ~\new_[12554]_ );
  assign \new_[2149]_  = ~\new_[2233]_  | (~\new_[2326]_  & ~\new_[12554]_ );
  assign \new_[2150]_  = ~\new_[2230]_  & (~\new_[7186]_  | ~\new_[5358]_ );
  assign \new_[2151]_  = ~\new_[2231]_  | (~\new_[2327]_  & ~\new_[12554]_ );
  assign \new_[2152]_  = \new_[2219]_ ;
  assign \new_[2153]_  = ~\new_[11829]_  & ~\new_[10964]_ ;
  assign \new_[2154]_  = ~\new_[11703]_  & ~\new_[10964]_ ;
  assign n1231 = ~\new_[3481]_  & (~\new_[2324]_  | ~\new_[3240]_ );
  assign \new_[2156]_  = ~\new_[2238]_  | (~\new_[5649]_  & ~\new_[2551]_ );
  assign \new_[2157]_  = ~\new_[2249]_  | ~\new_[6738]_ ;
  assign \new_[2158]_  = ~\new_[2251]_  | ~\new_[6738]_ ;
  assign \new_[2159]_  = ~\new_[2252]_  & (~\new_[2383]_  | ~\new_[4153]_ );
  assign \new_[2160]_  = ~\new_[6736]_  & ~\new_[2257]_ ;
  assign n1296 = ~\new_[2259]_  | ~\new_[2396]_ ;
  assign n1301 = ~\new_[2260]_  | ~\new_[2330]_ ;
  assign n1291 = ~\new_[2261]_  | ~\new_[2331]_ ;
  assign n1306 = ~\new_[2262]_  | ~\new_[2332]_ ;
  assign n1316 = ~\new_[2264]_  | ~\new_[2334]_ ;
  assign n1311 = ~\new_[2263]_  | ~\new_[2333]_ ;
  assign n1521 = ~\new_[2265]_  | ~\new_[2336]_ ;
  assign n1326 = ~\new_[2267]_  | ~\new_[2337]_ ;
  assign n1331 = ~\new_[2268]_  | ~\new_[2338]_ ;
  assign n1336 = ~\new_[2269]_  | ~\new_[2339]_ ;
  assign n1321 = ~\new_[2266]_  | ~\new_[2335]_ ;
  assign n1341 = ~\new_[2270]_  | ~\new_[2340]_ ;
  assign n1346 = ~\new_[2272]_  | ~\new_[2342]_ ;
  assign n1281 = ~\new_[2271]_  | ~\new_[2341]_ ;
  assign n1351 = ~\new_[2273]_  | ~\new_[2397]_ ;
  assign n1286 = ~\new_[2274]_  | ~\new_[2398]_ ;
  assign n1356 = ~\new_[2275]_  | ~\new_[2343]_ ;
  assign n1371 = ~\new_[2276]_  | ~\new_[2344]_ ;
  assign n1271 = ~\new_[11379]_  | ~\new_[2345]_ ;
  assign n1361 = ~\new_[2277]_  | ~\new_[2346]_ ;
  assign n1366 = ~\new_[2278]_  | ~\new_[2347]_ ;
  assign n1376 = ~\new_[2279]_  | ~\new_[2348]_ ;
  assign n1381 = ~\new_[2280]_  | ~\new_[2349]_ ;
  assign n1276 = ~\new_[2282]_  | ~\new_[2350]_ ;
  assign n1391 = ~\new_[2283]_  | ~\new_[2352]_ ;
  assign n1386 = ~\new_[2281]_  | ~\new_[2351]_ ;
  assign n1396 = ~\new_[2284]_  | ~\new_[2399]_ ;
  assign n1266 = ~\new_[2285]_  | ~\new_[2353]_ ;
  assign n1411 = ~\new_[2287]_  | ~\new_[2401]_ ;
  assign n1401 = ~\new_[2288]_  | ~\new_[2402]_ ;
  assign n1416 = ~\new_[2289]_  | ~\new_[2403]_ ;
  assign n1421 = ~\new_[2290]_  | ~\new_[2404]_ ;
  assign n1406 = ~\new_[2286]_  | ~\new_[2400]_ ;
  assign n1431 = ~\new_[2291]_  | ~\new_[2405]_ ;
  assign n1426 = ~\new_[2292]_  | ~\new_[2406]_ ;
  assign n1261 = ~\new_[2293]_  | ~\new_[2407]_ ;
  assign n1436 = ~\new_[2294]_  | ~\new_[2408]_ ;
  assign n1441 = ~\new_[2295]_  | ~\new_[2409]_ ;
  assign n1446 = ~\new_[2296]_  | ~\new_[2410]_ ;
  assign n1256 = ~\new_[2297]_  | ~\new_[2411]_ ;
  assign n1451 = ~\new_[2298]_  | ~\new_[2412]_ ;
  assign n1236 = ~\new_[2299]_  | ~\new_[2413]_ ;
  assign n1461 = ~\new_[2301]_  | ~\new_[2415]_ ;
  assign n1466 = ~\new_[2302]_  | ~\new_[2416]_ ;
  assign n1456 = ~\new_[2300]_  | ~\new_[2414]_ ;
  assign n1476 = ~\new_[2303]_  | ~\new_[2417]_ ;
  assign n1471 = ~\new_[2304]_  | ~\new_[2395]_ ;
  assign n1251 = ~\new_[2305]_  | ~\new_[2391]_ ;
  assign n1481 = ~\new_[2306]_  | ~\new_[2418]_ ;
  assign n1486 = ~\new_[2308]_  | ~\new_[2419]_ ;
  assign n1491 = ~\new_[2307]_  | ~\new_[2420]_ ;
  assign n1241 = ~\new_[2309]_  | ~\new_[2421]_ ;
  assign n1506 = ~\new_[2310]_  | ~\new_[2422]_ ;
  assign n1496 = ~\new_[2311]_  | ~\new_[2423]_ ;
  assign n1501 = ~\new_[2312]_  | ~\new_[2424]_ ;
  assign n1246 = ~\new_[2313]_  | ~\new_[2425]_ ;
  assign \new_[2217]_  = ~\new_[11736]_ ;
  assign \new_[2218]_  = ~\new_[2314]_  | ~\new_[10310]_ ;
  assign \new_[2219]_  = ~\new_[12519]_ ;
  assign \new_[2220]_  = ~\new_[10108]_  & (~\new_[4816]_  | ~\new_[2384]_ );
  assign \new_[2221]_  = ~\new_[2321]_  | ~\new_[12469]_ ;
  assign \new_[2222]_  = ~\new_[11823]_  & ~\new_[2323]_ ;
  assign \new_[2223]_  = ~\new_[7288]_  | ~\new_[2317]_  | ~\new_[11733]_ ;
  assign n1516 = ~\new_[3481]_  & (~\new_[2969]_  | ~\new_[2382]_ );
  assign n1511 = ~\new_[3481]_  & (~\new_[2883]_  | ~\new_[2382]_ );
  assign \new_[2226]_  = ~\new_[2329]_  | ~\new_[10108]_ ;
  assign \new_[2227]_  = ~\new_[12760]_  | ~\new_[7018]_ ;
  assign \new_[2228]_  = ~\new_[2328]_  & ~\new_[12384]_ ;
  assign \new_[2229]_  = ~\new_[7564]_  & ~\new_[12552]_ ;
  assign \new_[2230]_  = ~\new_[6122]_  & ~\new_[2371]_ ;
  assign \new_[2231]_  = ~\new_[2374]_  | ~\new_[9634]_ ;
  assign \new_[2232]_  = ~\new_[12424]_  | ~\new_[9634]_ ;
  assign \new_[2233]_  = ~\new_[2373]_  | ~\new_[9634]_ ;
  assign \new_[2234]_  = (~\new_[2435]_  | ~\new_[11833]_ ) & (~\new_[9580]_  | ~\new_[8070]_ );
  assign \new_[2235]_  = \new_[2376]_  | \new_[2426]_ ;
  assign \new_[2236]_  = \new_[2426]_  | \new_[2377]_ ;
  assign \new_[2237]_  = \new_[6812]_  | \new_[2375]_ ;
  assign \new_[2238]_  = ~\new_[2378]_  | ~\new_[11731]_ ;
  assign \new_[2239]_  = (~\new_[2436]_  | ~\new_[11833]_ ) & (~\new_[9260]_  | ~\new_[8490]_ );
  assign \new_[2240]_  = ~\new_[2483]_  & (~\new_[12760]_  | ~\new_[4153]_ );
  assign \new_[2241]_  = ~\new_[2379]_  & (~\new_[12762]_  | ~\new_[4153]_ );
  assign \new_[2242]_  = \new_[8392]_  ? \new_[12469]_  : \new_[2434]_ ;
  assign \new_[2243]_  = ~\new_[2383]_  & ~\new_[2431]_ ;
  assign \new_[2244]_  = ~\new_[6685]_  & ~\new_[12759]_ ;
  assign \new_[2245]_  = ~\new_[11416]_  & ~\new_[7300]_ ;
  assign \new_[2246]_  = ~\new_[6685]_  & ~\new_[12761]_ ;
  assign \new_[2247]_  = ~\new_[12217]_  & ~\new_[7300]_ ;
  assign \new_[2248]_  = \new_[11416]_  | \new_[6733]_ ;
  assign \new_[2249]_  = ~\new_[4547]_  | ~\new_[2384]_ ;
  assign \new_[2250]_  = \new_[12217]_  | \new_[6733]_ ;
  assign \new_[2251]_  = ~\new_[4560]_  | ~\new_[2384]_ ;
  assign \new_[2252]_  = ~\new_[11416]_  & ~\new_[11467]_ ;
  assign \new_[2253]_  = ~\new_[11569]_  & ~\new_[8707]_ ;
  assign \new_[2254]_  = \new_[3879]_  | \new_[2387]_ ;
  assign \new_[2255]_  = ~\new_[7186]_  | ~\new_[2389]_ ;
  assign \new_[2256]_  = ~\new_[11944]_  | ~\new_[2389]_ ;
  assign \new_[2257]_  = ~\new_[2329]_ ;
  assign \new_[2258]_  = \\u0_csc_reg[10] ;
  assign \new_[2259]_  = ~\new_[2496]_  & (~\new_[11381]_  | ~\new_[2451]_ );
  assign \new_[2260]_  = ~\new_[2497]_  & (~\new_[11381]_  | ~\new_[2452]_ );
  assign \new_[2261]_  = ~\new_[2498]_  & (~\new_[11381]_  | ~\new_[2453]_ );
  assign \new_[2262]_  = ~\new_[2499]_  & (~\new_[11381]_  | ~\new_[2454]_ );
  assign \new_[2263]_  = ~\new_[2500]_  & (~\new_[11381]_  | ~\new_[2455]_ );
  assign \new_[2264]_  = ~\new_[2501]_  & (~\new_[11381]_  | ~\new_[2456]_ );
  assign \new_[2265]_  = ~\new_[2503]_  & (~\new_[11381]_  | ~\new_[2458]_ );
  assign \new_[2266]_  = ~\new_[2502]_  & (~\new_[11381]_  | ~\new_[2457]_ );
  assign \new_[2267]_  = ~\new_[2504]_  & (~\new_[11381]_  | ~\new_[2459]_ );
  assign \new_[2268]_  = ~\new_[2505]_  & (~\new_[11381]_  | ~\new_[2460]_ );
  assign \new_[2269]_  = ~\new_[2506]_  & (~\new_[11381]_  | ~\new_[2461]_ );
  assign \new_[2270]_  = ~\new_[2507]_  & (~\new_[11381]_  | ~\new_[2462]_ );
  assign \new_[2271]_  = ~\new_[2508]_  & (~\new_[11381]_  | ~\new_[2463]_ );
  assign \new_[2272]_  = ~\new_[2509]_  & (~\new_[11381]_  | ~\new_[2464]_ );
  assign \new_[2273]_  = ~\new_[2510]_  & (~\new_[11381]_  | ~\new_[2465]_ );
  assign \new_[2274]_  = ~\new_[2511]_  & (~\new_[11381]_  | ~\new_[2466]_ );
  assign \new_[2275]_  = ~\new_[2512]_  & (~\new_[11381]_  | ~\new_[2467]_ );
  assign \new_[2276]_  = ~\new_[2513]_  & (~\new_[11381]_  | ~\new_[2468]_ );
  assign \new_[2277]_  = ~\new_[2514]_  & (~\new_[11381]_  | ~\new_[2469]_ );
  assign \new_[2278]_  = ~\new_[2515]_  & (~\new_[11381]_  | ~\new_[2470]_ );
  assign \new_[2279]_  = ~\new_[2516]_  & (~\new_[11381]_  | ~\new_[2471]_ );
  assign \new_[2280]_  = ~\new_[2517]_  & (~\new_[11381]_  | ~\new_[2472]_ );
  assign \new_[2281]_  = ~\new_[2519]_  & (~\new_[11381]_  | ~\new_[2474]_ );
  assign \new_[2282]_  = ~\new_[2518]_  & (~\new_[11381]_  | ~\new_[2473]_ );
  assign \new_[2283]_  = ~\new_[2520]_  & (~\new_[11381]_  | ~\new_[2475]_ );
  assign \new_[2284]_  = ~\new_[2521]_  & (~\new_[11381]_  | ~\new_[2476]_ );
  assign \new_[2285]_  = ~\new_[2522]_  & (~\new_[11381]_  | ~\new_[2477]_ );
  assign \new_[2286]_  = ~\new_[2523]_  & (~\new_[2451]_  | ~\new_[12601]_ );
  assign \new_[2287]_  = ~\new_[2524]_  & (~\new_[2452]_  | ~\new_[12601]_ );
  assign \new_[2288]_  = ~\new_[2525]_  & (~\new_[2453]_  | ~\new_[12601]_ );
  assign \new_[2289]_  = ~\new_[2526]_  & (~\new_[2454]_  | ~\new_[12601]_ );
  assign \new_[2290]_  = ~\new_[2527]_  & (~\new_[2455]_  | ~\new_[12601]_ );
  assign \new_[2291]_  = ~\new_[2528]_  & (~\new_[2456]_  | ~\new_[12601]_ );
  assign \new_[2292]_  = ~\new_[2529]_  & (~\new_[2457]_  | ~\new_[12601]_ );
  assign \new_[2293]_  = ~\new_[2530]_  & (~\new_[2458]_  | ~\new_[12601]_ );
  assign \new_[2294]_  = ~\new_[2531]_  & (~\new_[2459]_  | ~\new_[12601]_ );
  assign \new_[2295]_  = ~\new_[2532]_  & (~\new_[2460]_  | ~\new_[12601]_ );
  assign \new_[2296]_  = ~\new_[2533]_  & (~\new_[2461]_  | ~\new_[7727]_ );
  assign \new_[2297]_  = ~\new_[2534]_  & (~\new_[2462]_  | ~\new_[12601]_ );
  assign \new_[2298]_  = ~\new_[2535]_  & (~\new_[2463]_  | ~\new_[7727]_ );
  assign \new_[2299]_  = ~\new_[2536]_  & (~\new_[2464]_  | ~\new_[12601]_ );
  assign \new_[2300]_  = ~\new_[2537]_  & (~\new_[2465]_  | ~\new_[12601]_ );
  assign \new_[2301]_  = ~\new_[2538]_  & (~\new_[2466]_  | ~\new_[12601]_ );
  assign \new_[2302]_  = ~\new_[2539]_  & (~\new_[2467]_  | ~\new_[12601]_ );
  assign \new_[2303]_  = ~\new_[2540]_  & (~\new_[2468]_  | ~\new_[12601]_ );
  assign \new_[2304]_  = ~\new_[2541]_  & (~\new_[11380]_  | ~\new_[12601]_ );
  assign \new_[2305]_  = ~\new_[2542]_  & (~\new_[2469]_  | ~\new_[12601]_ );
  assign \new_[2306]_  = ~\new_[2543]_  & (~\new_[2470]_  | ~\new_[12601]_ );
  assign \new_[2307]_  = ~\new_[2545]_  & (~\new_[2472]_  | ~\new_[7727]_ );
  assign \new_[2308]_  = ~\new_[2544]_  & (~\new_[2471]_  | ~\new_[12601]_ );
  assign \new_[2309]_  = ~\new_[2546]_  & (~\new_[2473]_  | ~\new_[12601]_ );
  assign \new_[2310]_  = ~\new_[2547]_  & (~\new_[2474]_  | ~\new_[7727]_ );
  assign \new_[2311]_  = ~\new_[2548]_  & (~\new_[2475]_  | ~\new_[12601]_ );
  assign \new_[2312]_  = ~\new_[2549]_  & (~\new_[2476]_  | ~\new_[12601]_ );
  assign \new_[2313]_  = ~\new_[2550]_  & (~\new_[7727]_  | ~\new_[2477]_ );
  assign \new_[2314]_  = ~\new_[12552]_ ;
  assign \new_[2315]_  = \\u0_csc_reg[5] ;
  assign \new_[2316]_  = \\u0_csc_reg[4] ;
  assign \new_[2317]_  = ~\new_[2375]_ ;
  assign \new_[2318]_  = ~\new_[2429]_  & ~\new_[2430]_ ;
  assign \new_[2319]_  = \new_[11830]_  & \new_[7443]_ ;
  assign \new_[2320]_  = ~\new_[12674]_  | ~\new_[7018]_ ;
  assign \new_[2321]_  = ~\new_[2433]_  & ~\new_[10108]_ ;
  assign \new_[2322]_  = ~\new_[11830]_  | ~\new_[7018]_ ;
  assign \new_[2323]_  = ~\new_[11739]_ ;
  assign \new_[2324]_  = \new_[3879]_  | \new_[2433]_ ;
  assign \new_[2325]_  = ~\new_[2432]_  & (~\new_[6337]_  | ~\new_[10217]_ );
  assign \new_[2326]_  = ~\new_[2432]_  & (~\new_[12499]_  | ~\new_[10217]_ );
  assign \new_[2327]_  = ~\new_[2432]_  & (~\new_[6336]_  | ~\new_[10217]_ );
  assign \new_[2328]_  = ~\new_[2383]_ ;
  assign \new_[2329]_  = ~\new_[6076]_  | ~\new_[2437]_ ;
  assign \new_[2330]_  = ~\new_[11284]_  | ~\new_[11014]_ ;
  assign \new_[2331]_  = ~\new_[11284]_  | ~\new_[11122]_ ;
  assign \new_[2332]_  = ~\new_[11284]_  | ~\new_[11005]_ ;
  assign \new_[2333]_  = ~\new_[11284]_  | ~\new_[11136]_ ;
  assign \new_[2334]_  = ~\new_[11284]_  | ~\new_[11194]_ ;
  assign \new_[2335]_  = ~\new_[11284]_  | ~\new_[11137]_ ;
  assign \new_[2336]_  = ~\new_[11284]_  | ~\new_[11027]_ ;
  assign \new_[2337]_  = ~\new_[11284]_  | ~\new_[11002]_ ;
  assign \new_[2338]_  = ~\new_[11284]_  | ~\new_[11216]_ ;
  assign \new_[2339]_  = ~\new_[11284]_  | ~\new_[11035]_ ;
  assign \new_[2340]_  = ~\new_[11284]_  | ~\new_[2103]_ ;
  assign \new_[2341]_  = ~\new_[11284]_  | ~\new_[11076]_ ;
  assign \new_[2342]_  = ~\new_[11284]_  | ~\new_[11132]_ ;
  assign \new_[2343]_  = ~\new_[11284]_  | ~\new_[11128]_ ;
  assign \new_[2344]_  = ~\new_[11284]_  | ~\new_[11251]_ ;
  assign \new_[2345]_  = ~\new_[11284]_  | ~\new_[11044]_ ;
  assign \new_[2346]_  = ~\new_[11284]_  | ~\new_[11244]_ ;
  assign \new_[2347]_  = ~\new_[11284]_  | ~\new_[2108]_ ;
  assign \new_[2348]_  = ~\new_[11284]_  | ~\new_[11261]_ ;
  assign \new_[2349]_  = ~\new_[11284]_  | ~\new_[11006]_ ;
  assign \new_[2350]_  = ~\new_[11284]_  | ~\new_[11232]_ ;
  assign \new_[2351]_  = ~\new_[11284]_  | ~\new_[11143]_ ;
  assign \new_[2352]_  = ~\new_[11284]_  | ~\new_[11160]_ ;
  assign \new_[2353]_  = ~\new_[11284]_  | ~\new_[2085]_ ;
  assign \new_[2354]_  = ~u2_u0_bank0_open_reg;
  assign \new_[2355]_  = ~u2_u0_bank1_open_reg;
  assign \new_[2356]_  = ~u2_u0_bank3_open_reg;
  assign \new_[2357]_  = ~u2_u1_bank0_open_reg;
  assign \new_[2358]_  = ~u2_u1_bank1_open_reg;
  assign \new_[2359]_  = ~u2_u1_bank2_open_reg;
  assign \new_[2360]_  = ~\\u0_csc_reg[6] ;
  assign \new_[2361]_  = ~\\u0_csc_reg[7] ;
  assign \new_[2362]_  = ~\\u0_csc_reg[9] ;
  assign \new_[2363]_  = \\u0_sp_csc_reg[10] ;
  assign \new_[2364]_  = \\u0_sp_csc_reg[4] ;
  assign \new_[2365]_  = ~\\u0_sp_csc_reg[7] ;
  assign \new_[2366]_  = ~\\u0_sp_csc_reg[9] ;
  assign \new_[2367]_  = ~\\u0_sp_csc_reg[6] ;
  assign \new_[2368]_  = \\u0_sp_csc_reg[3] ;
  assign \new_[2369]_  = \\u0_sp_csc_reg[2] ;
  assign \new_[2370]_  = ~\\u0_csc_reg[11] ;
  assign \new_[2371]_  = ~\new_[8021]_  & (~\new_[2554]_  | ~\new_[9648]_ );
  assign \new_[2372]_  = ~u2_u1_bank3_open_reg;
  assign \new_[2373]_  = ~\new_[2481]_  | (~\new_[8817]_  & ~\new_[12469]_ );
  assign \new_[2374]_  = ~\new_[2482]_  | (~\new_[8484]_  & ~\new_[12469]_ );
  assign \new_[2375]_  = \new_[2551]_  | \new_[9902]_ ;
  assign \new_[2376]_  = ~\new_[2553]_  | ~\new_[2551]_ ;
  assign \new_[2377]_  = ~\new_[2576]_  | ~\new_[2551]_ ;
  assign \new_[2378]_  = ~\new_[7714]_  & ~\new_[2551]_ ;
  assign \new_[2379]_  = ~\new_[12675]_  & ~\new_[11474]_ ;
  assign \new_[2380]_  = ~\new_[9658]_  | ~\new_[2487]_  | ~\new_[12052]_ ;
  assign \new_[2381]_  = \\u0_sp_csc_reg[5] ;
  assign \new_[2382]_  = ~\new_[3878]_  | ~\new_[12218]_ ;
  assign \new_[2383]_  = \new_[7269]_  | \new_[12591]_ ;
  assign \new_[2384]_  = ~\new_[12218]_  | ~\new_[12469]_ ;
  assign \new_[2385]_  = ~\new_[2433]_ ;
  assign \new_[2386]_  = ~\new_[11706]_ ;
  assign \new_[2387]_  = ~\new_[2434]_ ;
  assign \new_[2388]_  = ~u2_u0_bank2_open_reg;
  assign \new_[2389]_  = ~\new_[2437]_ ;
  assign \new_[2390]_  = \\u0_sp_csc_reg[1] ;
  assign \new_[2391]_  = ~\new_[11282]_  | ~\new_[11101]_ ;
  assign n1536 = ~\new_[2568]_  | ~\new_[2573]_  | ~\new_[2579]_ ;
  assign n1531 = ~\new_[2569]_  | ~\new_[2588]_  | ~\new_[2580]_ ;
  assign n1526 = ~\new_[2567]_  | ~\new_[2574]_  | ~\new_[2578]_ ;
  assign \new_[2395]_  = ~\new_[11282]_  | ~\new_[11225]_ ;
  assign \new_[2396]_  = ~\new_[11284]_  | ~\new_[2094]_ ;
  assign \new_[2397]_  = ~\new_[11284]_  | ~\new_[11084]_ ;
  assign \new_[2398]_  = ~\new_[11284]_  | ~\new_[11090]_ ;
  assign \new_[2399]_  = ~\new_[11284]_  | ~\new_[11206]_ ;
  assign \new_[2400]_  = ~\new_[11280]_  | ~\new_[2116]_ ;
  assign \new_[2401]_  = ~\new_[11280]_  | ~\new_[11037]_ ;
  assign \new_[2402]_  = ~\new_[11284]_  | ~\new_[11064]_ ;
  assign \new_[2403]_  = ~\new_[11284]_  | ~\new_[11120]_ ;
  assign \new_[2404]_  = ~\new_[11284]_  | ~\new_[11106]_ ;
  assign \new_[2405]_  = ~\new_[11284]_  | ~\new_[11260]_ ;
  assign \new_[2406]_  = ~\new_[11284]_  | ~\new_[11001]_ ;
  assign \new_[2407]_  = ~\new_[11280]_  | ~\new_[10985]_ ;
  assign \new_[2408]_  = ~\new_[11282]_  | ~\new_[11024]_ ;
  assign \new_[2409]_  = ~\new_[11282]_  | ~\new_[11169]_ ;
  assign \new_[2410]_  = ~\new_[11280]_  | ~\new_[11103]_ ;
  assign \new_[2411]_  = ~\new_[11284]_  | ~\new_[2081]_ ;
  assign \new_[2412]_  = ~\new_[11280]_  | ~\new_[11047]_ ;
  assign \new_[2413]_  = ~\new_[11280]_  | ~\new_[11171]_ ;
  assign \new_[2414]_  = ~\new_[11282]_  | ~\new_[11215]_ ;
  assign \new_[2415]_  = ~\new_[11282]_  | ~\new_[11262]_ ;
  assign \new_[2416]_  = ~\new_[11280]_  | ~\new_[10993]_ ;
  assign \new_[2417]_  = ~\new_[11280]_  | ~\new_[11104]_ ;
  assign \new_[2418]_  = ~\new_[11284]_  | ~\new_[2131]_ ;
  assign \new_[2419]_  = ~\new_[11284]_  | ~\new_[11038]_ ;
  assign \new_[2420]_  = ~\new_[11282]_  | ~\new_[11142]_ ;
  assign \new_[2421]_  = ~\new_[11282]_  | ~\new_[11083]_ ;
  assign \new_[2422]_  = ~\new_[11284]_  | ~\new_[11170]_ ;
  assign \new_[2423]_  = ~\new_[11284]_  | ~\new_[11154]_ ;
  assign \new_[2424]_  = ~\new_[11284]_  | ~\new_[11155]_ ;
  assign \new_[2425]_  = ~\new_[11284]_  | ~\new_[2075]_ ;
  assign \new_[2426]_  = ~\new_[2552]_  | ~\new_[9658]_ ;
  assign \new_[2427]_  = ~\new_[2554]_  | ~\new_[7018]_ ;
  assign \new_[2428]_  = ~\new_[3879]_  & ~\new_[2551]_ ;
  assign \new_[2429]_  = ~\new_[2486]_ ;
  assign \new_[2430]_  = \new_[7124]_  | \new_[12218]_ ;
  assign \new_[2431]_  = \new_[7123]_  | \new_[12218]_ ;
  assign \new_[2432]_  = \new_[12218]_  & \new_[10326]_ ;
  assign \new_[2433]_  = ~\new_[7376]_  & ~\new_[12218]_ ;
  assign \new_[2434]_  = \new_[7375]_  | \new_[12218]_ ;
  assign \new_[2435]_  = \new_[7121]_  | \new_[12218]_ ;
  assign \new_[2436]_  = \new_[7120]_  | \new_[12218]_ ;
  assign \new_[2437]_  = ~\new_[12218]_ ;
  assign \new_[2438]_  = ~\new_[2601]_  | ~\new_[4135]_  | ~\new_[2772]_  | ~\new_[4167]_ ;
  assign n1571 = ~\new_[2561]_  | (~\new_[2617]_  & ~\new_[2360]_ );
  assign n1581 = ~\new_[2562]_  | (~\new_[2617]_  & ~\new_[2362]_ );
  assign n1576 = ~\new_[2563]_  | (~\new_[2631]_  & ~\new_[2361]_ );
  assign n1586 = ~\new_[2595]_  | ~\new_[2589]_  | ~\new_[2581]_ ;
  assign n1591 = ~\new_[2599]_  | ~\new_[2593]_  | ~\new_[2582]_ ;
  assign n1631 = ~\new_[2600]_  | ~\new_[2594]_  | ~\new_[2583]_ ;
  assign n1606 = ~\new_[2564]_  | (~\new_[2631]_  & ~\new_[2367]_ );
  assign n1596 = ~\new_[2565]_  | (~\new_[2631]_  & ~\new_[2365]_ );
  assign n1601 = ~\new_[2566]_  | (~\new_[2631]_  & ~\new_[2366]_ );
  assign n1616 = ~\new_[2586]_  | ~\new_[2591]_  | ~\new_[2597]_ ;
  assign n1641 = ~\new_[2585]_  | ~\new_[2590]_  | ~\new_[2596]_ ;
  assign n1611 = ~\new_[2587]_  | ~\new_[2592]_  | ~\new_[2598]_ ;
  assign \new_[2451]_  = ~\new_[11289]_  & ~\new_[11217]_ ;
  assign \new_[2452]_  = ~\new_[11286]_  & ~\new_[10982]_ ;
  assign \new_[2453]_  = ~\new_[11286]_  & ~\new_[7968]_ ;
  assign \new_[2454]_  = ~\new_[11286]_  & ~\new_[7943]_ ;
  assign \new_[2455]_  = ~\new_[11288]_  & ~\new_[7917]_ ;
  assign \new_[2456]_  = ~\new_[11286]_  & ~\new_[7969]_ ;
  assign \new_[2457]_  = ~\new_[11288]_  & ~\new_[7922]_ ;
  assign \new_[2458]_  = ~\new_[11289]_  & ~\new_[7936]_ ;
  assign \new_[2459]_  = ~\new_[11288]_  & ~\new_[7941]_ ;
  assign \new_[2460]_  = ~\new_[11286]_  & ~\new_[7950]_ ;
  assign \new_[2461]_  = ~\new_[11288]_  & ~\new_[7981]_ ;
  assign \new_[2462]_  = ~\new_[11286]_  & ~\new_[11152]_ ;
  assign \new_[2463]_  = ~\new_[11286]_  & ~\new_[7970]_ ;
  assign \new_[2464]_  = ~\new_[11288]_  & ~\new_[7985]_ ;
  assign \new_[2465]_  = ~\new_[11286]_  & ~\new_[7984]_ ;
  assign \new_[2466]_  = ~\new_[11286]_  & ~\new_[7939]_ ;
  assign \new_[2467]_  = ~\new_[11289]_  & ~\new_[11023]_ ;
  assign \new_[2468]_  = ~\new_[11286]_  & ~\new_[11118]_ ;
  assign \new_[2469]_  = ~\new_[11288]_  & ~\new_[11096]_ ;
  assign \new_[2470]_  = ~\new_[11286]_  & ~\new_[10981]_ ;
  assign \new_[2471]_  = ~\new_[11286]_  & ~\new_[11032]_ ;
  assign \new_[2472]_  = ~\new_[11288]_  & ~\new_[10999]_ ;
  assign \new_[2473]_  = ~\new_[11286]_  & ~\new_[11149]_ ;
  assign \new_[2474]_  = ~\new_[11288]_  & ~\new_[11172]_ ;
  assign \new_[2475]_  = ~\new_[11286]_  & ~\new_[11157]_ ;
  assign \new_[2476]_  = ~\new_[11289]_  & ~\new_[11163]_ ;
  assign \new_[2477]_  = ~\new_[11286]_  & ~\new_[11077]_ ;
  assign \new_[2478]_  = \\u0_csc_reg[1] ;
  assign \new_[2479]_  = \\u0_csc_reg[3] ;
  assign n1621 = ~\new_[2604]_  | (~\new_[2617]_  & ~\new_[2370]_ );
  assign \new_[2481]_  = ~\new_[12469]_  | ~\new_[2576]_ ;
  assign \new_[2482]_  = ~\new_[12469]_  | ~\new_[2575]_ ;
  assign \new_[2483]_  = ~\new_[11825]_  & ~\new_[11474]_ ;
  assign \new_[2484]_  = ~\new_[11740]_  | ~\new_[11944]_ ;
  assign \new_[2485]_  = ~\new_[7186]_  | ~\new_[11740]_  | ~\new_[6540]_ ;
  assign \new_[2486]_  = ~\new_[7603]_  & ~\new_[12591]_ ;
  assign \new_[2487]_  = ~\new_[2552]_ ;
  assign n1546 = ~\new_[2555]_  | ~\new_[7431]_ ;
  assign n1636 = ~\new_[2556]_  | ~\new_[7439]_ ;
  assign n1566 = ~\new_[2559]_  | ~\new_[7429]_ ;
  assign n1561 = ~\new_[2558]_  | ~\new_[7427]_ ;
  assign n1551 = ~\new_[2557]_  | ~\new_[7433]_ ;
  assign n1626 = ~\new_[2560]_  | ~\new_[7430]_ ;
  assign \new_[2494]_  = \\u0_csc_reg[2] ;
  assign \new_[2495]_  = \new_[2720]_  ? \new_[4262]_  : n1661;
  assign \new_[2496]_  = ~\new_[10705]_  & ~\new_[11281]_ ;
  assign \new_[2497]_  = ~\new_[10437]_  & ~\new_[11279]_ ;
  assign \new_[2498]_  = ~\new_[10721]_  & ~\new_[11279]_ ;
  assign \new_[2499]_  = ~\new_[10737]_  & ~\new_[11279]_ ;
  assign \new_[2500]_  = ~\new_[10423]_  & ~\new_[11279]_ ;
  assign \new_[2501]_  = ~\new_[10616]_  & ~\new_[11279]_ ;
  assign \new_[2502]_  = ~\new_[10667]_  & ~\new_[11279]_ ;
  assign \new_[2503]_  = ~\new_[10464]_  & ~\new_[11385]_ ;
  assign \new_[2504]_  = ~\new_[10782]_  & ~\new_[11279]_ ;
  assign \new_[2505]_  = ~\new_[10567]_  & ~\new_[11279]_ ;
  assign \new_[2506]_  = ~\new_[10492]_  & ~\new_[11385]_ ;
  assign \new_[2507]_  = ~\new_[10399]_  & ~\new_[11385]_ ;
  assign \new_[2508]_  = ~\new_[10462]_  & ~\new_[11281]_ ;
  assign \new_[2509]_  = ~\new_[10663]_  & ~\new_[11279]_ ;
  assign \new_[2510]_  = ~\new_[10751]_  & ~\new_[11279]_ ;
  assign \new_[2511]_  = ~\new_[10605]_  & ~\new_[11279]_ ;
  assign \new_[2512]_  = ~\new_[10465]_  & ~\new_[11385]_ ;
  assign \new_[2513]_  = ~\new_[10395]_  & ~\new_[11281]_ ;
  assign \new_[2514]_  = ~\new_[10489]_  & ~\new_[11385]_ ;
  assign \new_[2515]_  = ~\new_[10672]_  & ~\new_[11281]_ ;
  assign \new_[2516]_  = ~\new_[10622]_  & ~\new_[11279]_ ;
  assign \new_[2517]_  = ~\new_[10577]_  & ~\new_[11279]_ ;
  assign \new_[2518]_  = ~\new_[10719]_  & ~\new_[11279]_ ;
  assign \new_[2519]_  = ~\new_[10540]_  & ~\new_[11279]_ ;
  assign \new_[2520]_  = ~\new_[10410]_  & ~\new_[11385]_ ;
  assign \new_[2521]_  = ~\new_[10453]_  & ~\new_[11385]_ ;
  assign \new_[2522]_  = ~\new_[10674]_  & ~\new_[11279]_ ;
  assign \new_[2523]_  = ~\new_[7393]_  & ~\new_[11279]_ ;
  assign \new_[2524]_  = ~\new_[7394]_  & ~\new_[11279]_ ;
  assign \new_[2525]_  = ~\new_[7395]_  & ~\new_[11385]_ ;
  assign \new_[2526]_  = ~\new_[7396]_  & ~\new_[11385]_ ;
  assign \new_[2527]_  = ~\new_[7397]_  & ~\new_[11385]_ ;
  assign \new_[2528]_  = ~\new_[7392]_  & ~\new_[11279]_ ;
  assign \new_[2529]_  = ~\new_[7398]_  & ~\new_[11279]_ ;
  assign \new_[2530]_  = ~\new_[7399]_  & ~\new_[11385]_ ;
  assign \new_[2531]_  = ~\new_[7400]_  & ~\new_[11385]_ ;
  assign \new_[2532]_  = ~\new_[7401]_  & ~\new_[11385]_ ;
  assign \new_[2533]_  = ~\new_[7388]_  & ~\new_[11385]_ ;
  assign \new_[2534]_  = ~\new_[7402]_  & ~\new_[11279]_ ;
  assign \new_[2535]_  = ~\new_[7403]_  & ~\new_[11279]_ ;
  assign \new_[2536]_  = ~\new_[7405]_  & ~\new_[11385]_ ;
  assign \new_[2537]_  = ~\new_[7404]_  & ~\new_[11279]_ ;
  assign \new_[2538]_  = ~\new_[7406]_  & ~\new_[11279]_ ;
  assign \new_[2539]_  = ~\new_[7387]_  & ~\new_[11385]_ ;
  assign \new_[2540]_  = ~\new_[7407]_  & ~\new_[11385]_ ;
  assign \new_[2541]_  = ~\new_[7408]_  & ~\new_[11279]_ ;
  assign \new_[2542]_  = ~\new_[7409]_  & ~\new_[11385]_ ;
  assign \new_[2543]_  = ~\new_[7410]_  & ~\new_[11385]_ ;
  assign \new_[2544]_  = ~\new_[7411]_  & ~\new_[11385]_ ;
  assign \new_[2545]_  = ~\new_[7412]_  & ~\new_[11385]_ ;
  assign \new_[2546]_  = ~\new_[7413]_  & ~\new_[11279]_ ;
  assign \new_[2547]_  = ~\new_[7384]_  & ~\new_[11279]_ ;
  assign \new_[2548]_  = ~\new_[7414]_  & ~\new_[11385]_ ;
  assign \new_[2549]_  = ~\new_[7383]_  & ~\new_[11279]_ ;
  assign \new_[2550]_  = ~\new_[7415]_  & ~\new_[11385]_ ;
  assign \new_[2551]_  = ~\new_[2575]_ ;
  assign \new_[2552]_  = ~\new_[12466]_ ;
  assign \new_[2553]_  = ~\new_[2576]_ ;
  assign \new_[2554]_  = ~\new_[11825]_ ;
  assign \new_[2555]_  = ~\new_[11199]_  | ~\new_[6350]_  | ~\new_[12202]_ ;
  assign \new_[2556]_  = ~\new_[11109]_  | ~\new_[6351]_  | ~\new_[12202]_ ;
  assign \new_[2557]_  = ~\new_[11176]_  | ~\new_[6352]_  | ~\new_[12202]_ ;
  assign \new_[2558]_  = ~\new_[11111]_  | ~\new_[6353]_  | ~\new_[12209]_ ;
  assign \new_[2559]_  = ~\new_[11067]_  | ~\new_[6354]_  | ~\new_[12209]_ ;
  assign \new_[2560]_  = ~\new_[11178]_  | ~\new_[6355]_  | ~\new_[12209]_ ;
  assign \new_[2561]_  = (~\new_[2611]_  | ~\new_[7765]_ ) & (~\new_[2610]_  | ~\new_[7727]_ );
  assign \new_[2562]_  = (~\new_[2614]_  | ~\new_[7765]_ ) & (~\new_[2616]_  | ~\new_[7727]_ );
  assign \new_[2563]_  = (~\new_[2613]_  | ~\new_[7765]_ ) & (~\new_[2612]_  | ~\new_[7727]_ );
  assign \new_[2564]_  = (~\new_[10479]_  | ~\new_[2617]_ ) & (~\new_[2610]_  | ~\new_[11381]_ );
  assign \new_[2565]_  = (~\new_[10472]_  | ~\new_[2617]_ ) & (~\new_[2612]_  | ~\new_[11381]_ );
  assign \new_[2566]_  = (~\new_[10467]_  | ~\new_[2617]_ ) & (~\new_[2616]_  | ~\new_[11381]_ );
  assign \new_[2567]_  = ~\new_[7715]_  | ~\new_[7765]_  | ~\new_[2617]_ ;
  assign \new_[2568]_  = ~\new_[7594]_  | ~\new_[7765]_  | ~\new_[2617]_ ;
  assign \new_[2569]_  = ~\new_[7619]_  | ~\new_[7765]_  | ~\new_[2617]_ ;
  assign n1646 = \new_[2478]_  ? \new_[2617]_  : \new_[7127]_ ;
  assign n1656 = \new_[2494]_  ? \new_[2617]_  : \new_[7128]_ ;
  assign n1651 = \new_[2479]_  ? \new_[2617]_  : \new_[7129]_ ;
  assign \new_[2573]_  = ~\new_[2623]_  | ~\new_[2316]_ ;
  assign \new_[2574]_  = ~\new_[2623]_  | ~\new_[2258]_ ;
  assign \new_[2575]_  = ~\new_[11373]_ ;
  assign \new_[2576]_  = ~\new_[11372]_ ;
  assign \new_[2577]_  = u5_cmd_a10_r_reg;
  assign \new_[2578]_  = ~\new_[2607]_  | ~\new_[7727]_ ;
  assign \new_[2579]_  = ~\new_[2608]_  | ~\new_[7727]_ ;
  assign \new_[2580]_  = ~\new_[2609]_  | ~\new_[12601]_ ;
  assign \new_[2581]_  = ~\new_[2607]_  | ~\new_[11381]_ ;
  assign \new_[2582]_  = ~\new_[2608]_  | ~\new_[11381]_ ;
  assign \new_[2583]_  = ~\new_[2609]_  | ~\new_[11381]_ ;
  assign mc_ras_pad_o_ = u7_mc_ras__reg;
  assign \new_[2585]_  = ~\new_[11153]_  | ~\new_[2615]_  | ~\new_[7813]_ ;
  assign \new_[2586]_  = ~\new_[11153]_  | ~\new_[2615]_  | ~\new_[7828]_ ;
  assign \new_[2587]_  = ~\new_[11153]_  | ~\new_[2615]_  | ~\new_[7851]_ ;
  assign \new_[2588]_  = ~\new_[2623]_  | ~\new_[10956]_ ;
  assign \new_[2589]_  = ~\new_[2623]_  | ~\new_[2363]_ ;
  assign \new_[2590]_  = ~\new_[2623]_  | ~\new_[2390]_ ;
  assign \new_[2591]_  = ~\new_[2623]_  | ~\new_[2369]_ ;
  assign \new_[2592]_  = ~\new_[2623]_  | ~\new_[2368]_ ;
  assign \new_[2593]_  = ~\new_[2623]_  | ~\new_[2364]_ ;
  assign \new_[2594]_  = ~\new_[2623]_  | ~\new_[2381]_ ;
  assign \new_[2595]_  = ~\new_[10949]_  | ~\new_[2617]_  | ~\new_[7715]_ ;
  assign \new_[2596]_  = ~\new_[7618]_  | ~\new_[2617]_  | ~\new_[10949]_ ;
  assign \new_[2597]_  = ~\new_[7616]_  | ~\new_[2617]_  | ~\new_[10949]_ ;
  assign \new_[2598]_  = ~\new_[7732]_  | ~\new_[2617]_  | ~\new_[10949]_ ;
  assign \new_[2599]_  = ~\new_[10949]_  | ~\new_[2617]_  | ~\new_[7594]_ ;
  assign \new_[2600]_  = ~\new_[10949]_  | ~\new_[2617]_  | ~\new_[7619]_ ;
  assign \new_[2601]_  = ~\new_[2621]_  & (~\new_[7682]_  | ~\new_[9746]_ );
  assign mc_adsc_pad_o_ = u7_mc_adsc__reg;
  assign n1661 = \new_[2622]_  | \new_[3501]_ ;
  assign \new_[2604]_  = \new_[7270]_  | \new_[2623]_ ;
  assign \new_[2605]_  = (~\new_[2641]_  & ~\new_[9913]_  & ~\new_[10419]_ ) | (~\new_[9813]_  & ~\new_[5643]_  & ~\new_[11316]_ );
  assign \new_[2606]_  = u5_wr_cycle_reg;
  assign \new_[2607]_  = \new_[2631]_  & \new_[7716]_ ;
  assign \new_[2608]_  = \new_[2631]_  & \new_[7733]_ ;
  assign \new_[2609]_  = \new_[2631]_  & \new_[7722]_ ;
  assign \new_[2610]_  = \new_[2631]_  & \new_[7951]_ ;
  assign \new_[2611]_  = \new_[2631]_  & \new_[7625]_ ;
  assign \new_[2612]_  = \new_[2631]_  & \new_[7723]_ ;
  assign \new_[2613]_  = \new_[2631]_  & \new_[7595]_ ;
  assign \new_[2614]_  = \new_[2631]_  & \new_[7624]_ ;
  assign \new_[2615]_  = \new_[2631]_  & \new_[9136]_ ;
  assign \new_[2616]_  = \new_[2631]_  & \new_[7724]_ ;
  assign \new_[2617]_  = ~\new_[2623]_ ;
  assign \new_[2618]_  = ~\new_[2625]_ ;
  assign n1666 = \new_[2647]_  ? \new_[10283]_  : n1716;
  assign \new_[2620]_  = ~\new_[4107]_  | ~\new_[2965]_  | ~\new_[5314]_  | ~\new_[2665]_ ;
  assign \new_[2621]_  = ~\new_[2640]_  | (~\new_[8725]_  & ~\new_[11503]_ );
  assign \new_[2622]_  = ~\new_[4759]_  | ~\new_[5282]_  | ~\new_[3284]_  | ~\new_[2670]_ ;
  assign \new_[2623]_  = ~\new_[2631]_ ;
  assign n1671 = ~\new_[5378]_  | ~\new_[5418]_  | ~\new_[2644]_  | ~\new_[3729]_ ;
  assign \new_[2625]_  = ~\new_[2739]_  | ~\new_[6549]_  | ~\new_[2648]_  | ~\new_[4101]_ ;
  assign \new_[2626]_  = ~\new_[8013]_  | ~\new_[5075]_  | ~\new_[2729]_  | ~\new_[2668]_ ;
  assign \new_[2627]_  = ~\new_[2669]_  & ~\new_[11404]_ ;
  assign \new_[2628]_  = ~\new_[2669]_  & ~\new_[11403]_ ;
  assign \new_[2629]_  = ~\new_[2774]_  | ~\new_[5371]_  | ~\new_[4281]_  | ~\new_[6721]_ ;
  assign mc_coe_pad_coe_o = u7_mc_c_oe_reg;
  assign \new_[2631]_  = \new_[2642]_ ;
  assign \new_[2632]_  = ~\new_[2642]_ ;
  assign \new_[2633]_  = ~\new_[2806]_  | ~\new_[5993]_  | ~\new_[2705]_  | ~\new_[4117]_ ;
  assign \new_[2634]_  = n1681 & \new_[11113]_ ;
  assign \new_[2635]_  = ~\new_[2667]_  & ~\new_[2880]_ ;
  assign \new_[2636]_  = ~\new_[2740]_  | ~\new_[5609]_  | ~\new_[2920]_  | ~\new_[4602]_ ;
  assign n1676 = ~\new_[3633]_  | ~\new_[2743]_  | ~\new_[8712]_  | ~\new_[3632]_ ;
  assign n5766 = u5_cs_le_reg;
  assign \new_[2639]_  = ~\new_[2958]_  | ~\new_[5743]_  | ~\new_[2718]_  | ~\new_[4136]_ ;
  assign \new_[2640]_  = (~\new_[2773]_  | ~\new_[10001]_ ) & (~\new_[7260]_  | ~\new_[11453]_ );
  assign \new_[2641]_  = \new_[5019]_  & \new_[2722]_ ;
  assign \new_[2642]_  = n1686 & \new_[10948]_ ;
  assign \new_[2643]_  = ~\new_[2777]_  | ~\new_[4272]_  | ~\new_[5367]_ ;
  assign \new_[2644]_  = ~\new_[2723]_  & ~\new_[3867]_ ;
  assign \new_[2645]_  = ~\new_[2871]_  | ~\new_[4925]_  | ~\new_[2708]_  | ~\new_[4120]_ ;
  assign \new_[2646]_  = ~\new_[2873]_  | ~\new_[6620]_  | ~\new_[2714]_  | ~\new_[3865]_ ;
  assign \new_[2647]_  = \\u5_cmd_del_reg[2] ;
  assign \new_[2648]_  = ~\new_[2725]_  & (~\new_[7682]_  | ~\new_[10102]_ );
  assign \new_[2649]_  = (~\new_[3687]_  | ~\new_[2805]_ ) & (~\new_[4296]_  | ~\new_[6036]_ );
  assign \new_[2650]_  = ~\new_[2795]_  & ~\new_[2702]_ ;
  assign \new_[2651]_  = ~\new_[2796]_  & ~\new_[2704]_ ;
  assign \new_[2652]_  = ~\new_[3007]_  | ~\new_[5728]_  | ~\new_[2706]_  | ~\new_[4118]_ ;
  assign \new_[2653]_  = ~\new_[2888]_  | ~\new_[5729]_  | ~\new_[2707]_  | ~\new_[4119]_ ;
  assign \new_[2654]_  = ~\new_[3010]_  | ~\new_[5730]_  | ~\new_[2709]_  | ~\new_[4121]_ ;
  assign \new_[2655]_  = ~\new_[2893]_  | ~\new_[5731]_  | ~\new_[2710]_  | ~\new_[4122]_ ;
  assign \new_[2656]_  = ~\new_[2894]_  | ~\new_[5732]_  | ~\new_[2688]_  | ~\new_[4125]_ ;
  assign \new_[2657]_  = ~\new_[2896]_  | ~\new_[5736]_  | ~\new_[2715]_  | ~\new_[4130]_ ;
  assign \new_[2658]_  = ~\new_[2897]_  | ~\new_[5738]_  | ~\new_[2716]_  | ~\new_[4133]_ ;
  assign \new_[2659]_  = ~\new_[2890]_  | ~\new_[4067]_  | ~\new_[2717]_  | ~\new_[6680]_ ;
  assign \new_[2660]_  = ~\new_[2864]_  & ~\new_[2689]_ ;
  assign \new_[2661]_  = ~\new_[4216]_  | ~\new_[5024]_  | ~\new_[2730]_  | ~\new_[2961]_ ;
  assign \new_[2662]_  = ~\new_[4051]_  | ~\new_[5119]_  | ~\new_[2731]_  | ~\new_[2770]_ ;
  assign \new_[2663]_  = ~\new_[4217]_  | ~\new_[5124]_  | ~\new_[2732]_  | ~\new_[2771]_ ;
  assign \new_[2664]_  = ~\new_[2686]_  & ~\new_[2807]_ ;
  assign \new_[2665]_  = \new_[2692]_  & \new_[7323]_ ;
  assign \new_[2666]_  = ~\new_[2950]_  | ~\new_[4211]_  | ~\new_[6547]_  | ~\new_[5820]_ ;
  assign \new_[2667]_  = ~\new_[4556]_  | ~\new_[5965]_  | ~\new_[4050]_  | ~\new_[2856]_ ;
  assign \new_[2668]_  = ~\new_[2741]_  & (~\new_[12534]_  | ~\new_[9856]_ );
  assign \new_[2669]_  = (~\new_[2857]_  | ~\new_[9299]_ ) & (~\new_[4242]_  | ~\new_[9926]_ );
  assign \new_[2670]_  = ~\new_[12430]_  & (~\new_[6459]_  | ~\new_[10278]_ );
  assign \new_[2671]_  = ~\new_[4960]_  | ~\new_[4279]_  | ~\new_[2870]_ ;
  assign \new_[2672]_  = ~\new_[7669]_  | ~\new_[4048]_  | ~\new_[2869]_ ;
  assign \new_[2673]_  = ~\new_[5844]_  | ~\new_[6463]_  | ~\new_[4103]_  | ~\new_[2872]_ ;
  assign \new_[2674]_  = ~\new_[2778]_  & (~\new_[12534]_  | ~\new_[11787]_ );
  assign \new_[2675]_  = ~\new_[2779]_  & (~\new_[12534]_  | ~\new_[9985]_ );
  assign \new_[2676]_  = ~\new_[2780]_  & (~\new_[12534]_  | ~\new_[10244]_ );
  assign \new_[2677]_  = ~\new_[2781]_  & (~\new_[12534]_  | ~\new_[11452]_ );
  assign \new_[2678]_  = ~\new_[2782]_  & (~\new_[12534]_  | ~\new_[9606]_ );
  assign \new_[2679]_  = ~\new_[2783]_  & (~\new_[12534]_  | ~\new_[9970]_ );
  assign n1681 = u5_mc_c_oe_reg;
  assign \new_[2681]_  = ~\new_[7170]_  | ~\new_[2802]_  | ~\new_[4670]_ ;
  assign \new_[2682]_  = ~\new_[2790]_  & ~\new_[2745]_ ;
  assign \new_[2683]_  = ~\new_[3014]_  | ~\new_[5735]_  | ~\new_[2766]_  | ~\new_[4129]_ ;
  assign \new_[2684]_  = ~\new_[2899]_  & ~\new_[2799]_ ;
  assign \new_[2685]_  = ~\new_[4132]_  | ~\new_[2964]_  | ~\new_[5968]_  | ~\new_[6147]_ ;
  assign \new_[2686]_  = ~\new_[4555]_  | ~\new_[5962]_  | ~\new_[4049]_  | ~\new_[2948]_ ;
  assign \new_[2687]_  = ~\new_[4565]_  | ~\new_[5521]_  | ~\new_[2828]_  | ~\new_[5522]_ ;
  assign \new_[2688]_  = ~\new_[2737]_ ;
  assign \new_[2689]_  = ~\new_[4572]_  | ~\new_[5581]_  | ~\new_[6292]_  | ~\new_[2938]_ ;
  assign \new_[2690]_  = ~\new_[2825]_  & (~\new_[12534]_  | ~\new_[11504]_ );
  assign \new_[2691]_  = ~\new_[2826]_  & (~\new_[12534]_  | ~\new_[10045]_ );
  assign \new_[2692]_  = ~\new_[2824]_  & (~\new_[7588]_  | ~\new_[10818]_ );
  assign \new_[2693]_  = ~\new_[2827]_  & (~\new_[7599]_  | ~\new_[11356]_ );
  assign \new_[2694]_  = ~\new_[4845]_  | ~\new_[5511]_  | ~\new_[2834]_  | ~\new_[5512]_ ;
  assign \new_[2695]_  = ~\new_[4846]_  | ~\new_[5030]_  | ~\new_[2835]_  | ~\new_[5515]_ ;
  assign \new_[2696]_  = ~\new_[4564]_  | ~\new_[5518]_  | ~\new_[2836]_  | ~\new_[5519]_ ;
  assign \new_[2697]_  = ~\new_[4847]_  | ~\new_[5524]_  | ~\new_[2838]_  | ~\new_[5525]_ ;
  assign \new_[2698]_  = ~\new_[4852]_  | ~\new_[5537]_  | ~\new_[2844]_  | ~\new_[5538]_ ;
  assign \new_[2699]_  = ~\new_[4853]_  | ~\new_[5540]_  | ~\new_[2846]_  | ~\new_[5927]_ ;
  assign \new_[2700]_  = ~\new_[4854]_  | ~\new_[5543]_  | ~\new_[2847]_  | ~\new_[5544]_ ;
  assign \new_[2701]_  = ~\new_[4855]_  | ~\new_[5546]_  | ~\new_[2848]_  | ~\new_[5547]_ ;
  assign \new_[2702]_  = ~\new_[4567]_  | ~\new_[5059]_  | ~\new_[2850]_  | ~\new_[5060]_ ;
  assign \new_[2703]_  = ~\new_[4858]_  | ~\new_[5558]_  | ~\new_[2851]_  | ~\new_[5559]_ ;
  assign \new_[2704]_  = ~\new_[4568]_  | ~\new_[5069]_  | ~\new_[2852]_  | ~\new_[5071]_ ;
  assign \new_[2705]_  = ~\new_[2752]_ ;
  assign \new_[2706]_  = ~\new_[2753]_ ;
  assign \new_[2707]_  = ~\new_[2754]_ ;
  assign \new_[2708]_  = ~\new_[2755]_ ;
  assign \new_[2709]_  = ~\new_[2756]_ ;
  assign \new_[2710]_  = ~\new_[2757]_ ;
  assign \new_[2711]_  = ~\new_[4570]_  | ~\new_[5575]_  | ~\new_[2853]_  | ~\new_[5576]_ ;
  assign \new_[2712]_  = ~\new_[4868]_  | ~\new_[5573]_  | ~\new_[2854]_  | ~\new_[5578]_ ;
  assign \new_[2713]_  = ~\new_[2759]_ ;
  assign \new_[2714]_  = ~\new_[2760]_ ;
  assign \new_[2715]_  = ~\new_[2761]_ ;
  assign \new_[2716]_  = ~\new_[2762]_ ;
  assign \new_[2717]_  = ~\new_[2764]_ ;
  assign \new_[2718]_  = ~\new_[2765]_ ;
  assign \new_[2719]_  = ~\\u1_bank_adr_reg[0] ;
  assign \new_[2720]_  = \\u1_row_adr_reg[10] ;
  assign \new_[2721]_  = \\u1_row_adr_reg[11] ;
  assign \new_[2722]_  = \new_[2858]_  | \new_[11298]_ ;
  assign \new_[2723]_  = ~\new_[3340]_  | ~\new_[3103]_  | ~\new_[2859]_  | ~\new_[3079]_ ;
  assign n1691 = \\u5_cmd_r_reg[2] ;
  assign \new_[2725]_  = ~\new_[2868]_  | (~\new_[8709]_  & ~\new_[11503]_ );
  assign \new_[2726]_  = ~\new_[3799]_  | ~\new_[11846]_  | ~\new_[5763]_  | ~\new_[2968]_ ;
  assign \new_[2727]_  = ~\new_[4822]_  | ~\new_[5972]_  | ~\new_[2865]_  | ~\new_[3216]_ ;
  assign \new_[2728]_  = ~\new_[3525]_  | ~\new_[5949]_  | ~\new_[5890]_  | ~\new_[2898]_ ;
  assign \new_[2729]_  = ~\new_[4280]_  & ~\new_[2874]_ ;
  assign \new_[2730]_  = ~\new_[4282]_  & ~\new_[2875]_ ;
  assign \new_[2731]_  = ~\new_[4284]_  & ~\new_[2876]_ ;
  assign \new_[2732]_  = ~\new_[4285]_  & ~\new_[2877]_ ;
  assign \new_[2733]_  = ~\new_[5720]_  | ~\new_[4276]_  | ~\new_[2891]_ ;
  assign \new_[2734]_  = ~\new_[5722]_  | ~\new_[4277]_  | ~\new_[2892]_ ;
  assign \new_[2735]_  = ~\new_[3299]_  | ~\new_[5953]_  | ~\new_[2917]_  | ~\new_[4599]_ ;
  assign \new_[2736]_  = ~\new_[3148]_  | ~\new_[5586]_  | ~\new_[3131]_  | ~\new_[4258]_ ;
  assign \new_[2737]_  = ~\new_[4871]_  | ~\new_[5583]_  | ~\new_[2903]_  | ~\new_[5956]_ ;
  assign \new_[2738]_  = ~\new_[4580]_  | ~\new_[5614]_  | ~\new_[2904]_  | ~\new_[5615]_ ;
  assign \new_[2739]_  = ~\new_[2900]_  & (~\new_[7599]_  | ~\new_[10265]_ );
  assign \new_[2740]_  = ~\new_[2902]_  & (~\new_[7067]_  | ~\new_[9989]_ );
  assign \new_[2741]_  = ~\new_[2932]_  | ~\new_[5567]_ ;
  assign \new_[2742]_  = ~\new_[4841]_  | ~\new_[5507]_  | ~\new_[2923]_  | ~\new_[5508]_ ;
  assign \new_[2743]_  = ~\new_[10231]_  | ~\new_[2922]_  | ~\new_[10139]_ ;
  assign \new_[2744]_  = ~\new_[4843]_  | ~\new_[5509]_  | ~\new_[2924]_  | ~\new_[5917]_ ;
  assign \new_[2745]_  = ~\new_[4848]_  | ~\new_[5527]_  | ~\new_[2925]_  | ~\new_[5528]_ ;
  assign \new_[2746]_  = ~\new_[4849]_  | ~\new_[5036]_  | ~\new_[2901]_  | ~\new_[5529]_ ;
  assign \new_[2747]_  = ~\new_[4850]_  | ~\new_[5531]_  | ~\new_[2962]_  | ~\new_[5533]_ ;
  assign \new_[2748]_  = ~\new_[4851]_  | ~\new_[5536]_  | ~\new_[2926]_  | ~\new_[5040]_ ;
  assign \new_[2749]_  = ~\new_[4856]_  | ~\new_[5549]_  | ~\new_[2928]_  | ~\new_[5550]_ ;
  assign \new_[2750]_  = ~\new_[4857]_  | ~\new_[5063]_  | ~\new_[2929]_  | ~\new_[5555]_ ;
  assign \new_[2751]_  = ~\new_[4859]_  | ~\new_[5561]_  | ~\new_[2930]_  | ~\new_[5562]_ ;
  assign \new_[2752]_  = ~\new_[4860]_  | ~\new_[5565]_  | ~\new_[2931]_  | ~\new_[5938]_ ;
  assign \new_[2753]_  = ~\new_[4862]_  | ~\new_[5568]_  | ~\new_[2933]_  | ~\new_[5940]_ ;
  assign \new_[2754]_  = ~\new_[4864]_  | ~\new_[5941]_  | ~\new_[2934]_  | ~\new_[5942]_ ;
  assign \new_[2755]_  = ~\new_[4569]_  | ~\new_[5554]_  | ~\new_[2935]_  | ~\new_[5944]_ ;
  assign \new_[2756]_  = ~\new_[4866]_  | ~\new_[5946]_  | ~\new_[2936]_  | ~\new_[5947]_ ;
  assign \new_[2757]_  = ~\new_[4867]_  | ~\new_[5574]_  | ~\new_[2937]_  | ~\new_[5948]_ ;
  assign \new_[2758]_  = ~\new_[4872]_  | ~\new_[5587]_  | ~\new_[2939]_  | ~\new_[5588]_ ;
  assign \new_[2759]_  = ~\new_[4873]_  | ~\new_[5960]_  | ~\new_[2940]_  | ~\new_[5961]_ ;
  assign \new_[2760]_  = ~\new_[4574]_  | ~\new_[5963]_  | ~\new_[2941]_  | ~\new_[5964]_ ;
  assign \new_[2761]_  = ~\new_[4877]_  | ~\new_[5582]_  | ~\new_[2942]_  | ~\new_[5967]_ ;
  assign \new_[2762]_  = ~\new_[4842]_  | ~\new_[5599]_  | ~\new_[2943]_  | ~\new_[5970]_ ;
  assign \new_[2763]_  = ~\new_[4879]_  | ~\new_[5600]_  | ~\new_[2944]_  | ~\new_[5601]_ ;
  assign \new_[2764]_  = ~\new_[4883]_  | ~\new_[5506]_  | ~\new_[2945]_  | ~\new_[5971]_ ;
  assign \new_[2765]_  = ~\new_[4885]_  | ~\new_[5973]_  | ~\new_[2946]_  | ~\new_[5974]_ ;
  assign \new_[2766]_  = ~\new_[2831]_ ;
  assign \new_[2767]_  = ~\\u1_bank_adr_reg[1] ;
  assign \new_[2768]_  = \\u1_row_adr_reg[9] ;
  assign \new_[2769]_  = \\u1_row_adr_reg[12] ;
  assign \new_[2770]_  = ~\new_[2955]_  & (~\new_[12534]_  | ~\new_[10056]_ );
  assign \new_[2771]_  = ~\new_[2956]_  & (~\new_[12534]_  | ~\new_[10059]_ );
  assign \new_[2772]_  = ~\new_[2957]_  & (~\new_[12534]_  | ~\new_[10089]_ );
  assign \new_[2773]_  = ~\new_[7295]_  & (~\new_[3965]_  | ~\new_[3075]_ );
  assign \new_[2774]_  = ~\new_[10001]_  | ~\new_[2959]_  | ~\new_[12664]_ ;
  assign \new_[2775]_  = ~\new_[6545]_  | ~\new_[3219]_  | ~\new_[4263]_  | ~\new_[6092]_ ;
  assign \new_[2776]_  = ~\new_[6546]_  | ~\new_[3231]_  | ~\new_[4266]_  | ~\new_[6093]_ ;
  assign \new_[2777]_  = ~\new_[2960]_  | ~\new_[10553]_ ;
  assign \new_[2778]_  = ~\new_[3086]_  | ~\new_[6078]_  | ~\new_[3053]_  | ~\new_[4607]_ ;
  assign \new_[2779]_  = ~\new_[3088]_  | ~\new_[6079]_  | ~\new_[3055]_  | ~\new_[4610]_ ;
  assign \new_[2780]_  = ~\new_[3090]_  | ~\new_[6080]_  | ~\new_[2951]_  | ~\new_[4618]_ ;
  assign \new_[2781]_  = ~\new_[3094]_  | ~\new_[6082]_  | ~\new_[2952]_  | ~\new_[4628]_ ;
  assign \new_[2782]_  = ~\new_[3096]_  | ~\new_[6084]_  | ~\new_[2953]_  | ~\new_[4630]_ ;
  assign \new_[2783]_  = ~\new_[3097]_  | ~\new_[6085]_  | ~\new_[2954]_  | ~\new_[4632]_ ;
  assign \new_[2784]_  = ~\new_[4609]_  | ~\new_[3226]_  | ~\new_[6165]_  | ~\new_[6124]_ ;
  assign \new_[2785]_  = ~\new_[4634]_  | ~\new_[3229]_  | ~\new_[6192]_  | ~\new_[6144]_ ;
  assign \new_[2786]_  = ~\new_[4638]_  | ~\new_[3230]_  | ~\new_[6201]_  | ~\new_[6152]_ ;
  assign \new_[2787]_  = ~\new_[5716]_  | ~\new_[4265]_  | ~\new_[2994]_ ;
  assign \new_[2788]_  = ~\new_[5717]_  | ~\new_[4267]_  | ~\new_[2995]_ ;
  assign \new_[2789]_  = ~\new_[5365]_  | ~\new_[4268]_  | ~\new_[2996]_ ;
  assign \new_[2790]_  = ~\new_[5718]_  | ~\new_[4269]_  | ~\new_[2997]_ ;
  assign \new_[2791]_  = ~\new_[5719]_  | ~\new_[4270]_  | ~\new_[2999]_ ;
  assign \new_[2792]_  = ~\new_[5366]_  | ~\new_[4271]_  | ~\new_[3000]_ ;
  assign \new_[2793]_  = ~\new_[5368]_  | ~\new_[4274]_  | ~\new_[3001]_ ;
  assign \new_[2794]_  = ~\new_[5369]_  | ~\new_[4275]_  | ~\new_[3002]_ ;
  assign \new_[2795]_  = ~\new_[5721]_  | ~\new_[4111]_  | ~\new_[3003]_ ;
  assign \new_[2796]_  = ~\new_[5726]_  | ~\new_[4116]_  | ~\new_[3004]_ ;
  assign \new_[2797]_  = ~\new_[5374]_  | ~\new_[4283]_  | ~\new_[3017]_ ;
  assign \new_[2798]_  = ~\new_[5741]_  | ~\new_[4286]_  | ~\new_[3020]_ ;
  assign \new_[2799]_  = ~\new_[5376]_  | ~\new_[4139]_  | ~\new_[3023]_ ;
  assign \new_[2800]_  = ~\new_[5744]_  | ~\new_[4264]_  | ~\new_[3025]_ ;
  assign n1696 = ~\new_[3121]_  | ~\new_[3111]_  | ~\new_[3098]_  | ~\new_[2983]_ ;
  assign \new_[2802]_  = ~\new_[2963]_  & (~\new_[7682]_  | ~\new_[9842]_ );
  assign \new_[2803]_  = ~\new_[2966]_  & ~\new_[3092]_ ;
  assign \new_[2804]_  = ~\new_[2967]_  & ~\new_[3009]_ ;
  assign \new_[2805]_  = ~\new_[5763]_  | ~\new_[11846]_  | ~\new_[2968]_  | ~\new_[3775]_ ;
  assign \new_[2806]_  = (~\new_[3030]_  | ~\new_[10001]_ ) & (~\new_[7100]_  | ~\new_[6393]_ );
  assign \new_[2807]_  = \new_[2889]_  | \new_[4836]_ ;
  assign \new_[2808]_  = ~\new_[5589]_  | ~\new_[2895]_  | ~\new_[3150]_ ;
  assign \new_[2809]_  = ~\new_[2887]_  & ~\new_[3035]_ ;
  assign \new_[2810]_  = ~\new_[3670]_  | ~\new_[5928]_  | ~\new_[3294]_  | ~\new_[4177]_ ;
  assign \new_[2811]_  = ~\new_[3083]_  & ~\new_[3008]_ ;
  assign \new_[2812]_  = ~\new_[2985]_  & ~\new_[3012]_ ;
  assign \new_[2813]_  = ~\new_[3301]_  | ~\new_[5591]_  | ~\new_[3132]_  | ~\new_[4600]_ ;
  assign \new_[2814]_  = ~\new_[2986]_  & ~\new_[3015]_ ;
  assign \new_[2815]_  = ~\new_[2987]_  & ~\new_[2982]_ ;
  assign \new_[2816]_  = ~\new_[2989]_  & ~\new_[3021]_ ;
  assign \new_[2817]_  = ~\new_[2990]_  & ~\new_[3022]_ ;
  assign \new_[2818]_  = ~\new_[2993]_  & (~\new_[6826]_  | ~\new_[9391]_ );
  assign \new_[2819]_  = ~\new_[2992]_  & (~\new_[12385]_  | ~\new_[9938]_ );
  assign \new_[2820]_  = ~\new_[2884]_ ;
  assign n1701 = \new_[11080]_  ? n5766 : \new_[3136]_ ;
  assign n1706 = \new_[2720]_  ? n5766 : \new_[3137]_ ;
  assign n1711 = \new_[2721]_  ? n5766 : \new_[3174]_ ;
  assign \new_[2824]_  = ~\new_[6176]_  | ~\new_[3039]_  | ~\new_[5752]_ ;
  assign \new_[2825]_  = ~\new_[3051]_  | ~\new_[6182]_ ;
  assign \new_[2826]_  = ~\new_[3052]_  | ~\new_[6186]_ ;
  assign \new_[2827]_  = ~\new_[6194]_  | ~\new_[3040]_  | ~\new_[5383]_ ;
  assign \new_[2828]_  = ~\new_[3038]_  & (~\new_[12534]_  | ~\new_[10053]_ );
  assign \new_[2829]_  = \\u1_row_adr_reg[3] ;
  assign \new_[2830]_  = \\u1_row_adr_reg[7] ;
  assign \new_[2831]_  = ~\new_[4875]_  | ~\new_[5594]_  | ~\new_[3071]_  | ~\new_[5966]_ ;
  assign \new_[2832]_  = ~\new_[4895]_  | ~\new_[5603]_  | ~\new_[3072]_  | ~\new_[5604]_ ;
  assign \new_[2833]_  = \\u1_row_adr_reg[0] ;
  assign \new_[2834]_  = ~\new_[3054]_  & (~\new_[12534]_  | ~\new_[10054]_ );
  assign \new_[2835]_  = ~\new_[3056]_  & (~\new_[12534]_  | ~\new_[9912]_ );
  assign \new_[2836]_  = ~\new_[3057]_  & (~\new_[12534]_  | ~\new_[10065]_ );
  assign \new_[2837]_  = ~\\u1_acs_addr_reg[23] ;
  assign \new_[2838]_  = ~\new_[3058]_  & (~\new_[12534]_  | ~\new_[10046]_ );
  assign \new_[2839]_  = \\u1_row_adr_reg[1] ;
  assign \new_[2840]_  = \\u1_row_adr_reg[2] ;
  assign \new_[2841]_  = \\u1_row_adr_reg[4] ;
  assign \new_[2842]_  = \\u1_row_adr_reg[5] ;
  assign \new_[2843]_  = \\u1_row_adr_reg[6] ;
  assign \new_[2844]_  = ~\new_[3059]_  & (~\new_[12534]_  | ~\new_[9880]_ );
  assign \new_[2845]_  = \\u1_row_adr_reg[8] ;
  assign \new_[2846]_  = ~\new_[3060]_  & (~\new_[12534]_  | ~\new_[9849]_ );
  assign \new_[2847]_  = ~\new_[3061]_  & (~\new_[12534]_  | ~\new_[10081]_ );
  assign \new_[2848]_  = ~\new_[3062]_  & (~\new_[12534]_  | ~\new_[10130]_ );
  assign \new_[2849]_  = ~\new_[3063]_  & (~\new_[12534]_  | ~\new_[10061]_ );
  assign \new_[2850]_  = ~\new_[3064]_  & (~\new_[12534]_  | ~\new_[9668]_ );
  assign \new_[2851]_  = ~\new_[3065]_  & (~\new_[12534]_  | ~\new_[10071]_ );
  assign \new_[2852]_  = ~\new_[3066]_  & (~\new_[12534]_  | ~\new_[9649]_ );
  assign \new_[2853]_  = ~\new_[3067]_  & (~\new_[12534]_  | ~\new_[10153]_ );
  assign \new_[2854]_  = ~\new_[3068]_  & (~\new_[12534]_  | ~\new_[10118]_ );
  assign \new_[2855]_  = ~\new_[3069]_  & (~\new_[12534]_  | ~\new_[9904]_ );
  assign \new_[2856]_  = ~\new_[3070]_  & (~\new_[12534]_  | ~\new_[9871]_ );
  assign \new_[2857]_  = ~\new_[3073]_  & ~\new_[9341]_ ;
  assign \new_[2858]_  = ~\new_[3074]_  & (~\new_[6029]_  | ~\new_[11316]_ );
  assign \new_[2859]_  = ~\new_[3078]_  & ~\new_[3221]_ ;
  assign \new_[2860]_  = ~\new_[6721]_  | ~\new_[11503]_  | ~\new_[3099]_ ;
  assign \new_[2861]_  = ~\new_[4903]_  & ~\new_[3080]_ ;
  assign \new_[2862]_  = ~\new_[4904]_  & ~\new_[3081]_ ;
  assign \new_[2863]_  = ~\new_[6081]_  | ~\new_[4626]_  | ~\new_[3093]_ ;
  assign \new_[2864]_  = ~\new_[6083]_  | ~\new_[4629]_  | ~\new_[3095]_ ;
  assign \new_[2865]_  = ~\new_[4920]_  & ~\new_[3082]_ ;
  assign \new_[2866]_  = ~\new_[3289]_  | ~\new_[5526]_  | ~\new_[3026]_  | ~\new_[4253]_ ;
  assign n1716 = ~\new_[3775]_  | ~\new_[2970]_  | ~\new_[6367]_ ;
  assign \new_[2868]_  = (~\new_[3101]_  | ~\new_[10001]_ ) & (~\new_[7353]_  | ~\new_[11453]_ );
  assign \new_[2869]_  = (~\new_[3104]_  | ~\new_[10001]_ ) & (~\new_[7093]_  | ~\new_[11453]_ );
  assign \new_[2870]_  = (~\new_[3105]_  | ~\new_[10001]_ ) & (~\new_[7098]_  | ~\new_[11453]_ );
  assign \new_[2871]_  = (~\new_[3106]_  | ~\new_[10001]_ ) & (~\new_[7103]_  | ~\new_[6393]_ );
  assign \new_[2872]_  = (~\new_[3102]_  | ~\new_[10001]_ ) & (~\new_[7995]_  | ~\new_[12306]_ );
  assign \new_[2873]_  = (~\new_[3107]_  | ~\new_[10001]_ ) & (~\new_[7087]_  | ~\new_[6393]_ );
  assign \new_[2874]_  = \new_[3006]_  | \new_[5727]_ ;
  assign \new_[2875]_  = \new_[3016]_  | \new_[5737]_ ;
  assign \new_[2876]_  = \new_[3018]_  | \new_[5739]_ ;
  assign \new_[2877]_  = \new_[3019]_  | \new_[5740]_ ;
  assign \new_[2878]_  = ~\new_[5504]_  | ~\new_[5789]_  | ~\new_[3115]_ ;
  assign \new_[2879]_  = ~\new_[5930]_  | ~\new_[3142]_  | ~\new_[6734]_ ;
  assign \new_[2880]_  = \new_[3013]_  | \new_[4837]_ ;
  assign \new_[2881]_  = ~\new_[5952]_  | ~\new_[8002]_  | ~\new_[3147]_ ;
  assign \new_[2882]_  = ~\new_[3085]_  & (~\new_[6826]_  | ~\new_[8977]_ );
  assign \new_[2883]_  = ~\new_[3100]_  & (~\new_[3704]_  | ~\new_[5703]_ );
  assign \new_[2884]_  = ~\new_[3385]_  | ~\new_[5955]_  | ~\new_[3273]_  | ~\new_[4290]_ ;
  assign n1726 = \new_[2768]_  ? n5766 : \new_[3267]_ ;
  assign n1721 = \new_[11179]_  ? n5766 : \new_[3285]_ ;
  assign \new_[2887]_  = ~\new_[7463]_  | ~\new_[3133]_  | ~\new_[4978]_ ;
  assign \new_[2888]_  = ~\new_[6986]_  | ~\new_[3117]_ ;
  assign \new_[2889]_  = ~\new_[7156]_  & (~\new_[3463]_  | ~\new_[3307]_ );
  assign \new_[2890]_  = ~\new_[6985]_  | ~\new_[3122]_ ;
  assign \new_[2891]_  = ~\new_[3028]_ ;
  assign \new_[2892]_  = ~\new_[3029]_ ;
  assign \new_[2893]_  = ~\new_[3031]_ ;
  assign \new_[2894]_  = ~\new_[3032]_ ;
  assign \new_[2895]_  = ~\new_[3120]_  & (~\new_[4840]_  | ~\new_[9978]_ );
  assign \new_[2896]_  = ~\new_[3033]_ ;
  assign \new_[2897]_  = ~\new_[3034]_ ;
  assign \new_[2898]_  = ~\new_[3118]_  & (~\new_[7329]_  | ~\new_[9655]_ );
  assign \new_[2899]_  = ~\new_[4579]_  | ~\new_[5610]_  | ~\new_[5611]_  | ~\new_[3318]_ ;
  assign \new_[2900]_  = ~\new_[6105]_  | ~\new_[3468]_  | ~\new_[6106]_  | ~\new_[4821]_ ;
  assign \new_[2901]_  = ~\new_[3192]_  & (~\new_[12534]_  | ~\new_[9737]_ );
  assign \new_[2902]_  = ~\new_[3175]_  | ~\new_[5634]_ ;
  assign \new_[2903]_  = ~\new_[3168]_  & (~\new_[12534]_  | ~\new_[9846]_ );
  assign \new_[2904]_  = ~\new_[3154]_  & (~\new_[12534]_  | ~\new_[10063]_ );
  assign \new_[2905]_  = ~\new_[3155]_  & (~\new_[11864]_  | ~\new_[10039]_ );
  assign \new_[2906]_  = ~\new_[3156]_  & (~\new_[11864]_  | ~\new_[9401]_ );
  assign \new_[2907]_  = ~\new_[3157]_  & (~\new_[6652]_  | ~\new_[9661]_ );
  assign \new_[2908]_  = ~\new_[3158]_  & (~\new_[6652]_  | ~\new_[9963]_ );
  assign \new_[2909]_  = ~\new_[3159]_  & (~\new_[11864]_  | ~\new_[9995]_ );
  assign \new_[2910]_  = ~\new_[3160]_  & (~\new_[11864]_  | ~\new_[10237]_ );
  assign \new_[2911]_  = ~\new_[3161]_  & (~\new_[11864]_  | ~\new_[9660]_ );
  assign \new_[2912]_  = ~\new_[3162]_  & (~\new_[6652]_  | ~\new_[9641]_ );
  assign \new_[2913]_  = ~\new_[3163]_  & (~\new_[11864]_  | ~\new_[10111]_ );
  assign \new_[2914]_  = ~\new_[3164]_  & (~\new_[6652]_  | ~\new_[10052]_ );
  assign \new_[2915]_  = ~\new_[12298]_  & (~\new_[11864]_  | ~\new_[9388]_ );
  assign \new_[2916]_  = ~\new_[3165]_  & (~\new_[6652]_  | ~\new_[10019]_ );
  assign \new_[2917]_  = ~\new_[3166]_  & (~\new_[11864]_  | ~\new_[9657]_ );
  assign \new_[2918]_  = ~\new_[3170]_  & (~\new_[11864]_  | ~\new_[9599]_ );
  assign \new_[2919]_  = ~\new_[3171]_  & (~\new_[6652]_  | ~\new_[9407]_ );
  assign \new_[2920]_  = ~\new_[3172]_  & (~\new_[11864]_  | ~\new_[9990]_ );
  assign \new_[2921]_  = ~\new_[3173]_  & (~\new_[11864]_  | ~\new_[10037]_ );
  assign \new_[2922]_  = ~\new_[3868]_  & ~\new_[3188]_ ;
  assign \new_[2923]_  = ~\new_[3189]_  & (~\new_[12534]_  | ~\new_[9953]_ );
  assign \new_[2924]_  = ~\new_[3190]_  & (~\new_[12534]_  | ~\new_[12060]_ );
  assign \new_[2925]_  = ~\new_[3191]_  & (~\new_[12534]_  | ~\new_[9822]_ );
  assign \new_[2926]_  = ~\new_[3194]_  & (~\new_[12534]_  | ~\new_[10078]_ );
  assign \new_[2927]_  = u5_cnt_reg;
  assign \new_[2928]_  = ~\new_[3195]_  & (~\new_[12534]_  | ~\new_[10082]_ );
  assign \new_[2929]_  = ~\new_[3196]_  & (~\new_[12534]_  | ~\new_[9807]_ );
  assign \new_[2930]_  = ~\new_[3197]_  & (~\new_[12534]_  | ~\new_[9694]_ );
  assign \new_[2931]_  = ~\new_[3198]_  & (~\new_[12534]_  | ~\new_[9965]_ );
  assign \new_[2932]_  = ~\new_[3199]_  & (~\new_[5865]_  | ~\new_[9326]_ );
  assign \new_[2933]_  = ~\new_[3200]_  & (~\new_[12534]_  | ~\new_[10055]_ );
  assign \new_[2934]_  = ~\new_[3201]_  & (~\new_[12534]_  | ~\new_[9841]_ );
  assign \new_[2935]_  = ~\new_[3202]_  & (~\new_[12534]_  | ~\new_[9610]_ );
  assign \new_[2936]_  = ~\new_[3203]_  & (~\new_[12534]_  | ~\new_[9843]_ );
  assign \new_[2937]_  = ~\new_[3204]_  & (~\new_[12534]_  | ~\new_[10087]_ );
  assign \new_[2938]_  = ~\new_[3205]_  & (~\new_[7239]_  | ~\new_[9657]_ );
  assign \new_[2939]_  = ~\new_[3206]_  & (~\new_[12534]_  | ~\new_[9847]_ );
  assign \new_[2940]_  = ~\new_[3207]_  & (~\new_[12534]_  | ~\new_[9872]_ );
  assign \new_[2941]_  = ~\new_[3209]_  & (~\new_[12534]_  | ~\new_[10051]_ );
  assign \new_[2942]_  = ~\new_[3210]_  & (~\new_[12534]_  | ~\new_[10044]_ );
  assign \new_[2943]_  = ~\new_[3211]_  & (~\new_[12534]_  | ~\new_[10049]_ );
  assign \new_[2944]_  = ~\new_[3212]_  & (~\new_[12534]_  | ~\new_[10050]_ );
  assign \new_[2945]_  = ~\new_[3213]_  & (~\new_[12534]_  | ~\new_[10043]_ );
  assign \new_[2946]_  = ~\new_[3214]_  & (~\new_[12534]_  | ~\new_[10048]_ );
  assign \new_[2947]_  = ~\new_[3215]_  & (~\new_[12534]_  | ~\new_[10107]_ );
  assign \new_[2948]_  = ~\new_[3187]_  & (~\new_[12534]_  | ~\new_[9967]_ );
  assign n1731 = \new_[2769]_  ? n5766 : \new_[3232]_ ;
  assign \new_[2950]_  = ~\new_[5412]_  & ~\new_[3218]_ ;
  assign \new_[2951]_  = ~\new_[5413]_  & ~\new_[3220]_ ;
  assign \new_[2952]_  = ~\new_[4605]_  & ~\new_[3222]_ ;
  assign \new_[2953]_  = ~\new_[5414]_  & ~\new_[3223]_ ;
  assign \new_[2954]_  = ~\new_[4606]_  & ~\new_[3224]_ ;
  assign \new_[2955]_  = ~\new_[4312]_  | ~\new_[3349]_  | ~\new_[5493]_  | ~\new_[6698]_ ;
  assign \new_[2956]_  = ~\new_[4469]_  | ~\new_[3350]_  | ~\new_[6033]_  | ~\new_[6715]_ ;
  assign \new_[2957]_  = ~\new_[4466]_  | ~\new_[3351]_  | ~\new_[5496]_  | ~\new_[6716]_ ;
  assign \new_[2958]_  = ~\new_[6986]_  | ~\new_[3217]_ ;
  assign \new_[2959]_  = ~\new_[3327]_  | ~\new_[3771]_  | ~\new_[3923]_ ;
  assign \new_[2960]_  = ~\new_[12665]_  & (~\new_[3233]_  | ~\new_[10010]_ );
  assign \new_[2961]_  = ~\new_[3227]_  & (~\new_[12534]_  | ~\new_[9870]_ );
  assign \new_[2962]_  = ~\new_[3193]_  & (~\new_[12534]_  | ~\new_[9854]_ );
  assign \new_[2963]_  = ~\new_[3089]_  | ~\new_[6074]_ ;
  assign \new_[2964]_  = ~\new_[4838]_  & (~\new_[6985]_  | ~\new_[3261]_ );
  assign \new_[2965]_  = ~\new_[5746]_  & (~\new_[6985]_  | ~\new_[3253]_ );
  assign \new_[2966]_  = ~\new_[7456]_  | ~\new_[3109]_  | ~\new_[5471]_ ;
  assign \new_[2967]_  = ~\new_[7448]_  | ~\new_[3110]_  | ~\new_[5472]_ ;
  assign \new_[2968]_  = ~\new_[3348]_  & ~\new_[3084]_ ;
  assign \new_[2969]_  = ~\new_[3108]_  & (~\new_[3704]_  | ~\new_[5695]_ );
  assign \new_[2970]_  = ~\new_[3239]_  & ~\new_[12470]_ ;
  assign \new_[2971]_  = \\u3_byte1_reg[5] ;
  assign \new_[2972]_  = ~\new_[3236]_  & (~\new_[12780]_  | ~\new_[9937]_ );
  assign n1746 = \new_[2833]_  ? n5766 : \new_[3372]_ ;
  assign n1756 = \new_[2839]_  ? n5766 : \new_[3373]_ ;
  assign n1761 = \new_[2840]_  ? n5766 : \new_[3374]_ ;
  assign n1736 = \new_[2829]_  ? n5766 : \new_[3375]_ ;
  assign n1766 = \new_[2841]_  ? n5766 : \new_[3376]_ ;
  assign n1771 = \new_[2842]_  ? n5766 : \new_[3377]_ ;
  assign n1776 = \new_[2843]_  ? n5766 : \new_[3378]_ ;
  assign n1741 = \new_[2830]_  ? n5766 : \new_[3379]_ ;
  assign n1781 = \new_[2845]_  ? n5766 : \new_[3380]_ ;
  assign \new_[2982]_  = ~\new_[5632]_  | ~\new_[3560]_  | ~\new_[5503]_  | ~\new_[5623]_ ;
  assign \new_[2983]_  = ~\new_[3243]_  | ~\new_[12664]_ ;
  assign \new_[2984]_  = ~\new_[7461]_  | ~\new_[3270]_  | ~\new_[4965]_ ;
  assign \new_[2985]_  = ~\new_[7466]_  | ~\new_[3274]_  | ~\new_[5449]_ ;
  assign \new_[2986]_  = ~\new_[7469]_  | ~\new_[3276]_  | ~\new_[5488]_ ;
  assign \new_[2987]_  = ~\new_[7470]_  | ~\new_[3279]_  | ~\new_[5492]_ ;
  assign \new_[2988]_  = ~\new_[7473]_  | ~\new_[3280]_  | ~\new_[5494]_ ;
  assign \new_[2989]_  = ~\new_[7453]_  | ~\new_[3282]_  | ~\new_[4985]_ ;
  assign \new_[2990]_  = ~\new_[7474]_  | ~\new_[3283]_  | ~\new_[4984]_ ;
  assign \new_[2991]_  = ~\new_[5081]_  | ~\new_[3604]_  | ~\new_[5910]_  | ~\new_[5627]_ ;
  assign \new_[2992]_  = ~\new_[5843]_  | ~\new_[7447]_  | ~\new_[6162]_  | ~\new_[3415]_ ;
  assign \new_[2993]_  = ~\new_[5866]_  | ~\new_[7458]_  | ~\new_[5915]_  | ~\new_[3427]_ ;
  assign \new_[2994]_  = ~\new_[6984]_  | ~\new_[3244]_ ;
  assign \new_[2995]_  = ~\new_[6984]_  | ~\new_[3245]_ ;
  assign \new_[2996]_  = ~\new_[6985]_  | ~\new_[3246]_ ;
  assign \new_[2997]_  = ~\new_[6985]_  | ~\new_[3247]_ ;
  assign \new_[2998]_  = \new_[3290]_  & \new_[5923]_ ;
  assign \new_[2999]_  = ~\new_[6984]_  | ~\new_[3248]_ ;
  assign \new_[3000]_  = ~\new_[6984]_  | ~\new_[3250]_ ;
  assign \new_[3001]_  = ~\new_[6984]_  | ~\new_[3252]_ ;
  assign \new_[3002]_  = ~\new_[6985]_  | ~\new_[3254]_ ;
  assign \new_[3003]_  = ~\new_[6986]_  | ~\new_[3255]_ ;
  assign \new_[3004]_  = ~\new_[6986]_  | ~\new_[3256]_ ;
  assign \new_[3005]_  = ~\new_[5053]_  | ~\new_[3591]_  | ~\new_[5566]_  | ~\new_[6607]_ ;
  assign \new_[3006]_  = ~\new_[7156]_  & (~\new_[3762]_  | ~\new_[3424]_ );
  assign \new_[3007]_  = ~\new_[6985]_  | ~\new_[3257]_ ;
  assign \new_[3008]_  = ~\new_[5055]_  | ~\new_[3592]_  | ~\new_[5569]_  | ~\new_[6727]_ ;
  assign \new_[3009]_  = ~\new_[5056]_  | ~\new_[3593]_  | ~\new_[5943]_  | ~\new_[6611]_ ;
  assign \new_[3010]_  = ~\new_[6985]_  | ~\new_[3258]_ ;
  assign \new_[3011]_  = ~\new_[6985]_  | ~\new_[3259]_ ;
  assign \new_[3012]_  = ~\new_[5073]_  | ~\new_[3599]_  | ~\new_[5590]_  | ~\new_[6583]_ ;
  assign \new_[3013]_  = ~\new_[7156]_  & (~\new_[3464]_  | ~\new_[3430]_ );
  assign \new_[3014]_  = ~\new_[6985]_  | ~\new_[3260]_ ;
  assign \new_[3015]_  = ~\new_[5077]_  | ~\new_[3601]_  | ~\new_[5595]_  | ~\new_[6623]_ ;
  assign \new_[3016]_  = ~\new_[7156]_  & (~\new_[3783]_  | ~\new_[3432]_ );
  assign \new_[3017]_  = ~\new_[6984]_  | ~\new_[3262]_ ;
  assign \new_[3018]_  = ~\new_[7156]_  & (~\new_[3789]_  | ~\new_[3433]_ );
  assign \new_[3019]_  = ~\new_[7156]_  & (~\new_[3791]_  | ~\new_[3435]_ );
  assign \new_[3020]_  = ~\new_[6984]_  | ~\new_[3263]_ ;
  assign \new_[3021]_  = ~\new_[3570]_  | ~\new_[5633]_  | ~\new_[5606]_  | ~\new_[6630]_ ;
  assign \new_[3022]_  = ~\new_[5084]_  | ~\new_[3606]_  | ~\new_[5607]_  | ~\new_[6603]_ ;
  assign \new_[3023]_  = ~\new_[6986]_  | ~\new_[3264]_ ;
  assign \new_[3024]_  = ~\new_[6984]_  | ~\new_[3265]_ ;
  assign \new_[3025]_  = ~\new_[6985]_  | ~\new_[3266]_ ;
  assign \new_[3026]_  = ~\new_[12287]_  & (~\new_[11864]_  | ~\new_[10128]_ );
  assign \new_[3027]_  = ~\new_[3249]_  & (~\new_[6652]_  | ~\new_[10011]_ );
  assign \new_[3028]_  = ~\new_[7156]_  & (~\new_[3751]_  | ~\new_[3412]_ );
  assign \new_[3029]_  = ~\new_[7156]_  & (~\new_[3756]_  | ~\new_[3407]_ );
  assign \new_[3030]_  = ~\new_[7295]_  & (~\new_[3760]_  | ~\new_[3423]_ );
  assign \new_[3031]_  = ~\new_[7156]_  & (~\new_[3461]_  | ~\new_[3408]_ );
  assign \new_[3032]_  = ~\new_[7156]_  & (~\new_[3462]_  | ~\new_[3409]_ );
  assign \new_[3033]_  = ~\new_[7156]_  & (~\new_[3465]_  | ~\new_[3410]_ );
  assign \new_[3034]_  = ~\new_[7156]_  & (~\new_[3786]_  | ~\new_[3411]_ );
  assign \new_[3035]_  = ~\new_[4717]_  | ~\new_[3499]_  | ~\new_[4898]_  | ~\new_[5078]_ ;
  assign \new_[3036]_  = u5_wb_cycle_reg;
  assign \new_[3037]_  = ~\new_[3305]_  & (~\new_[7329]_  | ~\new_[10037]_ );
  assign \new_[3038]_  = ~\new_[6696]_  | ~\new_[3319]_  | ~\new_[5441]_ ;
  assign \new_[3039]_  = ~\new_[3320]_  & (~\new_[12786]_  | ~\new_[9975]_ );
  assign \new_[3040]_  = ~\new_[3323]_  & (~\new_[12786]_  | ~\new_[10062]_ );
  assign \new_[3041]_  = \\u1_acs_addr_reg[19] ;
  assign \new_[3042]_  = \\u1_acs_addr_reg[20] ;
  assign \new_[3043]_  = \\u3_byte1_reg[0] ;
  assign \new_[3044]_  = \\u3_byte1_reg[1] ;
  assign \new_[3045]_  = \\u3_byte1_reg[2] ;
  assign \new_[3046]_  = \\u3_byte1_reg[3] ;
  assign \new_[3047]_  = \\u3_byte1_reg[4] ;
  assign \new_[3048]_  = \\u3_byte1_reg[7] ;
  assign \new_[3049]_  = \\u3_byte1_reg[6] ;
  assign \new_[3050]_  = ~\\u1_col_adr_reg[8] ;
  assign \new_[3051]_  = ~\new_[3321]_  & (~\new_[5865]_  | ~\new_[10111]_ );
  assign \new_[3052]_  = ~\new_[3322]_  & (~\new_[5865]_  | ~\new_[11860]_ );
  assign \new_[3053]_  = ~\new_[5410]_  & ~\new_[3331]_ ;
  assign \new_[3054]_  = ~\new_[4304]_  | ~\new_[3476]_  | ~\new_[5438]_  | ~\new_[6498]_ ;
  assign \new_[3055]_  = ~\new_[5411]_  & ~\new_[3332]_ ;
  assign \new_[3056]_  = ~\new_[4656]_  | ~\new_[3478]_  | ~\new_[5845]_  | ~\new_[6499]_ ;
  assign \new_[3057]_  = ~\new_[4308]_  | ~\new_[3479]_  | ~\new_[5846]_  | ~\new_[6500]_ ;
  assign \new_[3058]_  = ~\new_[4659]_  | ~\new_[3480]_  | ~\new_[5847]_  | ~\new_[6501]_ ;
  assign \new_[3059]_  = ~\new_[4667]_  | ~\new_[3483]_  | ~\new_[5852]_  | ~\new_[6507]_ ;
  assign \new_[3060]_  = ~\new_[4315]_  | ~\new_[3484]_  | ~\new_[5448]_  | ~\new_[6508]_ ;
  assign \new_[3061]_  = ~\new_[4673]_  | ~\new_[3485]_  | ~\new_[5853]_  | ~\new_[6509]_ ;
  assign \new_[3062]_  = ~\new_[4320]_  | ~\new_[3486]_  | ~\new_[5854]_  | ~\new_[6510]_ ;
  assign \new_[3063]_  = ~\new_[4321]_  | ~\new_[3487]_  | ~\new_[5455]_  | ~\new_[6512]_ ;
  assign \new_[3064]_  = ~\new_[4323]_  | ~\new_[3488]_  | ~\new_[5458]_  | ~\new_[6700]_ ;
  assign \new_[3065]_  = ~\new_[4326]_  | ~\new_[3489]_  | ~\new_[5857]_  | ~\new_[6515]_ ;
  assign \new_[3066]_  = ~\new_[4330]_  | ~\new_[3490]_  | ~\new_[5468]_  | ~\new_[6701]_ ;
  assign \new_[3067]_  = ~\new_[4435]_  | ~\new_[3491]_  | ~\new_[5618]_  | ~\new_[6519]_ ;
  assign \new_[3068]_  = ~\new_[4700]_  | ~\new_[3492]_  | ~\new_[5862]_  | ~\new_[6520]_ ;
  assign \new_[3069]_  = ~\new_[4446]_  | ~\new_[3493]_  | ~\new_[5476]_  | ~\new_[6521]_ ;
  assign \new_[3070]_  = ~\new_[4460]_  | ~\new_[3495]_  | ~\new_[5872]_  | ~\new_[6525]_ ;
  assign \new_[3071]_  = ~\new_[3329]_  & (~\new_[12534]_  | ~\new_[10015]_ );
  assign \new_[3072]_  = ~\new_[3330]_  & (~\new_[12534]_  | ~\new_[10140]_ );
  assign \new_[3073]_  = ~\new_[11713]_  | ~\new_[3326]_  | ~\new_[9885]_ ;
  assign \new_[3074]_  = ~\new_[5878]_  | (~\new_[9744]_  & ~\new_[3470]_ );
  assign \new_[3075]_  = ~\new_[3328]_  & (~\new_[9632]_  | ~\new_[5247]_ );
  assign n1751 = \new_[3333]_  | \new_[5008]_ ;
  assign \new_[3077]_  = ~\\u1_acs_addr_reg[22] ;
  assign \new_[3078]_  = (~\new_[6632]_  & ~\new_[3500]_  & ~\new_[7292]_ ) | (~\new_[3653]_  & ~\new_[7063]_  & ~\new_[7662]_ );
  assign \new_[3079]_  = (~\new_[3338]_  | ~\new_[5621]_ ) & (~\new_[3337]_  | ~\new_[6208]_ );
  assign \new_[3080]_  = \new_[3234]_  | \new_[5723]_ ;
  assign \new_[3081]_  = \new_[3235]_  | \new_[5724]_ ;
  assign \new_[3082]_  = \new_[3237]_  | \new_[5742]_ ;
  assign \new_[3083]_  = ~\new_[7462]_  | ~\new_[3361]_  | ~\new_[4951]_ ;
  assign \new_[3084]_  = ~\new_[5833]_  | ~\new_[3959]_  | ~\new_[3533]_ ;
  assign \new_[3085]_  = ~\new_[5861]_  | ~\new_[7465]_  | ~\new_[5912]_  | ~\new_[3545]_ ;
  assign \new_[3086]_  = ~\new_[6985]_  | ~\new_[3355]_ ;
  assign \new_[3087]_  = \new_[3381]_  & \new_[5916]_ ;
  assign \new_[3088]_  = ~\new_[6985]_  | ~\new_[3356]_ ;
  assign \new_[3089]_  = ~\new_[6985]_  | ~\new_[3358]_ ;
  assign \new_[3090]_  = ~\new_[6985]_  | ~\new_[3359]_ ;
  assign \new_[3091]_  = \new_[3383]_  & \new_[5929]_ ;
  assign \new_[3092]_  = ~\new_[5054]_  | ~\new_[3805]_  | ~\new_[5939]_  | ~\new_[6609]_ ;
  assign \new_[3093]_  = ~\new_[6985]_  | ~\new_[12524]_ ;
  assign \new_[3094]_  = ~\new_[6985]_  | ~\new_[3366]_ ;
  assign \new_[3095]_  = ~\new_[6985]_  | ~\new_[3367]_ ;
  assign \new_[3096]_  = ~\new_[6985]_  | ~\new_[3368]_ ;
  assign \new_[3097]_  = ~\new_[6985]_  | ~\new_[3369]_ ;
  assign \new_[3098]_  = ~\new_[3348]_  & ~\new_[4559]_ ;
  assign \new_[3099]_  = ~\new_[3354]_  | ~\new_[12664]_ ;
  assign \new_[3100]_  = ~\new_[3353]_  & ~\new_[4152]_ ;
  assign \new_[3101]_  = ~\new_[7295]_  & (~\new_[3943]_  | ~\new_[3534]_ );
  assign \new_[3102]_  = ~\new_[7295]_  & (~\new_[3728]_  | ~\new_[3535]_ );
  assign \new_[3103]_  = ~\new_[7178]_  | ~\new_[3346]_  | ~\new_[5621]_ ;
  assign \new_[3104]_  = ~\new_[7295]_  & (~\new_[3750]_  | ~\new_[3538]_ );
  assign \new_[3105]_  = ~\new_[7295]_  & (~\new_[3757]_  | ~\new_[3540]_ );
  assign \new_[3106]_  = ~\new_[7295]_  & (~\new_[3767]_  | ~\new_[3543]_ );
  assign \new_[3107]_  = ~\new_[7295]_  & (~\new_[3779]_  | ~\new_[3531]_ );
  assign \new_[3108]_  = ~\new_[3352]_  & ~\new_[3556]_ ;
  assign \new_[3109]_  = ~\new_[3360]_  & (~\new_[6679]_  | ~\new_[9611]_ );
  assign \new_[3110]_  = ~\new_[3362]_  & (~\new_[6679]_  | ~\new_[9644]_ );
  assign \new_[3111]_  = ~\new_[7263]_  & ~\new_[3413]_ ;
  assign \new_[3112]_  = ~\\u1_acs_addr_reg[9] ;
  assign \new_[3113]_  = ~\\u1_acs_addr_reg[10] ;
  assign \new_[3114]_  = \\u1_acs_addr_reg[2] ;
  assign \new_[3115]_  = ~\new_[3420]_  & ~\new_[4893]_ ;
  assign \new_[3116]_  = ~\new_[3915]_  | ~\new_[3753]_  | ~\new_[3579]_ ;
  assign \new_[3117]_  = ~\new_[3920]_  | ~\new_[3460]_  | ~\new_[3766]_ ;
  assign \new_[3118]_  = ~\new_[6031]_  | ~\new_[7464]_  | ~\new_[3425]_  | ~\new_[5409]_ ;
  assign \new_[3119]_  = ~\new_[3924]_  | ~\new_[3772]_  | ~\new_[3580]_ ;
  assign \new_[3120]_  = ~\new_[3679]_  | ~\new_[7391]_  | ~\new_[4802]_  | ~\new_[7241]_ ;
  assign \new_[3121]_  = ~\new_[3431]_  & ~\new_[5800]_ ;
  assign \new_[3122]_  = ~\new_[3932]_  | ~\new_[3466]_  | ~\new_[3794]_ ;
  assign \new_[3123]_  = ~\new_[3436]_  & (~\new_[12776]_  | ~\new_[10099]_ );
  assign \new_[3124]_  = ~\new_[3437]_  & (~\new_[12776]_  | ~\new_[10104]_ );
  assign \new_[3125]_  = ~\new_[3416]_  & (~\new_[11864]_  | ~\new_[10099]_ );
  assign \new_[3126]_  = ~\new_[3417]_  & (~\new_[11864]_  | ~\new_[10104]_ );
  assign \new_[3127]_  = ~\new_[3418]_  & (~\new_[6652]_  | ~\new_[9680]_ );
  assign \new_[3128]_  = ~\new_[3419]_  & (~\new_[11864]_  | ~\new_[9845]_ );
  assign \new_[3129]_  = ~\new_[3421]_  & (~\new_[11864]_  | ~\new_[10126]_ );
  assign \new_[3130]_  = ~\new_[3422]_  & (~\new_[11864]_  | ~\new_[9987]_ );
  assign \new_[3131]_  = ~\new_[3428]_  & (~\new_[11864]_  | ~\new_[9595]_ );
  assign \new_[3132]_  = ~\new_[3429]_  & (~\new_[11864]_  | ~\new_[10083]_ );
  assign \new_[3133]_  = ~\new_[11968]_  & (~\new_[6679]_  | ~\new_[10115]_ );
  assign \new_[3134]_  = ~\new_[3434]_  & (~\new_[11864]_  | ~\new_[9604]_ );
  assign \new_[3135]_  = ~\new_[3390]_  & (~\new_[12775]_  | ~\new_[10039]_ );
  assign \new_[3136]_  = \new_[3892]_  ? \new_[6075]_  : \new_[3596]_ ;
  assign \new_[3137]_  = \new_[3608]_  ? \new_[6075]_  : \new_[3896]_ ;
  assign \new_[3138]_  = \\u1_acs_addr_reg[21] ;
  assign \new_[3139]_  = ~\new_[3391]_  & (~\new_[7067]_  | ~\new_[9680]_ );
  assign \new_[3140]_  = ~\new_[3392]_  & (~\new_[7067]_  | ~\new_[10237]_ );
  assign \new_[3141]_  = ~\new_[3393]_  & (~\new_[7067]_  | ~\new_[9660]_ );
  assign \new_[3142]_  = ~\new_[3394]_  & (~\new_[7067]_  | ~\new_[9418]_ );
  assign \new_[3143]_  = ~\new_[3395]_  & (~\new_[7067]_  | ~\new_[10126]_ );
  assign \new_[3144]_  = ~\new_[3396]_  & (~\new_[7067]_  | ~\new_[10111]_ );
  assign \new_[3145]_  = \\u1_acs_addr_reg[18] ;
  assign \new_[3146]_  = ~\new_[3399]_  & (~\new_[7067]_  | ~\new_[9987]_ );
  assign \new_[3147]_  = ~\new_[3400]_  & (~\new_[7067]_  | ~\new_[9168]_ );
  assign \new_[3148]_  = ~\new_[3401]_  & (~\new_[7329]_  | ~\new_[9595]_ );
  assign \new_[3149]_  = ~\new_[3402]_  & (~\new_[7067]_  | ~\new_[9374]_ );
  assign \new_[3150]_  = ~\new_[3403]_  & (~\new_[7067]_  | ~\new_[9978]_ );
  assign \new_[3151]_  = ~\new_[3404]_  & (~\new_[7329]_  | ~\new_[9599]_ );
  assign \new_[3152]_  = ~\new_[3406]_  & (~\new_[7067]_  | ~\new_[10136]_ );
  assign \new_[3153]_  = ~\\u1_acs_addr_reg[4] ;
  assign \new_[3154]_  = \new_[5417]_  | \new_[3442]_ ;
  assign \new_[3155]_  = ~\new_[3665]_  | ~\new_[4774]_  | ~\new_[6206]_  | ~\new_[7331]_ ;
  assign \new_[3156]_  = ~\new_[3666]_  | ~\new_[4775]_  | ~\new_[6573]_  | ~\new_[7550]_ ;
  assign \new_[3157]_  = ~\new_[3667]_  | ~\new_[4777]_  | ~\new_[6580]_  | ~\new_[7552]_ ;
  assign \new_[3158]_  = ~\new_[4778]_  | ~\new_[3668]_  | ~\new_[6581]_  | ~\new_[7554]_ ;
  assign \new_[3159]_  = ~\new_[3669]_  | ~\new_[4784]_  | ~\new_[6585]_  | ~\new_[7561]_ ;
  assign \new_[3160]_  = ~\new_[3671]_  | ~\new_[4787]_  | ~\new_[6587]_  | ~\new_[7565]_ ;
  assign \new_[3161]_  = ~\new_[3672]_  | ~\new_[4788]_  | ~\new_[6590]_  | ~\new_[7566]_ ;
  assign \new_[3162]_  = ~\new_[3673]_  | ~\new_[4791]_  | ~\new_[6592]_  | ~\new_[7333]_ ;
  assign \new_[3163]_  = ~\new_[3674]_  | ~\new_[4534]_  | ~\new_[5988]_  | ~\new_[7236]_ ;
  assign \new_[3164]_  = ~\new_[3675]_  | ~\new_[4792]_  | ~\new_[6595]_  | ~\new_[7334]_ ;
  assign \new_[3165]_  = ~\new_[3677]_  | ~\new_[4797]_  | ~\new_[6616]_  | ~\new_[7342]_ ;
  assign \new_[3166]_  = ~\new_[3678]_  | ~\new_[6244]_  | ~\new_[4799]_  | ~\new_[7575]_ ;
  assign \new_[3167]_  = ~\\u1_acs_addr_reg[7] ;
  assign \new_[3168]_  = ~\new_[4451]_  | ~\new_[3650]_  | ~\new_[5420]_  | ~\new_[11460]_ ;
  assign \new_[3169]_  = \\u1_acs_addr_reg[13] ;
  assign \new_[3170]_  = ~\new_[3680]_  | ~\new_[4808]_  | ~\new_[6626]_  | ~\new_[7576]_ ;
  assign \new_[3171]_  = ~\new_[3682]_  | ~\new_[4541]_  | ~\new_[6619]_  | ~\new_[7568]_ ;
  assign \new_[3172]_  = ~\new_[3683]_  | ~\new_[4542]_  | ~\new_[6266]_  | ~\new_[7350]_ ;
  assign \new_[3173]_  = ~\new_[3684]_  | ~\new_[4543]_  | ~\new_[6631]_  | ~\new_[7349]_ ;
  assign \new_[3174]_  = \new_[3473]_  ? \new_[6075]_  : \new_[3962]_ ;
  assign \new_[3175]_  = ~\new_[3443]_  & (~\new_[12771]_  | ~\new_[9989]_ );
  assign \new_[3176]_  = \\u1_acs_addr_reg[16] ;
  assign \new_[3177]_  = \\u1_acs_addr_reg[14] ;
  assign \new_[3178]_  = ~\\u1_acs_addr_reg[11] ;
  assign \new_[3179]_  = \\u1_acs_addr_reg[17] ;
  assign \new_[3180]_  = \\u1_acs_addr_reg[12] ;
  assign \new_[3181]_  = ~\\u1_acs_addr_reg[8] ;
  assign \new_[3182]_  = \\u1_acs_addr_reg[0] ;
  assign \new_[3183]_  = \\u1_acs_addr_reg[1] ;
  assign \new_[3184]_  = ~\\u1_acs_addr_reg[3] ;
  assign \new_[3185]_  = ~\\u1_acs_addr_reg[5] ;
  assign \new_[3186]_  = ~\\u1_acs_addr_reg[6] ;
  assign \new_[3187]_  = ~\new_[3494]_  | ~\new_[5381]_  | ~\new_[4713]_ ;
  assign \new_[3188]_  = ~\new_[7286]_  | ~\new_[3459]_  | ~\new_[8018]_ ;
  assign \new_[3189]_  = ~\new_[4297]_  | ~\new_[3631]_  | ~\new_[5841]_  | ~\new_[6495]_ ;
  assign \new_[3190]_  = ~\new_[4301]_  | ~\new_[3634]_  | ~\new_[5842]_  | ~\new_[6496]_ ;
  assign \new_[3191]_  = ~\new_[4661]_  | ~\new_[3635]_  | ~\new_[5848]_  | ~\new_[6502]_ ;
  assign \new_[3192]_  = ~\new_[4663]_  | ~\new_[3636]_  | ~\new_[5849]_  | ~\new_[6503]_ ;
  assign \new_[3193]_  = ~\new_[4665]_  | ~\new_[3637]_  | ~\new_[5850]_  | ~\new_[6505]_ ;
  assign \new_[3194]_  = ~\new_[4666]_  | ~\new_[3638]_  | ~\new_[5851]_  | ~\new_[6697]_ ;
  assign \new_[3195]_  = ~\new_[4676]_  | ~\new_[3639]_  | ~\new_[5855]_  | ~\new_[6511]_ ;
  assign \new_[3196]_  = ~\new_[4680]_  | ~\new_[3640]_  | ~\new_[5856]_  | ~\new_[6514]_ ;
  assign \new_[3197]_  = ~\new_[4328]_  | ~\new_[3641]_  | ~\new_[5858]_  | ~\new_[6516]_ ;
  assign \new_[3198]_  = ~\new_[4333]_  | ~\new_[3642]_  | ~\new_[5469]_  | ~\new_[6704]_ ;
  assign \new_[3199]_  = ~\new_[4337]_  | ~\new_[3643]_  | ~\new_[5860]_  | ~\new_[6705]_ ;
  assign \new_[3200]_  = ~\new_[4319]_  | ~\new_[3644]_  | ~\new_[5969]_  | ~\new_[6517]_ ;
  assign \new_[3201]_  = ~\new_[4207]_  | ~\new_[3645]_  | ~\new_[5747]_  | ~\new_[6706]_ ;
  assign \new_[3202]_  = ~\new_[4235]_  | ~\new_[3646]_  | ~\new_[5373]_  | ~\new_[6707]_ ;
  assign \new_[3203]_  = ~\new_[4363]_  | ~\new_[3647]_  | ~\new_[6030]_  | ~\new_[6708]_ ;
  assign \new_[3204]_  = ~\new_[4394]_  | ~\new_[3648]_  | ~\new_[5822]_  | ~\new_[6709]_ ;
  assign \new_[3205]_  = ~\new_[4702]_  | ~\new_[3649]_  | ~\new_[5863]_  | ~\new_[6522]_ ;
  assign \new_[3206]_  = ~\new_[4454]_  | ~\new_[3651]_  | ~\new_[5867]_  | ~\new_[6524]_ ;
  assign \new_[3207]_  = ~\new_[4457]_  | ~\new_[3652]_  | ~\new_[5446]_  | ~\new_[6504]_ ;
  assign n1786 = ~\new_[3335]_  | (~\new_[5624]_  & ~\new_[4087]_ );
  assign \new_[3209]_  = ~\new_[4459]_  | ~\new_[3654]_  | ~\new_[5484]_  | ~\new_[6532]_ ;
  assign \new_[3210]_  = ~\new_[4463]_  | ~\new_[3657]_  | ~\new_[5873]_  | ~\new_[6712]_ ;
  assign \new_[3211]_  = ~\new_[4306]_  | ~\new_[3659]_  | ~\new_[5874]_  | ~\new_[6506]_ ;
  assign \new_[3212]_  = ~\new_[4724]_  | ~\new_[3660]_  | ~\new_[5875]_  | ~\new_[6528]_ ;
  assign \new_[3213]_  = ~\new_[4456]_  | ~\new_[3661]_  | ~\new_[5868]_  | ~\new_[6531]_ ;
  assign \new_[3214]_  = ~\new_[4468]_  | ~\new_[3663]_  | ~\new_[5466]_  | ~\new_[6703]_ ;
  assign \new_[3215]_  = ~\new_[4732]_  | ~\new_[3664]_  | ~\new_[5877]_  | ~\new_[6534]_ ;
  assign \new_[3216]_  = ~\new_[3471]_  & (~\new_[12534]_  | ~\new_[9594]_ );
  assign \new_[3217]_  = ~\new_[3933]_  | ~\new_[3467]_  | ~\new_[3588]_ ;
  assign \new_[3218]_  = ~\new_[3339]_  | (~\new_[12693]_  & ~\new_[9190]_ );
  assign \new_[3219]_  = ~\new_[3336]_  | ~\new_[7291]_ ;
  assign \new_[3220]_  = ~\new_[4317]_  | ~\new_[3341]_ ;
  assign \new_[3221]_  = (~\new_[6632]_  & ~\new_[3656]_  & ~\new_[7063]_ ) | (~\new_[3653]_  & ~\new_[6805]_  & ~\new_[8957]_ );
  assign \new_[3222]_  = ~\new_[4444]_  | ~\new_[3342]_ ;
  assign \new_[3223]_  = ~\new_[4452]_  | ~\new_[3343]_ ;
  assign \new_[3224]_  = ~\new_[4331]_  | ~\new_[3344]_ ;
  assign \new_[3225]_  = \\u1_acs_addr_reg[15] ;
  assign \new_[3226]_  = ~\new_[5715]_  & (~\new_[6986]_  | ~\new_[3503]_ );
  assign \new_[3227]_  = ~\new_[6037]_  | ~\new_[6713]_  | ~\new_[3347]_  | ~\new_[4464]_ ;
  assign \new_[3228]_  = ~\new_[5725]_  & (~\new_[6985]_  | ~\new_[3504]_ );
  assign \new_[3229]_  = ~\new_[5733]_  & (~\new_[6986]_  | ~\new_[3507]_ );
  assign \new_[3230]_  = ~\new_[5745]_  & (~\new_[6986]_  | ~\new_[3509]_ );
  assign \new_[3231]_  = ~\new_[10934]_  | ~\new_[9772]_  | ~\new_[3357]_  | ~\new_[12664]_ ;
  assign \new_[3232]_  = ~\new_[3474]_  | (~\new_[4097]_  & ~\new_[6075]_ );
  assign \new_[3233]_  = ~\new_[3558]_  & (~\new_[3655]_  | ~\new_[10177]_ );
  assign \new_[3234]_  = ~\new_[7156]_  & (~\new_[3953]_  | ~\new_[3700]_ );
  assign \new_[3235]_  = ~\new_[7156]_  & (~\new_[3955]_  | ~\new_[3701]_ );
  assign \new_[3236]_  = ~\new_[5048]_  | ~\new_[3990]_  | ~\new_[6187]_  | ~\new_[6598]_ ;
  assign \new_[3237]_  = ~\new_[7156]_  & (~\new_[3967]_  | ~\new_[3702]_ );
  assign \new_[3238]_  = ~\new_[3498]_  & (~\new_[9063]_  | ~\new_[12792]_ );
  assign \new_[3239]_  = ~\new_[4975]_  | ~\new_[3894]_  | ~\new_[3959]_  | ~\new_[5415]_ ;
  assign \new_[3240]_  = \new_[8093]_  | \new_[11833]_  | \new_[3556]_  | \new_[3704]_ ;
  assign \new_[3241]_  = \new_[8092]_  | \new_[11833]_  | \new_[3556]_  | \new_[3704]_ ;
  assign \new_[3242]_  = ~\new_[3508]_  & (~\new_[4840]_  | ~\new_[9374]_ );
  assign \new_[3243]_  = ~\new_[10139]_  | ~\new_[10231]_  | ~\new_[3717]_ ;
  assign \new_[3244]_  = ~\new_[3908]_  | ~\new_[3730]_  | ~\new_[3731]_ ;
  assign \new_[3245]_  = ~\new_[3718]_  | ~\new_[3577]_  | ~\new_[3733]_ ;
  assign \new_[3246]_  = ~\new_[3910]_  | ~\new_[3734]_  | ~\new_[3735]_ ;
  assign \new_[3247]_  = ~\new_[3719]_  | ~\new_[3736]_  | ~\new_[3737]_ ;
  assign \new_[3248]_  = ~\new_[3911]_  | ~\new_[3738]_  | ~\new_[3739]_ ;
  assign \new_[3249]_  = ~\new_[4781]_  | ~\new_[5978]_  | ~\new_[6154]_  | ~\new_[3685]_ ;
  assign \new_[3250]_  = ~\new_[3720]_  | ~\new_[3740]_  | ~\new_[3741]_ ;
  assign \new_[3251]_  = ~\new_[4947]_  & ~\new_[3537]_ ;
  assign \new_[3252]_  = ~\new_[3721]_  | ~\new_[3742]_  | ~\new_[3743]_ ;
  assign \new_[3253]_  = ~\new_[3912]_  | ~\new_[3745]_  | ~\new_[3746]_ ;
  assign \new_[3254]_  = ~\new_[3913]_  | ~\new_[3747]_  | ~\new_[3748]_ ;
  assign \new_[3255]_  = ~\new_[3916]_  | ~\new_[3754]_  | ~\new_[3755]_ ;
  assign \new_[3256]_  = ~\new_[3918]_  | ~\new_[3758]_  | ~\new_[3759]_ ;
  assign \new_[3257]_  = ~\new_[3919]_  | ~\new_[3764]_  | ~\new_[3765]_ ;
  assign \new_[3258]_  = ~\new_[3921]_  | ~\new_[3768]_  | ~\new_[3769]_ ;
  assign \new_[3259]_  = ~\new_[3928]_  | ~\new_[3777]_  | ~\new_[3778]_ ;
  assign \new_[3260]_  = ~\new_[3929]_  | ~\new_[3781]_  | ~\new_[3782]_ ;
  assign \new_[3261]_  = ~\new_[3722]_  | ~\new_[3582]_  | ~\new_[3785]_ ;
  assign \new_[3262]_  = ~\new_[3930]_  | ~\new_[3787]_  | ~\new_[3788]_ ;
  assign \new_[3263]_  = ~\new_[3931]_  | ~\new_[3583]_  | ~\new_[3793]_ ;
  assign \new_[3264]_  = ~\new_[3723]_  | ~\new_[3584]_  | ~\new_[3795]_ ;
  assign \new_[3265]_  = ~\new_[3934]_  | ~\new_[3585]_  | ~\new_[3796]_ ;
  assign \new_[3266]_  = ~\new_[3935]_  | ~\new_[3797]_  | ~\new_[3798]_ ;
  assign \new_[3267]_  = ~\new_[3559]_  & (~\new_[3716]_  | ~\new_[6075]_ );
  assign \new_[3268]_  = ~\new_[3539]_  & (~\new_[11864]_  | ~\new_[9418]_ );
  assign \new_[3269]_  = ~\new_[3541]_  & (~\new_[11864]_  | ~\new_[9958]_ );
  assign \new_[3270]_  = ~\new_[3542]_  & (~\new_[11864]_  | ~\new_[9326]_ );
  assign \new_[3271]_  = ~\new_[3544]_  & (~\new_[11864]_  | ~\new_[9479]_ );
  assign \new_[3272]_  = ~\new_[3546]_  & (~\new_[11864]_  | ~\new_[9618]_ );
  assign \new_[3273]_  = ~\new_[3547]_  & (~\new_[11864]_  | ~\new_[9682]_ );
  assign \new_[3274]_  = ~\new_[3548]_  & (~\new_[6679]_  | ~\new_[10097]_ );
  assign \new_[3275]_  = ~\new_[3549]_  & (~\new_[11864]_  | ~\new_[9675]_ );
  assign \new_[3276]_  = ~\new_[3550]_  & (~\new_[6679]_  | ~\new_[9709]_ );
  assign \new_[3277]_  = ~\new_[3551]_  & (~\new_[11864]_  | ~\new_[9109]_ );
  assign \new_[3278]_  = ~\new_[3552]_  & (~\new_[11864]_  | ~\new_[9567]_ );
  assign \new_[3279]_  = ~\new_[3553]_  & (~\new_[6679]_  | ~\new_[9707]_ );
  assign \new_[3280]_  = ~\new_[11956]_  & (~\new_[6679]_  | ~\new_[9684]_ );
  assign \new_[3281]_  = ~\new_[3554]_  & (~\new_[11864]_  | ~\new_[9389]_ );
  assign \new_[3282]_  = ~\new_[3555]_  & (~\new_[6679]_  | ~\new_[10137]_ );
  assign \new_[3283]_  = ~\new_[11922]_  & (~\new_[6679]_  | ~\new_[9665]_ );
  assign \new_[3284]_  = ~\new_[3557]_  & (~\new_[6097]_  | ~\new_[10200]_ );
  assign \new_[3285]_  = \new_[3893]_  ? \new_[6075]_  : \new_[3808]_ ;
  assign \new_[3286]_  = ~\new_[3514]_  & (~\new_[7067]_  | ~\new_[9401]_ );
  assign \new_[3287]_  = ~\new_[3515]_  & (~\new_[7067]_  | ~\new_[9661]_ );
  assign \new_[3288]_  = ~\new_[3516]_  & (~\new_[7329]_  | ~\new_[9963]_ );
  assign \new_[3289]_  = ~\new_[3517]_  & (~\new_[7329]_  | ~\new_[10128]_ );
  assign \new_[3290]_  = ~\new_[3518]_  & (~\new_[7329]_  | ~\new_[8805]_ );
  assign \new_[3291]_  = ~\new_[3519]_  & (~\new_[7067]_  | ~\new_[10011]_ );
  assign \new_[3292]_  = ~\new_[3520]_  & (~\new_[7067]_  | ~\new_[10263]_ );
  assign \new_[3293]_  = ~\new_[3521]_  & (~\new_[7329]_  | ~\new_[9995]_ );
  assign \new_[3294]_  = ~\new_[3532]_  & (~\new_[7329]_  | ~\new_[11772]_ );
  assign \new_[3295]_  = ~\new_[3522]_  & (~\new_[7067]_  | ~\new_[9845]_ );
  assign \new_[3296]_  = ~\new_[3523]_  & (~\new_[7329]_  | ~\new_[9641]_ );
  assign \new_[3297]_  = ~\new_[3524]_  & (~\new_[7329]_  | ~\new_[10287]_ );
  assign \new_[3298]_  = ~\new_[3526]_  & (~\new_[7067]_  | ~\new_[10019]_ );
  assign \new_[3299]_  = ~\new_[3527]_  & (~\new_[7067]_  | ~\new_[9657]_ );
  assign n1801 = \new_[3513]_  | \new_[5005]_ ;
  assign \new_[3301]_  = ~\new_[3528]_  & (~\new_[7329]_  | ~\new_[9710]_ );
  assign \new_[3302]_  = ~\new_[3529]_  & (~\new_[7067]_  | ~\new_[9604]_ );
  assign \new_[3303]_  = ~\new_[3530]_  & (~\new_[7067]_  | ~\new_[9407]_ );
  assign n1851 = \new_[3536]_  | \new_[5007]_ ;
  assign \new_[3305]_  = ~\new_[4976]_  | ~\new_[5088]_  | ~\new_[3725]_ ;
  assign n1806 = \new_[3571]_  | \new_[5006]_ ;
  assign \new_[3307]_  = ~\new_[3581]_  & (~\new_[8913]_  | ~\new_[4758]_ );
  assign \new_[3308]_  = ~\\u1_col_adr_reg[9] ;
  assign n1811 = \new_[10845]_  ? \new_[8800]_  : \new_[3609]_ ;
  assign n1821 = \new_[10968]_  ? \new_[8800]_  : \new_[3611]_ ;
  assign n1816 = \new_[10844]_  ? \new_[8800]_  : \new_[3610]_ ;
  assign n1826 = \new_[10916]_  ? \new_[8800]_  : \new_[3612]_ ;
  assign n1831 = \new_[10869]_  ? \new_[8800]_  : \new_[3613]_ ;
  assign n1791 = \new_[10852]_  ? \new_[8800]_  : \new_[3614]_ ;
  assign n1841 = \new_[10819]_  ? \new_[8800]_  : \new_[3615]_ ;
  assign n1836 = \new_[10833]_  ? \new_[8800]_  : \new_[3616]_ ;
  assign \new_[3317]_  = ~\new_[4772]_  & ~\new_[3586]_ ;
  assign \new_[3318]_  = ~\new_[3607]_  & ~\new_[5416]_ ;
  assign \new_[3319]_  = ~\new_[3587]_  & ~\new_[12075]_ ;
  assign \new_[3320]_  = ~\new_[4950]_  | ~\new_[3832]_  | ~\new_[7143]_  | ~\new_[6994]_ ;
  assign \new_[3321]_  = ~\new_[4957]_  | ~\new_[3838]_  | ~\new_[6117]_  | ~\new_[6995]_ ;
  assign \new_[3322]_  = ~\new_[4962]_  | ~\new_[3840]_  | ~\new_[6118]_  | ~\new_[6996]_ ;
  assign \new_[3323]_  = ~\new_[4979]_  | ~\new_[3857]_  | ~\new_[6115]_  | ~\new_[6993]_ ;
  assign n1796 = ~\new_[8848]_  | (~\new_[7156]_  & ~\new_[11275]_ );
  assign n1846 = ~\new_[9576]_  | (~\new_[3686]_  & ~\new_[10125]_ );
  assign \new_[3326]_  = ~\new_[3578]_  & ~\new_[9249]_ ;
  assign \new_[3327]_  = \new_[3597]_  | \new_[11277]_ ;
  assign \new_[3328]_  = ~\new_[3598]_  & ~\new_[11277]_ ;
  assign \new_[3329]_  = ~\new_[6119]_  | ~\new_[6526]_  | ~\new_[3497]_  | ~\new_[4461]_ ;
  assign \new_[3330]_  = ~\new_[6692]_  | ~\new_[6530]_  | ~\new_[3502]_  | ~\new_[4465]_ ;
  assign \new_[3331]_  = ~\new_[4299]_  | ~\new_[3475]_ ;
  assign \new_[3332]_  = ~\new_[4305]_  | ~\new_[3477]_ ;
  assign \new_[3333]_  = ~\new_[3512]_  & ~\new_[10826]_ ;
  assign n1916 = ~\new_[3472]_ ;
  assign \new_[3335]_  = \new_[3869]_  ? \new_[5624]_  : \new_[4087]_ ;
  assign \new_[3336]_  = (~\new_[5783]_  & ~\new_[11277]_  & ~\new_[10325]_ ) | (~\new_[10698]_  & ~\new_[4149]_  & ~\new_[10325]_ );
  assign \new_[3337]_  = ~\new_[3656]_  & ~\new_[8394]_ ;
  assign \new_[3338]_  = ~\new_[3658]_  & ~\new_[6805]_ ;
  assign \new_[3339]_  = ~\new_[9658]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3340]_  = \new_[5436]_  | \new_[3658]_ ;
  assign \new_[3341]_  = ~\new_[11492]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3342]_  = ~\new_[10496]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3343]_  = ~\new_[10250]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3344]_  = ~\new_[12755]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3345]_  = ~\new_[11473]_  | ~\new_[4709]_  | ~\new_[3901]_ ;
  assign \new_[3346]_  = ~\new_[3500]_ ;
  assign \new_[3347]_  = ~\new_[11367]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3348]_  = ~\new_[12578]_  | ~\new_[7176]_  | ~\new_[3894]_ ;
  assign \new_[3349]_  = ~\new_[11313]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3350]_  = ~\new_[11361]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3351]_  = ~\new_[10933]_  | ~\new_[3872]_  | ~\new_[10511]_ ;
  assign \new_[3352]_  = ~\new_[7956]_  | ~\new_[3703]_ ;
  assign \new_[3353]_  = ~\new_[4245]_  | ~\new_[10018]_  | ~\new_[3703]_  | ~\new_[7886]_ ;
  assign \new_[3354]_  = ~\new_[4171]_  | ~\new_[11263]_  | ~\new_[10001]_  | ~\new_[6289]_ ;
  assign \new_[3355]_  = ~\new_[3906]_  | ~\new_[3726]_  | ~\new_[3941]_ ;
  assign \new_[3356]_  = ~\new_[3907]_  | ~\new_[3727]_  | ~\new_[3945]_ ;
  assign \new_[3357]_  = ~\new_[3909]_  | ~\new_[3732]_  | ~\new_[3947]_ ;
  assign \new_[3358]_  = ~\new_[4475]_  | ~\new_[3744]_  | ~\new_[3950]_ ;
  assign \new_[3359]_  = ~\new_[3914]_  | ~\new_[3749]_  | ~\new_[3951]_ ;
  assign \new_[3360]_  = ~\new_[6608]_  | ~\new_[4623]_  | ~\new_[4156]_  | ~\new_[7338]_ ;
  assign \new_[3361]_  = ~\new_[11847]_  & (~\new_[11864]_  | ~\new_[9853]_ );
  assign \new_[3362]_  = ~\new_[6610]_  | ~\new_[4624]_  | ~\new_[4157]_  | ~\new_[7339]_ ;
  assign n1881 = ~\new_[3505]_ ;
  assign \new_[3364]_  = ~\new_[3689]_  & (~\new_[11864]_  | ~\new_[9582]_ );
  assign n1921 = ~\new_[3506]_ ;
  assign \new_[3366]_  = ~\new_[3922]_  | ~\new_[3770]_  | ~\new_[3958]_ ;
  assign \new_[3367]_  = ~\new_[4477]_  | ~\new_[3773]_  | ~\new_[3960]_ ;
  assign \new_[3368]_  = ~\new_[3925]_  | ~\new_[3774]_  | ~\new_[3961]_ ;
  assign \new_[3369]_  = ~\new_[3927]_  | ~\new_[3776]_  | ~\new_[3963]_ ;
  assign n1951 = ~\new_[3510]_ ;
  assign \new_[3371]_  = ~\new_[3699]_  & (~\new_[11864]_  | ~\new_[9379]_ );
  assign \new_[3372]_  = \new_[3895]_  ? \new_[6075]_  : \new_[3892]_ ;
  assign \new_[3373]_  = \new_[3897]_  ? \new_[6075]_  : \new_[3893]_ ;
  assign \new_[3374]_  = \new_[3898]_  ? \new_[6075]_  : \new_[3895]_ ;
  assign \new_[3375]_  = \new_[3899]_  ? \new_[6075]_  : \new_[3897]_ ;
  assign \new_[3376]_  = \new_[3900]_  ? \new_[6075]_  : \new_[3898]_ ;
  assign \new_[3377]_  = \new_[3902]_  ? \new_[6075]_  : \new_[3899]_ ;
  assign \new_[3378]_  = \new_[3903]_  ? \new_[6075]_  : \new_[3900]_ ;
  assign \new_[3379]_  = \new_[3904]_  ? \new_[6075]_  : \new_[3902]_ ;
  assign \new_[3380]_  = \new_[3896]_  ? \new_[6075]_  : \new_[3903]_ ;
  assign \new_[3381]_  = ~\new_[3690]_  & (~\new_[7329]_  | ~\new_[9383]_ );
  assign \new_[3382]_  = ~\new_[3691]_  & (~\new_[7067]_  | ~\new_[10031]_ );
  assign \new_[3383]_  = ~\new_[3692]_  & (~\new_[7067]_  | ~\new_[9930]_ );
  assign \new_[3384]_  = ~\new_[3693]_  & (~\new_[7067]_  | ~\new_[8977]_ );
  assign \new_[3385]_  = ~\new_[3694]_  & (~\new_[7067]_  | ~\new_[9682]_ );
  assign \new_[3386]_  = ~\new_[3695]_  & (~\new_[7067]_  | ~\new_[9107]_ );
  assign \new_[3387]_  = ~\new_[3696]_  & (~\new_[7067]_  | ~\new_[9391]_ );
  assign \new_[3388]_  = \\u5_ack_cnt_reg[3] ;
  assign \new_[3389]_  = ~\new_[3827]_  | ~\new_[5028]_  | ~\new_[4650]_ ;
  assign \new_[3390]_  = ~\new_[3828]_  | ~\new_[5029]_  | ~\new_[4302]_ ;
  assign \new_[3391]_  = ~\new_[3831]_  | ~\new_[5034]_  | ~\new_[4311]_ ;
  assign \new_[3392]_  = ~\new_[3833]_  | ~\new_[5535]_  | ~\new_[4674]_ ;
  assign \new_[3393]_  = ~\new_[3834]_  | ~\new_[5039]_  | ~\new_[4675]_ ;
  assign \new_[3394]_  = ~\new_[3835]_  | ~\new_[5041]_  | ~\new_[4678]_ ;
  assign \new_[3395]_  = ~\new_[3836]_  | ~\new_[5042]_  | ~\new_[4322]_ ;
  assign \new_[3396]_  = ~\new_[3837]_  | ~\new_[5044]_  | ~\new_[4681]_ ;
  assign \new_[3397]_  = ~\new_[3839]_  | ~\new_[5046]_  | ~\new_[4682]_ ;
  assign \new_[3398]_  = \\u5_ack_cnt_reg[1] ;
  assign \new_[3399]_  = ~\new_[3841]_  | ~\new_[5049]_  | ~\new_[4329]_ ;
  assign \new_[3400]_  = ~\new_[3849]_  | ~\new_[5065]_  | ~\new_[4684]_ ;
  assign \new_[3401]_  = ~\new_[3850]_  | ~\new_[5067]_  | ~\new_[4708]_ ;
  assign \new_[3402]_  = ~\new_[3851]_  | ~\new_[5070]_  | ~\new_[4455]_ ;
  assign \new_[3403]_  = ~\new_[3852]_  | ~\new_[5072]_  | ~\new_[4711]_ ;
  assign \new_[3404]_  = ~\new_[3858]_  | ~\new_[5570]_  | ~\new_[4720]_ ;
  assign \new_[3405]_  = ~\new_[3862]_  | ~\new_[5083]_  | ~\new_[4727]_ ;
  assign \new_[3406]_  = ~\new_[3864]_  | ~\new_[5045]_  | ~\new_[4733]_ ;
  assign \new_[3407]_  = ~\new_[3802]_  & (~\new_[9144]_  | ~\new_[5247]_ );
  assign \new_[3408]_  = ~\new_[3807]_  & (~\new_[9110]_  | ~\new_[5247]_ );
  assign \new_[3409]_  = ~\new_[3810]_  & (~\new_[9317]_  | ~\new_[5247]_ );
  assign \new_[3410]_  = ~\new_[3814]_  & (~\new_[9312]_  | ~\new_[5247]_ );
  assign \new_[3411]_  = ~\new_[3816]_  & (~\new_[9371]_  | ~\new_[5247]_ );
  assign \new_[3412]_  = ~\new_[3752]_  & (~\new_[9309]_  | ~\new_[5247]_ );
  assign \new_[3413]_  = ~\new_[3533]_ ;
  assign \new_[3414]_  = ~\new_[4022]_  | ~\new_[5403]_  | ~\new_[6686]_  | ~\new_[6267]_ ;
  assign \new_[3415]_  = ~\new_[6153]_  & ~\new_[3712]_ ;
  assign \new_[3416]_  = ~\new_[4054]_  | ~\new_[6579]_  | ~\new_[4776]_  | ~\new_[7551]_ ;
  assign \new_[3417]_  = ~\new_[4055]_  | ~\new_[4779]_  | ~\new_[6212]_  | ~\new_[7558]_ ;
  assign \new_[3418]_  = ~\new_[4056]_  | ~\new_[4782]_  | ~\new_[6584]_  | ~\new_[7578]_ ;
  assign \new_[3419]_  = ~\new_[4057]_  | ~\new_[4785]_  | ~\new_[6586]_  | ~\new_[7562]_ ;
  assign \new_[3420]_  = ~\new_[4058]_  | ~\new_[4786]_  | ~\new_[6724]_  | ~\new_[7563]_ ;
  assign \new_[3421]_  = ~\new_[4059]_  | ~\new_[4790]_  | ~\new_[6224]_  | ~\new_[7347]_ ;
  assign \new_[3422]_  = ~\new_[4060]_  | ~\new_[4793]_  | ~\new_[6232]_  | ~\new_[7335]_ ;
  assign \new_[3423]_  = ~\new_[3761]_  & (~\new_[9320]_  | ~\new_[4758]_ );
  assign \new_[3424]_  = ~\new_[3763]_  & (~\new_[8918]_  | ~\new_[4758]_ );
  assign \new_[3425]_  = ~\new_[3713]_  & ~\new_[7874]_ ;
  assign \new_[3426]_  = ~\new_[6157]_  & ~\new_[3714]_ ;
  assign \new_[3427]_  = ~\new_[6158]_  & ~\new_[3715]_ ;
  assign \new_[3428]_  = ~\new_[4064]_  | ~\new_[5998]_  | ~\new_[4536]_  | ~\new_[7240]_ ;
  assign \new_[3429]_  = ~\new_[4065]_  | ~\new_[4804]_  | ~\new_[6237]_  | ~\new_[7553]_ ;
  assign \new_[3430]_  = ~\new_[3780]_  & (~\new_[9878]_  | ~\new_[5247]_ );
  assign \new_[3431]_  = ~\new_[4706]_  | ~\new_[7175]_  | ~\new_[3812]_  | ~\new_[7197]_ ;
  assign \new_[3432]_  = ~\new_[3784]_  & (~\new_[9633]_  | ~\new_[4758]_ );
  assign \new_[3433]_  = ~\new_[3790]_  & (~\new_[9748]_  | ~\new_[4758]_ );
  assign \new_[3434]_  = ~\new_[4066]_  | ~\new_[11520]_  | ~\new_[6628]_  | ~\new_[7585]_ ;
  assign \new_[3435]_  = ~\new_[3792]_  & (~\new_[9319]_  | ~\new_[4758]_ );
  assign \new_[3436]_  = ~\new_[4655]_  | ~\new_[4024]_  | ~\new_[5629]_  | ~\new_[6634]_ ;
  assign \new_[3437]_  = ~\new_[4658]_  | ~\new_[4028]_  | ~\new_[5630]_  | ~\new_[7006]_ ;
  assign \new_[3438]_  = u4_rfr_req_reg;
  assign \new_[3439]_  = \\u5_ack_cnt_reg[0] ;
  assign \new_[3440]_  = \\u5_ack_cnt_reg[2] ;
  assign \new_[3441]_  = ~\new_[6017]_  | ~\new_[5394]_  | ~\new_[3676]_  | ~\new_[7637]_ ;
  assign \new_[3442]_  = ~\new_[3822]_  & ~\new_[12689]_ ;
  assign \new_[3443]_  = ~\new_[5432]_  & (~\new_[3866]_  | ~\new_[7657]_ );
  assign n1926 = ~\new_[3561]_ ;
  assign n1861 = ~\new_[3562]_ ;
  assign n1931 = ~\new_[3563]_ ;
  assign n1866 = ~\new_[3564]_ ;
  assign n1936 = ~\new_[3565]_ ;
  assign n1941 = ~\new_[3566]_ ;
  assign n1946 = ~\new_[3567]_ ;
  assign n1856 = ~\new_[3568]_ ;
  assign n1901 = ~\new_[3569]_ ;
  assign n1871 = (~\new_[5635]_  & ~\new_[10759]_ ) | (~\new_[3949]_  & ~\new_[10826]_ );
  assign n1891 = ~\new_[3572]_ ;
  assign n1906 = ~\new_[3573]_ ;
  assign n1911 = ~\new_[3574]_ ;
  assign n1896 = ~\new_[3575]_ ;
  assign n1876 = ~\new_[3576]_ ;
  assign \new_[3459]_  = ~\new_[11275]_  & ~\new_[7777]_ ;
  assign \new_[3460]_  = ~\new_[12567]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3461]_  = ~\new_[10411]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3462]_  = ~\new_[9674]_  | ~\new_[12527]_  | ~\new_[10529]_ ;
  assign \new_[3463]_  = ~\new_[11337]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3464]_  = ~\new_[11323]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3465]_  = ~\new_[11328]_  | ~\new_[12527]_  | ~\new_[10529]_ ;
  assign \new_[3466]_  = ~\new_[9946]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3467]_  = ~\new_[10960]_  | ~\new_[11275]_  | ~\new_[10529]_ ;
  assign \new_[3468]_  = ~\new_[4652]_  & (~\new_[3871]_  | ~\new_[8920]_ );
  assign n1886 = ~\new_[3589]_ ;
  assign \new_[3470]_  = ~\new_[3820]_  & (~\new_[6327]_  | ~\new_[12093]_ );
  assign \new_[3471]_  = ~\new_[6638]_  | ~\new_[6533]_  | ~\new_[3662]_  | ~\new_[4335]_ ;
  assign \new_[3472]_  = ~\new_[4998]_  & (~\new_[4096]_  | ~\new_[10759]_ );
  assign \new_[3473]_  = ~\new_[5913]_  | ~\new_[3874]_  | ~\new_[4483]_ ;
  assign \new_[3474]_  = ~\new_[3873]_  | ~\new_[6075]_ ;
  assign \new_[3475]_  = ~\new_[10291]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3476]_  = ~\new_[10827]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3477]_  = ~\new_[10922]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3478]_  = ~\new_[11355]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3479]_  = ~\new_[11348]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3480]_  = ~\new_[9997]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3481]_  = \new_[11944]_  | \new_[6639]_ ;
  assign \new_[3482]_  = \new_[11944]_  & \new_[5358]_ ;
  assign \new_[3483]_  = ~\new_[11343]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3484]_  = ~\new_[10808]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3485]_  = ~\new_[11340]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3486]_  = ~\new_[10243]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3487]_  = ~\new_[10938]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3488]_  = ~\new_[11735]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3489]_  = ~\new_[11316]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3490]_  = ~\new_[10108]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3491]_  = ~\new_[12453]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3492]_  = ~\new_[9926]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3493]_  = ~\new_[10950]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3494]_  = ~\new_[11337]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3495]_  = ~\new_[11323]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3496]_  = ~\new_[3704]_  | ~\new_[5701]_ ;
  assign \new_[3497]_  = ~\new_[10955]_  | ~\new_[3871]_  | ~\new_[10511]_ ;
  assign \new_[3498]_  = ~\new_[4292]_  | ~\new_[4545]_  | ~\new_[5017]_  | ~\new_[7549]_ ;
  assign \new_[3499]_  = ~\new_[11367]_  | ~\new_[4240]_  | ~\new_[7628]_ ;
  assign \new_[3500]_  = ~\new_[3877]_  | ~\new_[12736]_ ;
  assign \new_[3501]_  = ~\new_[5881]_  | ~\new_[4505]_  | ~\new_[11434]_  | ~\new_[5766]_ ;
  assign \new_[3502]_  = ~\new_[11526]_  | ~\new_[3870]_  | ~\new_[10511]_ ;
  assign \new_[3503]_  = ~\new_[4473]_  | ~\new_[3942]_  | ~\new_[4161]_ ;
  assign \new_[3504]_  = ~\new_[4476]_  | ~\new_[3956]_  | ~\new_[4164]_ ;
  assign \new_[3505]_  = ~\new_[5011]_  & (~\new_[4159]_  | ~\new_[10759]_ );
  assign \new_[3506]_  = ~\new_[5015]_  & (~\new_[4160]_  | ~\new_[10759]_ );
  assign \new_[3507]_  = ~\new_[4478]_  | ~\new_[3964]_  | ~\new_[4165]_ ;
  assign \new_[3508]_  = ~\new_[4225]_  | ~\new_[4801]_  | ~\new_[7442]_  | ~\new_[7579]_ ;
  assign \new_[3509]_  = ~\new_[4493]_  | ~\new_[3968]_  | ~\new_[4169]_ ;
  assign \new_[3510]_  = ~\new_[5001]_  & (~\new_[4154]_  | ~\new_[10759]_ );
  assign n1956 = ~\new_[3688]_ ;
  assign \new_[3512]_  = ~\new_[3875]_  & (~\new_[11271]_  | ~\new_[11114]_ );
  assign \new_[3513]_  = ~\new_[3937]_  & ~\new_[10826]_ ;
  assign \new_[3514]_  = ~\new_[4023]_  | ~\new_[5516]_  | ~\new_[4653]_ ;
  assign \new_[3515]_  = ~\new_[4025]_  | ~\new_[5520]_  | ~\new_[4307]_ ;
  assign \new_[3516]_  = ~\new_[4026]_  | ~\new_[5031]_  | ~\new_[4309]_ ;
  assign \new_[3517]_  = ~\new_[4029]_  | ~\new_[5523]_  | ~\new_[4660]_ ;
  assign \new_[3518]_  = ~\new_[4032]_  | ~\new_[5032]_  | ~\new_[4662]_ ;
  assign \new_[3519]_  = ~\new_[4033]_  | ~\new_[5033]_  | ~\new_[4664]_ ;
  assign \new_[3520]_  = ~\new_[4034]_  | ~\new_[5035]_  | ~\new_[4314]_ ;
  assign \new_[3521]_  = ~\new_[4035]_  | ~\new_[5037]_  | ~\new_[4668]_ ;
  assign \new_[3522]_  = ~\new_[4037]_  | ~\new_[5532]_  | ~\new_[4316]_ ;
  assign \new_[3523]_  = ~\new_[4038]_  | ~\new_[5043]_  | ~\new_[4324]_ ;
  assign \new_[3524]_  = ~\new_[4039]_  | ~\new_[5541]_  | ~\new_[4325]_ ;
  assign \new_[3525]_  = ~\new_[4752]_  & ~\new_[3998]_ ;
  assign \new_[3526]_  = ~\new_[4041]_  | ~\new_[5064]_  | ~\new_[4445]_ ;
  assign \new_[3527]_  = ~\new_[4043]_  | ~\new_[5066]_  | ~\new_[4447]_ ;
  assign \new_[3528]_  = ~\new_[4044]_  | ~\new_[5074]_  | ~\new_[4336]_ ;
  assign \new_[3529]_  = ~\new_[4045]_  | ~\new_[5571]_  | ~\new_[4723]_ ;
  assign \new_[3530]_  = ~\new_[4046]_  | ~\new_[5085]_  | ~\new_[4470]_ ;
  assign \new_[3531]_  = ~\new_[4007]_  & (~\new_[9820]_  | ~\new_[4758]_ );
  assign \new_[3532]_  = ~\new_[4036]_  | ~\new_[5038]_  | ~\new_[4672]_ ;
  assign \new_[3533]_  = ~\new_[12769]_  & ~\new_[3890]_ ;
  assign \new_[3534]_  = ~\new_[3944]_  & (~\new_[9629]_  | ~\new_[5247]_ );
  assign \new_[3535]_  = ~\new_[3946]_  & (~\new_[9628]_  | ~\new_[4758]_ );
  assign \new_[3536]_  = ~\new_[3948]_  & ~\new_[10826]_ ;
  assign \new_[3537]_  = ~\new_[7325]_  | ~\new_[4273]_  | ~\new_[7332]_  | ~\new_[4783]_ ;
  assign \new_[3538]_  = ~\new_[3952]_  & (~\new_[9630]_  | ~\new_[5248]_ );
  assign \new_[3539]_  = ~\new_[4218]_  | ~\new_[4789]_  | ~\new_[6223]_  | ~\new_[7580]_ ;
  assign \new_[3540]_  = ~\new_[3954]_  & (~\new_[9635]_  | ~\new_[5248]_ );
  assign \new_[3541]_  = ~\new_[4219]_  | ~\new_[4794]_  | ~\new_[6600]_  | ~\new_[7336]_ ;
  assign \new_[3542]_  = ~\new_[4220]_  | ~\new_[6605]_  | ~\new_[4795]_  | ~\new_[7337]_ ;
  assign \new_[3543]_  = ~\new_[3957]_  & (~\new_[8807]_  | ~\new_[4758]_ );
  assign \new_[3544]_  = ~\new_[4221]_  | ~\new_[4796]_  | ~\new_[6574]_  | ~\new_[7340]_ ;
  assign \new_[3545]_  = ~\new_[6155]_  & ~\new_[3891]_ ;
  assign \new_[3546]_  = ~\new_[4223]_  | ~\new_[4798]_  | ~\new_[6243]_  | ~\new_[7574]_ ;
  assign \new_[3547]_  = ~\new_[4224]_  | ~\new_[4800]_  | ~\new_[6245]_  | ~\new_[7567]_ ;
  assign \new_[3548]_  = ~\new_[4226]_  | ~\new_[4803]_  | ~\new_[6205]_  | ~\new_[7557]_ ;
  assign \new_[3549]_  = ~\new_[4227]_  | ~\new_[4805]_  | ~\new_[6250]_  | ~\new_[7570]_ ;
  assign \new_[3550]_  = ~\new_[4228]_  | ~\new_[4806]_  | ~\new_[6251]_  | ~\new_[7581]_ ;
  assign \new_[3551]_  = ~\new_[4229]_  | ~\new_[4807]_  | ~\new_[6254]_  | ~\new_[7582]_ ;
  assign \new_[3552]_  = ~\new_[4230]_  | ~\new_[4537]_  | ~\new_[6257]_  | ~\new_[7583]_ ;
  assign \new_[3553]_  = ~\new_[4232]_  | ~\new_[4538]_  | ~\new_[6258]_  | ~\new_[7584]_ ;
  assign \new_[3554]_  = ~\new_[4233]_  | ~\new_[4539]_  | ~\new_[6602]_  | ~\new_[7346]_ ;
  assign \new_[3555]_  = ~\new_[4234]_  | ~\new_[4540]_  | ~\new_[6593]_  | ~\new_[7348]_ ;
  assign \new_[3556]_  = \new_[9060]_  | \new_[3905]_ ;
  assign \new_[3557]_  = ~\new_[6283]_  | ~\new_[3926]_  | ~\new_[5711]_ ;
  assign \new_[3558]_  = ~\new_[3939]_  & (~\new_[5826]_  | ~\new_[6215]_ );
  assign \new_[3559]_  = ~\new_[5626]_  & ~\new_[3962]_ ;
  assign \new_[3560]_  = ~\new_[7246]_  & ~\new_[4012]_ ;
  assign \new_[3561]_  = ~\new_[4735]_  & (~\new_[4079]_  | ~\new_[10759]_ );
  assign \new_[3562]_  = ~\new_[4996]_  & (~\new_[4080]_  | ~\new_[10759]_ );
  assign \new_[3563]_  = ~\new_[4736]_  & (~\new_[4081]_  | ~\new_[10691]_ );
  assign \new_[3564]_  = ~\new_[5009]_  & (~\new_[4082]_  | ~\new_[10759]_ );
  assign \new_[3565]_  = ~\new_[5010]_  & (~\new_[4083]_  | ~\new_[10691]_ );
  assign \new_[3566]_  = ~\new_[5012]_  & (~\new_[4084]_  | ~\new_[10759]_ );
  assign \new_[3567]_  = ~\new_[5013]_  & (~\new_[4085]_  | ~\new_[10759]_ );
  assign \new_[3568]_  = ~\new_[5016]_  & (~\new_[4086]_  | ~\new_[10759]_ );
  assign \new_[3569]_  = ~\new_[5000]_  & (~\new_[4158]_  | ~\new_[10759]_ );
  assign \new_[3570]_  = ~\new_[3966]_  & (~\new_[12775]_  | ~\new_[10137]_ );
  assign \new_[3571]_  = ~\new_[3830]_  & ~\new_[10826]_ ;
  assign \new_[3572]_  = ~\new_[4999]_  & (~\new_[4172]_  | ~\new_[10759]_ );
  assign \new_[3573]_  = ~\new_[4997]_  & (~\new_[4173]_  | ~\new_[10759]_ );
  assign \new_[3574]_  = ~\new_[5003]_  & (~\new_[4175]_  | ~\new_[10759]_ );
  assign \new_[3575]_  = ~\new_[5002]_  & (~\new_[4070]_  | ~\new_[10759]_ );
  assign \new_[3576]_  = ~\new_[5004]_  & (~\new_[4078]_  | ~\new_[10759]_ );
  assign \new_[3577]_  = ~\new_[10928]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3578]_  = (~\new_[9879]_  | ~\new_[4020]_ ) & (~\new_[6671]_  | ~\new_[10086]_ );
  assign \new_[3579]_  = \new_[5391]_  | \new_[11272]_ ;
  assign \new_[3580]_  = \new_[5401]_  | \new_[11272]_ ;
  assign \new_[3581]_  = ~\new_[11274]_  & (~\new_[5834]_  | ~\new_[5983]_ );
  assign \new_[3582]_  = ~\new_[11356]_  | ~\new_[11275]_  | ~\new_[10441]_ ;
  assign \new_[3583]_  = ~\new_[11526]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3584]_  = ~\new_[10509]_  | ~\new_[12527]_  | ~\new_[10441]_ ;
  assign \new_[3585]_  = ~\new_[10526]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3586]_  = (~\new_[12684]_  & ~\new_[7655]_  & ~\new_[7523]_ ) | (~\new_[4576]_  & ~\new_[7523]_  & ~\new_[10485]_ );
  assign \new_[3587]_  = ~\new_[4657]_  | ~\new_[3829]_ ;
  assign \new_[3588]_  = \new_[3823]_  | \new_[11276]_ ;
  assign \new_[3589]_  = ~\new_[5014]_  & (~\new_[4042]_  | ~\new_[10691]_ );
  assign \new_[3590]_  = \new_[4332]_  & \new_[3842]_ ;
  assign \new_[3591]_  = \new_[4334]_  & \new_[3843]_ ;
  assign \new_[3592]_  = \new_[4310]_  & \new_[3844]_ ;
  assign \new_[3593]_  = \new_[4507]_  & \new_[3845]_ ;
  assign \new_[3594]_  = \new_[4348]_  & \new_[3846]_ ;
  assign \new_[3595]_  = \new_[4367]_  & \new_[3847]_ ;
  assign \new_[3596]_  = ~\new_[5617]_  | ~\new_[6285]_  | ~\new_[3848]_  | ~\new_[6204]_ ;
  assign \new_[3597]_  = (~\new_[4030]_  | ~\new_[7286]_ ) & (~\new_[11306]_  | ~\new_[7517]_ );
  assign \new_[3598]_  = (~\new_[4027]_  | ~\new_[7116]_ ) & (~\new_[11306]_  | ~\new_[7768]_ );
  assign \new_[3599]_  = \new_[4458]_  & \new_[3853]_ ;
  assign \new_[3600]_  = \new_[4714]_  & \new_[3854]_ ;
  assign \new_[3601]_  = \new_[4462]_  & \new_[3855]_ ;
  assign \new_[3602]_  = \new_[4718]_  & \new_[3856]_ ;
  assign \new_[3603]_  = \new_[4721]_  & \new_[3859]_ ;
  assign \new_[3604]_  = \new_[4725]_  & \new_[3860]_ ;
  assign \new_[3605]_  = \new_[4318]_  & \new_[3861]_ ;
  assign \new_[3606]_  = \new_[4467]_  & \new_[3863]_ ;
  assign \new_[3607]_  = ~\new_[12693]_  & (~\new_[4099]_  | ~\new_[9178]_ );
  assign \new_[3608]_  = ~\new_[6202]_  | ~\new_[6286]_  | ~\new_[4238]_  | ~\new_[4098]_ ;
  assign \new_[3609]_  = \new_[10817]_  ? \new_[4255]_  : \new_[3043]_ ;
  assign \new_[3610]_  = \new_[10908]_  ? \new_[4255]_  : \new_[3044]_ ;
  assign \new_[3611]_  = \new_[10885]_  ? \new_[4255]_  : \new_[3045]_ ;
  assign \new_[3612]_  = \new_[10878]_  ? \new_[4255]_  : \new_[3046]_ ;
  assign \new_[3613]_  = \new_[10901]_  ? \new_[4255]_  : \new_[3047]_ ;
  assign \new_[3614]_  = \new_[10825]_  ? \new_[4255]_  : \new_[2971]_ ;
  assign \new_[3615]_  = \new_[10828]_  ? \new_[4255]_  : \new_[3049]_ ;
  assign \new_[3616]_  = \new_[10896]_  ? \new_[4255]_  : \new_[3048]_ ;
  assign \new_[3617]_  = \new_[2833]_  ? \new_[4262]_  : \new_[8893]_ ;
  assign \new_[3618]_  = \new_[2839]_  ? \new_[4262]_  : \new_[8973]_ ;
  assign \new_[3619]_  = \new_[2840]_  ? \new_[4262]_  : \new_[8966]_ ;
  assign \new_[3620]_  = \new_[2829]_  ? \new_[4262]_  : \new_[8971]_ ;
  assign \new_[3621]_  = \new_[2841]_  ? \new_[4262]_  : \new_[8969]_ ;
  assign \new_[3622]_  = \new_[2842]_  ? \new_[4262]_  : \new_[8940]_ ;
  assign \new_[3623]_  = \new_[2843]_  ? \new_[4262]_  : \new_[8951]_ ;
  assign \new_[3624]_  = \new_[2830]_  ? \new_[4262]_  : \new_[8939]_ ;
  assign \new_[3625]_  = \new_[2845]_  ? \new_[4262]_  : \new_[11227]_ ;
  assign \new_[3626]_  = \new_[2768]_  ? \new_[4262]_  : \new_[11059]_ ;
  assign n1976 = ~\new_[4090]_  & ~\new_[8230]_ ;
  assign n1966 = ~\new_[4091]_  & ~\new_[8230]_ ;
  assign n1981 = ~\new_[4088]_  & ~\new_[8230]_ ;
  assign n1961 = ~\new_[4089]_  & ~\new_[8230]_ ;
  assign \new_[3631]_  = ~\new_[10634]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3632]_  = ~\new_[4300]_  | ~\new_[8018]_  | ~\new_[4298]_ ;
  assign \new_[3633]_  = ~\new_[4300]_  | ~\new_[8018]_  | ~\new_[4648]_ ;
  assign \new_[3634]_  = ~\new_[10838]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3635]_  = ~\new_[11576]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3636]_  = ~\new_[9379]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3637]_  = ~\new_[11332]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3638]_  = ~\new_[10177]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3639]_  = ~\new_[11320]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3640]_  = ~\new_[9913]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3641]_  = ~\new_[9785]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3642]_  = ~\new_[10802]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3643]_  = ~\new_[12093]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3644]_  = ~n5021 | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3645]_  = ~\new_[12567]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3646]_  = ~\new_[10164]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3647]_  = ~\new_[11363]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3648]_  = ~\new_[10411]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3649]_  = ~\new_[12554]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3650]_  = ~\new_[12054]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3651]_  = ~\new_[12598]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3652]_  = ~\new_[12610]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3653]_  = \new_[4144]_  | \new_[6632]_ ;
  assign \new_[3654]_  = ~\new_[11353]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3655]_  = ~\new_[4149]_  & ~\new_[10549]_ ;
  assign \new_[3656]_  = \new_[4144]_  | \new_[7263]_ ;
  assign \new_[3657]_  = ~\new_[11328]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3658]_  = \new_[4144]_  | \new_[8740]_ ;
  assign \new_[3659]_  = ~\new_[11310]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3660]_  = ~\new_[10419]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3661]_  = ~\new_[9946]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3662]_  = ~\new_[12044]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3663]_  = ~\new_[10960]_  | ~\new_[4095]_  | ~\new_[10511]_ ;
  assign \new_[3664]_  = ~\new_[10526]_  | ~\new_[4093]_  | ~\new_[10511]_ ;
  assign \new_[3665]_  = ~\new_[4100]_  & (~\new_[7685]_  | ~\new_[10102]_ );
  assign \new_[3666]_  = ~\new_[4102]_  & (~\new_[12308]_  | ~\new_[9584]_ );
  assign \new_[3667]_  = ~\new_[4104]_  & (~\new_[7591]_  | ~\new_[9588]_ );
  assign \new_[3668]_  = ~\new_[4105]_  & (~\new_[12308]_  | ~\new_[9933]_ );
  assign \new_[3669]_  = ~\new_[4106]_  & (~\new_[7591]_  | ~\new_[9842]_ );
  assign \new_[3670]_  = ~\new_[4108]_  & (~\new_[12307]_  | ~\new_[9975]_ );
  assign \new_[3671]_  = ~\new_[4109]_  & (~\new_[7685]_  | ~\new_[9489]_ );
  assign \new_[3672]_  = ~\new_[4110]_  & (~\new_[7685]_  | ~\new_[9593]_ );
  assign \new_[3673]_  = ~\new_[4112]_  & (~\new_[7591]_  | ~\new_[9601]_ );
  assign \new_[3674]_  = ~\new_[4113]_  & (~\new_[12307]_  | ~\new_[10064]_ );
  assign \new_[3675]_  = ~\new_[4114]_  & (~\new_[7591]_  | ~\new_[9585]_ );
  assign \new_[3676]_  = ~\new_[4115]_  & (~\new_[12307]_  | ~\new_[9937]_ );
  assign \new_[3677]_  = ~\new_[4123]_  & (~\new_[7591]_  | ~\new_[9614]_ );
  assign \new_[3678]_  = ~\new_[4124]_  & (~\new_[7685]_  | ~\new_[9589]_ );
  assign \new_[3679]_  = ~\new_[4128]_  & (~\new_[7591]_  | ~\new_[9613]_ );
  assign \new_[3680]_  = ~\new_[4131]_  & (~\new_[7591]_  | ~\new_[9408]_ );
  assign \new_[3681]_  = ~\new_[4134]_  & (~\new_[12307]_  | ~\new_[10047]_ );
  assign \new_[3682]_  = ~\new_[4137]_  & (~\new_[12308]_  | ~\new_[9393]_ );
  assign \new_[3683]_  = ~\new_[4138]_  & (~\new_[7685]_  | ~\new_[9874]_ );
  assign \new_[3684]_  = ~\new_[4140]_  & (~\new_[7591]_  | ~\new_[9863]_ );
  assign \new_[3685]_  = ~\new_[4142]_  & (~\new_[12492]_  | ~\new_[9960]_ );
  assign \new_[3686]_  = (~\new_[4449]_  | ~\wb_addr_i[10] ) & (~\new_[5181]_  | ~\wb_addr_i[10] );
  assign \new_[3687]_  = ~\new_[4148]_  | (~\new_[6036]_  & ~\new_[5639]_ );
  assign \new_[3688]_  = ~\new_[4155]_  & (~\new_[10125]_  | ~\new_[11059]_ );
  assign \new_[3689]_  = ~\new_[7304]_  | ~\new_[4549]_  | ~\new_[5806]_  | ~\new_[4625]_ ;
  assign \new_[3690]_  = ~\new_[4193]_  | ~\new_[5918]_  | ~\new_[4928]_ ;
  assign \new_[3691]_  = ~\new_[4194]_  | ~\new_[5920]_  | ~\new_[4932]_ ;
  assign \new_[3692]_  = ~\new_[4196]_  | ~\new_[5925]_  | ~\new_[4954]_ ;
  assign \new_[3693]_  = ~\new_[4200]_  | ~\new_[5932]_  | ~\new_[4692]_ ;
  assign \new_[3694]_  = ~\new_[4201]_  | ~\new_[5934]_  | ~\new_[4704]_ ;
  assign \new_[3695]_  = ~\new_[4202]_  | ~\new_[5936]_  | ~\new_[4669]_ ;
  assign \new_[3696]_  = ~\new_[4203]_  | ~\new_[5937]_  | ~\new_[4707]_ ;
  assign \new_[3697]_  = \\u3_byte0_reg[1] ;
  assign \new_[3698]_  = ~\new_[7324]_  | ~\new_[4608]_  | ~\new_[7548]_  | ~\new_[4773]_ ;
  assign \new_[3699]_  = ~\new_[7526]_  | ~\new_[4614]_  | ~\new_[7559]_  | ~\new_[4780]_ ;
  assign \new_[3700]_  = ~\new_[4162]_  & (~\new_[9626]_  | ~\new_[5247]_ );
  assign \new_[3701]_  = ~\new_[4163]_  & (~\new_[9877]_  | ~\new_[5247]_ );
  assign \new_[3702]_  = ~\new_[4168]_  & (~\new_[9625]_  | ~\new_[5247]_ );
  assign \new_[3703]_  = ~\new_[3878]_ ;
  assign \new_[3704]_  = ~\new_[3879]_ ;
  assign \new_[3705]_  = \\u3_byte0_reg[0] ;
  assign \new_[3706]_  = \\u3_byte0_reg[2] ;
  assign \new_[3707]_  = \\u3_byte0_reg[4] ;
  assign \new_[3708]_  = \\u3_byte0_reg[3] ;
  assign \new_[3709]_  = \\u3_byte0_reg[5] ;
  assign \new_[3710]_  = \\u3_byte0_reg[6] ;
  assign \new_[3711]_  = \\u3_byte0_reg[7] ;
  assign \new_[3712]_  = ~\new_[6011]_  | ~\new_[5785]_  | ~\new_[4053]_  | ~\new_[7636]_ ;
  assign \new_[3713]_  = ~\new_[6018]_  | ~\new_[5795]_  | ~\new_[4061]_  | ~\new_[7640]_ ;
  assign \new_[3714]_  = ~\new_[6021]_  | ~\new_[5801]_  | ~\new_[4062]_  | ~\new_[7639]_ ;
  assign \new_[3715]_  = ~\new_[6023]_  | ~\new_[5790]_  | ~\new_[4063]_  | ~\new_[7642]_ ;
  assign \new_[3716]_  = ~\new_[3904]_ ;
  assign \new_[3717]_  = ~\new_[4166]_  & ~\new_[11045]_ ;
  assign \new_[3718]_  = ~\new_[10928]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3719]_  = ~\new_[11576]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3720]_  = ~\new_[11332]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3721]_  = ~\new_[11343]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3722]_  = ~\new_[11356]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3723]_  = ~\new_[10509]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign n1971 = ~\new_[10124]_  & (~\new_[4522]_  | ~\new_[10934]_ );
  assign \new_[3725]_  = \new_[4052]_  | \new_[12683]_ ;
  assign \new_[3726]_  = ~\new_[10291]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3727]_  = ~\new_[10922]_  | ~\new_[11274]_  | ~\new_[10441]_ ;
  assign \new_[3728]_  = ~\new_[10743]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3729]_  = ~\new_[4553]_  & ~\new_[4068]_ ;
  assign \new_[3730]_  = ~\new_[11355]_  | ~\new_[11272]_  | ~\new_[10441]_ ;
  assign \new_[3731]_  = \new_[5385]_  | \new_[11277]_ ;
  assign \new_[3732]_  = ~\new_[11348]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3733]_  = \new_[4890]_  | \new_[11272]_ ;
  assign \new_[3734]_  = ~\new_[9997]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3735]_  = \new_[5386]_  | \new_[11277]_ ;
  assign \new_[3736]_  = ~\new_[11576]_  | ~\new_[11275]_  | ~\new_[10441]_ ;
  assign \new_[3737]_  = \new_[5387]_  | \new_[11277]_ ;
  assign \new_[3738]_  = ~\new_[10962]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3739]_  = \new_[5388]_  | \new_[11272]_ ;
  assign \new_[3740]_  = ~\new_[11332]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3741]_  = \new_[4891]_  | \new_[11276]_ ;
  assign \new_[3742]_  = ~\new_[11343]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3743]_  = \new_[5389]_  | \new_[11276]_ ;
  assign \new_[3744]_  = ~\new_[10808]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3745]_  = ~\new_[10818]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3746]_  = \new_[5390]_  | \new_[11275]_ ;
  assign \new_[3747]_  = ~\new_[11340]_  | ~\new_[11275]_  | ~\new_[10441]_ ;
  assign \new_[3748]_  = \new_[4892]_  | \new_[11272]_ ;
  assign \new_[3749]_  = ~\new_[11492]_  | ~\new_[11274]_  | ~\new_[10441]_ ;
  assign \new_[3750]_  = ~\new_[10243]_  | ~\new_[11276]_  | ~\new_[10441]_ ;
  assign \new_[3751]_  = ~\new_[11320]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3752]_  = ~\new_[11277]_  & (~\new_[5828]_  | ~\new_[6222]_ );
  assign \new_[3753]_  = ~\new_[10938]_  | ~\new_[11275]_  | ~\new_[10529]_ ;
  assign \new_[3754]_  = ~\new_[11735]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3755]_  = \new_[5392]_  | \new_[11277]_ ;
  assign \new_[3756]_  = ~\new_[9913]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3757]_  = ~\new_[11316]_  | ~\new_[11276]_  | ~\new_[10441]_ ;
  assign \new_[3758]_  = ~\new_[10108]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3759]_  = \new_[5395]_  | \new_[11275]_ ;
  assign \new_[3760]_  = ~\new_[10802]_  | ~\new_[11276]_  | ~\new_[10529]_ ;
  assign \new_[3761]_  = ~\new_[11276]_  & (~\new_[5830]_  | ~\new_[6604]_ );
  assign \new_[3762]_  = ~\new_[12093]_  | ~\new_[11275]_  | ~\new_[10441]_ ;
  assign \new_[3763]_  = ~\new_[11275]_  & (~\new_[5831]_  | ~\new_[6236]_ );
  assign \new_[3764]_  = ~n5021 | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3765]_  = \new_[5396]_  | \new_[11276]_ ;
  assign \new_[3766]_  = \new_[5397]_  | \new_[11274]_ ;
  assign \new_[3767]_  = ~\new_[10164]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3768]_  = ~\new_[11363]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3769]_  = \new_[5399]_  | \new_[11276]_ ;
  assign \new_[3770]_  = ~\new_[10496]_  | ~\new_[11274]_  | ~\new_[10441]_ ;
  assign \new_[3771]_  = ~\new_[9926]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3772]_  = ~\new_[9903]_  | ~\new_[11275]_  | ~\new_[10529]_ ;
  assign \new_[3773]_  = ~\new_[12554]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3774]_  = ~\new_[10250]_  | ~\new_[11276]_  | ~\new_[10441]_ ;
  assign \new_[3775]_  = ~\new_[4812]_  & ~\new_[4021]_ ;
  assign \new_[3776]_  = ~\new_[12755]_  | ~\new_[11276]_  | ~\new_[10441]_ ;
  assign \new_[3777]_  = ~\new_[12610]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3778]_  = \new_[5402]_  | \new_[11276]_ ;
  assign \new_[3779]_  = ~\new_[11353]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3780]_  = ~\new_[11272]_  & (~\new_[5835]_  | ~\new_[6006]_ );
  assign \new_[3781]_  = ~\new_[10955]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3782]_  = \new_[5404]_  | \new_[11276]_ ;
  assign \new_[3783]_  = ~\new_[11367]_  | ~\new_[11276]_  | ~\new_[10529]_ ;
  assign \new_[3784]_  = ~\new_[11277]_  & (~\new_[5836]_  | ~\new_[6253]_ );
  assign \new_[3785]_  = \new_[4894]_  | \new_[11277]_ ;
  assign \new_[3786]_  = ~\new_[11310]_  | ~\new_[11274]_  | ~\new_[10529]_ ;
  assign \new_[3787]_  = ~\new_[10419]_  | ~\new_[12527]_  | ~\new_[10441]_ ;
  assign \new_[3788]_  = \new_[5405]_  | \new_[11276]_ ;
  assign \new_[3789]_  = ~\new_[11313]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3790]_  = ~\new_[11277]_  & (~\new_[5837]_  | ~\new_[6230]_ );
  assign \new_[3791]_  = ~\new_[11361]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3792]_  = ~\new_[11276]_  & (~\new_[5838]_  | ~\new_[6260]_ );
  assign \new_[3793]_  = \new_[5406]_  | \new_[11276]_ ;
  assign \new_[3794]_  = \new_[5407]_  | \new_[11276]_ ;
  assign \new_[3795]_  = \new_[4896]_  | \new_[11276]_ ;
  assign \new_[3796]_  = \new_[5408]_  | \new_[11272]_ ;
  assign \new_[3797]_  = ~\new_[10919]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3798]_  = \new_[4897]_  | \new_[11277]_ ;
  assign \new_[3799]_  = ~\new_[6101]_  & ~\new_[4021]_ ;
  assign \new_[3800]_  = ~\new_[11275]_  & (~\new_[7005]_  | ~\new_[7299]_ );
  assign \new_[3801]_  = ~\new_[10743]_  | ~\new_[12239]_  | ~\new_[11885]_ ;
  assign \new_[3802]_  = ~\new_[11277]_  & (~\new_[5987]_  | ~\new_[5419]_ );
  assign \new_[3803]_  = ~\new_[11298]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3804]_  = ~\new_[12089]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3805]_  = \new_[4338]_  & \new_[4040]_ ;
  assign \new_[3806]_  = ~\new_[10411]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3807]_  = ~\new_[12527]_  & (~\new_[5995]_  | ~\new_[5400]_ );
  assign \new_[3808]_  = ~\new_[4753]_  | ~\new_[5913]_  | ~\new_[4097]_  | ~\new_[4483]_ ;
  assign \new_[3809]_  = ~\new_[12554]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3810]_  = ~\new_[11274]_  & (~\new_[5996]_  | ~\new_[6381]_ );
  assign \new_[3811]_  = ~\new_[11323]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3812]_  = ~\new_[4551]_  & ~\new_[4092]_ ;
  assign \new_[3813]_  = ~\new_[11328]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3814]_  = ~\new_[11274]_  & (~\new_[6002]_  | ~\new_[6103]_ );
  assign \new_[3815]_  = ~\new_[11356]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3816]_  = ~\new_[11274]_  & (~\new_[6007]_  | ~\new_[6104]_ );
  assign \new_[3817]_  = ~\new_[10933]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3818]_  = ~\new_[9946]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3819]_  = ~\new_[12044]_  | ~\new_[12239]_  | ~\new_[4294]_ ;
  assign \new_[3820]_  = ~\new_[12093]_  & (~\new_[6328]_  | ~\new_[4206]_ );
  assign \new_[3821]_  = ~\new_[10509]_  | ~\new_[12239]_  | ~\new_[11885]_ ;
  assign \new_[3822]_  = ~\new_[10063]_  & (~\new_[4244]_  | ~\new_[10511]_ );
  assign \new_[3823]_  = (~\new_[11305]_  | ~\new_[7310]_ ) & (~\new_[4584]_  | ~\new_[7116]_ );
  assign \new_[3824]_  = \new_[4262]_  | \new_[11068]_ ;
  assign \new_[3825]_  = \new_[4262]_  | \new_[11133]_ ;
  assign \new_[3826]_  = ~\new_[11885]_  | ~\new_[10818]_ ;
  assign \new_[3827]_  = ~\new_[9998]_  | ~\new_[4240]_  | ~\new_[7628]_ ;
  assign \new_[3828]_  = ~\new_[12273]_  | ~\new_[4241]_  | ~\new_[7630]_ ;
  assign \new_[3829]_  = ~\new_[10928]_  | ~\new_[11495]_  | ~\new_[10511]_ ;
  assign \new_[3830]_  = ~\new_[4204]_  & (~\new_[11271]_  | ~\new_[3042]_ );
  assign \new_[3831]_  = ~\new_[10177]_  | ~\new_[4240]_  | ~\new_[7522]_ ;
  assign \new_[3832]_  = ~\new_[10818]_  | ~\new_[11495]_  | ~\new_[10511]_ ;
  assign \new_[3833]_  = ~\new_[10243]_  | ~\new_[4240]_  | ~\new_[7522]_ ;
  assign \new_[3834]_  = ~\new_[11320]_  | ~\new_[4240]_  | ~\new_[7522]_ ;
  assign \new_[3835]_  = ~\new_[10938]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3836]_  = ~\new_[11735]_  | ~\new_[4241]_  | ~\new_[7630]_ ;
  assign \new_[3837]_  = ~\new_[11298]_  | ~\new_[4240]_  | ~\new_[7628]_ ;
  assign \new_[3838]_  = ~\new_[11298]_  | ~\new_[11495]_  | ~\new_[10511]_ ;
  assign \new_[3839]_  = ~\new_[12089]_  | ~\new_[4240]_  | ~\new_[7628]_ ;
  assign \new_[3840]_  = ~\new_[12089]_  | ~\new_[11495]_  | ~\new_[10511]_ ;
  assign \new_[3841]_  = ~\new_[10108]_  | ~\new_[4241]_  | ~\new_[7630]_ ;
  assign \new_[3842]_  = ~\new_[10802]_  | ~\new_[4240]_  | ~\new_[7664]_ ;
  assign \new_[3843]_  = ~\new_[12093]_  | ~\new_[4240]_  | ~\new_[7664]_ ;
  assign \new_[3844]_  = ~\new_[12567]_  | ~\new_[4240]_  | ~\new_[7629]_ ;
  assign \new_[3845]_  = ~\new_[10164]_  | ~\new_[4240]_  | ~\new_[7664]_ ;
  assign \new_[3846]_  = ~\new_[11363]_  | ~\new_[4240]_  | ~\new_[7629]_ ;
  assign \new_[3847]_  = ~\new_[10411]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3848]_  = \new_[5467]_  & \new_[4238]_ ;
  assign \new_[3849]_  = ~\new_[9903]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3850]_  = ~\new_[12598]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3851]_  = ~\new_[12610]_  | ~\new_[4241]_  | ~\new_[7630]_ ;
  assign \new_[3852]_  = ~\new_[11337]_  | ~\new_[4240]_  | ~\new_[7664]_ ;
  assign \new_[3853]_  = ~\new_[11353]_  | ~\new_[4240]_  | ~\new_[7663]_ ;
  assign \new_[3854]_  = ~\new_[10955]_  | ~\new_[4240]_  | ~\new_[7663]_ ;
  assign \new_[3855]_  = ~\new_[11328]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3856]_  = ~\new_[11356]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3857]_  = ~\new_[11356]_  | ~\new_[11495]_  | ~\new_[10511]_ ;
  assign \new_[3858]_  = ~\new_[10419]_  | ~\new_[4240]_  | ~\new_[7522]_ ;
  assign \new_[3859]_  = ~\new_[11310]_  | ~\new_[4240]_  | ~\new_[7663]_ ;
  assign \new_[3860]_  = ~\new_[11361]_  | ~\new_[4240]_  | ~\new_[7663]_ ;
  assign \new_[3861]_  = ~\new_[10933]_  | ~\new_[4240]_  | ~\new_[7631]_ ;
  assign \new_[3862]_  = ~\new_[12044]_  | ~\new_[4240]_  | ~\new_[7628]_ ;
  assign \new_[3863]_  = ~\new_[10960]_  | ~\new_[4240]_  | ~\new_[7663]_ ;
  assign \new_[3864]_  = ~\new_[10634]_  | ~\new_[4240]_  | ~\new_[7628]_ ;
  assign \new_[3865]_  = ~\new_[4291]_  & (~\new_[11500]_  | ~\new_[10051]_ );
  assign \new_[3866]_  = ~\new_[4243]_  | ~\new_[7708]_ ;
  assign \new_[3867]_  = (~\new_[5619]_  & ~\new_[7292]_  & ~\new_[7069]_ ) | (~\new_[4654]_  & ~\new_[6786]_  & ~\new_[7662]_ );
  assign \new_[3868]_  = \new_[4648]_  | \new_[4300]_ ;
  assign \new_[3869]_  = \new_[4450]_  | \new_[2927]_ ;
  assign \new_[3870]_  = ~\new_[4094]_ ;
  assign \new_[3871]_  = ~\new_[4094]_ ;
  assign \new_[3872]_  = ~\new_[4094]_ ;
  assign \new_[3873]_  = ~\new_[4098]_ ;
  assign \new_[3874]_  = ~\new_[4141]_ ;
  assign \new_[3875]_  = ~\new_[4995]_  & ~\new_[4508]_ ;
  assign \new_[3876]_  = \\u3_byte2_reg[7] ;
  assign \new_[3877]_  = ~\new_[4144]_ ;
  assign \new_[3878]_  = ~\new_[12340]_ ;
  assign \new_[3879]_  = \new_[12340]_ ;
  assign n5451 = u5_lmr_ack_reg;
  assign \new_[3881]_  = \\u5_ir_cnt_reg[1] ;
  assign \new_[3882]_  = ~\\u5_ir_cnt_reg[2] ;
  assign \mc_addr_pad_o[14]  = \\u7_mc_addr_reg[14] ;
  assign \new_[3884]_  = \\u3_byte2_reg[0] ;
  assign \new_[3885]_  = \\u3_byte2_reg[1] ;
  assign \new_[3886]_  = \\u3_byte2_reg[2] ;
  assign \new_[3887]_  = \\u3_byte2_reg[4] ;
  assign \new_[3888]_  = \\u3_byte2_reg[5] ;
  assign \new_[3889]_  = \\u3_byte2_reg[6] ;
  assign \new_[3890]_  = ~\new_[4150]_ ;
  assign \new_[3891]_  = ~\new_[6019]_  | ~\new_[5797]_  | ~\new_[4222]_  | ~\new_[7641]_ ;
  assign \new_[3892]_  = ~\new_[4738]_  | ~\new_[4825]_  | ~\new_[4481]_ ;
  assign \new_[3893]_  = ~\new_[4739]_  | ~\new_[4826]_  | ~\new_[4482]_ ;
  assign \new_[3894]_  = ~\new_[6363]_  & ~\new_[4178]_ ;
  assign \new_[3895]_  = ~\new_[4741]_  | ~\new_[4827]_  | ~\new_[4484]_ ;
  assign \new_[3896]_  = ~\new_[4743]_  | ~\new_[4828]_  | ~\new_[4485]_ ;
  assign \new_[3897]_  = ~\new_[4745]_  | ~\new_[4829]_  | ~\new_[4479]_ ;
  assign \new_[3898]_  = ~\new_[4746]_  | ~\new_[4830]_  | ~\new_[4487]_ ;
  assign \new_[3899]_  = ~\new_[4747]_  | ~\new_[4831]_  | ~\new_[4492]_ ;
  assign \new_[3900]_  = ~\new_[4748]_  | ~\new_[4832]_  | ~\new_[4488]_ ;
  assign \new_[3901]_  = ~\new_[6975]_  | ~\new_[4525]_ ;
  assign \new_[3902]_  = ~\new_[4751]_  | ~\new_[4833]_  | ~\new_[4489]_ ;
  assign \new_[3903]_  = ~\new_[4749]_  | ~\new_[4834]_  | ~\new_[4490]_ ;
  assign \new_[3904]_  = ~\new_[4750]_  | ~\new_[4835]_  | ~\new_[4491]_ ;
  assign \new_[3905]_  = ~\new_[11467]_  | ~\new_[4245]_ ;
  assign \new_[3906]_  = ~\new_[10291]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3907]_  = ~\new_[10922]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3908]_  = ~\new_[11355]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3909]_  = ~\new_[11348]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3910]_  = ~\new_[9997]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3911]_  = ~\new_[10962]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3912]_  = ~\new_[10818]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3913]_  = ~\new_[11340]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3914]_  = ~\new_[11492]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3915]_  = ~\new_[10938]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3916]_  = ~\new_[11735]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3917]_  = \\u3_byte2_reg[3] ;
  assign \new_[3918]_  = ~\new_[10108]_  | ~\new_[5247]_  | ~\new_[11045]_ ;
  assign \new_[3919]_  = ~n5021 | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3920]_  = ~\new_[12567]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3921]_  = ~\new_[11363]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3922]_  = ~\new_[10496]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3923]_  = ~\new_[10902]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3924]_  = ~\new_[9903]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3925]_  = ~\new_[10250]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3926]_  = ~\new_[4524]_  | ~\new_[10278]_ ;
  assign \new_[3927]_  = ~\new_[12755]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[3928]_  = ~\new_[12610]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3929]_  = ~\new_[10955]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3930]_  = ~\new_[10419]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3931]_  = ~\new_[11526]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3932]_  = ~\new_[9946]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3933]_  = ~\new_[10960]_  | ~\new_[4758]_  | ~\new_[11045]_ ;
  assign \new_[3934]_  = ~\new_[10526]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \new_[3935]_  = ~\new_[10919]_  | ~\new_[5247]_  | ~\new_[11233]_ ;
  assign \mc_addr_pad_o[13]  = \\u7_mc_addr_reg[13] ;
  assign \new_[3937]_  = ~\new_[4513]_  & (~\new_[11271]_  | ~\new_[3041]_ );
  assign \new_[3938]_  = ~\new_[4520]_  & (~\new_[12492]_  | ~\new_[9864]_ );
  assign \new_[3939]_  = \new_[11277]_  | \new_[10549]_ ;
  assign \new_[3940]_  = ~\new_[11277]_  & (~\new_[6978]_  | ~\new_[7169]_ );
  assign \new_[3941]_  = \new_[5781]_  | \new_[12527]_ ;
  assign \new_[3942]_  = ~\new_[9998]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3943]_  = ~\new_[12273]_  | ~\new_[11275]_  | ~\new_[10529]_ ;
  assign \new_[3944]_  = ~\new_[12527]_  & (~\new_[5824]_  | ~\new_[6572]_ );
  assign \new_[3945]_  = \new_[5784]_  | \new_[11277]_ ;
  assign \new_[3946]_  = ~\new_[11277]_  & (~\new_[5825]_  | ~\new_[6577]_ );
  assign \new_[3947]_  = \new_[4889]_  | \new_[11276]_ ;
  assign \new_[3948]_  = ~\new_[4529]_  & (~\new_[11271]_  | ~\new_[11102]_ );
  assign \new_[3949]_  = ~\new_[4530]_  & (~\new_[4995]_  | ~\new_[3138]_ );
  assign \new_[3950]_  = \new_[5787]_  | \new_[11277]_ ;
  assign \new_[3951]_  = \new_[5788]_  | \new_[11276]_ ;
  assign \new_[3952]_  = ~\new_[11275]_  & (~\new_[5827]_  | ~\new_[6589]_ );
  assign \new_[3953]_  = ~\new_[11298]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3954]_  = ~\new_[11275]_  & (~\new_[5829]_  | ~\new_[6596]_ );
  assign \new_[3955]_  = ~\new_[12089]_  | ~\new_[11277]_  | ~\new_[10529]_ ;
  assign \new_[3956]_  = ~\new_[9785]_  | ~\new_[12527]_  | ~\new_[10529]_ ;
  assign \new_[3957]_  = ~\new_[11272]_  & (~\new_[5832]_  | ~\new_[6612]_ );
  assign \new_[3958]_  = \new_[5796]_  | \new_[11277]_ ;
  assign \new_[3959]_  = ~\new_[5329]_  & ~\new_[4239]_ ;
  assign \new_[3960]_  = \new_[5798]_  | \new_[11277]_ ;
  assign \new_[3961]_  = \new_[5799]_  | \new_[11277]_ ;
  assign \new_[3962]_  = ~\new_[4744]_  | ~\new_[4486]_  | ~\new_[4639]_ ;
  assign \new_[3963]_  = \new_[5803]_  | \new_[11277]_ ;
  assign \new_[3964]_  = ~\new_[12598]_  | ~\new_[12527]_  | ~\new_[10529]_ ;
  assign \new_[3965]_  = ~\new_[10933]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[3966]_  = ~\new_[5432]_  & (~\new_[4578]_  | ~\new_[7319]_ );
  assign \new_[3967]_  = ~\new_[12044]_  | ~\new_[11275]_  | ~\new_[10529]_ ;
  assign \new_[3968]_  = ~\new_[10634]_  | ~\new_[12527]_  | ~\new_[10529]_ ;
  assign \new_[3969]_  = ~\new_[10827]_  | ~\new_[5638]_  | ~\new_[4645]_ ;
  assign \new_[3970]_  = ~\new_[10922]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[3971]_  = ~\new_[11355]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3972]_  = ~\new_[11348]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[3973]_  = ~\new_[10928]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3974]_  = ~\new_[9997]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3975]_  = ~\new_[11576]_  | ~\new_[5638]_  | ~\new_[4646]_ ;
  assign \new_[3976]_  = ~\new_[10962]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[3977]_  = ~\new_[11332]_  | ~\new_[5638]_  | ~\new_[4645]_ ;
  assign \new_[3978]_  = ~\new_[10177]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3979]_  = ~\new_[11343]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3980]_  = ~\new_[10808]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3981]_  = ~\new_[11340]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3982]_  = ~\new_[11492]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[3983]_  = ~\new_[10243]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[3984]_  = ~\new_[11320]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[3985]_  = ~\new_[10938]_  | ~\new_[5638]_  | ~\new_[4926]_ ;
  assign \new_[3986]_  = ~\new_[11735]_  | ~\new_[5242]_  | ~\new_[4926]_ ;
  assign \new_[3987]_  = ~\new_[9913]_  | ~\new_[5638]_  | ~\new_[4645]_ ;
  assign \new_[3988]_  = ~\new_[11316]_  | ~\new_[5638]_  | ~\new_[4645]_ ;
  assign \new_[3989]_  = ~\new_[9785]_  | ~\new_[12239]_  | ~\new_[4926]_ ;
  assign \new_[3990]_  = \new_[4963]_  & \new_[4197]_ ;
  assign \new_[3991]_  = ~\new_[10108]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[3992]_  = ~\new_[10802]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[3993]_  = ~\new_[12093]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[3994]_  = ~n5021 | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3995]_  = ~\new_[12567]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[3996]_  = ~\new_[10164]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[3997]_  = ~\new_[11363]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[3998]_  = (~\new_[12684]_  & ~\new_[7654]_  & ~\new_[7772]_ ) | (~\new_[4576]_  & ~\new_[7521]_  & ~\new_[12454]_ );
  assign \new_[3999]_  = ~\new_[12453]_  | ~\new_[12239]_  | ~\new_[4926]_ ;
  assign \new_[4000]_  = ~\new_[10496]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[4001]_  = ~\new_[9926]_  | ~\new_[5638]_  | ~\new_[4645]_ ;
  assign \new_[4002]_  = ~\new_[9903]_  | ~\new_[5242]_  | ~\new_[4926]_ ;
  assign \new_[4003]_  = ~\new_[10250]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[4004]_  = ~\new_[12598]_  | ~\new_[12239]_  | ~\new_[4926]_ ;
  assign \new_[4005]_  = ~\new_[12610]_  | ~\new_[5638]_  | ~\new_[4646]_ ;
  assign \new_[4006]_  = ~\new_[11353]_  | ~\new_[5638]_  | ~\new_[4646]_ ;
  assign \new_[4007]_  = ~\new_[11272]_  & (~\new_[6247]_  | ~\new_[6383]_ );
  assign \new_[4008]_  = ~\new_[10955]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[4009]_  = ~\new_[11367]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[4010]_  = ~\new_[10419]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[4011]_  = ~\new_[11310]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[4012]_  = (~\new_[12683]_  & ~\new_[7661]_  & ~\new_[7772]_ ) | (~\new_[11478]_  & ~\new_[7772]_  & ~\new_[11314]_ );
  assign \new_[4013]_  = ~\new_[11313]_  | ~\new_[5242]_  | ~\new_[4646]_ ;
  assign \new_[4014]_  = ~\new_[11361]_  | ~\new_[5638]_  | ~\new_[4646]_ ;
  assign \new_[4015]_  = ~\new_[11526]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[4016]_  = ~\new_[10960]_  | ~\new_[5638]_  | ~\new_[4646]_ ;
  assign \new_[4017]_  = ~\new_[10526]_  | ~\new_[5638]_  | ~\new_[11884]_ ;
  assign \new_[4018]_  = ~\new_[10919]_  | ~\new_[12239]_  | ~\new_[11884]_ ;
  assign \new_[4019]_  = ~\new_[10634]_  | ~\new_[12239]_  | ~\new_[4926]_ ;
  assign \new_[4020]_  = \new_[4844]_  ? \new_[11355]_  : \new_[6671]_ ;
  assign \new_[4021]_  = ~\new_[6457]_  | ~\new_[4706]_  | ~\new_[7197]_ ;
  assign \new_[4022]_  = ~\new_[6164]_  & ~\new_[4573]_ ;
  assign \new_[4023]_  = ~\new_[10827]_  | ~\new_[11477]_  | ~\new_[7522]_ ;
  assign \new_[4024]_  = ~\new_[11355]_  | ~\new_[4577]_  | ~\new_[7630]_ ;
  assign \new_[4025]_  = ~\new_[11348]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4026]_  = ~\new_[10928]_  | ~\new_[11477]_  | ~\new_[7629]_ ;
  assign \new_[4027]_  = ~\new_[4562]_  & (~\new_[7994]_  | ~\new_[10348]_ );
  assign \new_[4028]_  = ~\new_[10963]_  | ~\new_[4577]_  | ~\new_[7630]_ ;
  assign \new_[4029]_  = ~\new_[11576]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4030]_  = ~\new_[4561]_  & (~\new_[7994]_  | ~\new_[10724]_ );
  assign \new_[4031]_  = ~\new_[4586]_  & (~\new_[7077]_  | ~\new_[9607]_ );
  assign \new_[4032]_  = ~\new_[9647]_  | ~\new_[4577]_  | ~\new_[7630]_ ;
  assign \new_[4033]_  = ~\new_[11332]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4034]_  = ~\new_[11343]_  | ~\new_[11477]_  | ~\new_[7629]_ ;
  assign \new_[4035]_  = ~\new_[10808]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4036]_  = ~\new_[10818]_  | ~\new_[4577]_  | ~\new_[7630]_ ;
  assign \new_[4037]_  = ~\new_[11340]_  | ~\new_[11477]_  | ~\new_[7522]_ ;
  assign \new_[4038]_  = ~\new_[9913]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4039]_  = ~\new_[11316]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4040]_  = ~n5021 | ~\new_[11477]_  | ~\new_[7664]_ ;
  assign \new_[4041]_  = ~\new_[10902]_  | ~\new_[11477]_  | ~\new_[7629]_ ;
  assign \new_[4042]_  = \new_[8366]_  ? \new_[11269]_  : \new_[11131]_ ;
  assign \new_[4043]_  = ~\new_[12554]_  | ~\new_[11477]_  | ~\new_[7629]_ ;
  assign \new_[4044]_  = ~\new_[11323]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4045]_  = ~\new_[11526]_  | ~\new_[4575]_  | ~\new_[7522]_ ;
  assign \new_[4046]_  = ~\new_[10526]_  | ~\new_[11477]_  | ~\new_[7522]_ ;
  assign \new_[4047]_  = ~\new_[4581]_  & (~\new_[11864]_  | ~\new_[9979]_ );
  assign \new_[4048]_  = ~\new_[4640]_  & (~\new_[11500]_  | ~\new_[10130]_ );
  assign \new_[4049]_  = ~\new_[4641]_  & (~\new_[11500]_  | ~\new_[9967]_ );
  assign \new_[4050]_  = ~\new_[4642]_  & (~\new_[11500]_  | ~\new_[9871]_ );
  assign \new_[4051]_  = ~\new_[4737]_  & (~\new_[5865]_  | ~\new_[9707]_ );
  assign \new_[4052]_  = ~\new_[7322]_  & (~\new_[11415]_  | ~\new_[4992]_ );
  assign \new_[4053]_  = ~\new_[4611]_  & (~\new_[12308]_  | ~\new_[9938]_ );
  assign \new_[4054]_  = ~\new_[4612]_  & (~\new_[7685]_  | ~\new_[9587]_ );
  assign \new_[4055]_  = ~\new_[4613]_  & (~\new_[7685]_  | ~\new_[9592]_ );
  assign \new_[4056]_  = ~\new_[4615]_  & (~\new_[12308]_  | ~\new_[9612]_ );
  assign \new_[4057]_  = ~\new_[4617]_  & (~\new_[7591]_  | ~\new_[9678]_ );
  assign \new_[4058]_  = ~\new_[4619]_  & (~\new_[12307]_  | ~\new_[10040]_ );
  assign \new_[4059]_  = ~\new_[4620]_  & (~\new_[7685]_  | ~\new_[9615]_ );
  assign \new_[4060]_  = ~\new_[4622]_  & (~\new_[7685]_  | ~\new_[9602]_ );
  assign \new_[4061]_  = ~\new_[4627]_  & (~\new_[12308]_  | ~\new_[10084]_ );
  assign \new_[4062]_  = ~\new_[4631]_  & (~\new_[12308]_  | ~\new_[11515]_ );
  assign \new_[4063]_  = ~\new_[4633]_  & (~\new_[12308]_  | ~\new_[9844]_ );
  assign \new_[4064]_  = ~\new_[4635]_  & (~\new_[7591]_  | ~\new_[9824]_ );
  assign \new_[4065]_  = ~\new_[4636]_  & (~\new_[7685]_  | ~\new_[9609]_ );
  assign \new_[4066]_  = ~\new_[4616]_  & (~\new_[7591]_  | ~\new_[11521]_ );
  assign \new_[4067]_  = ~\new_[4728]_  & (~\new_[6811]_  | ~\new_[6683]_ );
  assign \new_[4068]_  = (~\new_[5619]_  & ~\new_[6805]_  & ~\new_[6786]_ ) | (~\new_[6578]_  & ~\new_[5619]_  & ~\new_[7263]_ );
  assign n1991 = \new_[10845]_  ? \new_[4927]_  : \new_[3705]_ ;
  assign \new_[4070]_  = \new_[6527]_  ? \new_[11269]_  : \new_[3176]_ ;
  assign n1986 = \new_[10844]_  ? \new_[4927]_  : \new_[3697]_ ;
  assign n1996 = \new_[10968]_  ? \new_[4927]_  : \new_[3706]_ ;
  assign n2006 = \new_[10916]_  ? \new_[4927]_  : \new_[3708]_ ;
  assign n2001 = \new_[10869]_  ? \new_[4927]_  : \new_[3707]_ ;
  assign n2011 = \new_[10852]_  ? \new_[4927]_  : \new_[3709]_ ;
  assign n2016 = \new_[10819]_  ? \new_[4927]_  : \new_[3710]_ ;
  assign n2021 = \new_[10833]_  ? \new_[4927]_  : \new_[3711]_ ;
  assign \new_[4078]_  = \new_[5823]_  ? \new_[11269]_  : \new_[3145]_ ;
  assign \new_[4079]_  = \new_[10354]_  ? \new_[11269]_  : \new_[3182]_ ;
  assign \new_[4080]_  = \new_[8481]_  ? \new_[4995]_  : \new_[11026]_ ;
  assign \new_[4081]_  = \new_[10232]_  ? \new_[11269]_  : \new_[3183]_ ;
  assign \new_[4082]_  = \new_[9692]_  ? \new_[4995]_  : \new_[3114]_ ;
  assign \new_[4083]_  = \new_[9153]_  ? \new_[11269]_  : \new_[10710]_ ;
  assign \new_[4084]_  = \new_[8766]_  ? \new_[11269]_  : \new_[11100]_ ;
  assign \new_[4085]_  = \new_[8816]_  ? \new_[11269]_  : \new_[10820]_ ;
  assign \new_[4086]_  = \new_[8261]_  ? \new_[11269]_  : \new_[11051]_ ;
  assign \new_[4087]_  = \new_[4706]_  | \new_[2927]_ ;
  assign \new_[4088]_  = \new_[10297]_  ? \new_[6070]_  : \new_[5061]_ ;
  assign \new_[4089]_  = \new_[9994]_  ? \new_[6070]_  : \new_[5062]_ ;
  assign \new_[4090]_  = ~\new_[5641]_  & (~\new_[5239]_  | ~\new_[6070]_ );
  assign \new_[4091]_  = (~\new_[5026]_  | ~\new_[6070]_ ) & (~\new_[10685]_  | ~\new_[5651]_ );
  assign \new_[4092]_  = ~\new_[12486]_  | ~\new_[4703]_ ;
  assign \new_[4093]_  = \new_[11495]_ ;
  assign \new_[4094]_  = ~\new_[11495]_ ;
  assign \new_[4095]_  = \new_[11495]_ ;
  assign \new_[4096]_  = \new_[7872]_  ? \new_[11269]_  : \new_[3180]_ ;
  assign \new_[4097]_  = ~\new_[4740]_  & (~\new_[6806]_  | ~\wb_addr_i[24] );
  assign \new_[4098]_  = ~\new_[4742]_  & (~\new_[6806]_  | ~\wb_addr_i[22] );
  assign \new_[4099]_  = ~\new_[10511]_  | ~\new_[4730]_  | ~\new_[8311]_ ;
  assign \new_[4100]_  = ~\new_[5980]_  | (~\new_[12738]_  & ~\new_[10258]_ );
  assign \new_[4101]_  = ~\new_[4651]_  & (~\new_[7539]_  | ~\new_[10265]_ );
  assign \new_[4102]_  = ~\new_[6207]_  | (~\new_[12743]_  & ~\new_[9718]_ );
  assign \new_[4103]_  = ~\new_[4649]_  & (~\new_[11500]_  | ~\new_[9620]_ );
  assign \new_[4104]_  = ~\new_[6210]_  | (~\new_[12745]_  & ~\new_[9867]_ );
  assign \new_[4105]_  = ~\new_[6211]_  | (~\new_[12738]_  & ~\new_[10146]_ );
  assign \new_[4106]_  = ~\new_[6216]_  | (~\new_[12738]_  & ~\new_[10155]_ );
  assign \new_[4107]_  = ~\new_[4671]_  & (~\new_[11500]_  | ~\new_[9848]_ );
  assign \new_[4108]_  = ~\new_[5984]_  | (~\new_[12738]_  & ~\new_[10161]_ );
  assign \new_[4109]_  = ~\new_[6219]_  | (~\new_[12738]_  & ~\new_[9996]_ );
  assign \new_[4110]_  = ~\new_[6221]_  | (~\new_[12738]_  & ~\new_[9908]_ );
  assign \new_[4111]_  = ~\new_[4679]_  & (~\new_[11500]_  | ~\new_[9668]_ );
  assign \new_[4112]_  = ~\new_[6226]_  | (~\new_[12738]_  & ~\new_[9866]_ );
  assign \new_[4113]_  = ~\new_[5625]_  | (~\new_[12738]_  & ~\new_[9617]_ );
  assign \new_[4114]_  = ~\new_[6228]_  | (~\new_[12738]_  & ~\new_[10262]_ );
  assign \new_[4115]_  = ~\new_[5990]_  | (~\new_[12738]_  & ~\new_[9590]_ );
  assign \new_[4116]_  = ~\new_[4683]_  & (~\new_[11500]_  | ~\new_[9649]_ );
  assign \new_[4117]_  = ~\new_[4685]_  & (~\new_[11500]_  | ~\new_[9965]_ );
  assign \new_[4118]_  = ~\new_[4686]_  & (~\new_[11500]_  | ~\new_[10055]_ );
  assign \new_[4119]_  = ~\new_[4687]_  & (~\new_[11500]_  | ~\new_[9841]_ );
  assign \new_[4120]_  = ~\new_[4688]_  & (~\new_[11500]_  | ~\new_[9610]_ );
  assign \new_[4121]_  = ~\new_[4689]_  & (~\new_[11500]_  | ~\new_[9843]_ );
  assign \new_[4122]_  = ~\new_[4643]_  & (~\new_[11500]_  | ~\new_[10087]_ );
  assign \new_[4123]_  = ~\new_[6263]_  | (~\new_[12743]_  & ~\new_[10255]_ );
  assign \new_[4124]_  = ~\new_[6229]_  | (~\new_[12738]_  & ~\new_[9653]_ );
  assign \new_[4125]_  = ~\new_[4705]_  & (~\new_[11500]_  | ~\new_[9846]_ );
  assign \new_[4126]_  = ~\\u5_ir_cnt_reg[3] ;
  assign \new_[4127]_  = ~\new_[4710]_  & (~\new_[11500]_  | ~\new_[9872]_ );
  assign \new_[4128]_  = ~\new_[6248]_  | ~\new_[4712]_ ;
  assign \new_[4129]_  = ~\new_[4715]_  & (~\new_[11500]_  | ~\new_[10015]_ );
  assign \new_[4130]_  = ~\new_[4716]_  & (~\new_[11500]_  | ~\new_[10044]_ );
  assign \new_[4131]_  = ~\new_[6255]_  | (~\new_[12738]_  & ~\new_[9921]_ );
  assign \new_[4132]_  = ~\new_[4719]_  & (~\new_[11500]_  | ~\new_[10127]_ );
  assign \new_[4133]_  = ~\new_[4722]_  & (~\new_[11500]_  | ~\new_[10049]_ );
  assign \new_[4134]_  = ~\new_[5628]_  | (~\new_[12738]_  & ~\new_[12113]_ );
  assign \new_[4135]_  = ~\new_[4726]_  & (~\new_[7539]_  | ~\new_[10089]_ );
  assign \new_[4136]_  = ~\new_[4729]_  & (~\new_[11500]_  | ~\new_[10048]_ );
  assign \new_[4137]_  = ~\new_[6262]_  | (~\new_[12746]_  & ~\new_[9732]_ );
  assign \new_[4138]_  = ~\new_[6265]_  | (~\new_[12743]_  & ~\new_[10166]_ );
  assign \new_[4139]_  = ~\new_[4731]_  & (~\new_[11500]_  | ~\new_[9608]_ );
  assign \new_[4140]_  = ~\new_[6264]_  | (~\new_[12738]_  & ~\new_[10199]_ );
  assign \new_[4141]_  = ~\new_[6204]_  | ~\new_[5617]_  | ~\new_[6203]_  | ~\new_[5644]_ ;
  assign \new_[4142]_  = ~\new_[7527]_  | (~\new_[12742]_  & ~\new_[9922]_ );
  assign \new_[4143]_  = ~\new_[6690]_  | ~\new_[4922]_  | ~\new_[5283]_ ;
  assign \new_[4144]_  = \new_[4734]_  & \new_[9750]_ ;
  assign \new_[4145]_  = \\u5_ir_cnt_reg[0] ;
  assign \new_[4146]_  = ~u5_mc_adv_r1_reg;
  assign \new_[4147]_  = u5_tmr2_done_reg;
  assign \new_[4148]_  = ~\new_[4453]_ ;
  assign \new_[4149]_  = (~\new_[12528]_  | ~\new_[10529]_ ) & (~\new_[5642]_  | ~\new_[11045]_ );
  assign \new_[4150]_  = ~\new_[7011]_  & ~\new_[12470]_ ;
  assign \new_[4151]_  = ~\new_[11474]_  | ~\new_[4709]_ ;
  assign \new_[4152]_  = ~\new_[11474]_  | ~\new_[12337]_ ;
  assign \new_[4153]_  = \new_[11468]_  & \new_[4974]_ ;
  assign \new_[4154]_  = \new_[7002]_  ? \new_[11269]_  : \new_[3225]_ ;
  assign \new_[4155]_  = ~\new_[9895]_  & (~\new_[5648]_  | ~\new_[6034]_ );
  assign \new_[4156]_  = ~\new_[4756]_  & (~\new_[7683]_  | ~\new_[10210]_ );
  assign \new_[4157]_  = ~\new_[4757]_  & (~\new_[7683]_  | ~\new_[9969]_ );
  assign \new_[4158]_  = \new_[7341]_  ? \new_[11269]_  : \new_[3177]_ ;
  assign \new_[4159]_  = \new_[8409]_  ? \new_[4995]_  : \new_[10836]_ ;
  assign \new_[4160]_  = \new_[8483]_  ? \new_[4995]_  : \new_[11205]_ ;
  assign \new_[4161]_  = \new_[5782]_  | \new_[11276]_ ;
  assign \new_[4162]_  = ~\new_[12528]_  & (~\new_[6109]_  | ~\new_[6594]_ );
  assign \new_[4163]_  = ~\new_[11277]_  & (~\new_[6110]_  | ~\new_[6597]_ );
  assign \new_[4164]_  = \new_[5791]_  | \new_[11276]_ ;
  assign \new_[4165]_  = \new_[5804]_  | \new_[12527]_ ;
  assign \new_[4166]_  = ~\new_[4758]_ ;
  assign \new_[4167]_  = \new_[4557]_  & \new_[5605]_ ;
  assign \new_[4168]_  = ~\new_[12527]_  & (~\new_[6111]_  | ~\new_[6618]_ );
  assign \new_[4169]_  = \new_[5794]_  | \new_[11276]_ ;
  assign \new_[4170]_  = ~\new_[5463]_  | ~\new_[7459]_  | ~\new_[4603]_  | ~\new_[12382]_ ;
  assign \new_[4171]_  = ~\new_[12527]_  & (~\new_[7631]_  | ~\new_[12696]_ );
  assign \new_[4172]_  = \new_[7614]_  ? \new_[4995]_  : \new_[3169]_ ;
  assign \new_[4173]_  = \new_[7798]_  ? \new_[4995]_  : \new_[11235]_ ;
  assign \new_[4174]_  = ~\new_[11337]_  | ~\new_[12239]_  | ~\new_[4926]_ ;
  assign \new_[4175]_  = \new_[7374]_  ? \new_[11271]_  : \new_[3179]_ ;
  assign \new_[4176]_  = ~\new_[4817]_  & (~\new_[11976]_  | ~\new_[10047]_ );
  assign \new_[4177]_  = ~\new_[4820]_  & (~\new_[11976]_  | ~\new_[9975]_ );
  assign \new_[4178]_  = ~\new_[6364]_  | ~\new_[12785]_  | ~\new_[4968]_  | ~\new_[7183]_ ;
  assign \new_[4179]_  = ~\new_[4886]_  & (~\new_[12534]_  | ~\new_[9608]_ );
  assign \new_[4180]_  = \\u3_u0_r0_reg[16] ;
  assign \new_[4181]_  = \\u3_u0_r0_reg[22] ;
  assign \new_[4182]_  = \\u3_u0_r1_reg[26] ;
  assign \new_[4183]_  = \\u3_u0_r2_reg[25] ;
  assign n2036 = ~\new_[4899]_  | ~\new_[10722]_ ;
  assign \new_[4185]_  = \\u3_u0_r2_reg[3] ;
  assign \new_[4186]_  = \\u3_u0_r0_reg[1] ;
  assign \new_[4187]_  = ~\new_[4926]_  & ~\new_[11814]_ ;
  assign \new_[4188]_  = \\u3_u0_r0_reg[18] ;
  assign \new_[4189]_  = \\u3_u0_r0_reg[19] ;
  assign \new_[4190]_  = \\u3_u0_r0_reg[10] ;
  assign \new_[4191]_  = \\u3_u0_r2_reg[32] ;
  assign n2041 = ~\new_[4900]_  & ~\new_[10928]_ ;
  assign \new_[4193]_  = ~\new_[10291]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4194]_  = ~\new_[10922]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4195]_  = \\u3_u0_r2_reg[27] ;
  assign \new_[4196]_  = ~\new_[11492]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4197]_  = ~\new_[9785]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4198]_  = \\u3_u0_r2_reg[29] ;
  assign \new_[4199]_  = \\u3_u0_r0_reg[14] ;
  assign \new_[4200]_  = ~\new_[10496]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4201]_  = ~\new_[12054]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4202]_  = ~\new_[10250]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4203]_  = ~\new_[12755]_  | ~\new_[11477]_  | ~\new_[7628]_ ;
  assign \new_[4204]_  = ~\new_[4995]_  & ~\new_[5384]_ ;
  assign \new_[4205]_  = \\u3_u0_r2_reg[18] ;
  assign \new_[4206]_  = \new_[12557]_  | \new_[10839]_ ;
  assign \new_[4207]_  = ~\new_[12688]_  | ~\new_[9841]_ ;
  assign \new_[4208]_  = ~\new_[4888]_  & (~\new_[11864]_  | ~\new_[9383]_ );
  assign \new_[4209]_  = ~\new_[5022]_  & (~\new_[5865]_  | ~\new_[9383]_ );
  assign \new_[4210]_  = ~\new_[5025]_  & (~\new_[5865]_  | ~\new_[10031]_ );
  assign \new_[4211]_  = ~\new_[5514]_  & (~\new_[5865]_  | ~\new_[9388]_ );
  assign \new_[4212]_  = ~\new_[5050]_  & (~\new_[5865]_  | ~\new_[9930]_ );
  assign \new_[4213]_  = ~\new_[5086]_  & (~\new_[5865]_  | ~\new_[8977]_ );
  assign \new_[4214]_  = ~\new_[5121]_  & (~\new_[5865]_  | ~\new_[9107]_ );
  assign \new_[4215]_  = ~\new_[5068]_  & (~\new_[5865]_  | ~\new_[9391]_ );
  assign \new_[4216]_  = ~\new_[4923]_  & (~\new_[6384]_  | ~\new_[10115]_ );
  assign \new_[4217]_  = ~\new_[4924]_  & (~\new_[6384]_  | ~\new_[9684]_ );
  assign \new_[4218]_  = ~\new_[4902]_  & (~\new_[7685]_  | ~\new_[9621]_ );
  assign \new_[4219]_  = ~\new_[4905]_  & (~\new_[7750]_  | ~\new_[9855]_ );
  assign \new_[4220]_  = ~\new_[4906]_  & (~\new_[7750]_  | ~\new_[9598]_ );
  assign \new_[4221]_  = ~\new_[4907]_  & (~\new_[7750]_  | ~\new_[9837]_ );
  assign \new_[4222]_  = ~\new_[4908]_  & (~\new_[12307]_  | ~\new_[9616]_ );
  assign \new_[4223]_  = ~\new_[4909]_  & (~\new_[7685]_  | ~\new_[9586]_ );
  assign \new_[4224]_  = ~\new_[4901]_  & (~\new_[7750]_  | ~\new_[9857]_ );
  assign \new_[4225]_  = ~\new_[4910]_  & (~\new_[7685]_  | ~\new_[9663]_ );
  assign \new_[4226]_  = ~\new_[4911]_  & (~\new_[12308]_  | ~\new_[9581]_ );
  assign \new_[4227]_  = ~\new_[4912]_  & (~\new_[12308]_  | ~\new_[9862]_ );
  assign \new_[4228]_  = ~\new_[4913]_  & (~\new_[12308]_  | ~\new_[9840]_ );
  assign \new_[4229]_  = ~\new_[4914]_  & (~\new_[7684]_  | ~\new_[10062]_ );
  assign \new_[4230]_  = ~\new_[4915]_  & (~\new_[7684]_  | ~\new_[9818]_ );
  assign \new_[4231]_  = \\u3_u0_r2_reg[21] ;
  assign \new_[4232]_  = ~\new_[4916]_  & (~\new_[12308]_  | ~\new_[9659]_ );
  assign \new_[4233]_  = ~\new_[4918]_  & (~\new_[7684]_  | ~\new_[9746]_ );
  assign \new_[4234]_  = ~\new_[4919]_  & (~\new_[7683]_  | ~\new_[9850]_ );
  assign \new_[4235]_  = ~\new_[12688]_  | ~\new_[9610]_ ;
  assign \new_[4236]_  = ~\\u3_u0_wr_adr_reg[1] ;
  assign \new_[4237]_  = ~\\u3_u0_wr_adr_reg[3] ;
  assign \new_[4238]_  = \new_[5911]_  & \new_[5018]_ ;
  assign \new_[4239]_  = \new_[7012]_  | \new_[4970]_ ;
  assign \new_[4240]_  = ~\new_[4576]_ ;
  assign \new_[4241]_  = ~\new_[11478]_ ;
  assign \new_[4242]_  = u5_rfr_ack_r_reg;
  assign \new_[4243]_  = ~\new_[11510]_  | ~\new_[4989]_ ;
  assign \new_[4244]_  = \new_[4992]_  | n3951;
  assign \new_[4245]_  = ~\new_[4974]_  & ~\new_[10964]_ ;
  assign n2086 = ~\new_[5243]_  | (~\new_[6739]_  & ~\new_[7600]_ );
  assign n2046 = ~\new_[5244]_  | (~\new_[6740]_  & ~\new_[7600]_ );
  assign \new_[4248]_  = ~\new_[4930]_  & (~\new_[8282]_  | ~\new_[11485]_ );
  assign \new_[4249]_  = \\u3_u0_r2_reg[14] ;
  assign \new_[4250]_  = ~\new_[4934]_  & (~\new_[8416]_  | ~\new_[11485]_ );
  assign \new_[4251]_  = ~\new_[4936]_  & (~\new_[8397]_  | ~\new_[11485]_ );
  assign \new_[4252]_  = ~\new_[4938]_  & (~\new_[8264]_  | ~\new_[11485]_ );
  assign \new_[4253]_  = ~\new_[4941]_  & (~\new_[8265]_  | ~\new_[11485]_ );
  assign \new_[4254]_  = ~\new_[4944]_  & (~\new_[8266]_  | ~\new_[11485]_ );
  assign \new_[4255]_  = \new_[4927]_  | \new_[10665]_ ;
  assign \new_[4256]_  = ~\new_[4952]_  & (~\new_[8269]_  | ~\new_[11485]_ );
  assign \new_[4257]_  = ~\new_[4958]_  & (~\new_[8273]_  | ~\new_[11485]_ );
  assign \new_[4258]_  = ~\new_[4973]_  & (~\new_[8262]_  | ~\new_[11485]_ );
  assign \new_[4259]_  = ~\new_[4982]_  & (~\new_[8283]_  | ~\new_[11485]_ );
  assign \new_[4260]_  = ~\new_[4988]_  & (~\new_[8278]_  | ~\new_[11485]_ );
  assign \new_[4261]_  = ~\new_[4991]_  & (~\new_[8275]_  | ~\new_[11485]_ );
  assign \new_[4262]_  = \new_[4933]_  & \new_[7987]_ ;
  assign \new_[4263]_  = ~\new_[4931]_  & (~\new_[11500]_  | ~\new_[10054]_ );
  assign \new_[4264]_  = ~\new_[4993]_  & (~\new_[11500]_  | ~\new_[10063]_ );
  assign \new_[4265]_  = ~\new_[4935]_  & (~\new_[11500]_  | ~\new_[9912]_ );
  assign \new_[4266]_  = ~\new_[4937]_  & (~\new_[11500]_  | ~\new_[10065]_ );
  assign \new_[4267]_  = ~\new_[4939]_  & (~\new_[11500]_  | ~\new_[10053]_ );
  assign \new_[4268]_  = ~\new_[4940]_  & (~\new_[11500]_  | ~\new_[10046]_ );
  assign \new_[4269]_  = ~\new_[4942]_  & (~\new_[11500]_  | ~\new_[9822]_ );
  assign \new_[4270]_  = ~\new_[4943]_  & (~\new_[11500]_  | ~\new_[9737]_ );
  assign \new_[4271]_  = ~\new_[4945]_  & (~\new_[11500]_  | ~\new_[9854]_ );
  assign \new_[4272]_  = ~\new_[4946]_  & (~\new_[11500]_  | ~\new_[10078]_ );
  assign \new_[4273]_  = ~\new_[4948]_  & (~\new_[12749]_  | ~\new_[9880]_ );
  assign \new_[4274]_  = ~\new_[4949]_  & (~\new_[11500]_  | ~\new_[9880]_ );
  assign \new_[4275]_  = ~\new_[4953]_  & (~\new_[11500]_  | ~\new_[10081]_ );
  assign \new_[4276]_  = ~\new_[4955]_  & (~\new_[11500]_  | ~\new_[10082]_ );
  assign \new_[4277]_  = ~\new_[4956]_  & (~\new_[11500]_  | ~\new_[9807]_ );
  assign \new_[4278]_  = \\u3_u0_r2_reg[10] ;
  assign \new_[4279]_  = ~\new_[4959]_  & (~\new_[11500]_  | ~\new_[10071]_ );
  assign \new_[4280]_  = ~\new_[6969]_  | (~\new_[6267]_  & ~\new_[9691]_ );
  assign \new_[4281]_  = ~\new_[4967]_  & (~\new_[11500]_  | ~\new_[10118]_ );
  assign \new_[4282]_  = ~\new_[6982]_  | (~\new_[6267]_  & ~\new_[10172]_ );
  assign \new_[4283]_  = ~\new_[4981]_  & (~\new_[11500]_  | ~\new_[10050]_ );
  assign \new_[4284]_  = ~\new_[6987]_  | (~\new_[6267]_  & ~\new_[9955]_ );
  assign \new_[4285]_  = ~\new_[6976]_  | (~\new_[6267]_  & ~\new_[9911]_ );
  assign \new_[4286]_  = ~\new_[4977]_  & (~\new_[11500]_  | ~\new_[10140]_ );
  assign \new_[4287]_  = ~\new_[4990]_  & (~\new_[11500]_  | ~\new_[10107]_ );
  assign \new_[4288]_  = ~\new_[4983]_  & (~\new_[12749]_  | ~\new_[9953]_ );
  assign \new_[4289]_  = \\u3_u0_r2_reg[12] ;
  assign \new_[4290]_  = ~\new_[4971]_  & (~\new_[8524]_  | ~\new_[11485]_ );
  assign \new_[4291]_  = ~\new_[7234]_  | (~\new_[6267]_  & ~\new_[9623]_ );
  assign \new_[4292]_  = ~\new_[4929]_  & (~\new_[7873]_  | ~\new_[9591]_ );
  assign \new_[4293]_  = \new_[4994]_  | \new_[7295]_ ;
  assign \new_[4294]_  = ~\new_[4644]_ ;
  assign \new_[4295]_  = \\u3_u0_r1_reg[9] ;
  assign \new_[4296]_  = ~\new_[5639]_  & ~\new_[7023]_ ;
  assign \new_[4297]_  = ~\new_[12690]_  | ~\new_[9953]_ ;
  assign \new_[4298]_  = ~\new_[4648]_ ;
  assign \new_[4299]_  = ~\new_[12688]_  | ~\new_[11787]_ ;
  assign \new_[4300]_  = ~\new_[12683]_  | ~\new_[12689]_ ;
  assign \new_[4301]_  = ~\new_[12690]_  | ~\new_[12060]_ ;
  assign \new_[4302]_  = ~\new_[7629]_  | ~\new_[12682]_  | ~\new_[7649]_ ;
  assign \new_[4303]_  = \\u3_u0_r1_reg[7] ;
  assign \new_[4304]_  = ~\new_[12692]_  | ~\new_[10054]_ ;
  assign \new_[4305]_  = ~\new_[12688]_  | ~\new_[9985]_ ;
  assign \new_[4306]_  = ~\new_[12688]_  | ~\new_[10049]_ ;
  assign \new_[4307]_  = ~\new_[7631]_  | ~\new_[12679]_  | ~\new_[7483]_ ;
  assign \new_[4308]_  = ~\new_[12692]_  | ~\new_[10065]_ ;
  assign \new_[4309]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7311]_ ;
  assign \new_[4310]_  = ~\new_[7663]_  | ~\new_[12682]_  | ~\new_[7506]_ ;
  assign \new_[4311]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7487]_ ;
  assign \new_[4312]_  = ~\new_[12688]_  | ~\new_[10056]_ ;
  assign \new_[4313]_  = \\u3_u0_r1_reg[3] ;
  assign \new_[4314]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7314]_ ;
  assign \new_[4315]_  = ~\new_[12688]_  | ~\new_[9849]_ ;
  assign \new_[4316]_  = ~\new_[7663]_  | ~\new_[12679]_  | ~\new_[7489]_ ;
  assign \new_[4317]_  = ~\new_[12688]_  | ~\new_[10244]_ ;
  assign \new_[4318]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7768]_ ;
  assign \new_[4319]_  = ~\new_[12688]_  | ~\new_[10055]_ ;
  assign \new_[4320]_  = ~\new_[12692]_  | ~\new_[10130]_ ;
  assign \new_[4321]_  = ~\new_[12692]_  | ~\new_[10061]_ ;
  assign \new_[4322]_  = ~\new_[7629]_  | ~\new_[12678]_  | ~\new_[7494]_ ;
  assign \new_[4323]_  = ~\new_[12690]_  | ~\new_[9668]_ ;
  assign \new_[4324]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7495]_ ;
  assign \new_[4325]_  = ~\new_[7663]_  | ~\new_[12679]_  | ~\new_[7497]_ ;
  assign \new_[4326]_  = ~\new_[12692]_  | ~\new_[10071]_ ;
  assign \new_[4327]_  = ~\new_[12738]_  & ~\new_[11865]_ ;
  assign \new_[4328]_  = ~\new_[12690]_  | ~\new_[9694]_ ;
  assign \new_[4329]_  = ~\new_[7629]_  | ~\new_[12678]_  | ~\new_[7502]_ ;
  assign \new_[4330]_  = ~\new_[12688]_  | ~\new_[9649]_ ;
  assign \new_[4331]_  = ~\new_[12688]_  | ~\new_[9970]_ ;
  assign \new_[4332]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7503]_ ;
  assign \new_[4333]_  = ~\new_[12688]_  | ~\new_[9965]_ ;
  assign \new_[4334]_  = ~\new_[7629]_  | ~\new_[12678]_  | ~\new_[7514]_ ;
  assign \new_[4335]_  = ~\new_[12688]_  | ~\new_[9594]_ ;
  assign \new_[4336]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7315]_ ;
  assign \new_[4337]_  = ~\new_[12690]_  | ~\new_[9856]_ ;
  assign \new_[4338]_  = ~\new_[7629]_  | ~\new_[12678]_  | ~\new_[7488]_ ;
  assign \new_[4339]_  = \\u3_u0_r1_reg[32] ;
  assign \new_[4340]_  = ~\\u3_u0_wr_adr_reg[0] ;
  assign \new_[4341]_  = ~\\u3_u0_wr_adr_reg[2] ;
  assign \new_[4342]_  = \\u3_u0_r0_reg[0] ;
  assign \new_[4343]_  = \\u3_u0_r0_reg[11] ;
  assign \new_[4344]_  = \\u3_u0_r0_reg[12] ;
  assign \new_[4345]_  = \\u3_u0_r0_reg[13] ;
  assign \new_[4346]_  = \\u3_u0_r0_reg[15] ;
  assign \new_[4347]_  = \\u3_u0_r0_reg[17] ;
  assign \new_[4348]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7485]_ ;
  assign \new_[4349]_  = \\u3_u0_r0_reg[20] ;
  assign \new_[4350]_  = \\u3_u0_r0_reg[21] ;
  assign \new_[4351]_  = \\u3_u0_r0_reg[23] ;
  assign \new_[4352]_  = \\u3_u0_r0_reg[24] ;
  assign \new_[4353]_  = \\u3_u0_r0_reg[26] ;
  assign \new_[4354]_  = \\u3_u0_r0_reg[27] ;
  assign \new_[4355]_  = \\u3_u0_r0_reg[28] ;
  assign \new_[4356]_  = \\u3_u0_r0_reg[2] ;
  assign \new_[4357]_  = \\u3_u0_r0_reg[30] ;
  assign \new_[4358]_  = \\u3_u0_r0_reg[31] ;
  assign \new_[4359]_  = \\u3_u0_r0_reg[33] ;
  assign \new_[4360]_  = \\u3_u0_r0_reg[34] ;
  assign \new_[4361]_  = \\u3_u0_r0_reg[35] ;
  assign \new_[4362]_  = \\u3_u0_r0_reg[4] ;
  assign \new_[4363]_  = ~\new_[12688]_  | ~\new_[9843]_ ;
  assign \new_[4364]_  = \\u3_u0_r0_reg[9] ;
  assign \new_[4365]_  = \\u3_u0_r1_reg[0] ;
  assign \new_[4366]_  = \\u3_u0_r1_reg[11] ;
  assign \new_[4367]_  = ~\new_[7629]_  | ~\new_[12685]_  | ~\new_[7508]_ ;
  assign \new_[4368]_  = \\u3_u0_r1_reg[10] ;
  assign \new_[4369]_  = \\u3_u0_r1_reg[12] ;
  assign \new_[4370]_  = \\u3_u0_r1_reg[13] ;
  assign \new_[4371]_  = \\u3_u0_r1_reg[15] ;
  assign \new_[4372]_  = \\u3_u0_r1_reg[16] ;
  assign \new_[4373]_  = \\u3_u0_r1_reg[17] ;
  assign \new_[4374]_  = \\u3_u0_r1_reg[19] ;
  assign \new_[4375]_  = \\u3_u0_r1_reg[1] ;
  assign \new_[4376]_  = \\u3_u0_r1_reg[20] ;
  assign \new_[4377]_  = \\u3_u0_r1_reg[23] ;
  assign \new_[4378]_  = \\u3_u0_r1_reg[22] ;
  assign \new_[4379]_  = \\u3_u0_r1_reg[24] ;
  assign \new_[4380]_  = \\u3_u0_r1_reg[25] ;
  assign \new_[4381]_  = \\u3_u0_r1_reg[27] ;
  assign \new_[4382]_  = \\u3_u0_r1_reg[28] ;
  assign \new_[4383]_  = \\u3_u0_r1_reg[2] ;
  assign \new_[4384]_  = \\u3_u0_r1_reg[30] ;
  assign \new_[4385]_  = \\u3_u0_r1_reg[31] ;
  assign \new_[4386]_  = \\u3_u0_r1_reg[33] ;
  assign \new_[4387]_  = \\u3_u0_r1_reg[34] ;
  assign \new_[4388]_  = \\u3_u0_r1_reg[35] ;
  assign \new_[4389]_  = \\u3_u0_r1_reg[4] ;
  assign \new_[4390]_  = \\u3_u0_r1_reg[5] ;
  assign \new_[4391]_  = \\u3_u0_r1_reg[6] ;
  assign \new_[4392]_  = \\u3_u0_r1_reg[8] ;
  assign \new_[4393]_  = \\u3_u0_r2_reg[0] ;
  assign \new_[4394]_  = ~\new_[12688]_  | ~\new_[10087]_ ;
  assign \new_[4395]_  = \\u3_u0_r2_reg[11] ;
  assign \new_[4396]_  = \\u3_u0_r2_reg[13] ;
  assign \new_[4397]_  = \\u3_u0_r2_reg[15] ;
  assign \new_[4398]_  = \\u3_u0_r2_reg[16] ;
  assign \new_[4399]_  = \\u3_u0_r2_reg[17] ;
  assign \new_[4400]_  = \\u3_u0_r2_reg[19] ;
  assign \new_[4401]_  = \\u3_u0_r2_reg[1] ;
  assign \new_[4402]_  = \\u3_u0_r2_reg[20] ;
  assign \new_[4403]_  = \\u3_u0_r2_reg[22] ;
  assign \new_[4404]_  = \\u3_u0_r2_reg[23] ;
  assign \new_[4405]_  = \\u3_u0_r2_reg[24] ;
  assign \new_[4406]_  = \\u3_u0_r2_reg[26] ;
  assign \new_[4407]_  = \\u3_u0_r2_reg[28] ;
  assign \new_[4408]_  = \\u3_u0_r2_reg[2] ;
  assign \new_[4409]_  = \\u3_u0_r2_reg[30] ;
  assign \new_[4410]_  = \\u3_u0_r2_reg[31] ;
  assign \new_[4411]_  = \\u3_u0_r2_reg[33] ;
  assign \new_[4412]_  = \\u3_u0_r2_reg[34] ;
  assign \new_[4413]_  = \\u3_u0_r2_reg[35] ;
  assign \new_[4414]_  = \\u3_u0_r2_reg[4] ;
  assign \new_[4415]_  = \\u3_u0_r2_reg[5] ;
  assign \new_[4416]_  = \\u3_u0_r2_reg[6] ;
  assign \new_[4417]_  = \\u3_u0_r2_reg[8] ;
  assign \new_[4418]_  = \\u3_u0_r3_reg[0] ;
  assign \new_[4419]_  = \\u3_u0_r3_reg[11] ;
  assign \new_[4420]_  = \\u3_u0_r3_reg[12] ;
  assign \new_[4421]_  = \\u3_u0_r3_reg[13] ;
  assign \new_[4422]_  = \\u3_u0_r3_reg[15] ;
  assign \new_[4423]_  = \\u3_u0_r3_reg[16] ;
  assign \new_[4424]_  = \\u3_u0_r3_reg[17] ;
  assign \new_[4425]_  = \\u3_u0_r3_reg[19] ;
  assign \new_[4426]_  = \\u3_u0_r3_reg[1] ;
  assign \new_[4427]_  = \\u3_u0_r3_reg[20] ;
  assign \new_[4428]_  = \\u3_u0_r3_reg[22] ;
  assign \new_[4429]_  = \\u3_u0_r3_reg[23] ;
  assign \new_[4430]_  = \\u3_u0_r3_reg[24] ;
  assign \new_[4431]_  = \\u3_u0_r3_reg[26] ;
  assign \new_[4432]_  = \\u3_u0_r3_reg[28] ;
  assign \new_[4433]_  = \\u3_u0_r3_reg[2] ;
  assign \new_[4434]_  = \\u3_u0_r3_reg[31] ;
  assign \new_[4435]_  = ~\new_[12692]_  | ~\new_[10153]_ ;
  assign \new_[4436]_  = \\u3_u0_r3_reg[33] ;
  assign \new_[4437]_  = \\u3_u0_r3_reg[34] ;
  assign \new_[4438]_  = \\u3_u0_r3_reg[35] ;
  assign \new_[4439]_  = \\u3_u0_r3_reg[4] ;
  assign \new_[4440]_  = \\u3_u0_r3_reg[5] ;
  assign \new_[4441]_  = \\u3_u0_r3_reg[6] ;
  assign \new_[4442]_  = \\u3_u0_r3_reg[9] ;
  assign \new_[4443]_  = \\u3_u0_r3_reg[8] ;
  assign \new_[4444]_  = ~\new_[12688]_  | ~\new_[11452]_ ;
  assign \new_[4445]_  = ~\new_[7663]_  | ~\new_[12679]_  | ~\new_[7517]_ ;
  assign \new_[4446]_  = ~\new_[12688]_  | ~\new_[9904]_ ;
  assign \new_[4447]_  = ~\new_[7522]_  | ~\new_[12678]_  | ~\new_[7499]_ ;
  assign \new_[4448]_  = \\u3_u0_r1_reg[29] ;
  assign \new_[4449]_  = ~\new_[6322]_  | ~\new_[6034]_  | ~\new_[6654]_ ;
  assign \new_[4450]_  = ~\new_[4706]_ ;
  assign \new_[4451]_  = ~\new_[12688]_  | ~\new_[9846]_ ;
  assign \new_[4452]_  = ~\new_[12688]_  | ~\new_[9606]_ ;
  assign \new_[4453]_  = ~\new_[7077]_  & ~\new_[12239]_ ;
  assign \new_[4454]_  = ~\new_[12690]_  | ~\new_[9847]_ ;
  assign \new_[4455]_  = ~\new_[7629]_  | ~\new_[12679]_  | ~\new_[7500]_ ;
  assign \new_[4456]_  = ~\new_[12688]_  | ~\new_[10043]_ ;
  assign \new_[4457]_  = ~\new_[12690]_  | ~\new_[9872]_ ;
  assign \new_[4458]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7660]_ ;
  assign \new_[4459]_  = ~\new_[12688]_  | ~\new_[10051]_ ;
  assign \new_[4460]_  = ~\new_[12690]_  | ~\new_[9871]_ ;
  assign \new_[4461]_  = ~\new_[12692]_  | ~\new_[10015]_ ;
  assign \new_[4462]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7498]_ ;
  assign \new_[4463]_  = ~\new_[12688]_  | ~\new_[10044]_ ;
  assign \new_[4464]_  = ~\new_[12692]_  | ~\new_[9870]_ ;
  assign \new_[4465]_  = ~\new_[12690]_  | ~\new_[10140]_ ;
  assign \new_[4466]_  = ~\new_[12688]_  | ~\new_[10089]_ ;
  assign \new_[4467]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7310]_ ;
  assign \new_[4468]_  = ~\new_[12688]_  | ~\new_[10048]_ ;
  assign \new_[4469]_  = ~\new_[12688]_  | ~\new_[10059]_ ;
  assign \new_[4470]_  = ~\new_[7663]_  | ~\new_[12685]_  | ~\new_[7321]_ ;
  assign \new_[4471]_  = \new_[5285]_  & \new_[11450]_ ;
  assign n2031 = ~\new_[8357]_  | ~\new_[5287]_ ;
  assign \new_[4473]_  = ~\new_[9998]_  | ~\new_[5248]_  | ~\new_[11045]_ ;
  assign \new_[4474]_  = \\u3_u0_r1_reg[21] ;
  assign \new_[4475]_  = ~\new_[10808]_  | ~\new_[5248]_  | ~\new_[11045]_ ;
  assign \new_[4476]_  = ~\new_[9785]_  | ~\new_[5248]_  | ~\new_[11233]_ ;
  assign \new_[4477]_  = ~\new_[9968]_  | ~\new_[5248]_  | ~\new_[11045]_ ;
  assign \new_[4478]_  = ~\new_[12598]_  | ~\new_[5248]_  | ~\new_[11045]_ ;
  assign \new_[4479]_  = (~\new_[6290]_  | ~\wb_addr_i[15] ) & (~\new_[6666]_  | ~\wb_addr_i[14] );
  assign \new_[4480]_  = \\u3_u0_r0_reg[7] ;
  assign \new_[4481]_  = (~\new_[6290]_  | ~\wb_addr_i[12] ) & (~\new_[6063]_  | ~\wb_addr_i[11] );
  assign \new_[4482]_  = (~\new_[5646]_  | ~\wb_addr_i[13] ) & (~\new_[6063]_  | ~\wb_addr_i[12] );
  assign \new_[4483]_  = (~\new_[6290]_  | ~\wb_addr_i[25] ) & (~\new_[11725]_  | ~\wb_addr_i[23] );
  assign \new_[4484]_  = (~\new_[6290]_  | ~\wb_addr_i[14] ) & (~\new_[6666]_  | ~\wb_addr_i[13] );
  assign \new_[4485]_  = (~\new_[5646]_  | ~\wb_addr_i[22] ) & (~\new_[6063]_  | ~\wb_addr_i[21] );
  assign \new_[4486]_  = (~\new_[6290]_  | ~\wb_addr_i[23] ) & (~\new_[6063]_  | ~\wb_addr_i[22] );
  assign \new_[4487]_  = (~\new_[6290]_  | ~\wb_addr_i[16] ) & (~\new_[6666]_  | ~\wb_addr_i[15] );
  assign \new_[4488]_  = (~\new_[5646]_  | ~\wb_addr_i[18] ) & (~\new_[6666]_  | ~\wb_addr_i[17] );
  assign \new_[4489]_  = (~\new_[5646]_  | ~\wb_addr_i[19] ) & (~\new_[6063]_  | ~\wb_addr_i[18] );
  assign \new_[4490]_  = (~\new_[5646]_  | ~\wb_addr_i[20] ) & (~\new_[6666]_  | ~\wb_addr_i[19] );
  assign \new_[4491]_  = (~\new_[5646]_  | ~\wb_addr_i[21] ) & (~\new_[6666]_  | ~\wb_addr_i[20] );
  assign \new_[4492]_  = (~\new_[6290]_  | ~\wb_addr_i[17] ) & (~\new_[6063]_  | ~\wb_addr_i[16] );
  assign \new_[4493]_  = ~\new_[10634]_  | ~\new_[5248]_  | ~\new_[11045]_ ;
  assign \new_[4494]_  = \\u3_u0_r1_reg[18] ;
  assign \new_[4495]_  = \\u3_u0_r3_reg[7] ;
  assign n2051 = \new_[10845]_  ? \new_[5640]_  : \new_[3884]_ ;
  assign n2056 = \new_[10844]_  ? \new_[5640]_  : \new_[3885]_ ;
  assign n2061 = \new_[10968]_  ? \new_[5640]_  : \new_[3886]_ ;
  assign n2081 = \new_[10916]_  ? \new_[5640]_  : \new_[3917]_ ;
  assign n2066 = \new_[10869]_  ? \new_[5640]_  : \new_[3887]_ ;
  assign n2071 = \new_[10852]_  ? \new_[5640]_  : \new_[3888]_ ;
  assign n2076 = \new_[10819]_  ? \new_[5640]_  : \new_[3889]_ ;
  assign n2026 = \new_[10833]_  ? \new_[5640]_  : \new_[3876]_ ;
  assign \new_[4504]_  = \\u3_u0_r3_reg[3] ;
  assign \new_[4505]_  = ~\new_[5245]_  & (~\new_[6674]_  | ~\new_[10200]_ );
  assign \new_[4506]_  = \\u3_u0_r3_reg[30] ;
  assign \new_[4507]_  = ~\new_[7629]_  | ~\new_[12678]_  | ~\new_[7507]_ ;
  assign \new_[4508]_  = \new_[11114]_  ^ \new_[5645]_ ;
  assign \new_[4509]_  = \\u3_u0_r3_reg[32] ;
  assign \new_[4510]_  = \\u3_u0_r1_reg[14] ;
  assign \new_[4511]_  = \\u3_u0_r3_reg[25] ;
  assign \new_[4512]_  = \\u3_u0_r3_reg[29] ;
  assign \new_[4513]_  = ~\new_[4995]_  & ~\new_[5350]_ ;
  assign \new_[4514]_  = \\u3_u0_r0_reg[8] ;
  assign \new_[4515]_  = \\u3_u0_r3_reg[27] ;
  assign \new_[4516]_  = \\u3_u0_r0_reg[5] ;
  assign \new_[4517]_  = \\u3_u0_r3_reg[14] ;
  assign \new_[4518]_  = \\u3_u0_r3_reg[21] ;
  assign \new_[4519]_  = \\u3_u0_r0_reg[6] ;
  assign \new_[4520]_  = ~\new_[5393]_  | ~\new_[7306]_  | ~\new_[6016]_ ;
  assign \new_[4521]_  = \\u3_u0_r2_reg[7] ;
  assign \new_[4522]_  = ~u4_rfr_clr_reg;
  assign \new_[4523]_  = \\u3_u0_r0_reg[3] ;
  assign \new_[4524]_  = ~\new_[12740]_  | ~\new_[4813]_ ;
  assign \new_[4525]_  = ~\new_[7159]_  & ~\new_[11277]_ ;
  assign \new_[4526]_  = ~\new_[6729]_  | ~\new_[4813]_ ;
  assign \new_[4527]_  = \\u3_u0_r3_reg[18] ;
  assign \new_[4528]_  = \\u3_u0_r0_reg[32] ;
  assign \new_[4529]_  = ~\new_[4995]_  & ~\new_[4839]_ ;
  assign \new_[4530]_  = ~\new_[11271]_  & ~\new_[7114]_ ;
  assign \new_[4531]_  = \\u3_u0_r0_reg[29] ;
  assign \new_[4532]_  = \\u3_u0_r0_reg[25] ;
  assign \new_[4533]_  = \\u3_u0_r2_reg[9] ;
  assign \new_[4534]_  = ~\new_[4811]_  & (~\new_[11976]_  | ~\new_[10064]_ );
  assign \new_[4535]_  = \\u3_u0_r3_reg[10] ;
  assign \new_[4536]_  = ~\new_[4814]_  & (~\new_[11976]_  | ~\new_[9824]_ );
  assign \new_[4537]_  = ~\new_[5340]_  & (~\new_[11976]_  | ~\new_[9818]_ );
  assign \new_[4538]_  = ~\new_[5341]_  & (~\new_[11976]_  | ~\new_[9659]_ );
  assign \new_[4539]_  = ~\new_[5342]_  & (~\new_[11976]_  | ~\new_[9746]_ );
  assign \new_[4540]_  = ~\new_[5343]_  & (~\new_[11976]_  | ~\new_[9850]_ );
  assign \new_[4541]_  = ~\new_[5344]_  & (~\new_[11976]_  | ~\new_[9393]_ );
  assign \new_[4542]_  = ~\new_[5345]_  & (~\new_[11976]_  | ~\new_[9874]_ );
  assign \new_[4543]_  = ~\new_[5346]_  & (~\new_[11976]_  | ~\new_[9863]_ );
  assign \new_[4544]_  = ~\new_[5347]_  & (~\new_[11976]_  | ~\new_[9596]_ );
  assign \new_[4545]_  = (~\new_[5749]_  | ~\new_[8408]_ ) & (~\new_[8215]_  | ~\new_[12657]_ );
  assign n2101 = (~n2921 & ~\new_[10072]_ ) | (~\new_[4146]_  & ~n5306);
  assign \new_[4547]_  = ~\new_[8022]_  & (~\new_[5695]_  | ~\new_[12469]_ );
  assign n2091 = ~\new_[10928]_  & (~\new_[5859]_  | ~\new_[5871]_ );
  assign \new_[4549]_  = ~\new_[5398]_  & (~\new_[8218]_  | ~\new_[12655]_ );
  assign n2096 = ~\new_[5431]_  & ~\new_[10928]_ ;
  assign \new_[4551]_  = ~\new_[7534]_  | ~\new_[6283]_  | ~\new_[6466]_  | ~\new_[5994]_ ;
  assign \mc_addr_pad_o[23]  = \\u7_mc_addr_reg[23] ;
  assign \new_[4553]_  = (~\new_[6805]_  & ~\new_[8394]_  & ~\new_[6722]_ ) | (~\new_[5981]_  & ~\new_[6722]_  & ~\new_[8740]_ );
  assign \mc_addr_pad_o[17]  = \\u7_mc_addr_reg[17] ;
  assign \new_[4555]_  = ~\new_[5585]_  & (~\new_[5865]_  | ~\new_[9978]_ );
  assign \new_[4556]_  = ~\new_[5592]_  & (~\new_[5865]_  | ~\new_[10083]_ );
  assign \new_[4557]_  = ~\new_[5584]_  & (~\new_[5865]_  | ~\new_[9389]_ );
  assign n2106 = ~\new_[4823]_ ;
  assign \new_[4559]_  = ~\new_[6116]_  | ~\new_[7296]_  | ~\new_[11503]_  | ~\new_[7863]_ ;
  assign \new_[4560]_  = ~\new_[8044]_  & (~\new_[5703]_  | ~\new_[12469]_ );
  assign \new_[4561]_  = ~\new_[7994]_  & (~\new_[5879]_  | ~\new_[6376]_ );
  assign \new_[4562]_  = ~\new_[7994]_  & (~\new_[5879]_  | ~\new_[6677]_ );
  assign \new_[4563]_  = \new_[5513]_  & \new_[12736]_ ;
  assign \new_[4564]_  = ~\new_[5865]_  | ~\new_[9661]_ ;
  assign \new_[4565]_  = ~\new_[5865]_  | ~\new_[9963]_ ;
  assign \new_[4566]_  = ~\new_[5865]_  | ~\new_[9418]_ ;
  assign \new_[4567]_  = ~\new_[5865]_  | ~\new_[10126]_ ;
  assign \new_[4568]_  = ~\new_[5865]_  | ~\new_[9987]_ ;
  assign \new_[4569]_  = ~\new_[5865]_  | ~\new_[9644]_ ;
  assign \new_[4570]_  = ~\new_[5865]_  | ~\new_[9655]_ ;
  assign \new_[4571]_  = ~\new_[5865]_  | ~\new_[9168]_ ;
  assign \new_[4572]_  = ~\new_[5865]_  | ~\new_[9657]_ ;
  assign \new_[4573]_  = \new_[5475]_  | \new_[6688]_ ;
  assign \new_[4574]_  = ~\new_[5865]_  | ~\new_[10097]_ ;
  assign \new_[4575]_  = \new_[11477]_ ;
  assign \new_[4576]_  = ~\new_[11479]_ ;
  assign \new_[4577]_  = \new_[11477]_ ;
  assign \new_[4578]_  = ~\new_[5977]_  | ~\new_[7708]_  | ~\new_[7988]_ ;
  assign \new_[4579]_  = ~\new_[5865]_  | ~\new_[9990]_ ;
  assign \new_[4580]_  = ~\new_[5865]_  | ~\new_[10037]_ ;
  assign \new_[4581]_  = ~\new_[7446]_  | (~\new_[6640]_  & ~\new_[9851]_ );
  assign \new_[4582]_  = ~\new_[5437]_  & (~\new_[8414]_  | ~\new_[11485]_ );
  assign \new_[4583]_  = ~\new_[5440]_  & (~\new_[8144]_  | ~\new_[11485]_ );
  assign \new_[4584]_  = ~\new_[7760]_  | (~\new_[5879]_  & ~\new_[7823]_ );
  assign \new_[4585]_  = ~\new_[5442]_  & (~\new_[8418]_  | ~\new_[11485]_ );
  assign \new_[4586]_  = ~\new_[7452]_  | (~\new_[6640]_  & ~\new_[9894]_ );
  assign \new_[4587]_  = ~\new_[5445]_  & (~\new_[8267]_  | ~\new_[11485]_ );
  assign \new_[4588]_  = ~\new_[5447]_  & (~\new_[8268]_  | ~\new_[11485]_ );
  assign \new_[4589]_  = ~\new_[7457]_  | (~\new_[6641]_  & ~\new_[10161]_ );
  assign \new_[4590]_  = ~\new_[5452]_  & (~\new_[8270]_  | ~\new_[11485]_ );
  assign \new_[4591]_  = ~\new_[5453]_  & (~\new_[8271]_  | ~\new_[11485]_ );
  assign \new_[4592]_  = ~\new_[5454]_  & (~\new_[8276]_  | ~\new_[11485]_ );
  assign \new_[4593]_  = ~\new_[5457]_  & (~\new_[8421]_  | ~\new_[11485]_ );
  assign \new_[4594]_  = ~\new_[5459]_  & (~\new_[8272]_  | ~\new_[11485]_ );
  assign \new_[4595]_  = ~\new_[5460]_  & (~\new_[8146]_  | ~\new_[11485]_ );
  assign \new_[4596]_  = ~\new_[5465]_  & (~\new_[8419]_  | ~\new_[11485]_ );
  assign \new_[4597]_  = ~\new_[5474]_  & (~\new_[8279]_  | ~\new_[11485]_ );
  assign \new_[4598]_  = ~\new_[5497]_  & (~\new_[8280]_  | ~\new_[11485]_ );
  assign \new_[4599]_  = ~\new_[5477]_  & (~\new_[8420]_  | ~\new_[11485]_ );
  assign \new_[4600]_  = ~\new_[5486]_  & (~\new_[8277]_  | ~\new_[11485]_ );
  assign \new_[4601]_  = ~\new_[5490]_  & (~\new_[8281]_  | ~\new_[11485]_ );
  assign \new_[4602]_  = ~\new_[5483]_  & (~\new_[8417]_  | ~\new_[11485]_ );
  assign \new_[4603]_  = ~\new_[5501]_  & (~\new_[11864]_  | ~\new_[9340]_ );
  assign \new_[4604]_  = ~\new_[5500]_  & (~\new_[6809]_  | ~\new_[10263]_ );
  assign \new_[4605]_  = ~\new_[6710]_  | (~\new_[7176]_  & ~\new_[9177]_ );
  assign \new_[4606]_  = ~\new_[6702]_  | (~\new_[7176]_  & ~\new_[9715]_ );
  assign \new_[4607]_  = ~\new_[5433]_  & (~\new_[11500]_  | ~\new_[11787]_ );
  assign \new_[4608]_  = ~\new_[5434]_  & (~\new_[12751]_  | ~\new_[11787]_ );
  assign \new_[4609]_  = ~\new_[5435]_  & (~\new_[11500]_  | ~\new_[12060]_ );
  assign \new_[4610]_  = ~\new_[5439]_  & (~\new_[11500]_  | ~\new_[9985]_ );
  assign \new_[4611]_  = ~\new_[6220]_  | (~\new_[12741]_  & ~\new_[10208]_ );
  assign \new_[4612]_  = ~\new_[6209]_  | (~\new_[12741]_  & ~\new_[10229]_ );
  assign \new_[4613]_  = ~\new_[6213]_  | (~\new_[12742]_  & ~\new_[10234]_ );
  assign \new_[4614]_  = ~\new_[5443]_  & (~\new_[12747]_  | ~\new_[9737]_ );
  assign \new_[4615]_  = ~\new_[6214]_  | (~\new_[12742]_  & ~\new_[9838]_ );
  assign \new_[4616]_  = ~\new_[6217]_  | (~\new_[12741]_  & ~\new_[9925]_ );
  assign \new_[4617]_  = ~\new_[6218]_  | (~\new_[12738]_  & ~\new_[10254]_ );
  assign \new_[4618]_  = ~\new_[5451]_  & (~\new_[11500]_  | ~\new_[10244]_ );
  assign \new_[4619]_  = ~\new_[5985]_  | (~\new_[12742]_  & ~\new_[10057]_ );
  assign \new_[4620]_  = ~\new_[6225]_  | ~\new_[5456]_ ;
  assign \new_[4621]_  = ~\new_[5462]_  & (~\new_[11500]_  | ~\new_[9694]_ );
  assign \new_[4622]_  = ~\new_[6233]_  | ~\new_[5464]_ ;
  assign \new_[4623]_  = ~\new_[5470]_  & (~\new_[12748]_  | ~\new_[10055]_ );
  assign \new_[4624]_  = ~\new_[5650]_  & (~\new_[12750]_  | ~\new_[9610]_ );
  assign \new_[4625]_  = ~\new_[5354]_  & (~\new_[12751]_  | ~\new_[9843]_ );
  assign \new_[4626]_  = ~\new_[5375]_  & (~\new_[11500]_  | ~\new_[10153]_ );
  assign \new_[4627]_  = ~\new_[6615]_  | (~\new_[12745]_  & ~\new_[10150]_ );
  assign \new_[4628]_  = ~\new_[5505]_  & (~\new_[11500]_  | ~\new_[11452]_ );
  assign \new_[4629]_  = ~\new_[5478]_  & (~\new_[11500]_  | ~\new_[9839]_ );
  assign \new_[4630]_  = ~\new_[5479]_  & (~\new_[11500]_  | ~\new_[9606]_ );
  assign \new_[4631]_  = ~\new_[6241]_  | (~\new_[12738]_  & ~\new_[9305]_ );
  assign \new_[4632]_  = ~\new_[5444]_  & (~\new_[11500]_  | ~\new_[9970]_ );
  assign \new_[4633]_  = ~\new_[6227]_  | (~\new_[12740]_  & ~\new_[9715]_ );
  assign \new_[4634]_  = ~\new_[5480]_  & (~\new_[11500]_  | ~\new_[9847]_ );
  assign \new_[4635]_  = ~\new_[6231]_  | (~\new_[12738]_  & ~\new_[9743]_ );
  assign \new_[4636]_  = ~\new_[6249]_  | ~\new_[5485]_ ;
  assign \new_[4637]_  = ~\new_[6003]_  | (~\new_[12742]_  & ~\new_[10172]_ );
  assign \new_[4638]_  = ~\new_[5499]_  & (~\new_[11500]_  | ~\new_[9953]_ );
  assign \new_[4639]_  = (~\new_[11715]_  | ~\wb_addr_i[22] ) & (~\new_[5997]_  | ~\wb_addr_i[21] );
  assign \new_[4640]_  = ~\new_[7530]_  | (~\new_[6267]_  & ~\new_[9996]_ );
  assign \new_[4641]_  = \new_[7536]_  | \new_[5482]_ ;
  assign \new_[4642]_  = \new_[7542]_  | \new_[5487]_ ;
  assign \new_[4643]_  = ~\new_[6267]_  & ~\new_[9954]_ ;
  assign \new_[4644]_  = ~\new_[11885]_ ;
  assign \new_[4645]_  = ~\new_[12549]_ ;
  assign \new_[4646]_  = ~\new_[12549]_ ;
  assign \new_[4647]_  = ~\new_[7186]_  | ~\new_[11943]_ ;
  assign \new_[4648]_  = \new_[12683]_  & \new_[12665]_ ;
  assign \new_[4649]_  = ~\new_[6267]_  & ~\new_[9861]_ ;
  assign \new_[4650]_  = ~\new_[7628]_  | ~\new_[12682]_  | ~\new_[7648]_ ;
  assign \new_[4651]_  = ~\new_[6267]_  & ~\new_[10258]_ ;
  assign \new_[4652]_  = \new_[12690]_  & \new_[10265]_ ;
  assign \new_[4653]_  = ~\new_[7631]_  | ~\new_[12679]_  | ~\new_[7766]_ ;
  assign \new_[4654]_  = \new_[5619]_  | \new_[12735]_ ;
  assign \new_[4655]_  = ~\new_[7630]_  | ~\new_[12682]_  | ~\new_[7482]_ ;
  assign \new_[4656]_  = ~\new_[12688]_  | ~\new_[9912]_ ;
  assign \new_[4657]_  = ~\new_[12692]_  | ~\new_[10053]_ ;
  assign \new_[4658]_  = ~\new_[7630]_  | ~\new_[12679]_  | ~\new_[7484]_ ;
  assign \new_[4659]_  = ~\new_[12692]_  | ~\new_[10046]_ ;
  assign \new_[4660]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7486]_ ;
  assign \new_[4661]_  = ~\new_[12692]_  | ~\new_[9822]_ ;
  assign \new_[4662]_  = ~\new_[7630]_  | ~\new_[12682]_  | ~\new_[7312]_ ;
  assign \new_[4663]_  = ~\new_[12690]_  | ~\new_[9737]_ ;
  assign \new_[4664]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7313]_ ;
  assign \new_[4665]_  = ~\new_[12688]_  | ~\new_[9854]_ ;
  assign \new_[4666]_  = ~\new_[12692]_  | ~\new_[10078]_ ;
  assign \new_[4667]_  = ~\new_[12690]_  | ~\new_[9880]_ ;
  assign \new_[4668]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7767]_ ;
  assign \new_[4669]_  = ~\new_[7664]_  | ~\new_[12679]_  | ~\new_[7658]_ ;
  assign \new_[4670]_  = \new_[6267]_  | \new_[10155]_ ;
  assign \new_[4671]_  = ~\new_[6267]_  & ~\new_[10161]_ ;
  assign \new_[4672]_  = ~\new_[7630]_  | ~\new_[12678]_  | ~\new_[7651]_ ;
  assign \new_[4673]_  = ~\new_[12690]_  | ~\new_[10081]_ ;
  assign \new_[4674]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7491]_ ;
  assign \new_[4675]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7492]_ ;
  assign \new_[4676]_  = ~\new_[12688]_  | ~\new_[10082]_ ;
  assign \new_[4677]_  = ~\new_[6267]_  & ~\new_[9924]_ ;
  assign \new_[4678]_  = ~\new_[7628]_  | ~\new_[12679]_  | ~\new_[7493]_ ;
  assign \new_[4679]_  = ~\new_[6267]_  & ~\new_[9941]_ ;
  assign \new_[4680]_  = ~\new_[12688]_  | ~\new_[9807]_ ;
  assign \new_[4681]_  = ~\new_[7628]_  | ~\new_[12679]_  | ~\new_[7496]_ ;
  assign \new_[4682]_  = ~\new_[7628]_  | ~\new_[12682]_  | ~\new_[7501]_ ;
  assign \new_[4683]_  = ~\new_[6267]_  & ~\new_[9738]_ ;
  assign \new_[4684]_  = ~\new_[7628]_  | ~\new_[12679]_  | ~\new_[7511]_ ;
  assign \new_[4685]_  = ~\new_[6267]_  & ~\new_[9345]_ ;
  assign \new_[4686]_  = ~\new_[6267]_  & ~\new_[9956]_ ;
  assign \new_[4687]_  = ~\new_[6267]_  & ~\new_[10101]_ ;
  assign \new_[4688]_  = ~\new_[6267]_  & ~\new_[9836]_ ;
  assign \new_[4689]_  = ~\new_[6267]_  & ~\new_[9927]_ ;
  assign mc_bg_pad_o = u7_mc_bg_reg;
  assign \new_[4691]_  = u5_susp_sel_r_reg;
  assign \new_[4692]_  = ~\new_[7664]_  | ~\new_[12679]_  | ~\new_[7656]_ ;
  assign \mc_addr_pad_o[22]  = \\u7_mc_addr_reg[22] ;
  assign \mc_addr_pad_o[21]  = \\u7_mc_addr_reg[21] ;
  assign \mc_addr_pad_o[19]  = \\u7_mc_addr_reg[19] ;
  assign \mc_addr_pad_o[20]  = \\u7_mc_addr_reg[20] ;
  assign \mc_addr_pad_o[18]  = \\u7_mc_addr_reg[18] ;
  assign \mc_addr_pad_o[16]  = \\u7_mc_addr_reg[16] ;
  assign \mc_addr_pad_o[15]  = \\u7_mc_addr_reg[15] ;
  assign \new_[4700]_  = ~\new_[12690]_  | ~\new_[10118]_ ;
  assign \new_[4701]_  = ~\new_[6267]_  & ~\new_[9742]_ ;
  assign \new_[4702]_  = ~\new_[12690]_  | ~\new_[9839]_ ;
  assign \new_[4703]_  = ~\new_[4970]_ ;
  assign \new_[4704]_  = ~\new_[7664]_  | ~\new_[12682]_  | ~\new_[7317]_ ;
  assign \new_[4705]_  = ~\new_[6267]_  & ~\new_[9860]_ ;
  assign \new_[4706]_  = \new_[7564]_  & \new_[5637]_ ;
  assign \new_[4707]_  = ~\new_[7664]_  | ~\new_[12679]_  | ~\new_[7659]_ ;
  assign \new_[4708]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7652]_ ;
  assign \new_[4709]_  = ~\new_[4974]_ ;
  assign \new_[4710]_  = ~\new_[6267]_  & ~\new_[9717]_ ;
  assign \new_[4711]_  = ~\new_[7628]_  | ~\new_[12679]_  | ~\new_[7513]_ ;
  assign \new_[4712]_  = ~\new_[12744]_  | ~\new_[9978]_ ;
  assign \new_[4713]_  = ~\new_[12692]_  | ~\new_[9967]_ ;
  assign \new_[4714]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7519]_ ;
  assign \new_[4715]_  = ~\new_[6267]_  & ~\new_[9918]_ ;
  assign \new_[4716]_  = ~\new_[6267]_  & ~\new_[9905]_ ;
  assign \new_[4717]_  = ~\new_[7628]_  | ~\new_[12678]_  | ~\new_[7515]_ ;
  assign \new_[4718]_  = ~\new_[7663]_  | ~\new_[12685]_  | ~\new_[7480]_ ;
  assign \new_[4719]_  = ~\new_[6267]_  & ~\new_[9714]_ ;
  assign \new_[4720]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7318]_ ;
  assign \new_[4721]_  = ~\new_[7631]_  | ~\new_[12685]_  | ~\new_[7504]_ ;
  assign \new_[4722]_  = ~\new_[6267]_  & ~\new_[9859]_ ;
  assign \new_[4723]_  = ~\new_[7631]_  | ~\new_[12678]_  | ~\new_[7320]_ ;
  assign \new_[4724]_  = ~\new_[12692]_  | ~\new_[10050]_ ;
  assign \new_[4725]_  = ~\new_[7663]_  | ~\new_[12678]_  | ~\new_[7518]_ ;
  assign \new_[4726]_  = ~\new_[6267]_  & ~\new_[9739]_ ;
  assign \new_[4727]_  = ~\new_[7628]_  | ~\new_[12682]_  | ~\new_[7505]_ ;
  assign \new_[4728]_  = ~\new_[6267]_  & (~\new_[1433]_  | ~\new_[10767]_ );
  assign \new_[4729]_  = ~\new_[6267]_  & ~\new_[9899]_ ;
  assign \new_[4730]_  = ~\new_[4989]_ ;
  assign \new_[4731]_  = ~\new_[6267]_  & ~\new_[10166]_ ;
  assign \new_[4732]_  = ~\new_[12692]_  | ~\new_[10107]_ ;
  assign \new_[4733]_  = ~\new_[7628]_  | ~\new_[12678]_  | ~\new_[7647]_ ;
  assign \new_[4734]_  = ~\new_[11558]_  & ~\new_[11263]_ ;
  assign \new_[4735]_  = ~\new_[10759]_  & (~\new_[7364]_  | ~\new_[6038]_ );
  assign \new_[4736]_  = ~\new_[10691]_  & (~\new_[6319]_  | ~\new_[6039]_ );
  assign \new_[4737]_  = ~\new_[6012]_  | ~\new_[5647]_ ;
  assign \new_[4738]_  = (~\new_[6035]_  | ~\wb_addr_i[12] ) & (~\new_[11725]_  | ~\wb_addr_i[10] );
  assign \new_[4739]_  = (~\new_[6035]_  | ~\wb_addr_i[13] ) & (~\new_[11725]_  | ~\wb_addr_i[11] );
  assign \new_[4740]_  = ~\new_[5020]_ ;
  assign \new_[4741]_  = (~\new_[6035]_  | ~\wb_addr_i[14] ) & (~\new_[11725]_  | ~\wb_addr_i[12] );
  assign \new_[4742]_  = ~\new_[5021]_ ;
  assign \new_[4743]_  = (~\new_[6035]_  | ~\wb_addr_i[22] ) & (~\new_[11725]_  | ~\wb_addr_i[20] );
  assign \new_[4744]_  = (~\new_[6035]_  | ~\wb_addr_i[23] ) & (~\new_[11725]_  | ~\wb_addr_i[21] );
  assign \new_[4745]_  = (~\new_[6035]_  | ~\wb_addr_i[15] ) & (~\new_[11725]_  | ~\wb_addr_i[13] );
  assign \new_[4746]_  = (~\new_[6035]_  | ~\wb_addr_i[16] ) & (~\new_[11725]_  | ~\wb_addr_i[14] );
  assign \new_[4747]_  = (~\new_[6035]_  | ~\wb_addr_i[17] ) & (~\new_[11725]_  | ~\wb_addr_i[15] );
  assign \new_[4748]_  = (~\new_[6035]_  | ~\wb_addr_i[18] ) & (~\new_[11725]_  | ~\wb_addr_i[16] );
  assign \new_[4749]_  = (~\new_[6035]_  | ~\wb_addr_i[20] ) & (~\new_[11725]_  | ~\wb_addr_i[18] );
  assign \new_[4750]_  = (~\new_[6035]_  | ~\wb_addr_i[21] ) & (~\new_[11725]_  | ~\wb_addr_i[19] );
  assign \new_[4751]_  = (~\new_[6035]_  | ~\wb_addr_i[19] ) & (~\new_[11725]_  | ~\wb_addr_i[17] );
  assign \new_[4752]_  = ~\new_[5631]_  | (~\new_[12778]_  & ~\new_[10150]_ );
  assign \new_[4753]_  = \new_[6286]_  & \new_[5644]_ ;
  assign \new_[4754]_  = (~\new_[5780]_  | ~\new_[11560]_ ) & (~\new_[12533]_  | ~\new_[1643]_ );
  assign \new_[4755]_  = \new_[10522]_  ? \new_[11062]_  : \new_[5712]_ ;
  assign \new_[4756]_  = ~\new_[5792]_  | ~\new_[7476]_  | ~\new_[6274]_ ;
  assign \new_[4757]_  = ~\new_[5793]_  | ~\new_[7477]_  | ~\new_[6275]_ ;
  assign \new_[4758]_  = ~\new_[5249]_ ;
  assign \new_[4759]_  = ~\new_[10200]_  | (~\new_[5765]_  & ~\new_[6723]_ );
  assign \new_[4760]_  = ~\new_[5349]_  & (~\new_[7226]_  | ~\new_[9979]_ );
  assign \new_[4761]_  = ~\new_[5351]_  & (~\new_[7226]_  | ~\new_[11772]_ );
  assign \new_[4762]_  = ~\new_[5352]_  & (~\new_[7226]_  | ~\new_[9418]_ );
  assign \new_[4763]_  = ~\new_[5353]_  & (~\new_[7226]_  | ~\new_[9340]_ );
  assign \new_[4764]_  = ~\new_[5355]_  & (~\new_[7226]_  | ~\new_[9618]_ );
  assign \new_[4765]_  = ~\new_[5356]_  & (~\new_[7226]_  | ~\new_[9682]_ );
  assign \new_[4766]_  = ~\new_[5357]_  & (~\new_[7226]_  | ~\new_[9980]_ );
  assign \new_[4767]_  = ~\new_[5362]_  & (~\new_[7226]_  | ~\new_[9567]_ );
  assign \new_[4768]_  = ~\new_[5359]_  & (~\new_[7226]_  | ~\new_[9707]_ );
  assign \new_[4769]_  = ~\new_[5360]_  & (~\new_[7226]_  | ~\new_[9389]_ );
  assign \new_[4770]_  = ~\new_[5361]_  & (~\new_[7226]_  | ~\new_[9665]_ );
  assign \new_[4771]_  = ~\new_[5363]_  & (~\new_[7226]_  | ~\new_[10136]_ );
  assign \new_[4772]_  = ~\new_[7130]_  | ~\new_[5620]_  | ~\new_[6675]_ ;
  assign \new_[4773]_  = ~\new_[5301]_  & (~\new_[11976]_  | ~\new_[12000]_ );
  assign \new_[4774]_  = ~\new_[5302]_  & (~\new_[11976]_  | ~\new_[10102]_ );
  assign \new_[4775]_  = ~\new_[5303]_  & (~\new_[11976]_  | ~\new_[9584]_ );
  assign \new_[4776]_  = ~\new_[5304]_  & (~\new_[11976]_  | ~\new_[9587]_ );
  assign \new_[4777]_  = ~\new_[5305]_  & (~\new_[11976]_  | ~\new_[9588]_ );
  assign \new_[4778]_  = ~\new_[5306]_  & (~\new_[11976]_  | ~\new_[9933]_ );
  assign \new_[4779]_  = ~\new_[5307]_  & (~\new_[11976]_  | ~\new_[9592]_ );
  assign \new_[4780]_  = ~\new_[5309]_  & (~\new_[11976]_  | ~\new_[9929]_ );
  assign \new_[4781]_  = ~\new_[5310]_  & (~\new_[7873]_  | ~\new_[9960]_ );
  assign \new_[4782]_  = ~\new_[5311]_  & (~\new_[11976]_  | ~\new_[9612]_ );
  assign \new_[4783]_  = ~\new_[5312]_  & (~\new_[11976]_  | ~\new_[9603]_ );
  assign \new_[4784]_  = ~\new_[5313]_  & (~\new_[11976]_  | ~\new_[9842]_ );
  assign \new_[4785]_  = ~\new_[5315]_  & (~\new_[11976]_  | ~\new_[9678]_ );
  assign \new_[4786]_  = ~\new_[5316]_  & (~\new_[11976]_  | ~\new_[10040]_ );
  assign \new_[4787]_  = ~\new_[5317]_  & (~\new_[11976]_  | ~\new_[9489]_ );
  assign \new_[4788]_  = ~\new_[5318]_  & (~\new_[11976]_  | ~\new_[9593]_ );
  assign \new_[4789]_  = ~\new_[5319]_  & (~\new_[11976]_  | ~\new_[9621]_ );
  assign \new_[4790]_  = ~\new_[5320]_  & (~\new_[11976]_  | ~\new_[9615]_ );
  assign \new_[4791]_  = ~\new_[5321]_  & (~\new_[11976]_  | ~\new_[9601]_ );
  assign \new_[4792]_  = ~\new_[5322]_  & (~\new_[11976]_  | ~\new_[9585]_ );
  assign \new_[4793]_  = ~\new_[5323]_  & (~\new_[11976]_  | ~\new_[9602]_ );
  assign \new_[4794]_  = ~\new_[5324]_  & (~\new_[11976]_  | ~\new_[9855]_ );
  assign \new_[4795]_  = ~\new_[5325]_  & (~\new_[11976]_  | ~\new_[9598]_ );
  assign \new_[4796]_  = ~\new_[5326]_  & (~\new_[11976]_  | ~\new_[9837]_ );
  assign \new_[4797]_  = ~\new_[5327]_  & (~\new_[11976]_  | ~\new_[9614]_ );
  assign \new_[4798]_  = ~\new_[5328]_  & (~\new_[11976]_  | ~\new_[9586]_ );
  assign \new_[4799]_  = ~\new_[5330]_  & (~\new_[11976]_  | ~\new_[9589]_ );
  assign \new_[4800]_  = ~\new_[5331]_  & (~\new_[11976]_  | ~\new_[9857]_ );
  assign \new_[4801]_  = ~\new_[5332]_  & (~\new_[11976]_  | ~\new_[9663]_ );
  assign \new_[4802]_  = ~\new_[5333]_  & (~\new_[11976]_  | ~\new_[9613]_ );
  assign \new_[4803]_  = ~\new_[5334]_  & (~\new_[11976]_  | ~\new_[9581]_ );
  assign \new_[4804]_  = ~\new_[5335]_  & (~\new_[11976]_  | ~\new_[9609]_ );
  assign \new_[4805]_  = ~\new_[5336]_  & (~\new_[11976]_  | ~\new_[9862]_ );
  assign \new_[4806]_  = ~\new_[5337]_  & (~\new_[11976]_  | ~\new_[9840]_ );
  assign \new_[4807]_  = ~\new_[5338]_  & (~\new_[11976]_  | ~\new_[10062]_ );
  assign \new_[4808]_  = ~\new_[5339]_  & (~\new_[11976]_  | ~\new_[9408]_ );
  assign \new_[4809]_  = \new_[6642]_  | \new_[5748]_ ;
  assign \new_[4810]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10485]_ ) | (~\new_[12710]_  & ~\new_[12672]_  & ~\new_[10485]_ );
  assign \new_[4811]_  = (~\new_[12651]_  & ~\new_[8408]_  & ~\new_[11299]_ ) | (~\new_[12704]_  & ~\new_[12672]_  & ~\new_[11299]_ );
  assign \new_[4812]_  = \new_[5800]_  | \new_[7109]_ ;
  assign \new_[4813]_  = \new_[5802]_  & \new_[12486]_ ;
  assign \new_[4814]_  = (~\new_[12650]_  & ~\new_[8408]_  & ~\new_[12599]_ ) | (~\new_[12714]_  & ~\new_[12672]_  & ~\new_[12599]_ );
  assign \new_[4815]_  = ~\new_[5818]_  & ~\new_[6997]_ ;
  assign \new_[4816]_  = ~\new_[5701]_  | ~\new_[12469]_ ;
  assign \new_[4817]_  = (~\new_[12651]_  & ~\new_[8408]_  & ~\new_[12045]_ ) | (~\new_[12710]_  & ~\new_[12672]_  & ~\new_[12045]_ );
  assign \new_[4818]_  = ~\new_[5786]_  & (~\new_[7226]_  | ~\new_[10128]_ );
  assign \new_[4819]_  = ~\new_[5358]_ ;
  assign \new_[4820]_  = (~\new_[12654]_  & ~\new_[8408]_  & ~\new_[10551]_ ) | (~\new_[7862]_  & ~\new_[7297]_  & ~\new_[12654]_ );
  assign \new_[4821]_  = ~\new_[5819]_  & (~\new_[6384]_  | ~\new_[10039]_ );
  assign \new_[4822]_  = ~\new_[5821]_  & (~\new_[6384]_  | ~\new_[12110]_ );
  assign \new_[4823]_  = ~\new_[8192]_  | ~\new_[7426]_  | ~\new_[6733]_  | ~\new_[6738]_ ;
  assign \new_[4824]_  = ~\new_[5751]_  & (~\new_[7226]_  | ~\new_[9388]_ );
  assign \new_[4825]_  = (~\new_[6041]_  | ~\wb_addr_i[10] ) & (~\new_[11715]_  | ~\wb_addr_i[11] );
  assign \new_[4826]_  = (~\new_[6041]_  | ~\wb_addr_i[11] ) & (~\new_[11715]_  | ~\wb_addr_i[12] );
  assign \new_[4827]_  = (~\new_[6041]_  | ~\wb_addr_i[12] ) & (~\new_[11715]_  | ~\wb_addr_i[13] );
  assign \new_[4828]_  = (~\new_[6041]_  | ~\wb_addr_i[20] ) & (~\new_[11715]_  | ~\wb_addr_i[21] );
  assign \new_[4829]_  = (~\new_[6041]_  | ~\wb_addr_i[13] ) & (~\new_[11715]_  | ~\wb_addr_i[14] );
  assign \new_[4830]_  = (~\new_[6041]_  | ~\wb_addr_i[14] ) & (~\new_[11715]_  | ~\wb_addr_i[15] );
  assign \new_[4831]_  = (~\new_[6041]_  | ~\wb_addr_i[15] ) & (~\new_[11715]_  | ~\wb_addr_i[16] );
  assign \new_[4832]_  = (~\new_[6041]_  | ~\wb_addr_i[16] ) & (~\new_[11715]_  | ~\wb_addr_i[17] );
  assign \new_[4833]_  = (~\new_[6041]_  | ~\wb_addr_i[17] ) & (~\new_[11715]_  | ~\wb_addr_i[18] );
  assign \new_[4834]_  = (~\new_[6041]_  | ~\wb_addr_i[18] ) & (~\new_[11715]_  | ~\wb_addr_i[19] );
  assign \new_[4835]_  = (~\new_[6041]_  | ~\wb_addr_i[19] ) & (~\new_[11715]_  | ~\wb_addr_i[20] );
  assign \new_[4836]_  = ~\new_[5982]_  | ~\new_[6099]_ ;
  assign \new_[4837]_  = ~\new_[6032]_  | ~\new_[6100]_ ;
  assign \new_[4838]_  = ~\new_[7189]_  | ~\new_[5773]_ ;
  assign \new_[4839]_  = \new_[11102]_  ^ \new_[6107]_ ;
  assign \new_[4840]_  = ~\new_[7182]_  | ~\new_[5833]_ ;
  assign \new_[4841]_  = ~\new_[5865]_  | ~\new_[10136]_ ;
  assign \new_[4842]_  = ~\new_[5865]_  | ~\new_[9567]_ ;
  assign \new_[4843]_  = ~\new_[5865]_  | ~\new_[9979]_ ;
  assign \new_[4844]_  = (~\new_[7131]_  & ~\new_[11348]_  & ~\new_[10722]_ ) | (~\new_[11327]_  & ~\new_[6636]_  & ~\new_[11348]_ );
  assign \new_[4845]_  = ~\new_[5865]_  | ~\new_[9401]_ ;
  assign \new_[4846]_  = ~\new_[5865]_  | ~\new_[10099]_ ;
  assign \new_[4847]_  = ~\new_[5865]_  | ~\new_[10104]_ ;
  assign \new_[4848]_  = ~\new_[5865]_  | ~\new_[10128]_ ;
  assign \new_[4849]_  = ~\new_[5865]_  | ~\new_[8805]_ ;
  assign \new_[4850]_  = ~\new_[5865]_  | ~\new_[10011]_ ;
  assign \new_[4851]_  = ~\new_[5865]_  | ~\new_[9680]_ ;
  assign \new_[4852]_  = ~\new_[5865]_  | ~\new_[10263]_ ;
  assign \new_[4853]_  = ~\new_[5865]_  | ~\new_[9995]_ ;
  assign \new_[4854]_  = ~\new_[5865]_  | ~\new_[9845]_ ;
  assign \new_[4855]_  = ~\new_[5865]_  | ~\new_[10237]_ ;
  assign \new_[4856]_  = ~\new_[5865]_  | ~\new_[9660]_ ;
  assign \new_[4857]_  = ~\new_[5865]_  | ~\new_[9641]_ ;
  assign \new_[4858]_  = ~\new_[5865]_  | ~\new_[10052]_ ;
  assign \new_[4859]_  = ~\new_[5865]_  | ~\new_[9340]_ ;
  assign \new_[4860]_  = ~\new_[5865]_  | ~\new_[9958]_ ;
  assign \new_[4861]_  = \new_[6555]_  & \new_[5885]_ ;
  assign \new_[4862]_  = ~\new_[5865]_  | ~\new_[9611]_ ;
  assign \new_[4863]_  = \new_[6556]_  & \new_[5886]_ ;
  assign \new_[4864]_  = ~\new_[5865]_  | ~\new_[9853]_ ;
  assign \new_[4865]_  = \new_[6557]_  & \new_[5887]_ ;
  assign \new_[4866]_  = ~\new_[5865]_  | ~\new_[9582]_ ;
  assign \new_[4867]_  = ~\new_[5865]_  | ~\new_[9104]_ ;
  assign \new_[4868]_  = ~\new_[5865]_  | ~\new_[10019]_ ;
  assign \new_[4869]_  = \new_[5954]_  & \new_[5894]_ ;
  assign \new_[4870]_  = \new_[6560]_  & \new_[5895]_ ;
  assign \new_[4871]_  = ~\new_[5865]_  | ~\new_[9682]_ ;
  assign \new_[4872]_  = ~\new_[5865]_  | ~\new_[9595]_ ;
  assign \new_[4873]_  = ~\new_[5865]_  | ~\new_[9374]_ ;
  assign \new_[4874]_  = \new_[6563]_  & \new_[5897]_ ;
  assign \new_[4875]_  = ~\new_[5865]_  | ~\new_[9675]_ ;
  assign \new_[4876]_  = \new_[6565]_  & \new_[5900]_ ;
  assign \new_[4877]_  = ~\new_[5865]_  | ~\new_[9709]_ ;
  assign \new_[4878]_  = \new_[6566]_  & \new_[5901]_ ;
  assign \new_[4879]_  = ~\new_[5865]_  | ~\new_[9599]_ ;
  assign \new_[4880]_  = \new_[6568]_  & \new_[5903]_ ;
  assign \new_[4881]_  = \new_[6197]_  & \new_[5892]_ ;
  assign \new_[4882]_  = ~\new_[6280]_  | ~\new_[6198]_  | ~\new_[6731]_ ;
  assign \new_[4883]_  = ~\new_[5865]_  | ~\new_[10137]_ ;
  assign \new_[4884]_  = \new_[6199]_  & \new_[5906]_ ;
  assign \new_[4885]_  = ~\new_[5865]_  | ~\new_[9665]_ ;
  assign \new_[4886]_  = ~\new_[6281]_  | ~\new_[6200]_  | ~\new_[6732]_ ;
  assign \new_[4887]_  = ~\new_[5865]_  | ~\new_[9407]_ ;
  assign \new_[4888]_  = ~\new_[7445]_  | (~\new_[6284]_  & ~\new_[12003]_ );
  assign \new_[4889]_  = (~\new_[6747]_  | ~\new_[7825]_ ) & (~\new_[11306]_  | ~\new_[7483]_ );
  assign \new_[4890]_  = (~\new_[6748]_  | ~\new_[7776]_ ) & (~\new_[11305]_  | ~\new_[7311]_ );
  assign \new_[4891]_  = (~\new_[6752]_  | ~\new_[7776]_ ) & (~\new_[11305]_  | ~\new_[7313]_ );
  assign \new_[4892]_  = (~\new_[6756]_  | ~\new_[7776]_ ) & (~\new_[11303]_  | ~\new_[7489]_ );
  assign \new_[4893]_  = ~\new_[11484]_  | (~\new_[6283]_  & ~\new_[10057]_ );
  assign \new_[4894]_  = (~\new_[6769]_  | ~\new_[7776]_ ) & (~\new_[11304]_  | ~\new_[7480]_ );
  assign \new_[4895]_  = ~\new_[5876]_  | ~\new_[9604]_ ;
  assign \new_[4896]_  = (~\new_[6775]_  | ~\new_[7776]_ ) & (~\new_[11305]_  | ~\new_[7512]_ );
  assign \new_[4897]_  = (~\new_[6761]_  | ~\new_[7776]_ ) & (~\new_[11303]_  | ~\new_[7322]_ );
  assign \new_[4898]_  = ~\new_[5909]_  & (~\new_[7329]_  | ~\new_[10115]_ );
  assign \new_[4899]_  = ~\new_[5869]_  & (~\new_[3881]_  | ~\new_[6621]_ );
  assign \new_[4900]_  = ~\new_[5870]_  & (~\new_[11033]_  | ~\new_[6621]_ );
  assign \new_[4901]_  = ~\new_[6246]_  | (~\new_[12745]_  & ~\new_[9860]_ );
  assign \new_[4902]_  = ~\new_[5986]_  | (~\new_[12738]_  & ~\new_[9924]_ );
  assign \new_[4903]_  = ~\new_[11499]_  | (~\new_[6267]_  & ~\new_[9617]_ );
  assign \new_[4904]_  = ~\new_[6968]_  | (~\new_[6267]_  & ~\new_[11865]_ );
  assign \new_[4905]_  = ~\new_[6234]_  | (~\new_[12742]_  & ~\new_[9345]_ );
  assign \new_[4906]_  = ~\new_[6235]_  | (~\new_[12743]_  & ~\new_[9691]_ );
  assign \new_[4907]_  = ~\new_[6239]_  | (~\new_[12742]_  & ~\new_[9954]_ );
  assign \new_[4908]_  = ~\new_[6242]_  | (~\new_[12738]_  & ~\new_[9177]_ );
  assign \new_[4909]_  = ~\new_[5991]_  | (~\new_[12738]_  & ~\new_[9742]_ );
  assign \new_[4910]_  = ~\new_[5999]_  | (~\new_[12745]_  & ~\new_[9717]_ );
  assign \new_[4911]_  = ~\new_[6001]_  | (~\new_[12738]_  & ~\new_[9623]_ );
  assign \new_[4912]_  = ~\new_[6000]_  | (~\new_[12738]_  & ~\new_[9918]_ );
  assign \new_[4913]_  = ~\new_[6252]_  | (~\new_[12738]_  & ~\new_[9905]_ );
  assign \new_[4914]_  = ~\new_[6240]_  | (~\new_[12746]_  & ~\new_[9714]_ );
  assign \new_[4915]_  = ~\new_[6238]_  | (~\new_[12746]_  & ~\new_[9859]_ );
  assign \new_[4916]_  = ~\new_[6259]_  | (~\new_[12738]_  & ~\new_[9955]_ );
  assign \new_[4917]_  = ~\new_[6004]_  | (~\new_[12738]_  & ~\new_[9911]_ );
  assign \new_[4918]_  = ~\new_[6261]_  | (~\new_[12738]_  & ~\new_[9739]_ );
  assign \new_[4919]_  = ~\new_[5992]_  | (~\new_[12738]_  & ~\new_[9713]_ );
  assign \new_[4920]_  = ~\new_[6971]_  | (~\new_[6267]_  & ~\new_[12113]_ );
  assign \new_[4921]_  = ~\new_[5979]_  | (~\new_[12742]_  & ~\new_[9899]_ );
  assign \new_[4922]_  = ~\new_[5430]_ ;
  assign \new_[4923]_  = ~\new_[6024]_  | (~\new_[12070]_  & ~\new_[10172]_ );
  assign \new_[4924]_  = ~\new_[6025]_  | (~\new_[12070]_  & ~\new_[9911]_ );
  assign \new_[4925]_  = \new_[6027]_  | \new_[7863]_ ;
  assign \new_[4926]_  = ~\new_[12549]_ ;
  assign \new_[4927]_  = ~u5_pack_le0_reg;
  assign \new_[4928]_  = ~\new_[7628]_  | ~\new_[12679]_  | ~\new_[7481]_ ;
  assign \new_[4929]_  = ~\new_[12738]_  & (~\new_[10517]_  | ~\new_[10747]_ );
  assign \new_[4930]_  = ~\new_[6640]_  & ~\new_[9718]_ ;
  assign \new_[4931]_  = ~\new_[6267]_  & ~\new_[9718]_ ;
  assign \new_[4932]_  = ~\new_[7664]_  | ~\new_[12678]_  | ~\new_[7650]_ ;
  assign \new_[4933]_  = \new_[5977]_  | \new_[10348]_ ;
  assign \new_[4934]_  = ~\new_[6640]_  & ~\new_[10229]_ ;
  assign \new_[4935]_  = ~\new_[6267]_  & ~\new_[10229]_ ;
  assign \new_[4936]_  = ~\new_[6640]_  & ~\new_[9867]_ ;
  assign \new_[4937]_  = ~\new_[6267]_  & ~\new_[9867]_ ;
  assign \new_[4938]_  = ~\new_[6640]_  & ~\new_[10146]_ ;
  assign \new_[4939]_  = ~\new_[6267]_  & ~\new_[10146]_ ;
  assign \new_[4940]_  = ~\new_[6267]_  & ~\new_[10234]_ ;
  assign \new_[4941]_  = ~\new_[6640]_  & ~\new_[10256]_ ;
  assign \new_[4942]_  = ~\new_[6267]_  & ~\new_[10256]_ ;
  assign \new_[4943]_  = ~\new_[6267]_  & ~\new_[9894]_ ;
  assign \new_[4944]_  = ~\new_[6640]_  & ~\new_[9922]_ ;
  assign \new_[4945]_  = ~\new_[6267]_  & ~\new_[9922]_ ;
  assign \new_[4946]_  = ~\new_[6267]_  & ~\new_[9838]_ ;
  assign \new_[4947]_  = ~\new_[6640]_  & (~\new_[1433]_  | ~\new_[11344]_ );
  assign \new_[4948]_  = ~\new_[12741]_  & ~\new_[10340]_ ;
  assign \new_[4949]_  = ~\new_[6267]_  & ~\new_[10340]_ ;
  assign \new_[4950]_  = ~\new_[12690]_  | ~\new_[9848]_ ;
  assign \new_[4951]_  = \new_[6641]_  | \new_[10101]_ ;
  assign \new_[4952]_  = ~\new_[6640]_  & ~\new_[10254]_ ;
  assign \new_[4953]_  = ~\new_[6267]_  & ~\new_[10254]_ ;
  assign \new_[4954]_  = ~\new_[7628]_  | ~\new_[12679]_  | ~\new_[7490]_ ;
  assign \new_[4955]_  = ~\new_[6267]_  & ~\new_[9908]_ ;
  assign \new_[4956]_  = ~\new_[6267]_  & ~\new_[9866]_ ;
  assign \new_[4957]_  = ~\new_[12690]_  | ~\new_[11504]_ ;
  assign \new_[4958]_  = ~\new_[6640]_  & ~\new_[10262]_ ;
  assign \new_[4959]_  = ~\new_[6267]_  & ~\new_[10262]_ ;
  assign \new_[4960]_  = \new_[6026]_  | \new_[7863]_ ;
  assign n2196 = ~\new_[11845]_  | ~\new_[12725]_  | ~\new_[12322]_ ;
  assign \new_[4962]_  = ~\new_[12690]_  | ~\new_[10045]_ ;
  assign \new_[4963]_  = ~\new_[7628]_  | ~\new_[12681]_  | ~\new_[7653]_ ;
  assign \new_[4964]_  = \new_[6641]_  | \new_[9345]_ ;
  assign \new_[4965]_  = \new_[6641]_  | \new_[9691]_ ;
  assign \new_[4966]_  = \new_[6641]_  | \new_[9927]_ ;
  assign \new_[4967]_  = ~\new_[6267]_  & ~\new_[10255]_ ;
  assign \new_[4968]_  = ~\new_[5475]_ ;
  assign mc_adv_pad_o_ = u7_mc_adv__reg;
  assign \new_[4970]_  = ~\new_[12652]_  | ~\new_[12738]_ ;
  assign \new_[4971]_  = ~\new_[6641]_  & ~\new_[9860]_ ;
  assign \new_[4972]_  = \new_[6640]_  | \new_[10167]_ ;
  assign \new_[4973]_  = ~\new_[6640]_  & ~\new_[9743]_ ;
  assign \new_[4974]_  = ~\new_[7180]_  & ~\new_[5977]_ ;
  assign \new_[4975]_  = ~\new_[6268]_  | ~\new_[5977]_ ;
  assign \new_[4976]_  = ~\new_[12679]_  | ~\new_[7418]_ ;
  assign \new_[4977]_  = ~\new_[6267]_  & ~\new_[9925]_ ;
  assign \new_[4978]_  = \new_[6641]_  | \new_[10172]_ ;
  assign \new_[4979]_  = ~\new_[12690]_  | ~\new_[10127]_ ;
  assign n2236 = ~\new_[11410]_  | ~\new_[9986]_  | ~\new_[6065]_ ;
  assign \new_[4981]_  = ~\new_[6267]_  & ~\new_[9921]_ ;
  assign \new_[4982]_  = ~\new_[6640]_  & ~\new_[9925]_ ;
  assign \new_[4983]_  = ~\new_[12741]_  & ~\new_[10167]_ ;
  assign \new_[4984]_  = \new_[6641]_  | \new_[9899]_ ;
  assign \new_[4985]_  = \new_[6641]_  | \new_[9713]_ ;
  assign n2241 = ~\new_[12507]_  & (~\new_[6066]_  | ~\new_[6068]_ );
  assign n2191 = ~\new_[12507]_  & (~\new_[6067]_  | ~\new_[6069]_ );
  assign \new_[4988]_  = ~\new_[6640]_  & ~\new_[9732]_ ;
  assign \new_[4989]_  = \new_[5977]_  & \new_[10754]_ ;
  assign \new_[4990]_  = ~\new_[6267]_  & ~\new_[9732]_ ;
  assign \new_[4991]_  = ~\new_[6640]_  & ~\new_[10199]_ ;
  assign \new_[4992]_  = \new_[5977]_  & \new_[10919]_ ;
  assign \new_[4993]_  = ~\new_[6267]_  & ~\new_[10199]_ ;
  assign \new_[4994]_  = \new_[10325]_  | \new_[7992]_  | \new_[11278]_  | \new_[7302]_ ;
  assign \new_[4995]_  = \new_[10259]_  & \new_[6008]_ ;
  assign \new_[4996]_  = ~\new_[10691]_  & (~\new_[6040]_  | ~\new_[6295]_ );
  assign \new_[4997]_  = ~\new_[10691]_  & (~\new_[6047]_  | ~\new_[6298]_ );
  assign \new_[4998]_  = ~\new_[10691]_  & (~\new_[6060]_  | ~\new_[6299]_ );
  assign \new_[4999]_  = ~\new_[10759]_  & (~\new_[6048]_  | ~\new_[6314]_ );
  assign \new_[5000]_  = ~\new_[10759]_  & (~\new_[6049]_  | ~\new_[6300]_ );
  assign \new_[5001]_  = ~\new_[10759]_  & (~\new_[6051]_  | ~\new_[6301]_ );
  assign \new_[5002]_  = ~\new_[10691]_  & (~\new_[6050]_  | ~\new_[6296]_ );
  assign \new_[5003]_  = ~\new_[10691]_  & (~\new_[6046]_  | ~\new_[6302]_ );
  assign \new_[5004]_  = ~\new_[10691]_  & (~\new_[6057]_  | ~\new_[6303]_ );
  assign \new_[5005]_  = ~\new_[10759]_  & (~\new_[6052]_  | ~\new_[6297]_ );
  assign \new_[5006]_  = ~\new_[10759]_  & (~\new_[6053]_  | ~\new_[6304]_ );
  assign \new_[5007]_  = ~\new_[10759]_  & (~\new_[6054]_  | ~\new_[6306]_ );
  assign \new_[5008]_  = ~\new_[10759]_  & (~\new_[6055]_  | ~\new_[6307]_ );
  assign \new_[5009]_  = ~\new_[10691]_  & (~\new_[6056]_  | ~\new_[6311]_ );
  assign \new_[5010]_  = ~\new_[10691]_  & (~\new_[6045]_  | ~\new_[6294]_ );
  assign \new_[5011]_  = ~\new_[10691]_  & (~\new_[6058]_  | ~\new_[6308]_ );
  assign \new_[5012]_  = ~\new_[10691]_  & (~\new_[6042]_  | ~\new_[6293]_ );
  assign \new_[5013]_  = ~\new_[10691]_  & (~\new_[6044]_  | ~\new_[6309]_ );
  assign \new_[5014]_  = ~\new_[10759]_  & (~\new_[6043]_  | ~\new_[6310]_ );
  assign \new_[5015]_  = ~\new_[10691]_  & (~\new_[6062]_  | ~\new_[6313]_ );
  assign \new_[5016]_  = ~\new_[10759]_  & (~\new_[6059]_  | ~\new_[6312]_ );
  assign \new_[5017]_  = (~\new_[12307]_  | ~\new_[9591]_ ) & (~\new_[12747]_  | ~\new_[12060]_ );
  assign \new_[5018]_  = (~\new_[6290]_  | ~\wb_addr_i[24] ) & (~\new_[6666]_  | ~\wb_addr_i[23] );
  assign \new_[5019]_  = ~\new_[11298]_  | ~\new_[6029]_  | ~\new_[11317]_ ;
  assign \new_[5020]_  = (~\new_[6291]_  | ~\wb_addr_i[26] ) & (~\new_[11716]_  | ~\wb_addr_i[25] );
  assign \new_[5021]_  = (~\new_[6291]_  | ~\wb_addr_i[24] ) & (~\new_[11716]_  | ~\wb_addr_i[23] );
  assign \new_[5022]_  = ~\new_[6009]_  | (~\new_[6320]_  & ~\new_[9096]_ );
  assign \new_[5023]_  = (~\new_[12783]_  | ~\new_[12000]_ ) & (~\new_[7344]_  | ~\new_[9383]_ );
  assign \new_[5024]_  = (~\new_[12784]_  | ~\new_[11973]_ ) & (~\new_[7344]_  | ~\new_[10115]_ );
  assign \new_[5025]_  = ~\new_[6010]_  | (~\new_[6320]_  & ~\new_[9322]_ );
  assign \new_[5026]_  = \new_[3398]_  ? \new_[6071]_  : \new_[10416]_ ;
  assign \new_[5027]_  = (~\new_[12783]_  | ~\new_[9938]_ ) & (~\new_[7344]_  | ~\new_[10031]_ );
  assign \new_[5028]_  = (~\new_[6086]_  | ~\new_[9998]_ ) & (~\new_[12775]_  | ~\new_[9979]_ );
  assign \new_[5029]_  = (~\new_[6088]_  | ~\new_[12273]_ ) & (~\new_[7008]_  | ~\new_[10265]_ );
  assign \new_[5030]_  = (~\new_[7059]_  | ~\new_[9912]_ ) & (~\new_[11553]_  | ~\new_[8871]_ );
  assign \new_[5031]_  = (~\new_[6090]_  | ~\new_[10928]_ ) & (~\new_[12775]_  | ~\new_[9963]_ );
  assign \new_[5032]_  = (~\new_[6089]_  | ~\new_[9647]_ ) & (~\new_[12777]_  | ~\new_[9607]_ );
  assign \new_[5033]_  = (~\new_[6088]_  | ~\new_[11331]_ ) & (~\new_[12768]_  | ~\new_[10011]_ );
  assign \new_[5034]_  = (~\new_[6088]_  | ~\new_[10177]_ ) & (~\new_[12771]_  | ~\new_[9680]_ );
  assign \new_[5035]_  = (~\new_[6090]_  | ~\new_[11343]_ ) & (~\new_[12776]_  | ~\new_[10263]_ );
  assign \new_[5036]_  = (~\new_[7059]_  | ~\new_[9737]_ ) & (~\new_[11553]_  | ~\new_[9099]_ );
  assign \new_[5037]_  = (~\new_[6088]_  | ~\new_[10808]_ ) & (~\new_[12775]_  | ~\new_[9995]_ );
  assign \new_[5038]_  = (~\new_[6089]_  | ~\new_[10818]_ ) & (~\new_[12775]_  | ~\new_[9627]_ );
  assign \new_[5039]_  = (~\new_[6087]_  | ~\new_[11320]_ ) & (~\new_[12768]_  | ~\new_[9660]_ );
  assign \new_[5040]_  = (~\new_[12784]_  | ~\new_[9612]_ ) & (~\new_[7239]_  | ~\new_[9680]_ );
  assign \new_[5041]_  = (~\new_[6088]_  | ~\new_[10938]_ ) & (~\new_[12768]_  | ~\new_[9418]_ );
  assign \new_[5042]_  = (~\new_[6088]_  | ~\new_[11735]_ ) & (~\new_[12775]_  | ~\new_[10126]_ );
  assign \new_[5043]_  = (~\new_[6088]_  | ~\new_[9913]_ ) & (~\new_[12768]_  | ~\new_[9641]_ );
  assign \new_[5044]_  = (~\new_[6086]_  | ~\new_[11298]_ ) & (~\new_[12777]_  | ~\new_[10111]_ );
  assign \new_[5045]_  = (~\new_[6086]_  | ~\new_[10634]_ ) & (~\new_[12777]_  | ~\new_[10136]_ );
  assign \new_[5046]_  = (~\new_[6086]_  | ~\new_[12089]_ ) & (~\new_[12775]_  | ~\new_[11860]_ );
  assign \new_[5047]_  = \new_[6641]_  | \new_[9954]_ ;
  assign \new_[5048]_  = (~\new_[6089]_  | ~\new_[9785]_ ) & (~\new_[12774]_  | ~\new_[9936]_ );
  assign \new_[5049]_  = (~\new_[6088]_  | ~\new_[10108]_ ) & (~\new_[12773]_  | ~\new_[9987]_ );
  assign \new_[5050]_  = ~\new_[6013]_  | (~\new_[6320]_  & ~\new_[9568]_ );
  assign \new_[5051]_  = (~\new_[12783]_  | ~\new_[10040]_ ) & (~\new_[7344]_  | ~\new_[9930]_ );
  assign \new_[5052]_  = (~\new_[6086]_  | ~\new_[10802]_ ) & (~\new_[12771]_  | ~\new_[9958]_ );
  assign \new_[5053]_  = (~\new_[6086]_  | ~\new_[12093]_ ) & (~\new_[12769]_  | ~\new_[9326]_ );
  assign \new_[5054]_  = (~\new_[6087]_  | ~n5021) & (~\new_[12779]_  | ~\new_[9611]_ );
  assign \new_[5055]_  = (~\new_[12593]_  | ~\new_[12567]_ ) & (~\new_[12773]_  | ~\new_[9853]_ );
  assign \new_[5056]_  = (~\new_[6087]_  | ~\new_[10164]_ ) & (~\new_[12779]_  | ~\new_[9644]_ );
  assign \new_[5057]_  = (~\new_[6087]_  | ~\new_[11363]_ ) & (~\new_[12774]_  | ~\new_[9582]_ );
  assign \new_[5058]_  = (~\new_[6086]_  | ~\new_[10411]_ ) & (~\new_[12775]_  | ~\new_[9479]_ );
  assign \new_[5059]_  = (~\new_[7059]_  | ~\new_[9668]_ ) & (~\new_[11553]_  | ~\new_[8909]_ );
  assign \new_[5060]_  = (~\new_[12784]_  | ~\new_[9615]_ ) & (~\new_[7239]_  | ~\new_[10126]_ );
  assign \new_[5061]_  = \new_[11148]_  ? \new_[6071]_  : \new_[10013]_ ;
  assign \new_[5062]_  = \new_[10855]_  ? \new_[6071]_  : \new_[9670]_ ;
  assign \new_[5063]_  = (~\new_[7059]_  | ~\new_[9807]_ ) & (~\new_[11553]_  | ~\new_[8922]_ );
  assign \new_[5064]_  = (~\new_[6087]_  | ~\new_[10902]_ ) & (~\new_[12777]_  | ~\new_[10019]_ );
  assign \new_[5065]_  = (~\new_[6088]_  | ~\new_[9903]_ ) & (~\new_[12770]_  | ~\new_[9618]_ );
  assign \new_[5066]_  = (~\new_[6090]_  | ~\new_[9648]_ ) & (~\new_[12768]_  | ~\new_[9950]_ );
  assign \new_[5067]_  = (~\new_[6088]_  | ~\new_[12598]_ ) & (~\new_[12776]_  | ~\new_[9980]_ );
  assign \new_[5068]_  = ~\new_[6022]_  | (~\new_[6320]_  & ~\new_[9296]_ );
  assign \new_[5069]_  = (~\new_[7059]_  | ~\new_[9649]_ ) & (~\new_[11553]_  | ~\new_[8901]_ );
  assign \new_[5070]_  = (~\new_[6090]_  | ~\new_[12610]_ ) & (~\new_[12774]_  | ~\new_[9374]_ );
  assign \new_[5071]_  = (~\new_[12784]_  | ~\new_[9602]_ ) & (~\new_[7239]_  | ~\new_[9987]_ );
  assign \new_[5072]_  = (~\new_[6088]_  | ~\new_[11337]_ ) & (~\new_[12769]_  | ~\new_[9978]_ );
  assign \new_[5073]_  = (~\new_[12593]_  | ~\new_[11353]_ ) & (~\new_[12779]_  | ~\new_[10097]_ );
  assign \new_[5074]_  = (~\new_[6087]_  | ~\new_[11323]_ ) & (~\new_[12768]_  | ~\new_[10083]_ );
  assign \new_[5075]_  = (~\new_[12784]_  | ~\new_[9598]_ ) & (~\new_[7344]_  | ~\new_[9326]_ );
  assign \new_[5076]_  = (~\new_[6086]_  | ~\new_[10955]_ ) & (~\new_[12775]_  | ~\new_[9675]_ );
  assign \new_[5077]_  = (~\new_[6086]_  | ~\new_[11328]_ ) & (~\new_[12773]_  | ~\new_[9709]_ );
  assign \new_[5078]_  = (~\new_[6087]_  | ~\new_[11367]_ ) & (~\new_[12771]_  | ~\new_[10115]_ );
  assign \new_[5079]_  = (~\new_[12593]_  | ~\new_[11356]_ ) & (~\new_[12776]_  | ~\new_[9619]_ );
  assign \new_[5080]_  = (~\new_[12593]_  | ~\new_[11310]_ ) & (~\new_[12775]_  | ~\new_[9567]_ );
  assign \new_[5081]_  = ~\new_[7229]_  & (~\new_[6087]_  | ~\new_[11361]_ );
  assign \new_[5082]_  = (~\new_[6086]_  | ~\new_[10933]_ ) & (~\new_[12776]_  | ~\new_[9389]_ );
  assign \new_[5083]_  = (~\new_[6086]_  | ~\new_[12044]_ ) & (~\new_[12775]_  | ~\new_[12110]_ );
  assign \new_[5084]_  = (~\new_[6086]_  | ~\new_[10960]_ ) & (~\new_[12773]_  | ~\new_[9665]_ );
  assign \new_[5085]_  = (~\new_[6090]_  | ~\new_[10526]_ ) & (~\new_[12779]_  | ~\new_[9407]_ );
  assign \new_[5086]_  = ~\new_[6014]_  | (~\new_[6320]_  & ~\new_[9101]_ );
  assign \new_[5087]_  = (~\new_[12783]_  | ~\new_[9616]_ ) & (~\new_[7344]_  | ~\new_[8977]_ );
  assign \new_[5088]_  = (~\new_[6090]_  | ~\new_[10919]_ ) & (~\new_[12774]_  | ~\new_[10037]_ );
  assign n2246 = \new_[10845]_  ? \new_[12504]_  : \new_[4342]_ ;
  assign n2151 = \new_[10885]_  ? \new_[12504]_  : \new_[4190]_ ;
  assign n2251 = \new_[10878]_  ? \new_[12504]_  : \new_[4343]_ ;
  assign n2256 = \new_[10901]_  ? \new_[12504]_  : \new_[4344]_ ;
  assign \new_[5093]_  = (~\new_[12784]_  | ~\new_[11515]_ ) & (~\new_[7344]_  | ~\new_[9107]_ );
  assign n2261 = \new_[10825]_  ? \new_[12504]_  : \new_[4345]_ ;
  assign n2171 = \new_[10828]_  ? \new_[12504]_  : \new_[4199]_ ;
  assign \new_[5096]_  = (~\new_[12784]_  | ~\new_[9844]_ ) & (~\new_[7344]_  | ~\new_[9391]_ );
  assign n2266 = \new_[10896]_  ? \new_[12504]_  : \new_[4346]_ ;
  assign n2111 = \new_[10943]_  ? \new_[12504]_  : \new_[4180]_ ;
  assign n2271 = \new_[10860]_  ? \new_[12504]_  : \new_[4347]_ ;
  assign n2141 = \new_[10868]_  ? \new_[12504]_  : \new_[4188]_ ;
  assign n2276 = \new_[10972]_  ? \new_[12504]_  : \new_[4349]_ ;
  assign n2146 = \new_[10847]_  ? \new_[12504]_  : \new_[4189]_ ;
  assign n2281 = \new_[10832]_  ? \new_[12504]_  : \new_[4350]_ ;
  assign n2136 = \new_[10844]_  ? \new_[12504]_  : \new_[4186]_ ;
  assign n2116 = \new_[10843]_  ? \new_[12504]_  : \new_[4181]_ ;
  assign n2286 = \new_[10814]_  ? \new_[12504]_  : \new_[4351]_ ;
  assign n2291 = \new_[10942]_  ? \new_[12504]_  : \new_[4352]_ ;
  assign n2846 = \new_[10923]_  ? \new_[12504]_  : \new_[4532]_ ;
  assign n2296 = \new_[10939]_  ? \new_[12504]_  : \new_[4353]_ ;
  assign n2301 = \new_[10879]_  ? \new_[12504]_  : \new_[4354]_ ;
  assign n2306 = \new_[10835]_  ? \new_[12504]_  : \new_[4355]_ ;
  assign n2841 = \new_[10867]_  ? \new_[12504]_  : \new_[4531]_ ;
  assign n2311 = \new_[10968]_  ? \new_[12504]_  : \new_[4356]_ ;
  assign n2321 = \new_[10935]_  ? \new_[12504]_  : \new_[4358]_ ;
  assign n2316 = \new_[10947]_  ? \new_[12504]_  : \new_[4357]_ ;
  assign n2836 = \new_[10970]_  ? \new_[12504]_  : \new_[4528]_ ;
  assign n2326 = \new_[10911]_  ? \new_[12504]_  : \new_[4359]_ ;
  assign n2331 = \new_[10900]_  ? \new_[12504]_  : \new_[4360]_ ;
  assign \new_[5119]_  = (~\new_[12784]_  | ~\new_[9659]_ ) & (~\new_[7344]_  | ~\new_[9707]_ );
  assign n2336 = \new_[10831]_  ? \new_[12504]_  : \new_[4361]_ ;
  assign \new_[5121]_  = ~\new_[6020]_  | (~\new_[6320]_  & ~\new_[9030]_ );
  assign n2826 = \new_[10916]_  ? \new_[12504]_  : \new_[4523]_ ;
  assign n2341 = \new_[10869]_  ? \new_[12504]_  : \new_[4362]_ ;
  assign \new_[5124]_  = (~\new_[12784]_  | ~\new_[11962]_ ) & (~\new_[7344]_  | ~\new_[9684]_ );
  assign n2796 = \new_[10852]_  ? \new_[12504]_  : \new_[4516]_ ;
  assign n2811 = \new_[10819]_  ? \new_[12504]_  : \new_[4519]_ ;
  assign n2741 = \new_[10833]_  ? \new_[12504]_  : \new_[4480]_ ;
  assign n2786 = \new_[10817]_  ? \new_[12504]_  : \new_[4514]_ ;
  assign n2351 = \new_[10845]_  ? \new_[6068]_  : \new_[4365]_ ;
  assign n2346 = \new_[10908]_  ? \new_[12504]_  : \new_[4364]_ ;
  assign n2361 = \new_[10885]_  ? \new_[6068]_  : \new_[4368]_ ;
  assign n2356 = \new_[10878]_  ? \new_[6068]_  : \new_[4366]_ ;
  assign n2366 = \new_[10901]_  ? \new_[6068]_  : \new_[4369]_ ;
  assign n2371 = \new_[10825]_  ? \new_[6068]_  : \new_[4370]_ ;
  assign n2376 = \new_[10896]_  ? \new_[6068]_  : \new_[4371]_ ;
  assign n2771 = \new_[10828]_  ? \new_[6068]_  : \new_[4510]_ ;
  assign n2381 = \new_[10943]_  ? \new_[6068]_  : \new_[4372]_ ;
  assign n2386 = \new_[10860]_  ? \new_[6068]_  : \new_[4373]_ ;
  assign n2746 = \new_[10868]_  ? \new_[6068]_  : \new_[4494]_ ;
  assign n2391 = \new_[10847]_  ? \new_[6068]_  : \new_[4374]_ ;
  assign n2396 = \new_[10844]_  ? \new_[6068]_  : \new_[4375]_ ;
  assign n2401 = \new_[10972]_  ? \new_[6068]_  : \new_[4376]_ ;
  assign n2736 = \new_[10832]_  ? \new_[6068]_  : \new_[4474]_ ;
  assign n2411 = \new_[10843]_  ? \new_[6068]_  : \new_[4378]_ ;
  assign n2406 = \new_[10814]_  ? \new_[6068]_  : \new_[4377]_ ;
  assign n2416 = \new_[10942]_  ? \new_[6068]_  : \new_[4379]_ ;
  assign n2421 = \new_[10923]_  ? \new_[6068]_  : \new_[4380]_ ;
  assign n2121 = \new_[10939]_  ? \new_[6068]_  : \new_[4182]_ ;
  assign n2426 = \new_[10879]_  ? \new_[6068]_  : \new_[4381]_ ;
  assign n2431 = \new_[10835]_  ? \new_[6068]_  : \new_[4382]_ ;
  assign n2731 = \new_[10867]_  ? \new_[6068]_  : \new_[4448]_ ;
  assign n2436 = \new_[10968]_  ? \new_[6068]_  : \new_[4383]_ ;
  assign n2441 = \new_[10947]_  ? \new_[6068]_  : \new_[4384]_ ;
  assign n2446 = \new_[10935]_  ? \new_[6068]_  : \new_[4385]_ ;
  assign n2231 = \new_[10970]_  ? \new_[6068]_  : \new_[4339]_ ;
  assign n2451 = \new_[10911]_  ? \new_[6068]_  : \new_[4386]_ ;
  assign n2456 = \new_[10900]_  ? \new_[6068]_  : \new_[4387]_ ;
  assign n2461 = \new_[10831]_  ? \new_[6068]_  : \new_[4388]_ ;
  assign n2226 = \new_[10916]_  ? \new_[6068]_  : \new_[4313]_ ;
  assign n2466 = \new_[10869]_  ? \new_[6068]_  : \new_[4389]_ ;
  assign n2471 = \new_[10852]_  ? \new_[6068]_  : \new_[4390]_ ;
  assign n2476 = \new_[10819]_  ? \new_[6068]_  : \new_[4391]_ ;
  assign n2221 = \new_[10833]_  ? \new_[6068]_  : \new_[4303]_ ;
  assign n2481 = \new_[10817]_  ? \new_[6068]_  : \new_[4392]_ ;
  assign n2216 = \new_[10908]_  ? \new_[6068]_  : \new_[4295]_ ;
  assign n2486 = \new_[10845]_  ? \new_[6069]_  : \new_[4393]_ ;
  assign n2206 = \new_[10885]_  ? \new_[6069]_  : \new_[4278]_ ;
  assign n2491 = \new_[10878]_  ? \new_[6069]_  : \new_[4395]_ ;
  assign n2211 = \new_[10901]_  ? \new_[6069]_  : \new_[4289]_ ;
  assign n2496 = \new_[10825]_  ? \new_[6069]_  : \new_[4396]_ ;
  assign n2201 = \new_[10828]_  ? \new_[6069]_  : \new_[4249]_ ;
  assign n2501 = \new_[10896]_  ? \new_[6069]_  : \new_[4397]_ ;
  assign n2506 = \new_[10943]_  ? \new_[6069]_  : \new_[4398]_ ;
  assign n2511 = \new_[10860]_  ? \new_[6069]_  : \new_[4399]_ ;
  assign n2176 = \new_[10868]_  ? \new_[6069]_  : \new_[4205]_ ;
  assign n2516 = \new_[10847]_  ? \new_[6069]_  : \new_[4400]_ ;
  assign n2521 = \new_[10844]_  ? \new_[6069]_  : \new_[4401]_ ;
  assign n2526 = \new_[10972]_  ? \new_[6069]_  : \new_[4402]_ ;
  assign n2181 = \new_[10832]_  ? \new_[6069]_  : \new_[4231]_ ;
  assign n2531 = \new_[10843]_  ? \new_[6069]_  : \new_[4403]_ ;
  assign \new_[5181]_  = \new_[6035]_  | \new_[11716]_ ;
  assign n2536 = \new_[10814]_  ? \new_[6069]_  : \new_[4404]_ ;
  assign n2541 = \new_[10942]_  ? \new_[6069]_  : \new_[4405]_ ;
  assign n2126 = \new_[10923]_  ? \new_[6069]_  : \new_[4183]_ ;
  assign n2546 = \new_[10939]_  ? \new_[6069]_  : \new_[4406]_ ;
  assign n2161 = \new_[10879]_  ? \new_[6069]_  : \new_[4195]_ ;
  assign n2551 = \new_[10835]_  ? \new_[6069]_  : \new_[4407]_ ;
  assign n2166 = \new_[10867]_  ? \new_[6069]_  : \new_[4198]_ ;
  assign n2556 = \new_[10968]_  ? \new_[6069]_  : \new_[4408]_ ;
  assign n2561 = \new_[10947]_  ? \new_[6069]_  : \new_[4409]_ ;
  assign n2566 = \new_[10935]_  ? \new_[6069]_  : \new_[4410]_ ;
  assign n2156 = \new_[10970]_  ? \new_[6069]_  : \new_[4191]_ ;
  assign n2571 = \new_[10911]_  ? \new_[6069]_  : \new_[4411]_ ;
  assign n2576 = \new_[10900]_  ? \new_[6069]_  : \new_[4412]_ ;
  assign n2581 = \new_[10831]_  ? \new_[6069]_  : \new_[4413]_ ;
  assign n2131 = \new_[10916]_  ? \new_[6069]_  : \new_[4185]_ ;
  assign n2586 = \new_[10869]_  ? \new_[6069]_  : \new_[4414]_ ;
  assign n2591 = \new_[10852]_  ? \new_[6069]_  : \new_[4415]_ ;
  assign n2596 = \new_[10819]_  ? \new_[6069]_  : \new_[4416]_ ;
  assign n2816 = \new_[10833]_  ? \new_[6069]_  : \new_[4521]_ ;
  assign n2601 = \new_[10817]_  ? \new_[6069]_  : \new_[4417]_ ;
  assign n2851 = \new_[10908]_  ? \new_[6069]_  : \new_[4533]_ ;
  assign n2606 = \new_[10845]_  ? \new_[11410]_  : \new_[4418]_ ;
  assign n2856 = \new_[10885]_  ? \new_[11410]_  : \new_[4535]_ ;
  assign n2611 = \new_[10878]_  ? \new_[11410]_  : \new_[4419]_ ;
  assign n2616 = \new_[10901]_  ? \new_[11410]_  : \new_[4420]_ ;
  assign n2621 = \new_[10825]_  ? \new_[11410]_  : \new_[4421]_ ;
  assign n2801 = \new_[10828]_  ? \new_[11410]_  : \new_[4517]_ ;
  assign n2626 = \new_[10896]_  ? \new_[11410]_  : \new_[4422]_ ;
  assign n2631 = \new_[10943]_  ? \new_[11410]_  : \new_[4423]_ ;
  assign n2636 = \new_[10860]_  ? \new_[11410]_  : \new_[4424]_ ;
  assign n2831 = \new_[10868]_  ? \new_[11410]_  : \new_[4527]_ ;
  assign n2641 = \new_[10847]_  ? \new_[11410]_  : \new_[4425]_ ;
  assign n2646 = \new_[10844]_  ? \new_[11410]_  : \new_[4426]_ ;
  assign n2651 = \new_[10972]_  ? \new_[11410]_  : \new_[4427]_ ;
  assign n2806 = \new_[10832]_  ? \new_[11410]_  : \new_[4518]_ ;
  assign n2656 = \new_[10843]_  ? \new_[11410]_  : \new_[4428]_ ;
  assign n2661 = \new_[10814]_  ? \new_[11410]_  : \new_[4429]_ ;
  assign n2666 = \new_[10942]_  ? \new_[11410]_  : \new_[4430]_ ;
  assign n2776 = \new_[10923]_  ? \new_[11410]_  : \new_[4511]_ ;
  assign n2671 = \new_[10939]_  ? \new_[11410]_  : \new_[4431]_ ;
  assign n2791 = \new_[10879]_  ? \new_[11410]_  : \new_[4515]_ ;
  assign n2676 = \new_[10835]_  ? \new_[11410]_  : \new_[4432]_ ;
  assign n2781 = \new_[10867]_  ? \new_[11410]_  : \new_[4512]_ ;
  assign n2681 = \new_[10968]_  ? \new_[11410]_  : \new_[4433]_ ;
  assign n2761 = \new_[10947]_  ? \new_[11410]_  : \new_[4506]_ ;
  assign n2686 = \new_[10935]_  ? \new_[11410]_  : \new_[4434]_ ;
  assign n2766 = \new_[10970]_  ? \new_[11410]_  : \new_[4509]_ ;
  assign n2691 = \new_[10911]_  ? \new_[11410]_  : \new_[4436]_ ;
  assign n2696 = \new_[10900]_  ? \new_[11410]_  : \new_[4437]_ ;
  assign n2701 = \new_[10831]_  ? \new_[11410]_  : \new_[4438]_ ;
  assign n2756 = \new_[10916]_  ? \new_[11410]_  : \new_[4504]_ ;
  assign n2706 = \new_[10869]_  ? \new_[11410]_  : \new_[4439]_ ;
  assign n2711 = \new_[10852]_  ? \new_[11410]_  : \new_[4440]_ ;
  assign n2716 = \new_[10819]_  ? \new_[11410]_  : \new_[4441]_ ;
  assign n2751 = \new_[10833]_  ? \new_[11410]_  : \new_[4495]_ ;
  assign n2726 = \new_[10817]_  ? \new_[11410]_  : \new_[4443]_ ;
  assign n2721 = \new_[10908]_  ? \new_[11410]_  : \new_[4442]_ ;
  assign \new_[5239]_  = \new_[3439]_  ^ \new_[6071]_ ;
  assign \new_[5240]_  = ~\new_[5662]_  & (~\new_[8914]_  | ~\new_[7065]_ );
  assign \new_[5241]_  = ~\new_[5668]_  & (~\new_[9111]_  | ~\new_[7226]_ );
  assign \new_[5242]_  = ~\new_[12240]_ ;
  assign \new_[5243]_  = (~\new_[3169]_  | ~\new_[7366]_ ) & (~\new_[11080]_  | ~\new_[6064]_ );
  assign \new_[5244]_  = (~\new_[3177]_  | ~\new_[7366]_ ) & (~\new_[11179]_  | ~\new_[7286]_ );
  assign \new_[5245]_  = ~\new_[12677]_  & ~\new_[5713]_ ;
  assign \new_[5246]_  = ~\new_[5693]_  & ~\new_[7864]_ ;
  assign \new_[5247]_  = \new_[5642]_ ;
  assign \new_[5248]_  = \new_[5642]_ ;
  assign \new_[5249]_  = ~\new_[5642]_ ;
  assign \new_[5250]_  = ~\new_[5657]_  & (~\new_[7577]_  | ~\new_[8919]_ );
  assign \new_[5251]_  = ~\new_[5653]_  & (~\new_[7226]_  | ~\new_[9383]_ );
  assign \new_[5252]_  = ~\new_[5655]_  & (~\new_[7226]_  | ~\new_[9401]_ );
  assign \new_[5253]_  = ~\new_[5656]_  & (~\new_[7226]_  | ~\new_[10031]_ );
  assign \new_[5254]_  = ~\new_[5658]_  & (~\new_[7226]_  | ~\new_[10099]_ );
  assign \new_[5255]_  = ~\new_[5659]_  & (~\new_[7226]_  | ~\new_[9661]_ );
  assign \new_[5256]_  = ~\new_[5660]_  & (~\new_[7226]_  | ~\new_[9963]_ );
  assign \new_[5257]_  = ~\new_[5661]_  & (~\new_[7226]_  | ~\new_[10104]_ );
  assign \new_[5258]_  = ~\new_[5663]_  & (~\new_[7226]_  | ~\new_[9607]_ );
  assign \new_[5259]_  = ~\new_[5664]_  & (~\new_[7226]_  | ~\new_[10011]_ );
  assign \new_[5260]_  = ~\new_[5665]_  & (~\new_[7226]_  | ~\new_[9680]_ );
  assign \new_[5261]_  = ~\new_[5666]_  & (~\new_[7226]_  | ~\new_[10263]_ );
  assign \new_[5262]_  = ~\new_[5667]_  & (~\new_[7226]_  | ~\new_[9995]_ );
  assign \new_[5263]_  = ~\new_[5669]_  & (~\new_[7226]_  | ~\new_[9930]_ );
  assign \new_[5264]_  = ~\new_[5670]_  & (~\new_[7226]_  | ~\new_[10237]_ );
  assign \new_[5265]_  = ~\new_[5671]_  & (~\new_[7226]_  | ~\new_[9660]_ );
  assign \new_[5266]_  = ~\new_[5673]_  & (~\new_[7226]_  | ~\new_[9641]_ );
  assign \new_[5267]_  = ~\new_[5675]_  & (~\new_[7226]_  | ~\new_[10111]_ );
  assign \new_[5268]_  = ~\new_[5676]_  & (~\new_[7226]_  | ~\new_[10287]_ );
  assign \new_[5269]_  = ~\new_[5677]_  & (~\new_[7226]_  | ~\new_[11860]_ );
  assign \new_[5270]_  = ~\new_[5679]_  & (~\new_[7226]_  | ~\new_[9958]_ );
  assign \new_[5271]_  = ~\new_[5680]_  & (~\new_[7226]_  | ~\new_[9326]_ );
  assign \new_[5272]_  = ~\new_[5681]_  & (~\new_[7226]_  | ~\new_[9611]_ );
  assign \new_[5273]_  = ~\new_[5682]_  & (~\new_[7226]_  | ~\new_[9853]_ );
  assign \new_[5274]_  = ~\new_[5683]_  & (~\new_[7226]_  | ~\new_[9644]_ );
  assign \new_[5275]_  = ~\new_[5684]_  & (~\new_[7226]_  | ~\new_[9582]_ );
  assign \new_[5276]_  = ~\new_[5685]_  & (~\new_[7226]_  | ~\new_[9479]_ );
  assign \new_[5277]_  = ~\new_[5686]_  & (~\new_[7226]_  | ~\new_[9655]_ );
  assign \new_[5278]_  = ~\new_[5687]_  & (~\new_[7226]_  | ~\new_[8977]_ );
  assign \new_[5279]_  = ~\new_[5688]_  & (~\new_[7226]_  | ~\new_[10019]_ );
  assign \new_[5280]_  = ~\new_[5689]_  & (~\new_[7226]_  | ~\new_[9657]_ );
  assign \new_[5281]_  = ~\new_[5690]_  & (~\new_[7226]_  | ~\new_[9107]_ );
  assign \new_[5282]_  = ~\new_[5714]_  & (~\new_[6719]_  | ~\new_[10278]_ );
  assign \new_[5283]_  = ~\new_[6689]_  & ~\new_[12568]_ ;
  assign \new_[5284]_  = ~\new_[5692]_  & (~\new_[7226]_  | ~\new_[9374]_ );
  assign \new_[5285]_  = ~\new_[12512]_  | ~\new_[12233]_  | ~\new_[12514]_ ;
  assign \new_[5286]_  = ~\new_[5694]_  & (~\new_[7226]_  | ~\new_[10097]_ );
  assign \new_[5287]_  = ~\new_[9914]_  | ~\new_[9902]_  | ~\new_[5710]_  | ~\new_[9885]_ ;
  assign \new_[5288]_  = ~\new_[5696]_  & (~\new_[7226]_  | ~\new_[9675]_ );
  assign \new_[5289]_  = ~\new_[5697]_  & (~\new_[7226]_  | ~\new_[9709]_ );
  assign \new_[5290]_  = ~\new_[5698]_  & (~\new_[7226]_  | ~\new_[10115]_ );
  assign \new_[5291]_  = ~\new_[5699]_  & (~\new_[7226]_  | ~\new_[9109]_ );
  assign \new_[5292]_  = ~\new_[5700]_  & (~\new_[7226]_  | ~\new_[9599]_ );
  assign \new_[5293]_  = ~\new_[5702]_  & (~\new_[7226]_  | ~\new_[9684]_ );
  assign \new_[5294]_  = ~\new_[5704]_  & (~\new_[7226]_  | ~\new_[9604]_ );
  assign \new_[5295]_  = ~\new_[5705]_  & (~\new_[7226]_  | ~\new_[10137]_ );
  assign \new_[5296]_  = ~\new_[5706]_  & (~\new_[7226]_  | ~\new_[12110]_ );
  assign \new_[5297]_  = ~\new_[5707]_  & (~\new_[7226]_  | ~\new_[9989]_ );
  assign \new_[5298]_  = ~\new_[5708]_  & (~\new_[7226]_  | ~\new_[9407]_ );
  assign \new_[5299]_  = ~\new_[5709]_  & (~\new_[7226]_  | ~\new_[10037]_ );
  assign n2821 = ~\new_[7918]_  | ~\new_[7721]_  | ~\new_[5674]_  | ~\new_[7705]_ ;
  assign \new_[5301]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10402]_ ) | (~\new_[12700]_  & ~\new_[12672]_  & ~\new_[10402]_ );
  assign \new_[5302]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[12274]_ ) | (~\new_[12700]_  & ~\new_[12672]_  & ~\new_[12274]_ );
  assign \new_[5303]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10698]_ ) | (~\new_[12701]_  & ~\new_[12672]_  & ~\new_[10698]_ );
  assign \new_[5304]_  = (~\new_[12652]_  & ~\new_[8499]_  & ~\new_[12184]_ ) | (~\new_[12699]_  & ~\new_[12672]_  & ~\new_[12184]_ );
  assign \new_[5305]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[11349]_ ) | (~\new_[12709]_  & ~\new_[12672]_  & ~\new_[11349]_ );
  assign \new_[5306]_  = (~\new_[12654]_  & ~\new_[8499]_  & ~\new_[10722]_ ) | (~\new_[12713]_  & ~\new_[12672]_  & ~\new_[10722]_ );
  assign \new_[5307]_  = (~\new_[12651]_  & ~\new_[8499]_  & ~\new_[11737]_ ) | (~\new_[12705]_  & ~\new_[12672]_  & ~\new_[11737]_ );
  assign \new_[5308]_  = (~\new_[12654]_  & ~\new_[8408]_  & ~\new_[11575]_ ) | (~\new_[12711]_  & ~\new_[12672]_  & ~\new_[11575]_ );
  assign \new_[5309]_  = (~\new_[12652]_  & ~\new_[8408]_  & ~\new_[10809]_ ) | (~\new_[12709]_  & ~\new_[12672]_  & ~\new_[10809]_ );
  assign \new_[5310]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[11334]_ ) | (~\new_[12710]_  & ~\new_[12672]_  & ~\new_[11334]_ );
  assign \new_[5311]_  = (~\new_[12651]_  & ~\new_[8499]_  & ~\new_[10752]_ ) | (~\new_[12706]_  & ~\new_[12672]_  & ~\new_[10752]_ );
  assign \new_[5312]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[11344]_ ) | (~\new_[12710]_  & ~\new_[12672]_  & ~\new_[11344]_ );
  assign \new_[5313]_  = (~\new_[12656]_  & ~\new_[11525]_  & ~\new_[10920]_ ) | (~\new_[12700]_  & ~\new_[12672]_  & ~\new_[10920]_ );
  assign \new_[5314]_  = ~\new_[6102]_  & (~\new_[7344]_  | ~\new_[9627]_ );
  assign \new_[5315]_  = (~\new_[12652]_  & ~\new_[11525]_  & ~\new_[11341]_ ) | (~\new_[12698]_  & ~\new_[12672]_  & ~\new_[11341]_ );
  assign \new_[5316]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[11493]_ ) | (~\new_[12699]_  & ~\new_[12672]_  & ~\new_[11493]_ );
  assign \new_[5317]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[10673]_ ) | (~\new_[12709]_  & ~\new_[12672]_  & ~\new_[10673]_ );
  assign \new_[5318]_  = (~\new_[12651]_  & ~\new_[8408]_  & ~\new_[11321]_ ) | (~\new_[12707]_  & ~\new_[12672]_  & ~\new_[11321]_ );
  assign \new_[5319]_  = (~\new_[12654]_  & ~\new_[11525]_  & ~\new_[11012]_ ) | (~\new_[12698]_  & ~\new_[12672]_  & ~\new_[11012]_ );
  assign \new_[5320]_  = (~\new_[12650]_  & ~\new_[8408]_  & ~\new_[11881]_ ) | (~\new_[12711]_  & ~\new_[12672]_  & ~\new_[11881]_ );
  assign \new_[5321]_  = (~\new_[12651]_  & ~\new_[8408]_  & ~\new_[10872]_ ) | (~\new_[12710]_  & ~\new_[12672]_  & ~\new_[10872]_ );
  assign \new_[5322]_  = (~\new_[12652]_  & ~\new_[11525]_  & ~\new_[11317]_ ) | (~\new_[12701]_  & ~\new_[12672]_  & ~\new_[11317]_ );
  assign \new_[5323]_  = (~\new_[12654]_  & ~\new_[8408]_  & ~\new_[10591]_ ) | (~\new_[12705]_  & ~\new_[12672]_  & ~\new_[10591]_ );
  assign \new_[5324]_  = (~\new_[12652]_  & ~\new_[8499]_  & ~\new_[10897]_ ) | (~\new_[12705]_  & ~\new_[12672]_  & ~\new_[10897]_ );
  assign \new_[5325]_  = (~\new_[12650]_  & ~\new_[8499]_  & ~\new_[12094]_ ) | (~\new_[12716]_  & ~\new_[12672]_  & ~\new_[12094]_ );
  assign \new_[5326]_  = (~\new_[12650]_  & ~\new_[8499]_  & ~\new_[10676]_ ) | (~\new_[12704]_  & ~\new_[12672]_  & ~\new_[10676]_ );
  assign \new_[5327]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[10724]_ ) | (~\new_[12709]_  & ~\new_[12672]_  & ~\new_[10724]_ );
  assign \new_[5328]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10704]_ ) | (~\new_[12698]_  & ~\new_[12672]_  & ~\new_[10704]_ );
  assign \new_[5329]_  = \new_[12614]_  | \new_[12495]_  | \new_[7864]_  | \new_[12496]_ ;
  assign \new_[5330]_  = (~\new_[12651]_  & ~\new_[8408]_  & ~\new_[12555]_ ) | (~\new_[12707]_  & ~\new_[12672]_  & ~\new_[12555]_ );
  assign \new_[5331]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[12052]_ ) | (~\new_[12706]_  & ~\new_[12672]_  & ~\new_[12052]_ );
  assign \new_[5332]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[12611]_ ) | (~\new_[12709]_  & ~\new_[12672]_  & ~\new_[12611]_ );
  assign \new_[5333]_  = (~\new_[12651]_  & ~\new_[8408]_  & ~\new_[11338]_ ) | (~\new_[12714]_  & ~\new_[12672]_  & ~\new_[11338]_ );
  assign \new_[5334]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[11393]_ ) | (~\new_[12701]_  & ~\new_[12672]_  & ~\new_[11393]_ );
  assign \new_[5335]_  = (~\new_[12652]_  & ~\new_[8408]_  & ~\new_[11324]_ ) | (~\new_[12699]_  & ~\new_[12672]_  & ~\new_[11324]_ );
  assign \new_[5336]_  = (~\new_[12650]_  & ~\new_[8499]_  & ~\new_[10579]_ ) | (~\new_[12709]_  & ~\new_[12672]_  & ~\new_[10579]_ );
  assign \new_[5337]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[11329]_ ) | (~\new_[12700]_  & ~\new_[12281]_  & ~\new_[11329]_ );
  assign \new_[5338]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[12400]_ ) | (~\new_[12698]_  & ~\new_[12672]_  & ~\new_[12400]_ );
  assign \new_[5339]_  = (~\new_[12654]_  & ~\new_[8499]_  & ~\new_[10771]_ ) | (~\new_[12706]_  & ~\new_[12672]_  & ~\new_[10771]_ );
  assign \new_[5340]_  = (~\new_[12650]_  & ~\new_[8499]_  & ~\new_[11311]_ ) | (~\new_[12711]_  & ~\new_[12672]_  & ~\new_[11311]_ );
  assign \new_[5341]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[11314]_ ) | (~\new_[12701]_  & ~\new_[12672]_  & ~\new_[11314]_ );
  assign \new_[5342]_  = (~\new_[12650]_  & ~\new_[8499]_  & ~\new_[10348]_ ) | (~\new_[12711]_  & ~\new_[12672]_  & ~\new_[10348]_ );
  assign \new_[5343]_  = (~\new_[12656]_  & ~\new_[8499]_  & ~\new_[10767]_ ) | (~\new_[12700]_  & ~\new_[12672]_  & ~\new_[10767]_ );
  assign \new_[5344]_  = (~\new_[12654]_  & ~\new_[8408]_  & ~\new_[10715]_ ) | (~\new_[12713]_  & ~\new_[12672]_  & ~\new_[10715]_ );
  assign \new_[5345]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10754]_ ) | (~\new_[12700]_  & ~\new_[12672]_  & ~\new_[10754]_ );
  assign \new_[5346]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10783]_ ) | (~\new_[12707]_  & ~\new_[12672]_  & ~\new_[10783]_ );
  assign \new_[5347]_  = (~\new_[12656]_  & ~\new_[8408]_  & ~\new_[10328]_ ) | (~\new_[12707]_  & ~\new_[12672]_  & ~\new_[10328]_ );
  assign \new_[5348]_  = ~\new_[12508]_ ;
  assign \new_[5349]_  = ~\new_[6316]_  & (~\new_[6395]_  | ~\new_[9851]_ );
  assign \new_[5350]_  = \new_[3041]_  ^ \new_[6359]_ ;
  assign \new_[5351]_  = ~\new_[6316]_  & (~\new_[6399]_  | ~\new_[10161]_ );
  assign \new_[5352]_  = ~\new_[6316]_  & (~\new_[6400]_  | ~\new_[9924]_ );
  assign \new_[5353]_  = ~\new_[6316]_  & (~\new_[6402]_  | ~\new_[9590]_ );
  assign \new_[5354]_  = ~\new_[12741]_  & ~\new_[9927]_ ;
  assign \new_[5355]_  = ~\new_[6316]_  & (~\new_[6449]_  | ~\new_[9742]_ );
  assign \new_[5356]_  = ~\new_[6316]_  & (~\new_[6456]_  | ~\new_[9860]_ );
  assign \new_[5357]_  = ~\new_[6316]_  & (~\new_[6462]_  | ~\new_[9743]_ );
  assign \new_[5358]_  = \new_[11120]_  ? \new_[12622]_  : \new_[11005]_ ;
  assign \new_[5359]_  = ~\new_[6317]_  & (~\new_[6432]_  | ~\new_[9955]_ );
  assign \new_[5360]_  = ~\new_[6316]_  & (~\new_[6406]_  | ~\new_[9739]_ );
  assign \new_[5361]_  = ~\new_[6316]_  & (~\new_[6469]_  | ~\new_[9899]_ );
  assign \new_[5362]_  = ~\new_[6316]_  & (~\new_[6468]_  | ~\new_[9859]_ );
  assign \new_[5363]_  = ~\new_[6316]_  & (~\new_[6470]_  | ~\new_[10167]_ );
  assign n2876 = ~\new_[6820]_  | (~\new_[6391]_  & ~\new_[11113]_ );
  assign \new_[5365]_  = (~\new_[7083]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9592]_ );
  assign \new_[5366]_  = (~\new_[7088]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9960]_ );
  assign \new_[5367]_  = (~\new_[7089]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9612]_ );
  assign \new_[5368]_  = (~\new_[7090]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9603]_ );
  assign \new_[5369]_  = (~\new_[7092]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9678]_ );
  assign \new_[5370]_  = ~\new_[7200]_  | ~\new_[6094]_ ;
  assign \new_[5371]_  = (~\new_[7105]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9614]_ );
  assign \new_[5372]_  = ~\new_[7214]_  | ~\new_[6096]_ ;
  assign \new_[5373]_  = ~\new_[11894]_  | ~\new_[9644]_ ;
  assign \new_[5374]_  = (~\new_[6816]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9408]_ );
  assign \new_[5375]_  = ~\new_[6267]_  & ~\new_[10150]_ ;
  assign \new_[5376]_  = (~\new_[6817]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9874]_ );
  assign \new_[5377]_  = (~\new_[6818]_  | ~\new_[6393]_ ) & (~\new_[7995]_  | ~\new_[9393]_ );
  assign \new_[5378]_  = \new_[6113]_  | \new_[7063]_ ;
  assign \new_[5379]_  = \new_[6171]_  & \new_[6130]_ ;
  assign \new_[5380]_  = \new_[6190]_  & \new_[6145]_ ;
  assign \new_[5381]_  = ~\new_[6714]_  & (~\new_[11894]_  | ~\new_[9978]_ );
  assign \new_[5382]_  = \new_[6193]_  & \new_[6146]_ ;
  assign \new_[5383]_  = ~\new_[5865]_  | ~\new_[9619]_ ;
  assign \new_[5384]_  = \new_[3042]_  ^ \new_[6398]_ ;
  assign \new_[5385]_  = (~\new_[6746]_  | ~\new_[7776]_ ) & (~\new_[11304]_  | ~\new_[7482]_ );
  assign \new_[5386]_  = (~\new_[6749]_  | ~\new_[7776]_ ) & (~\new_[11304]_  | ~\new_[7484]_ );
  assign \new_[5387]_  = (~\new_[6750]_  | ~\new_[7825]_ ) & (~\new_[11304]_  | ~\new_[7486]_ );
  assign \new_[5388]_  = (~\new_[6751]_  | ~\new_[7825]_ ) & (~\new_[11304]_  | ~\new_[7312]_ );
  assign \new_[5389]_  = (~\new_[6753]_  | ~\new_[7776]_ ) & (~\new_[11304]_  | ~\new_[7314]_ );
  assign \new_[5390]_  = (~\new_[6754]_  | ~\new_[7825]_ ) & (~\new_[11305]_  | ~\new_[7651]_ );
  assign \new_[5391]_  = (~\new_[6758]_  | ~\new_[7777]_ ) & (~\new_[11302]_  | ~\new_[7493]_ );
  assign \new_[5392]_  = (~\new_[6759]_  | ~\new_[7823]_ ) & (~\new_[11304]_  | ~\new_[7494]_ );
  assign \new_[5393]_  = \new_[12709]_  | \new_[7423]_ ;
  assign \new_[5394]_  = \new_[12710]_  | \new_[7165]_ ;
  assign \new_[5395]_  = (~\new_[6763]_  | ~\new_[7823]_ ) & (~\new_[11301]_  | ~\new_[7502]_ );
  assign \new_[5396]_  = (~\new_[6764]_  | ~\new_[7823]_ ) & (~\new_[11301]_  | ~\new_[7488]_ );
  assign \new_[5397]_  = (~\new_[6765]_  | ~\new_[7823]_ ) & (~\new_[11306]_  | ~\new_[7506]_ );
  assign \new_[5398]_  = ~\new_[12700]_  & ~\new_[7425]_ ;
  assign \new_[5399]_  = (~\new_[6766]_  | ~\new_[7823]_ ) & (~\new_[11306]_  | ~\new_[7485]_ );
  assign \new_[5400]_  = ~\new_[7007]_  & (~\new_[11305]_  | ~\new_[7508]_ );
  assign \new_[5401]_  = (~\new_[6768]_  | ~\new_[7777]_ ) & (~\new_[11305]_  | ~\new_[7511]_ );
  assign \new_[5402]_  = (~\new_[6772]_  | ~\new_[7823]_ ) & (~\new_[11302]_  | ~\new_[7500]_ );
  assign \new_[5403]_  = ~\new_[6277]_  & ~\new_[7141]_ ;
  assign \new_[5404]_  = (~\new_[6745]_  | ~\new_[7777]_ ) & (~\new_[11305]_  | ~\new_[7519]_ );
  assign \new_[5405]_  = (~\new_[6773]_  | ~\new_[7776]_ ) & (~\new_[11303]_  | ~\new_[7318]_ );
  assign \new_[5406]_  = (~\new_[6774]_  | ~\new_[7825]_ ) & (~\new_[11303]_  | ~\new_[7320]_ );
  assign \new_[5407]_  = (~\new_[6744]_  | ~\new_[7823]_ ) & (~\new_[11305]_  | ~\new_[7516]_ );
  assign \new_[5408]_  = (~\new_[6760]_  | ~\new_[7776]_ ) & (~\new_[11304]_  | ~\new_[7321]_ );
  assign \new_[5409]_  = ~\new_[6156]_  & (~\new_[11864]_  | ~\new_[9655]_ );
  assign \new_[5410]_  = ~\new_[6693]_  | (~\new_[7176]_  & ~\new_[12003]_ );
  assign \new_[5411]_  = ~\new_[6694]_  | (~\new_[7176]_  & ~\new_[10208]_ );
  assign \new_[5412]_  = ~\new_[6695]_  | (~\new_[7176]_  & ~\new_[9861]_ );
  assign \new_[5413]_  = ~\new_[6699]_  | (~\new_[7176]_  & ~\new_[10057]_ );
  assign \new_[5414]_  = ~\new_[6711]_  | (~\new_[7176]_  & ~\new_[9305]_ );
  assign \new_[5415]_  = ~\new_[5807]_ ;
  assign \new_[5416]_  = ~\new_[6717]_  | (~\new_[7176]_  & ~\new_[10166]_ );
  assign \new_[5417]_  = ~\new_[6536]_  | (~\new_[7176]_  & ~\new_[10199]_ );
  assign \new_[5418]_  = ~\new_[6114]_  | ~\new_[6396]_ ;
  assign \new_[5419]_  = (~\new_[11305]_  | ~\new_[7495]_ ) & (~\new_[7662]_  | ~\new_[7366]_ );
  assign \new_[5420]_  = (~\new_[11894]_  | ~\new_[9682]_ ) & (~\new_[7289]_  | ~\new_[8524]_ );
  assign n2906 = ~\new_[5809]_ ;
  assign n2866 = ~\new_[5810]_ ;
  assign n2901 = ~\new_[5811]_ ;
  assign n2891 = ~\new_[5812]_ ;
  assign n2886 = ~\new_[5813]_ ;
  assign n2881 = ~\new_[5814]_ ;
  assign n2861 = ~\new_[5815]_ ;
  assign n2911 = ~\new_[5816]_ ;
  assign n2896 = ~\new_[5817]_ ;
  assign \new_[5430]_  = ~\new_[8001]_  | ~\new_[8003]_  | ~\new_[11774]_  | ~\new_[12746]_ ;
  assign \new_[5431]_  = \new_[4145]_  ^ \new_[6621]_ ;
  assign \new_[5432]_  = \new_[12683]_  | \new_[7191]_ ;
  assign \new_[5433]_  = ~\new_[6267]_  & ~\new_[12003]_ ;
  assign \new_[5434]_  = ~\new_[12741]_  & ~\new_[12003]_ ;
  assign \new_[5435]_  = ~\new_[6267]_  & ~\new_[9851]_ ;
  assign \new_[5436]_  = ~\new_[6208]_  | ~\new_[7167]_ ;
  assign \new_[5437]_  = ~\new_[6284]_  & ~\new_[10258]_ ;
  assign \new_[5438]_  = ~\new_[11894]_  | ~\new_[9401]_ ;
  assign \new_[5439]_  = ~\new_[6267]_  & ~\new_[10208]_ ;
  assign \new_[5440]_  = ~\new_[6284]_  & ~\new_[9861]_ ;
  assign \new_[5441]_  = ~\new_[11894]_  | ~\new_[9963]_ ;
  assign \new_[5442]_  = ~\new_[6284]_  & ~\new_[10234]_ ;
  assign \new_[5443]_  = ~\new_[12738]_  & ~\new_[9894]_ ;
  assign \new_[5444]_  = ~\new_[6267]_  & ~\new_[9715]_ ;
  assign \new_[5445]_  = ~\new_[6284]_  & ~\new_[9838]_ ;
  assign \new_[5446]_  = ~\new_[11894]_  | ~\new_[9374]_ ;
  assign \new_[5447]_  = ~\new_[6284]_  & ~\new_[10155]_ ;
  assign \new_[5448]_  = ~\new_[11894]_  | ~\new_[9995]_ ;
  assign \new_[5449]_  = \new_[6283]_  | \new_[9623]_ ;
  assign \new_[5450]_  = \new_[6283]_  | \new_[9918]_ ;
  assign \new_[5451]_  = ~\new_[6267]_  & ~\new_[10057]_ ;
  assign \new_[5452]_  = ~\new_[6284]_  & ~\new_[9996]_ ;
  assign \new_[5453]_  = ~\new_[6284]_  & ~\new_[9908]_ ;
  assign \new_[5454]_  = ~\new_[6284]_  & ~\new_[9924]_ ;
  assign \new_[5455]_  = ~\new_[11894]_  | ~\new_[9418]_ ;
  assign \new_[5456]_  = ~\new_[12744]_  | ~\new_[10126]_ ;
  assign \new_[5457]_  = ~\new_[6284]_  & ~\new_[9941]_ ;
  assign \new_[5458]_  = ~\new_[11894]_  | ~\new_[10126]_ ;
  assign \new_[5459]_  = ~\new_[6284]_  & ~\new_[9866]_ ;
  assign \new_[5460]_  = ~\new_[6284]_  & ~\new_[9617]_ ;
  assign \new_[5461]_  = ~\new_[6284]_  & ~\new_[11865]_ ;
  assign \new_[5462]_  = ~\new_[6267]_  & ~\new_[9590]_ ;
  assign \new_[5463]_  = \new_[6284]_  | \new_[9590]_ ;
  assign \new_[5464]_  = ~\new_[12744]_  | ~\new_[9987]_ ;
  assign \new_[5465]_  = ~\new_[6284]_  & ~\new_[9738]_ ;
  assign \new_[5466]_  = ~\new_[11894]_  | ~\new_[9665]_ ;
  assign \new_[5467]_  = \new_[6202]_  & \new_[6203]_ ;
  assign \new_[5468]_  = ~\new_[11894]_  | ~\new_[9987]_ ;
  assign \new_[5469]_  = ~\new_[11894]_  | ~\new_[9958]_ ;
  assign \new_[5470]_  = ~\new_[12741]_  & ~\new_[9956]_ ;
  assign \new_[5471]_  = \new_[6283]_  | \new_[9956]_ ;
  assign \new_[5472]_  = \new_[6283]_  | \new_[9836]_ ;
  assign \new_[5473]_  = ~\new_[12738]_  & ~\new_[10101]_ ;
  assign \new_[5474]_  = ~\new_[6284]_  & ~\new_[10255]_ ;
  assign \new_[5475]_  = ~\new_[12693]_  | ~\new_[7326]_ ;
  assign \new_[5476]_  = ~\new_[11894]_  | ~\new_[9618]_ ;
  assign \new_[5477]_  = ~\new_[6284]_  & ~\new_[9304]_ ;
  assign \new_[5478]_  = ~\new_[6267]_  & ~\new_[9304]_ ;
  assign \new_[5479]_  = ~\new_[6267]_  & ~\new_[9305]_ ;
  assign \new_[5480]_  = ~\new_[6267]_  & ~\new_[9743]_ ;
  assign \new_[5481]_  = \new_[6256]_  & \new_[11434]_ ;
  assign \new_[5482]_  = ~\new_[6267]_  & ~\new_[9816]_ ;
  assign \new_[5483]_  = ~\new_[6284]_  & ~\new_[10166]_ ;
  assign \new_[5484]_  = ~\new_[11894]_  | ~\new_[10097]_ ;
  assign \new_[5485]_  = ~\new_[12739]_  | ~\new_[10083]_ ;
  assign \new_[5486]_  = ~\new_[6284]_  & ~\new_[9868]_ ;
  assign \new_[5487]_  = ~\new_[6267]_  & ~\new_[9868]_ ;
  assign \new_[5488]_  = \new_[6283]_  | \new_[9905]_ ;
  assign \new_[5489]_  = \new_[6283]_  | \new_[9714]_ ;
  assign \new_[5490]_  = ~\new_[6284]_  & ~\new_[9921]_ ;
  assign \new_[5491]_  = \new_[6283]_  | \new_[9859]_ ;
  assign \new_[5492]_  = \new_[6283]_  | \new_[9955]_ ;
  assign \new_[5493]_  = ~\new_[11894]_  | ~\new_[9707]_ ;
  assign \new_[5494]_  = \new_[6283]_  | \new_[9911]_ ;
  assign \new_[5495]_  = \new_[6283]_  | \new_[9739]_ ;
  assign \new_[5496]_  = ~\new_[11894]_  | ~\new_[9389]_ ;
  assign \new_[5497]_  = ~\new_[6284]_  & ~\new_[9742]_ ;
  assign \new_[5498]_  = ~\new_[6284]_  & ~\new_[12113]_ ;
  assign \new_[5499]_  = ~\new_[6267]_  & ~\new_[10167]_ ;
  assign \new_[5500]_  = ~\new_[7455]_  | (~\new_[12109]_  & ~\new_[10340]_ );
  assign \new_[5501]_  = ~\new_[7243]_  | (~\new_[7020]_  & ~\new_[9590]_ );
  assign \new_[5502]_  = ~\new_[6637]_  | (~\new_[6827]_  & ~\new_[9590]_ );
  assign \new_[5503]_  = (~\new_[6660]_  | ~\new_[10056]_ ) & (~\new_[7067]_  | ~\new_[9707]_ );
  assign \new_[5504]_  = (~\new_[12780]_  | ~\new_[10040]_ ) & (~\new_[11864]_  | ~\new_[9930]_ );
  assign \new_[5505]_  = ~\new_[6267]_  & ~\new_[9177]_ ;
  assign \new_[5506]_  = (~\new_[7059]_  | ~\new_[10043]_ ) & (~\new_[6321]_  | ~\new_[9294]_ );
  assign \new_[5507]_  = (~\new_[7059]_  | ~\new_[9953]_ ) & (~\new_[11553]_  | ~\new_[9118]_ );
  assign \new_[5508]_  = (~\new_[12783]_  | ~\new_[9596]_ ) & (~\new_[7571]_  | ~\new_[10136]_ );
  assign \new_[5509]_  = (~\new_[7059]_  | ~\new_[12060]_ ) & (~\new_[11553]_  | ~\new_[9089]_ );
  assign \new_[5510]_  = ~\new_[6777]_  & (~\new_[6657]_  | ~\new_[10054]_ );
  assign \new_[5511]_  = (~\new_[7059]_  | ~\new_[10054]_ ) & (~\new_[6321]_  | ~\new_[8873]_ );
  assign \new_[5512]_  = (~\new_[12784]_  | ~\new_[9584]_ ) & (~\new_[7571]_  | ~\new_[9401]_ );
  assign \new_[5513]_  = ~\new_[6789]_  & (~\new_[6656]_  | ~\new_[9620]_ );
  assign \new_[5514]_  = (~\new_[7213]_  & ~\new_[9190]_ ) | (~\new_[6720]_  & ~\new_[9159]_ );
  assign \new_[5515]_  = (~\new_[12784]_  | ~\new_[9587]_ ) & (~\new_[7571]_  | ~\new_[10099]_ );
  assign \new_[5516]_  = (~\new_[6346]_  | ~\new_[10827]_ ) & (~\new_[12774]_  | ~\new_[9401]_ );
  assign \new_[5517]_  = ~\new_[6779]_  & (~\new_[6657]_  | ~\new_[10065]_ );
  assign \new_[5518]_  = (~\new_[7059]_  | ~\new_[10065]_ ) & (~\new_[6321]_  | ~\new_[8897]_ );
  assign \new_[5519]_  = (~\new_[12784]_  | ~\new_[9588]_ ) & (~\new_[7571]_  | ~\new_[9661]_ );
  assign \new_[5520]_  = (~\new_[6346]_  | ~\new_[11348]_ ) & (~\new_[12777]_  | ~\new_[9661]_ );
  assign \new_[5521]_  = (~\new_[7059]_  | ~\new_[10053]_ ) & (~\new_[11553]_  | ~\new_[9330]_ );
  assign \new_[5522]_  = (~\new_[12783]_  | ~\new_[9933]_ ) & (~\new_[7571]_  | ~\new_[9963]_ );
  assign \new_[5523]_  = (~\new_[6346]_  | ~\new_[11576]_ ) & (~\new_[12768]_  | ~\new_[10128]_ );
  assign \new_[5524]_  = (~\new_[7059]_  | ~\new_[10046]_ ) & (~\new_[6664]_  | ~\new_[8863]_ );
  assign \new_[5525]_  = (~\new_[12784]_  | ~\new_[9592]_ ) & (~\new_[7239]_  | ~\new_[10104]_ );
  assign \new_[5526]_  = ~\new_[6782]_  & (~\new_[6657]_  | ~\new_[9822]_ );
  assign \new_[5527]_  = (~\new_[7059]_  | ~\new_[9822]_ ) & (~\new_[6664]_  | ~\new_[9082]_ );
  assign \new_[5528]_  = (~\new_[12784]_  | ~\new_[12293]_ ) & (~\new_[7571]_  | ~\new_[10128]_ );
  assign \new_[5529]_  = (~\new_[12783]_  | ~\new_[9929]_ ) & (~\new_[7239]_  | ~\new_[9607]_ );
  assign \new_[5530]_  = ~\new_[6783]_  & (~\new_[6657]_  | ~\new_[9854]_ );
  assign \new_[5531]_  = (~\new_[7059]_  | ~\new_[9854]_ ) & (~\new_[6664]_  | ~\new_[9077]_ );
  assign \new_[5532]_  = (~\new_[6346]_  | ~\new_[11340]_ ) & (~\new_[12779]_  | ~\new_[9845]_ );
  assign \new_[5533]_  = (~\new_[12784]_  | ~\new_[9960]_ ) & (~\new_[7239]_  | ~\new_[10011]_ );
  assign \new_[5534]_  = ~\new_[6784]_  & (~\new_[6657]_  | ~\new_[10078]_ );
  assign \new_[5535]_  = (~\new_[6346]_  | ~\new_[10243]_ ) & (~\new_[12773]_  | ~\new_[10237]_ );
  assign \new_[5536]_  = (~\new_[7059]_  | ~\new_[10078]_ ) & (~\new_[6664]_  | ~\new_[8898]_ );
  assign \new_[5537]_  = (~\new_[7059]_  | ~\new_[9880]_ ) & (~\new_[6664]_  | ~\new_[8902]_ );
  assign \new_[5538]_  = (~\new_[12784]_  | ~\new_[9603]_ ) & (~\new_[7571]_  | ~\new_[10263]_ );
  assign \new_[5539]_  = ~\new_[6787]_  & (~\new_[6657]_  | ~\new_[9849]_ );
  assign \new_[5540]_  = (~\new_[7059]_  | ~\new_[9849]_ ) & (~\new_[11553]_  | ~\new_[9324]_ );
  assign \new_[5541]_  = (~\new_[6346]_  | ~\new_[11316]_ ) & (~\new_[12770]_  | ~\new_[10287]_ );
  assign \new_[5542]_  = ~\new_[6788]_  & (~\new_[6657]_  | ~\new_[10081]_ );
  assign \new_[5543]_  = (~\new_[7059]_  | ~\new_[10081]_ ) & (~\new_[6664]_  | ~\new_[8943]_ );
  assign \new_[5544]_  = (~\new_[12783]_  | ~\new_[9678]_ ) & (~\new_[7571]_  | ~\new_[9845]_ );
  assign \new_[5545]_  = ~\new_[6790]_  & (~\new_[6657]_  | ~\new_[10130]_ );
  assign \new_[5546]_  = (~\new_[7059]_  | ~\new_[10130]_ ) & (~\new_[6321]_  | ~\new_[8895]_ );
  assign \new_[5547]_  = (~\new_[12784]_  | ~\new_[9489]_ ) & (~\new_[7239]_  | ~\new_[10237]_ );
  assign \new_[5548]_  = ~\new_[6791]_  & (~\new_[6657]_  | ~\new_[10082]_ );
  assign \new_[5549]_  = (~\new_[7059]_  | ~\new_[10082]_ ) & (~\new_[6664]_  | ~\new_[8868]_ );
  assign \new_[5550]_  = (~\new_[12784]_  | ~\new_[9593]_ ) & (~\new_[7571]_  | ~\new_[9660]_ );
  assign \new_[5551]_  = (~\new_[7059]_  | ~\new_[10061]_ ) & (~\new_[11553]_  | ~\new_[9092]_ );
  assign \new_[5552]_  = ~\new_[7201]_  & (~\new_[6660]_  | ~\new_[9668]_ );
  assign \new_[5553]_  = ~\new_[6793]_  & (~\new_[6657]_  | ~\new_[9807]_ );
  assign \new_[5554]_  = (~\new_[7059]_  | ~\new_[9610]_ ) & (~\new_[6664]_  | ~\new_[9579]_ );
  assign \new_[5555]_  = (~\new_[12784]_  | ~\new_[9601]_ ) & (~\new_[7571]_  | ~\new_[9641]_ );
  assign \new_[5556]_  = ~\new_[7055]_  & (~\new_[6656]_  | ~\new_[11504]_ );
  assign \new_[5557]_  = ~\new_[6792]_  & (~\new_[6657]_  | ~\new_[10071]_ );
  assign \new_[5558]_  = (~\new_[7059]_  | ~\new_[10071]_ ) & (~\new_[6321]_  | ~\new_[8904]_ );
  assign \new_[5559]_  = (~\new_[12784]_  | ~\new_[9585]_ ) & (~\new_[7239]_  | ~\new_[10287]_ );
  assign \new_[5560]_  = ~\new_[7203]_  & (~\new_[6659]_  | ~\new_[10089]_ );
  assign \new_[5561]_  = (~\new_[7059]_  | ~\new_[9694]_ ) & (~\new_[6321]_  | ~\new_[9114]_ );
  assign \new_[5562]_  = (~\new_[12786]_  | ~\new_[9937]_ ) & (~\new_[7344]_  | ~\new_[9340]_ );
  assign \new_[5563]_  = ~\new_[7057]_  & (~\new_[6660]_  | ~\new_[9649]_ );
  assign \new_[5564]_  = ~\new_[7205]_  & (~\new_[6659]_  | ~\new_[9965]_ );
  assign \new_[5565]_  = (~\new_[7059]_  | ~\new_[9965]_ ) & (~\new_[6664]_  | ~\new_[9358]_ );
  assign \new_[5566]_  = ~\new_[7206]_  & (~\new_[6659]_  | ~\new_[9856]_ );
  assign \new_[5567]_  = (~\new_[7059]_  | ~\new_[9856]_ ) & (~\new_[11553]_  | ~\new_[8906]_ );
  assign \new_[5568]_  = (~\new_[7059]_  | ~\new_[10055]_ ) & (~\new_[6321]_  | ~\new_[9823]_ );
  assign \new_[5569]_  = ~\new_[7208]_  & (~\new_[6659]_  | ~\new_[9841]_ );
  assign \new_[5570]_  = (~\new_[6346]_  | ~\new_[10419]_ ) & (~\new_[12768]_  | ~\new_[9599]_ );
  assign \new_[5571]_  = (~\new_[6346]_  | ~\new_[11526]_ ) & (~\new_[12771]_  | ~\new_[9604]_ );
  assign \new_[5572]_  = ~\new_[7210]_  & (~\new_[6659]_  | ~\new_[10087]_ );
  assign \new_[5573]_  = (~\new_[7059]_  | ~\new_[10118]_ ) & (~\new_[6321]_  | ~\new_[8907]_ );
  assign \new_[5574]_  = (~\new_[7059]_  | ~\new_[10087]_ ) & (~\new_[6664]_  | ~\new_[9338]_ );
  assign \new_[5575]_  = (~\new_[7059]_  | ~\new_[10153]_ ) & (~\new_[11553]_  | ~\new_[9646]_ );
  assign \new_[5576]_  = (~\new_[12784]_  | ~\new_[10084]_ ) & (~\new_[7239]_  | ~\new_[9655]_ );
  assign \new_[5577]_  = ~\new_[6801]_  & (~\new_[6657]_  | ~\new_[10118]_ );
  assign \new_[5578]_  = (~\new_[12783]_  | ~\new_[9614]_ ) & (~\new_[7239]_  | ~\new_[10019]_ );
  assign \new_[5579]_  = (~\new_[12783]_  | ~\new_[9586]_ ) & (~\new_[7239]_  | ~\new_[9618]_ );
  assign \new_[5580]_  = (~\new_[7059]_  | ~\new_[9904]_ ) & (~\new_[11553]_  | ~\new_[9123]_ );
  assign \new_[5581]_  = (~\new_[7059]_  | ~\new_[9839]_ ) & (~\new_[6664]_  | ~\new_[9093]_ );
  assign \new_[5582]_  = (~\new_[7059]_  | ~\new_[10044]_ ) & (~\new_[6321]_  | ~\new_[9293]_ );
  assign \new_[5583]_  = (~\new_[7059]_  | ~\new_[9846]_ ) & (~\new_[6321]_  | ~\new_[9085]_ );
  assign \new_[5584]_  = ~\new_[6279]_  | (~\new_[6720]_  & ~\new_[9291]_ );
  assign \new_[5585]_  = ~\new_[6276]_  | (~\new_[6720]_  & ~\new_[9049]_ );
  assign \new_[5586]_  = ~\new_[6798]_  & (~\new_[6656]_  | ~\new_[9847]_ );
  assign \new_[5587]_  = (~\new_[7059]_  | ~\new_[9847]_ ) & (~\new_[11553]_  | ~\new_[9295]_ );
  assign \new_[5588]_  = (~\new_[12783]_  | ~\new_[9824]_ ) & (~\new_[7571]_  | ~\new_[9980]_ );
  assign \new_[5589]_  = ~\new_[6797]_  & (~\new_[6656]_  | ~\new_[9967]_ );
  assign \new_[5590]_  = ~\new_[7232]_  & (~\new_[6658]_  | ~\new_[10051]_ );
  assign \new_[5591]_  = ~\new_[6799]_  & (~\new_[6657]_  | ~\new_[9871]_ );
  assign \new_[5592]_  = ~\new_[6278]_  | (~\new_[6720]_  & ~\new_[9084]_ );
  assign \new_[5593]_  = ~\new_[7223]_  & (~\new_[6658]_  | ~\new_[10015]_ );
  assign \new_[5594]_  = (~\new_[7059]_  | ~\new_[10015]_ ) & (~\new_[6321]_  | ~\new_[9292]_ );
  assign \new_[5595]_  = ~\new_[7224]_  & (~\new_[6658]_  | ~\new_[10044]_ );
  assign \new_[5596]_  = ~\new_[7218]_  & (~\new_[6658]_  | ~\new_[10127]_ );
  assign \new_[5597]_  = ~\new_[6800]_  & (~\new_[6657]_  | ~\new_[10050]_ );
  assign \new_[5598]_  = ~\new_[7228]_  & (~\new_[6659]_  | ~\new_[10049]_ );
  assign \new_[5599]_  = (~\new_[7059]_  | ~\new_[10049]_ ) & (~\new_[6321]_  | ~\new_[9378]_ );
  assign \new_[5600]_  = (~\new_[7059]_  | ~\new_[10050]_ ) & (~\new_[6664]_  | ~\new_[8931]_ );
  assign \new_[5601]_  = (~\new_[12784]_  | ~\new_[9408]_ ) & (~\new_[7571]_  | ~\new_[9599]_ );
  assign \new_[5602]_  = ~\new_[6794]_  & (~\new_[6657]_  | ~\new_[10140]_ );
  assign \new_[5603]_  = (~\new_[7059]_  | ~\new_[10140]_ ) & (~\new_[6664]_  | ~\new_[8923]_ );
  assign \new_[5604]_  = (~\new_[12784]_  | ~\new_[11521]_ ) & (~\new_[7239]_  | ~\new_[9604]_ );
  assign \new_[5605]_  = (~\new_[12783]_  | ~\new_[9746]_ ) & (~\new_[7571]_  | ~\new_[9389]_ );
  assign \new_[5606]_  = ~\new_[7230]_  & (~\new_[6659]_  | ~\new_[10043]_ );
  assign \new_[5607]_  = ~\new_[7231]_  & (~\new_[6659]_  | ~\new_[10048]_ );
  assign \new_[5608]_  = ~\new_[6803]_  & (~\new_[6657]_  | ~\new_[10107]_ );
  assign \new_[5609]_  = ~\new_[7068]_  & (~\new_[6660]_  | ~\new_[9608]_ );
  assign \new_[5610]_  = (~\new_[7059]_  | ~\new_[9608]_ ) & (~\new_[11553]_  | ~\new_[9349]_ );
  assign \new_[5611]_  = (~\new_[12784]_  | ~\new_[9874]_ ) & (~\new_[7571]_  | ~\new_[9989]_ );
  assign \new_[5612]_  = (~\new_[7059]_  | ~\new_[10107]_ ) & (~\new_[6664]_  | ~\new_[8908]_ );
  assign \new_[5613]_  = (~\new_[12784]_  | ~\new_[9393]_ ) & (~\new_[7571]_  | ~\new_[9407]_ );
  assign \new_[5614]_  = (~\new_[7059]_  | ~\new_[10063]_ ) & (~\new_[6321]_  | ~\new_[9323]_ );
  assign \new_[5615]_  = (~\new_[12784]_  | ~\new_[9863]_ ) & (~\new_[7571]_  | ~\new_[10037]_ );
  assign \new_[5616]_  = ~\new_[7070]_  & (~\new_[6656]_  | ~\new_[9953]_ );
  assign \new_[5617]_  = ~\new_[6291]_  | ~\wb_addr_i[25] ;
  assign \new_[5618]_  = ~\new_[11894]_  | ~\new_[9655]_ ;
  assign \new_[5619]_  = ~\new_[12171]_  | ~\new_[12665]_  | ~\new_[6317]_ ;
  assign \new_[5620]_  = ~\new_[12771]_  | ~\new_[9388]_ ;
  assign \new_[5621]_  = ~\new_[6663]_  & ~\new_[6786]_ ;
  assign \new_[5622]_  = ~\new_[12747]_  | ~\new_[9620]_ ;
  assign \new_[5623]_  = ~\new_[12775]_  | ~\new_[9707]_ ;
  assign \new_[5624]_  = ~\new_[6809]_  & ~\new_[7235]_ ;
  assign \new_[5625]_  = ~\new_[12747]_  | ~\new_[11504]_ ;
  assign \new_[5626]_  = ~\new_[6374]_  | ~\new_[6285]_ ;
  assign \new_[5627]_  = ~\new_[12771]_  | ~\new_[9684]_ ;
  assign \new_[5628]_  = ~\new_[12747]_  | ~\new_[9594]_ ;
  assign \new_[5629]_  = ~\new_[6088]_  | ~\new_[11355]_ ;
  assign \new_[5630]_  = ~\new_[6088]_  | ~\new_[10963]_ ;
  assign \new_[5631]_  = ~\new_[6088]_  | ~\new_[12453]_ ;
  assign \new_[5632]_  = ~\new_[6087]_  | ~\new_[11313]_ ;
  assign \new_[5633]_  = ~\new_[6087]_  | ~\new_[9946]_ ;
  assign \new_[5634]_  = ~\new_[6088]_  | ~\new_[10509]_ ;
  assign \new_[5635]_  = ~\new_[6305]_  & (~\new_[7288]_  | ~\wb_addr_i[21] );
  assign n2871 = (~\new_[6377]_  & ~\new_[8707]_  & ~\new_[8720]_ ) | (~\new_[10305]_  & ~\new_[8231]_  & ~\new_[10501]_ );
  assign \new_[5637]_  = ~\new_[5242]_ ;
  assign \new_[5638]_  = \new_[5242]_ ;
  assign \new_[5639]_  = ~\new_[12239]_ ;
  assign \new_[5640]_  = ~u5_pack_le2_reg;
  assign \new_[5641]_  = ~\new_[6070]_  & ~\new_[3439]_ ;
  assign \new_[5642]_  = ~\new_[12532]_  & ~\new_[10957]_ ;
  assign \new_[5643]_  = ~\new_[6029]_ ;
  assign \new_[5644]_  = ~\new_[6666]_  | ~\wb_addr_i[24] ;
  assign \new_[5645]_  = ~\new_[3138]_  | ~\new_[11102]_  | ~\new_[6095]_  | ~\new_[10877]_ ;
  assign \new_[5646]_  = ~\new_[6034]_ ;
  assign \new_[5647]_  = ~\new_[10846]_  | ~\new_[11553]_  | ~\new_[9659]_ ;
  assign \new_[5648]_  = ~\new_[6035]_ ;
  assign \new_[5649]_  = ~\new_[6063]_  & (~\new_[11731]_  | ~\new_[7827]_ );
  assign \new_[5650]_  = ~\new_[12741]_  & ~\new_[9836]_ ;
  assign \new_[5651]_  = ~\new_[6070]_ ;
  assign \new_[5652]_  = ~\new_[6072]_ ;
  assign \new_[5653]_  = ~\new_[6317]_  & (~\new_[6950]_  | ~\new_[12003]_ );
  assign \new_[5654]_  = ~\new_[6316]_  & (~\new_[6951]_  | ~\new_[10258]_ );
  assign \new_[5655]_  = ~\new_[6316]_  & (~\new_[7137]_  | ~\new_[9718]_ );
  assign \new_[5656]_  = ~\new_[6317]_  & (~\new_[6952]_  | ~\new_[10208]_ );
  assign \new_[5657]_  = ~\new_[6317]_  & (~\new_[6953]_  | ~\new_[9861]_ );
  assign \new_[5658]_  = ~\new_[6317]_  & (~\new_[6954]_  | ~\new_[10229]_ );
  assign \new_[5659]_  = ~\new_[6316]_  & (~\new_[7138]_  | ~\new_[9867]_ );
  assign \new_[5660]_  = ~\new_[6317]_  & (~\new_[7139]_  | ~\new_[10146]_ );
  assign \new_[5661]_  = ~\new_[6317]_  & (~\new_[6956]_  | ~\new_[10234]_ );
  assign \new_[5662]_  = ~\new_[6316]_  & (~\new_[6957]_  | ~\new_[10256]_ );
  assign \new_[5663]_  = ~\new_[6316]_  & (~\new_[6958]_  | ~\new_[9894]_ );
  assign \new_[5664]_  = ~\new_[6316]_  & (~\new_[6959]_  | ~\new_[9922]_ );
  assign \new_[5665]_  = ~\new_[6316]_  & (~\new_[6960]_  | ~\new_[9838]_ );
  assign \new_[5666]_  = ~\new_[6317]_  & (~\new_[6961]_  | ~\new_[10340]_ );
  assign \new_[5667]_  = ~\new_[6316]_  & (~\new_[7142]_  | ~\new_[10155]_ );
  assign \new_[5668]_  = ~\new_[6317]_  & (~\new_[6963]_  | ~\new_[10254]_ );
  assign \new_[5669]_  = ~\new_[6317]_  & (~\new_[6964]_  | ~\new_[10057]_ );
  assign \new_[5670]_  = ~\new_[6317]_  & (~\new_[7144]_  | ~\new_[9996]_ );
  assign \new_[5671]_  = ~\new_[6316]_  & (~\new_[6965]_  | ~\new_[9908]_ );
  assign \new_[5672]_  = \new_[6379]_  | \new_[6316]_ ;
  assign \new_[5673]_  = ~\new_[6316]_  & (~\new_[7145]_  | ~\new_[9866]_ );
  assign \new_[5674]_  = ~\new_[6349]_  & (~\new_[7608]_  | ~\new_[10793]_ );
  assign \new_[5675]_  = ~\new_[6317]_  & (~\new_[6966]_  | ~\new_[9617]_ );
  assign \new_[5676]_  = ~\new_[6316]_  & (~\new_[7146]_  | ~\new_[10262]_ );
  assign \new_[5677]_  = ~\new_[6317]_  & (~\new_[6967]_  | ~\new_[11865]_ );
  assign \new_[5678]_  = \new_[6380]_  | \new_[6316]_ ;
  assign \new_[5679]_  = ~\new_[6317]_  & (~\new_[7147]_  | ~\new_[9345]_ );
  assign \new_[5680]_  = ~\new_[6317]_  & (~\new_[7148]_  | ~\new_[9691]_ );
  assign \new_[5681]_  = ~\new_[6316]_  & (~\new_[7149]_  | ~\new_[9956]_ );
  assign \new_[5682]_  = ~\new_[6316]_  & (~\new_[6894]_  | ~\new_[10101]_ );
  assign \new_[5683]_  = ~\new_[6316]_  & (~\new_[6979]_  | ~\new_[9836]_ );
  assign \new_[5684]_  = ~\new_[6316]_  & (~\new_[6955]_  | ~\new_[9927]_ );
  assign \new_[5685]_  = ~\new_[6317]_  & (~\new_[7133]_  | ~\new_[9954]_ );
  assign \new_[5686]_  = ~\new_[6316]_  & (~\new_[7046]_  | ~\new_[10150]_ );
  assign \new_[5687]_  = ~\new_[6317]_  & (~\new_[7071]_  | ~\new_[9177]_ );
  assign \new_[5688]_  = ~\new_[6316]_  & (~\new_[7162]_  | ~\new_[10255]_ );
  assign \new_[5689]_  = ~\new_[6317]_  & (~\new_[6970]_  | ~\new_[9653]_ );
  assign \new_[5690]_  = ~\new_[6317]_  & (~\new_[6973]_  | ~\new_[9305]_ );
  assign \new_[5691]_  = ~\new_[6317]_  & (~\new_[6974]_  | ~\new_[9372]_ );
  assign \new_[5692]_  = ~\new_[6316]_  & (~\new_[7153]_  | ~\new_[9717]_ );
  assign \new_[5693]_  = ~\new_[11808]_  | ~\new_[12727]_  | ~\new_[6465]_  | ~\new_[12650]_ ;
  assign \new_[5694]_  = ~\new_[6316]_  & (~\new_[6977]_  | ~\new_[9623]_ );
  assign \new_[5695]_  = ~\new_[6339]_  | (~\new_[2136]_  & ~\new_[12619]_ );
  assign \new_[5696]_  = ~\new_[6316]_  & (~\new_[7122]_  | ~\new_[9918]_ );
  assign \new_[5697]_  = ~\new_[6316]_  & (~\new_[6980]_  | ~\new_[9905]_ );
  assign \new_[5698]_  = ~\new_[6316]_  & (~\new_[6981]_  | ~\new_[10172]_ );
  assign \new_[5699]_  = ~\new_[6316]_  & (~\new_[6962]_  | ~\new_[9714]_ );
  assign \new_[5700]_  = ~\new_[6316]_  & (~\new_[6983]_  | ~\new_[9921]_ );
  assign \new_[5701]_  = ~\new_[6340]_  | ~\new_[6673]_ ;
  assign \new_[5702]_  = ~\new_[6317]_  & (~\new_[7140]_  | ~\new_[9911]_ );
  assign \new_[5703]_  = ~\new_[6338]_  | (~\new_[2134]_  & ~\new_[12622]_ );
  assign \new_[5704]_  = ~\new_[6316]_  & (~\new_[6988]_  | ~\new_[9925]_ );
  assign \new_[5705]_  = ~\new_[6316]_  & (~\new_[7158]_  | ~\new_[9713]_ );
  assign \new_[5706]_  = ~\new_[6317]_  & (~\new_[6989]_  | ~\new_[12113]_ );
  assign \new_[5707]_  = ~\new_[6317]_  & (~\new_[6990]_  | ~\new_[10166]_ );
  assign \new_[5708]_  = ~\new_[6316]_  & (~\new_[6991]_  | ~\new_[9732]_ );
  assign \new_[5709]_  = ~\new_[6316]_  & (~\new_[6992]_  | ~\new_[10199]_ );
  assign \new_[5710]_  = ~\new_[6077]_ ;
  assign \new_[5711]_  = ~\new_[6365]_  & (~\new_[7874]_  | ~\new_[2055]_ );
  assign \new_[5712]_  = (~\new_[6687]_  | ~\new_[11778]_ ) & (~\new_[2055]_  | ~\new_[11779]_ );
  assign \new_[5713]_  = (~\new_[6687]_  | ~\new_[7772]_ ) & (~\new_[10278]_  | ~\new_[7992]_ );
  assign \new_[5714]_  = (~\new_[11450]_  & ~\new_[10522]_ ) | (~\new_[12240]_  & ~\new_[11505]_ );
  assign \new_[5715]_  = ~\new_[6348]_  | (~\new_[7863]_  & ~\new_[9302]_ );
  assign \new_[5716]_  = (~\new_[7081]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[9587]_ );
  assign \new_[5717]_  = (~\new_[7082]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[9933]_ );
  assign \new_[5718]_  = (~\new_[7084]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[12293]_ );
  assign \new_[5719]_  = (~\new_[7085]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[9929]_ );
  assign \new_[5720]_  = (~\new_[7094]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[9593]_ );
  assign \new_[5721]_  = (~\new_[7096]_  | ~\new_[6683]_ ) & (~\new_[7995]_  | ~\new_[9615]_ );
  assign \new_[5722]_  = (~\new_[7097]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[9601]_ );
  assign \new_[5723]_  = ~\new_[7533]_  | ~\new_[6356]_ ;
  assign \new_[5724]_  = ~\new_[7535]_  | ~\new_[6357]_ ;
  assign \new_[5725]_  = ~\new_[7389]_  | ~\new_[6358]_ ;
  assign \new_[5726]_  = (~\new_[7251]_  | ~\new_[6683]_ ) & (~\new_[7995]_  | ~\new_[9602]_ );
  assign \new_[5727]_  = ~\new_[7209]_  | ~\new_[6360]_ ;
  assign \new_[5728]_  = (~\new_[7252]_  | ~\new_[6682]_ ) & (~\new_[7682]_  | ~\new_[10210]_ );
  assign \new_[5729]_  = (~\new_[7253]_  | ~\new_[6682]_ ) & (~\new_[7682]_  | ~\new_[9865]_ );
  assign \new_[5730]_  = (~\new_[7254]_  | ~\new_[6683]_ ) & (~\new_[7682]_  | ~\new_[9906]_ );
  assign \new_[5731]_  = (~\new_[7255]_  | ~\new_[6683]_ ) & (~\new_[7682]_  | ~\new_[9837]_ );
  assign \new_[5732]_  = (~\new_[7257]_  | ~\new_[6682]_ ) & (~\new_[7682]_  | ~\new_[9857]_ );
  assign \new_[5733]_  = ~\new_[7529]_  | ~\new_[6361]_ ;
  assign \new_[5734]_  = (~\new_[7250]_  | ~\new_[6682]_ ) & (~\new_[7682]_  | ~\new_[9663]_ );
  assign \new_[5735]_  = (~\new_[7108]_  | ~\new_[6682]_ ) & (~\new_[7682]_  | ~\new_[9862]_ );
  assign \new_[5736]_  = (~\new_[6813]_  | ~\new_[6682]_ ) & (~\new_[7995]_  | ~\new_[9840]_ );
  assign \new_[5737]_  = ~\new_[7225]_  | ~\new_[6369]_ ;
  assign \new_[5738]_  = (~\new_[7099]_  | ~\new_[6682]_ ) & (~\new_[7995]_  | ~\new_[9818]_ );
  assign \new_[5739]_  = ~\new_[7198]_  | ~\new_[6371]_ ;
  assign \new_[5740]_  = ~\new_[7217]_  | ~\new_[6372]_ ;
  assign \new_[5741]_  = (~\new_[7086]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[11521]_ );
  assign \new_[5742]_  = ~\new_[7544]_  | ~\new_[6373]_ ;
  assign \new_[5743]_  = (~\new_[7248]_  | ~\new_[6682]_ ) & (~\new_[7682]_  | ~\new_[11928]_ );
  assign \new_[5744]_  = (~\new_[6819]_  | ~\new_[6684]_ ) & (~\new_[7995]_  | ~\new_[9863]_ );
  assign \new_[5745]_  = ~\new_[7546]_  | ~\new_[6375]_ ;
  assign \new_[5746]_  = \new_[7528]_  | \new_[6347]_ ;
  assign \new_[5747]_  = ~\new_[11894]_  | ~\new_[9853]_ ;
  assign \new_[5748]_  = ~\new_[6540]_  | ~\new_[6733]_ ;
  assign \new_[5749]_  = ~\new_[7627]_  & ~\new_[12656]_ ;
  assign \new_[5750]_  = ~\new_[12064]_  | ~\new_[9985]_ ;
  assign \new_[5751]_  = ~\new_[6394]_  & ~\new_[9190]_ ;
  assign \new_[5752]_  = ~\new_[6384]_  | ~\new_[11772]_ ;
  assign \new_[5753]_  = ~\new_[12064]_  | ~\new_[10244]_ ;
  assign \new_[5754]_  = ~\new_[12064]_  | ~\new_[9694]_ ;
  assign \new_[5755]_  = ~\new_[12064]_  | ~\new_[9965]_ ;
  assign \new_[5756]_  = ~\new_[12064]_  | ~\new_[9856]_ ;
  assign \new_[5757]_  = ~\new_[12064]_  | ~\new_[10055]_ ;
  assign \new_[5758]_  = ~\new_[12064]_  | ~\new_[9841]_ ;
  assign \new_[5759]_  = ~\new_[12064]_  | ~\new_[9610]_ ;
  assign \new_[5760]_  = ~\new_[12064]_  | ~\new_[9843]_ ;
  assign \new_[5761]_  = ~\new_[12064]_  | ~\new_[10087]_ ;
  assign \new_[5762]_  = ~\new_[12064]_  | ~\new_[9846]_ ;
  assign \new_[5763]_  = ~\new_[11439]_  & ~\new_[6972]_ ;
  assign \new_[5764]_  = ~\new_[12064]_  | ~\new_[9606]_ ;
  assign \new_[5765]_  = ~\new_[6457]_  | ~\new_[7175]_ ;
  assign \new_[5766]_  = ~\new_[6461]_  | ~\new_[10200]_ ;
  assign \new_[5767]_  = ~\new_[12064]_  | ~\new_[9872]_ ;
  assign \new_[5768]_  = ~\new_[12064]_  | ~\new_[10051]_ ;
  assign \new_[5769]_  = ~\new_[12064]_  | ~\new_[10015]_ ;
  assign \new_[5770]_  = ~\new_[12064]_  | ~\new_[10044]_ ;
  assign \new_[5771]_  = ~\new_[12064]_  | ~\new_[9870]_ ;
  assign \new_[5772]_  = ~\new_[12064]_  | ~\new_[10127]_ ;
  assign \new_[5773]_  = ~\new_[7091]_  | ~\new_[6393]_ ;
  assign \new_[5774]_  = ~\new_[12064]_  | ~\new_[10049]_ ;
  assign \new_[5775]_  = ~\new_[12064]_  | ~\new_[10056]_ ;
  assign \new_[5776]_  = ~\new_[12064]_  | ~\new_[10059]_ ;
  assign \new_[5777]_  = ~\new_[12064]_  | ~\new_[10089]_ ;
  assign \new_[5778]_  = ~\new_[12064]_  | ~\new_[10043]_ ;
  assign \new_[5779]_  = ~\new_[12064]_  | ~\new_[10048]_ ;
  assign \new_[5780]_  = ~\new_[8219]_  & ~\new_[6535]_ ;
  assign \new_[5781]_  = (~\new_[6741]_  | ~\new_[7825]_ ) & (~\new_[11306]_  | ~\new_[7481]_ );
  assign \new_[5782]_  = (~\new_[7049]_  | ~\new_[7823]_ ) & (~\new_[11306]_  | ~\new_[7648]_ );
  assign \new_[5783]_  = (~\new_[6743]_  | ~\new_[7777]_ ) & (~\new_[11306]_  | ~\new_[7766]_ );
  assign \new_[5784]_  = (~\new_[6755]_  | ~\new_[7825]_ ) & (~\new_[11306]_  | ~\new_[7650]_ );
  assign \new_[5785]_  = \new_[12700]_  | \new_[7752]_ ;
  assign \new_[5786]_  = \new_[6397]_  & \new_[9822]_ ;
  assign \new_[5787]_  = (~\new_[7048]_  | ~\new_[7777]_ ) & (~\new_[11306]_  | ~\new_[7767]_ );
  assign \new_[5788]_  = (~\new_[6757]_  | ~\new_[7777]_ ) & (~\new_[11306]_  | ~\new_[7490]_ );
  assign \new_[5789]_  = ~\new_[6541]_  & (~\new_[12385]_  | ~\new_[10040]_ );
  assign \new_[5790]_  = \new_[12701]_  | \new_[7753]_ ;
  assign \new_[5791]_  = (~\new_[7050]_  | ~\new_[7994]_ ) & (~\new_[11306]_  | ~\new_[7653]_ );
  assign \new_[5792]_  = \new_[12700]_  | \new_[7754]_ ;
  assign \new_[5793]_  = \new_[12700]_  | \new_[7755]_ ;
  assign \new_[5794]_  = (~\new_[7051]_  | ~\new_[7823]_ ) & (~\new_[11306]_  | ~\new_[7647]_ );
  assign \new_[5795]_  = \new_[12705]_  | \new_[7756]_ ;
  assign \new_[5796]_  = (~\new_[6762]_  | ~\new_[7777]_ ) & (~\new_[11306]_  | ~\new_[7656]_ );
  assign \new_[5797]_  = \new_[12701]_  | \new_[7757]_ ;
  assign \new_[5798]_  = (~\new_[6770]_  | ~\new_[7777]_ ) & (~\new_[11306]_  | ~\new_[7499]_ );
  assign \new_[5799]_  = (~\new_[6742]_  | ~\new_[7825]_ ) & (~\new_[11306]_  | ~\new_[7658]_ );
  assign \new_[5800]_  = ~\new_[8001]_  | ~\new_[11449]_  | ~\new_[6735]_ ;
  assign \new_[5801]_  = \new_[12709]_  | \new_[7758]_ ;
  assign \new_[5802]_  = ~\new_[12376]_  & ~\new_[12613]_ ;
  assign \new_[5803]_  = (~\new_[6771]_  | ~\new_[7825]_ ) & (~\new_[11306]_  | ~\new_[7659]_ );
  assign \new_[5804]_  = (~\new_[7047]_  | ~\new_[7823]_ ) & (~\new_[11306]_  | ~\new_[7652]_ );
  assign n2921 = (~\new_[6737]_  | ~\new_[12780]_ ) & (~\new_[7066]_  | ~\new_[12606]_ );
  assign \new_[5806]_  = ~\new_[6539]_  & (~\new_[7540]_  | ~\new_[9906]_ );
  assign \new_[5807]_  = ~\new_[6463]_  | (~\new_[7174]_  & ~\new_[7807]_ );
  assign \new_[5808]_  = ~\new_[6691]_  & (~\new_[6663]_  | ~\new_[9978]_ );
  assign \new_[5809]_  = ~\new_[6475]_  & (~\new_[3176]_  | ~\new_[6832]_ );
  assign \new_[5810]_  = ~\new_[6476]_  & (~\new_[3179]_  | ~\new_[7366]_ );
  assign \new_[5811]_  = ~\new_[6477]_  & (~\new_[3145]_  | ~\new_[7366]_ );
  assign \new_[5812]_  = ~\new_[6478]_  & (~\new_[3041]_  | ~\new_[7366]_ );
  assign \new_[5813]_  = ~\new_[6481]_  & (~\new_[3138]_  | ~\new_[6832]_ );
  assign \new_[5814]_  = ~\new_[6482]_  & (~\new_[11102]_  | ~\new_[6832]_ );
  assign \new_[5815]_  = ~\new_[6483]_  & (~\new_[11114]_  | ~\new_[6832]_ );
  assign \new_[5816]_  = ~\new_[6492]_  & (~\new_[3225]_  | ~\new_[6832]_ );
  assign \new_[5817]_  = ~\new_[6480]_  & (~\new_[3042]_  | ~\new_[6832]_ );
  assign \new_[5818]_  = ~\new_[7326]_  | ~\new_[12782]_  | ~\new_[11895]_  | ~\new_[12694]_ ;
  assign \new_[5819]_  = (~\new_[12070]_  & ~\new_[10258]_ ) | (~\new_[6720]_  & ~\new_[9642]_ );
  assign \new_[5820]_  = (~\new_[12455]_  | ~\new_[8919]_ ) & (~\new_[12783]_  | ~\new_[12306]_ );
  assign \new_[5821]_  = (~\new_[12070]_  & ~\new_[12113]_ ) | (~\new_[6720]_  & ~\new_[9664]_ );
  assign \new_[5822]_  = ~\new_[11894]_  | ~\new_[9479]_ ;
  assign \new_[5823]_  = \new_[3145]_  ^ \new_[6718]_ ;
  assign \new_[5824]_  = ~\new_[11302]_  | ~\new_[7649]_ ;
  assign \new_[5825]_  = ~\new_[11305]_  | ~\new_[7510]_ ;
  assign \new_[5826]_  = ~\new_[11305]_  | ~\new_[7487]_ ;
  assign \new_[5827]_  = ~\new_[11306]_  | ~\new_[7491]_ ;
  assign \new_[5828]_  = ~\new_[11305]_  | ~\new_[7492]_ ;
  assign \new_[5829]_  = ~\new_[11302]_  | ~\new_[7497]_ ;
  assign \new_[5830]_  = ~\new_[11306]_  | ~\new_[7503]_ ;
  assign \new_[5831]_  = ~\new_[11305]_  | ~\new_[7514]_ ;
  assign \new_[5832]_  = ~\new_[11306]_  | ~\new_[7507]_ ;
  assign \new_[5833]_  = \new_[6641]_  & \new_[12109]_ ;
  assign \new_[5834]_  = ~\new_[11305]_  | ~\new_[7513]_ ;
  assign \new_[5835]_  = ~\new_[11305]_  | ~\new_[7315]_ ;
  assign \new_[5836]_  = ~\new_[11303]_  | ~\new_[7515]_ ;
  assign \new_[5837]_  = ~\new_[11305]_  | ~\new_[7769]_ ;
  assign \new_[5838]_  = ~\new_[11303]_  | ~\new_[7518]_ ;
  assign \new_[5839]_  = \new_[6639]_  & \new_[12499]_ ;
  assign \new_[5840]_  = \new_[6639]_  & \new_[6337]_ ;
  assign \new_[5841]_  = ~\new_[11894]_  | ~\new_[10136]_ ;
  assign \new_[5842]_  = ~\new_[11894]_  | ~\new_[9979]_ ;
  assign \new_[5843]_  = \new_[6640]_  | \new_[10208]_ ;
  assign \new_[5844]_  = ~\new_[7102]_  | ~\new_[7298]_ ;
  assign \new_[5845]_  = ~\new_[11894]_  | ~\new_[10099]_ ;
  assign \new_[5846]_  = ~\new_[11894]_  | ~\new_[9661]_ ;
  assign \new_[5847]_  = ~\new_[11894]_  | ~\new_[10104]_ ;
  assign \new_[5848]_  = ~\new_[11894]_  | ~\new_[10128]_ ;
  assign \new_[5849]_  = ~\new_[11894]_  | ~\new_[8805]_ ;
  assign \new_[5850]_  = ~\new_[11894]_  | ~\new_[10011]_ ;
  assign \new_[5851]_  = ~\new_[11894]_  | ~\new_[9680]_ ;
  assign \new_[5852]_  = ~\new_[11894]_  | ~\new_[10263]_ ;
  assign \new_[5853]_  = ~\new_[11894]_  | ~\new_[9845]_ ;
  assign \new_[5854]_  = ~\new_[11894]_  | ~\new_[10237]_ ;
  assign \new_[5855]_  = ~\new_[11894]_  | ~\new_[9660]_ ;
  assign \new_[5856]_  = ~\new_[11894]_  | ~\new_[9641]_ ;
  assign \new_[5857]_  = ~\new_[11894]_  | ~\new_[10287]_ ;
  assign \new_[5858]_  = ~\new_[11894]_  | ~\new_[9936]_ ;
  assign \new_[5859]_  = ~\new_[11053]_  | ~\new_[6621]_ ;
  assign \new_[5860]_  = ~\new_[11894]_  | ~\new_[9326]_ ;
  assign \new_[5861]_  = \new_[6640]_  | \new_[9177]_ ;
  assign \new_[5862]_  = ~\new_[11894]_  | ~\new_[10019]_ ;
  assign \new_[5863]_  = ~\new_[11894]_  | ~\new_[9950]_ ;
  assign \new_[5864]_  = \new_[6640]_  | \new_[9305]_ ;
  assign \new_[5865]_  = ~\new_[6460]_ ;
  assign \new_[5866]_  = \new_[6640]_  | \new_[9715]_ ;
  assign \new_[5867]_  = ~\new_[11894]_  | ~\new_[9595]_ ;
  assign \new_[5868]_  = ~\new_[11894]_  | ~\new_[10137]_ ;
  assign \new_[5869]_  = ~\new_[10349]_  & ~\new_[6621]_ ;
  assign \new_[5870]_  = ~\new_[10003]_  & ~\new_[6621]_ ;
  assign \new_[5871]_  = \new_[10121]_  | \new_[6621]_ ;
  assign \new_[5872]_  = ~\new_[11894]_  | ~\new_[10083]_ ;
  assign \new_[5873]_  = ~\new_[11894]_  | ~\new_[9709]_ ;
  assign \new_[5874]_  = ~\new_[11894]_  | ~\new_[9567]_ ;
  assign \new_[5875]_  = ~\new_[11894]_  | ~\new_[9599]_ ;
  assign \new_[5876]_  = ~\new_[7176]_  | ~\new_[12070]_ ;
  assign \new_[5877]_  = ~\new_[11894]_  | ~\new_[9407]_ ;
  assign \new_[5878]_  = ~\new_[11335]_  | ~\new_[12094]_  | ~\new_[6327]_  | ~\new_[10456]_ ;
  assign \new_[5879]_  = ~\new_[6376]_  | ~\new_[7181]_ ;
  assign \new_[5880]_  = ~\new_[11062]_  | ~\new_[12691]_  | ~\new_[8413]_ ;
  assign \new_[5881]_  = ~\new_[6617]_  | ~\new_[10200]_ ;
  assign \new_[5882]_  = (~\new_[9817]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[9108]_ );
  assign \new_[5883]_  = (~\new_[9160]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9958]_ );
  assign \new_[5884]_  = (~\new_[8894]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9326]_ );
  assign \new_[5885]_  = (~\new_[9062]_  | ~\new_[7109]_ ) & (~\new_[7215]_  | ~\new_[9611]_ );
  assign \new_[5886]_  = (~\new_[9280]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9853]_ );
  assign \new_[5887]_  = (~\new_[8801]_  | ~\new_[7560]_ ) & (~\new_[7215]_  | ~\new_[9644]_ );
  assign \new_[5888]_  = (~\new_[9067]_  | ~\new_[7560]_ ) & (~\new_[7215]_  | ~\new_[9582]_ );
  assign \new_[5889]_  = (~\new_[8888]_  | ~\new_[7560]_ ) & (~\new_[7060]_  | ~\new_[9479]_ );
  assign \new_[5890]_  = (~\new_[9072]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[9655]_ );
  assign \new_[5891]_  = (~\new_[8803]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[8977]_ );
  assign \new_[5892]_  = (~\new_[9075]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[10137]_ );
  assign \new_[5893]_  = (~\new_[8885]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[9168]_ );
  assign \new_[5894]_  = (~\new_[8792]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9657]_ );
  assign \new_[5895]_  = (~\new_[9165]_  | ~\new_[7109]_ ) & (~\new_[7215]_  | ~\new_[9682]_ );
  assign \new_[5896]_  = (~\new_[9066]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9374]_ );
  assign \new_[5897]_  = (~\new_[9892]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[10097]_ );
  assign \new_[5898]_  = ~\new_[6730]_  & (~\new_[6663]_  | ~\new_[10083]_ );
  assign \new_[5899]_  = (~\new_[9273]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9675]_ );
  assign \new_[5900]_  = (~\new_[9086]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9709]_ );
  assign \new_[5901]_  = (~\new_[9274]_  | ~\new_[7109]_ ) & (~\new_[7215]_  | ~\new_[10115]_ );
  assign \new_[5902]_  = (~\new_[9070]_  | ~\new_[7109]_ ) & (~\new_[7215]_  | ~\new_[9567]_ );
  assign \new_[5903]_  = (~\new_[9390]_  | ~\new_[7109]_ ) & (~\new_[7215]_  | ~\new_[9707]_ );
  assign \new_[5904]_  = (~\new_[9348]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9684]_ );
  assign \new_[5905]_  = (~\new_[9282]_  | ~\new_[7109]_ ) & (~\new_[7215]_  | ~\new_[9389]_ );
  assign \new_[5906]_  = (~\new_[9276]_  | ~\new_[7560]_ ) & (~\new_[7060]_  | ~\new_[9665]_ );
  assign \new_[5907]_  = (~\new_[9821]_  | ~\new_[7109]_ ) & (~\new_[6826]_  | ~\new_[10031]_ );
  assign \new_[5908]_  = ~\new_[6159]_ ;
  assign \new_[5909]_  = ~\new_[6624]_  | ~\new_[7073]_ ;
  assign \new_[5910]_  = (~\new_[6810]_  | ~\new_[10059]_ ) & (~\new_[7067]_  | ~\new_[9684]_ );
  assign \new_[5911]_  = (~\new_[11719]_  | ~\wb_addr_i[23] ) & (~\new_[11725]_  | ~\wb_addr_i[22] );
  assign \new_[5912]_  = (~\new_[12780]_  | ~\new_[9616]_ ) & (~\new_[11864]_  | ~\new_[8977]_ );
  assign \new_[5913]_  = (~\new_[11719]_  | ~\wb_addr_i[24] ) & (~\new_[6804]_  | ~\wb_addr_i[23] );
  assign \new_[5914]_  = (~\new_[12780]_  | ~\new_[11515]_ ) & (~\new_[11864]_  | ~\new_[9107]_ );
  assign \new_[5915]_  = (~\new_[12385]_  | ~\new_[9844]_ ) & (~\new_[11864]_  | ~\new_[9391]_ );
  assign \new_[5916]_  = ~\new_[7188]_  & (~\new_[6810]_  | ~\new_[11787]_ );
  assign \new_[5917]_  = (~\new_[12783]_  | ~\new_[9591]_ ) & (~\new_[7571]_  | ~\new_[9979]_ );
  assign \new_[5918]_  = (~\new_[12592]_  | ~\new_[10291]_ ) & (~\new_[12773]_  | ~\new_[9383]_ );
  assign \new_[5919]_  = (~\new_[11997]_  | ~\new_[9587]_ ) & (~\new_[6665]_  | ~\new_[10099]_ );
  assign \new_[5920]_  = (~\new_[12592]_  | ~\new_[10922]_ ) & (~\new_[12779]_  | ~\new_[10031]_ );
  assign \new_[5921]_  = ~\new_[6780]_  & (~\new_[7008]_  | ~\new_[10053]_ );
  assign \new_[5922]_  = ~\new_[6781]_  & (~\new_[7008]_  | ~\new_[10046]_ );
  assign \new_[5923]_  = ~\new_[7193]_  & (~\new_[6810]_  | ~\new_[9737]_ );
  assign \new_[5924]_  = (~\new_[11997]_  | ~\new_[9929]_ ) & (~\new_[6665]_  | ~\new_[8805]_ );
  assign \new_[5925]_  = (~\new_[12592]_  | ~\new_[11492]_ ) & (~\new_[12779]_  | ~\new_[9930]_ );
  assign \new_[5926]_  = ~\new_[6785]_  & (~\new_[7008]_  | ~\new_[9880]_ );
  assign \new_[5927]_  = (~\new_[12784]_  | ~\new_[9842]_ ) & (~\new_[7571]_  | ~\new_[9995]_ );
  assign \new_[5928]_  = ~\new_[7195]_  & (~\new_[6810]_  | ~\new_[9848]_ );
  assign \new_[5929]_  = ~\new_[7196]_  & (~\new_[6810]_  | ~\new_[10244]_ );
  assign \new_[5930]_  = ~\new_[6776]_  & (~\new_[7008]_  | ~\new_[10061]_ );
  assign \new_[5931]_  = (~\new_[12783]_  | ~\new_[9621]_ ) & (~\new_[7239]_  | ~\new_[9418]_ );
  assign \new_[5932]_  = (~\new_[12592]_  | ~\new_[10496]_ ) & (~\new_[12779]_  | ~\new_[8977]_ );
  assign \new_[5933]_  = (~\new_[12786]_  | ~\new_[10064]_ ) & (~\new_[7571]_  | ~\new_[10111]_ );
  assign \new_[5934]_  = (~\new_[12592]_  | ~\new_[12054]_ ) & (~\new_[12774]_  | ~\new_[9682]_ );
  assign \new_[5935]_  = (~\new_[12786]_  | ~\new_[9864]_ ) & (~\new_[7571]_  | ~\new_[11860]_ );
  assign \new_[5936]_  = (~\new_[12592]_  | ~\new_[10250]_ ) & (~\new_[12779]_  | ~\new_[9107]_ );
  assign \new_[5937]_  = (~\new_[12593]_  | ~\new_[12755]_ ) & (~\new_[12779]_  | ~\new_[9391]_ );
  assign \new_[5938]_  = (~\new_[12783]_  | ~\new_[9855]_ ) & (~\new_[7344]_  | ~\new_[9958]_ );
  assign \new_[5939]_  = ~\new_[7207]_  & (~\new_[6810]_  | ~\new_[10055]_ );
  assign \new_[5940]_  = (~\new_[12783]_  | ~\new_[10210]_ ) & (~\new_[7344]_  | ~\new_[9611]_ );
  assign \new_[5941]_  = (~\new_[7059]_  | ~\new_[9841]_ ) & (~\new_[6664]_  | ~\new_[9321]_ );
  assign \new_[5942]_  = (~\new_[12783]_  | ~\new_[9865]_ ) & (~\new_[7571]_  | ~\new_[9853]_ );
  assign \new_[5943]_  = ~\new_[7233]_  & (~\new_[6810]_  | ~\new_[9610]_ );
  assign \new_[5944]_  = (~\new_[12783]_  | ~\new_[9969]_ ) & (~\new_[7344]_  | ~\new_[9644]_ );
  assign \new_[5945]_  = ~\new_[7192]_  & (~\new_[6810]_  | ~\new_[9843]_ );
  assign \new_[5946]_  = (~\new_[7059]_  | ~\new_[9843]_ ) & (~\new_[6664]_  | ~\new_[9329]_ );
  assign \new_[5947]_  = (~\new_[12783]_  | ~\new_[9906]_ ) & (~\new_[7344]_  | ~\new_[9582]_ );
  assign \new_[5948]_  = (~\new_[12783]_  | ~\new_[9837]_ ) & (~\new_[7344]_  | ~\new_[9479]_ );
  assign \new_[5949]_  = ~\new_[6795]_  & (~\new_[7008]_  | ~\new_[10153]_ );
  assign \new_[5950]_  = ~\new_[7211]_  & (~\new_[6810]_  | ~\new_[9985]_ );
  assign \new_[5951]_  = ~\new_[7212]_  & (~\new_[6810]_  | ~\new_[11452]_ );
  assign \new_[5952]_  = ~\new_[6796]_  & (~\new_[7008]_  | ~\new_[9904]_ );
  assign \new_[5953]_  = ~\new_[7064]_  & (~\new_[7008]_  | ~\new_[9839]_ );
  assign \new_[5954]_  = (~\new_[11997]_  | ~\new_[9589]_ ) & (~\new_[6665]_  | ~\new_[9657]_ );
  assign \new_[5955]_  = ~\new_[7199]_  & (~\new_[6810]_  | ~\new_[9846]_ );
  assign \new_[5956]_  = (~\new_[12783]_  | ~\new_[9857]_ ) & (~\new_[7344]_  | ~\new_[9682]_ );
  assign \new_[5957]_  = ~\new_[7194]_  & (~\new_[6810]_  | ~\new_[9606]_ );
  assign \new_[5958]_  = ~\new_[7202]_  & (~\new_[6810]_  | ~\new_[9970]_ );
  assign \new_[5959]_  = ~\new_[7221]_  & (~\new_[6810]_  | ~\new_[9872]_ );
  assign \new_[5960]_  = (~\new_[7059]_  | ~\new_[9872]_ ) & (~\new_[6664]_  | ~\new_[9102]_ );
  assign \new_[5961]_  = (~\new_[12784]_  | ~\new_[9663]_ ) & (~\new_[7571]_  | ~\new_[9374]_ );
  assign \new_[5962]_  = (~\new_[12784]_  | ~\new_[9613]_ ) & (~\new_[7571]_  | ~\new_[9978]_ );
  assign \new_[5963]_  = (~\new_[7059]_  | ~\new_[10051]_ ) & (~\new_[6664]_  | ~\new_[9117]_ );
  assign \new_[5964]_  = (~\new_[12783]_  | ~\new_[9581]_ ) & (~\new_[7344]_  | ~\new_[10097]_ );
  assign \new_[5965]_  = (~\new_[12784]_  | ~\new_[9609]_ ) & (~\new_[7571]_  | ~\new_[9710]_ );
  assign \new_[5966]_  = (~\new_[12783]_  | ~\new_[9862]_ ) & (~\new_[7344]_  | ~\new_[9675]_ );
  assign \new_[5967]_  = (~\new_[12784]_  | ~\new_[9840]_ ) & (~\new_[7571]_  | ~\new_[9709]_ );
  assign \new_[5968]_  = (~\new_[11997]_  | ~\new_[10062]_ ) & (~\new_[6665]_  | ~\new_[9619]_ );
  assign \new_[5969]_  = ~\new_[11894]_  | ~\new_[9611]_ ;
  assign \new_[5970]_  = (~\new_[12784]_  | ~\new_[9818]_ ) & (~\new_[7571]_  | ~\new_[9567]_ );
  assign \new_[5971]_  = (~\new_[12783]_  | ~\new_[9850]_ ) & (~\new_[7344]_  | ~\new_[10137]_ );
  assign \new_[5972]_  = (~\new_[12784]_  | ~\new_[10047]_ ) & (~\new_[7571]_  | ~\new_[12110]_ );
  assign \new_[5973]_  = (~\new_[7059]_  | ~\new_[10048]_ ) & (~\new_[6664]_  | ~\new_[9346]_ );
  assign \new_[5974]_  = (~\new_[12783]_  | ~\new_[11928]_ ) & (~\new_[7344]_  | ~\new_[9665]_ );
  assign \new_[5975]_  = ~\new_[6802]_  & (~\new_[7008]_  | ~\new_[10063]_ );
  assign \new_[5976]_  = (~\new_[11997]_  | ~\new_[9393]_ ) & (~\new_[6665]_  | ~\new_[9407]_ );
  assign \new_[5977]_  = u5_wb_wait_r_reg;
  assign \new_[5978]_  = ~\new_[12751]_  | (~\new_[8831]_  & ~\new_[9854]_ );
  assign \new_[5979]_  = ~\new_[12748]_  | ~\new_[10048]_ ;
  assign \new_[5980]_  = ~\new_[12751]_  | ~\new_[10265]_ ;
  assign \new_[5981]_  = \new_[7263]_  | \new_[7063]_ ;
  assign \new_[5982]_  = ~\new_[7263]_  | ~\new_[7662]_ ;
  assign \new_[5983]_  = ~\new_[11337]_  | ~\new_[7777]_  | ~\new_[6670]_ ;
  assign \new_[5984]_  = ~\new_[12747]_  | ~\new_[9848]_ ;
  assign \new_[5985]_  = ~\new_[12751]_  | ~\new_[10244]_ ;
  assign \new_[5986]_  = ~\new_[12747]_  | ~\new_[10061]_ ;
  assign \new_[5987]_  = ~\new_[9913]_  | ~\new_[7823]_  | ~\new_[6670]_ ;
  assign \new_[5988]_  = ~\new_[7077]_  | ~\new_[10111]_ ;
  assign \new_[5989]_  = ~\new_[7077]_  | ~\new_[11860]_ ;
  assign \new_[5990]_  = ~\new_[12751]_  | ~\new_[9694]_ ;
  assign \new_[5991]_  = ~\new_[12747]_  | ~\new_[9904]_ ;
  assign \new_[5992]_  = ~\new_[12751]_  | ~\new_[10043]_ ;
  assign \new_[5993]_  = \new_[6655]_  | \new_[7863]_ ;
  assign \new_[5994]_  = ~\new_[12751]_  & ~\new_[11864]_ ;
  assign \new_[5995]_  = ~\new_[10411]_  | ~\new_[7777]_  | ~\new_[7286]_ ;
  assign \new_[5996]_  = ~\new_[12054]_  | ~\new_[7777]_  | ~\new_[7286]_ ;
  assign \new_[5997]_  = ~\new_[7074]_  | ~\new_[6837]_ ;
  assign \new_[5998]_  = ~\new_[7077]_  | ~\new_[9980]_ ;
  assign \new_[5999]_  = ~\new_[12748]_  | ~\new_[9872]_ ;
  assign \new_[6000]_  = ~\new_[12751]_  | ~\new_[10015]_ ;
  assign \new_[6001]_  = ~\new_[10051]_  | ~\new_[12751]_ ;
  assign \new_[6002]_  = ~\new_[11328]_  | ~\new_[7777]_  | ~\new_[7286]_ ;
  assign \new_[6003]_  = ~\new_[12751]_  | ~\new_[9870]_ ;
  assign \new_[6004]_  = ~\new_[12749]_  | ~\new_[10059]_ ;
  assign \new_[6005]_  = ~\new_[7077]_  | ~\new_[12110]_ ;
  assign \new_[6006]_  = ~\new_[11323]_  | ~\new_[7777]_  | ~\new_[6670]_ ;
  assign \new_[6007]_  = ~\new_[11310]_  | ~\new_[7777]_  | ~\new_[7286]_ ;
  assign \new_[6008]_  = ~\new_[10212]_  | ~\new_[6833]_  | ~\new_[4147]_  | ~\new_[10468]_ ;
  assign \new_[6009]_  = ~\new_[7059]_  | ~\new_[11787]_ ;
  assign \new_[6010]_  = ~\new_[7059]_  | ~\new_[9985]_ ;
  assign \new_[6011]_  = ~\new_[10922]_  | ~\new_[12653]_  | ~\new_[8748]_ ;
  assign \new_[6012]_  = ~\new_[7059]_  | ~\new_[10056]_ ;
  assign \new_[6013]_  = ~\new_[7059]_  | ~\new_[10244]_ ;
  assign \new_[6014]_  = ~\new_[7059]_  | ~\new_[11452]_ ;
  assign \new_[6015]_  = ~\new_[12528]_  & ~\new_[7295]_ ;
  assign \new_[6016]_  = ~\new_[12089]_  | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6017]_  = ~\new_[9785]_  | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6018]_  = ~\new_[12453]_  | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6019]_  = ~\new_[10496]_  | ~\new_[12653]_  | ~\new_[8748]_ ;
  assign \new_[6020]_  = ~\new_[7059]_  | ~\new_[9606]_ ;
  assign \new_[6021]_  = ~\new_[10250]_  | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6022]_  = ~\new_[7059]_  | ~\new_[9970]_ ;
  assign \new_[6023]_  = ~\new_[12755]_  | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6024]_  = ~\new_[7059]_  | ~\new_[9870]_ ;
  assign \new_[6025]_  = ~\new_[7059]_  | ~\new_[10059]_ ;
  assign \new_[6026]_  = ~\new_[9585]_  & (~\new_[11727]_  | ~\new_[6662]_ );
  assign \new_[6027]_  = ~\new_[9969]_  & (~\new_[6836]_  | ~\new_[6662]_ );
  assign n2916 = ~\new_[6315]_  | (~\new_[7695]_  & ~\new_[7915]_ );
  assign \new_[6029]_  = \new_[9202]_  & \new_[6327]_ ;
  assign \new_[6030]_  = ~\new_[11894]_  | ~\new_[9582]_ ;
  assign \new_[6031]_  = \new_[6641]_  | \new_[10150]_ ;
  assign \new_[6032]_  = ~\new_[7263]_  | ~n3451;
  assign \new_[6033]_  = \new_[6720]_  | \new_[8896]_ ;
  assign \new_[6034]_  = ~\new_[6290]_ ;
  assign \new_[6035]_  = \new_[6291]_ ;
  assign \new_[6036]_  = ~\new_[6809]_ ;
  assign \new_[6037]_  = ~\new_[8983]_  | ~\new_[11553]_ ;
  assign \new_[6038]_  = (~\wb_addr_i[0]  | ~\new_[7288]_ ) & (~\wb_addr_i[1]  | ~\new_[6836]_ );
  assign \new_[6039]_  = (~\wb_addr_i[1]  | ~\new_[7288]_ ) & (~\new_[11264]_  | ~\wb_addr_i[3] );
  assign \new_[6040]_  = ~\new_[7288]_  | ~\wb_addr_i[10] ;
  assign \new_[6041]_  = ~\new_[6834]_  | ~\new_[7074]_  | ~\new_[6837]_ ;
  assign \new_[6042]_  = ~\new_[7288]_  | ~\wb_addr_i[5] ;
  assign \new_[6043]_  = ~\new_[6672]_  | ~\wb_addr_i[7] ;
  assign \new_[6044]_  = ~\new_[6672]_  | ~\wb_addr_i[6] ;
  assign \new_[6045]_  = ~\new_[6672]_  | ~\wb_addr_i[3] ;
  assign \new_[6046]_  = ~\new_[6672]_  | ~\wb_addr_i[17] ;
  assign \new_[6047]_  = ~\new_[7288]_  | ~\wb_addr_i[11] ;
  assign \new_[6048]_  = ~\new_[6672]_  | ~\wb_addr_i[13] ;
  assign \new_[6049]_  = ~\new_[6672]_  | ~\wb_addr_i[14] ;
  assign \new_[6050]_  = ~\new_[6672]_  | ~\wb_addr_i[16] ;
  assign \new_[6051]_  = ~\new_[6672]_  | ~\wb_addr_i[15] ;
  assign \new_[6052]_  = ~\new_[7288]_  | ~\wb_addr_i[19] ;
  assign \new_[6053]_  = ~\new_[7288]_  | ~\wb_addr_i[20] ;
  assign \new_[6054]_  = ~\new_[6672]_  | ~\wb_addr_i[22] ;
  assign \new_[6055]_  = ~\new_[6672]_  | ~\wb_addr_i[23] ;
  assign \new_[6056]_  = ~\new_[6672]_  | ~\wb_addr_i[2] ;
  assign \new_[6057]_  = ~\new_[6672]_  | ~\wb_addr_i[18] ;
  assign \new_[6058]_  = ~\new_[6672]_  | ~\wb_addr_i[4] ;
  assign \new_[6059]_  = ~\new_[7288]_  | ~\wb_addr_i[9] ;
  assign \new_[6060]_  = ~\new_[6672]_  | ~\wb_addr_i[12] ;
  assign n2926 = \new_[7288]_  & \new_[10164]_ ;
  assign \new_[6062]_  = ~\new_[7288]_  | ~\wb_addr_i[8] ;
  assign \new_[6063]_  = ~\new_[6322]_ ;
  assign \new_[6064]_  = ~\new_[6835]_ ;
  assign \new_[6065]_  = n2936 | \new_[4340]_ ;
  assign \new_[6066]_  = n2936 | \new_[4341]_ ;
  assign \new_[6067]_  = n2936 | \new_[4237]_ ;
  assign \new_[6068]_  = ~\new_[12506]_  | ~\new_[11162]_ ;
  assign \new_[6069]_  = ~\new_[12506]_  | ~\new_[11081]_ ;
  assign \new_[6070]_  = ~n2936 | ~\new_[7632]_ ;
  assign \new_[6071]_  = ~n2936 & ~\new_[7632]_ ;
  assign \new_[6072]_  = (~\new_[11418]_  & ~\new_[3036]_ ) | (~\new_[12516]_  & ~\new_[12515]_ );
  assign \new_[6073]_  = ~\new_[6676]_  & ~\new_[12075]_ ;
  assign \new_[6074]_  = (~\new_[7245]_  | ~\new_[11453]_ ) & (~\new_[8806]_  | ~\new_[7539]_ );
  assign \new_[6075]_  = ~\new_[6374]_ ;
  assign \new_[6076]_  = \new_[2115]_  ? \new_[12622]_  : \new_[2093]_ ;
  assign \new_[6077]_  = ~\new_[11713]_  | ~\new_[8875]_  | ~\new_[7000]_ ;
  assign \new_[6078]_  = (~\new_[7080]_  | ~\new_[11453]_ ) & (~\new_[7682]_  | ~\new_[12000]_ );
  assign \new_[6079]_  = (~\new_[7354]_  | ~\new_[11453]_ ) & (~\new_[7682]_  | ~\new_[9938]_ );
  assign \new_[6080]_  = (~\new_[7355]_  | ~\new_[11453]_ ) & (~\new_[7995]_  | ~\new_[10040]_ );
  assign \new_[6081]_  = (~\new_[7104]_  | ~\new_[11453]_ ) & (~\new_[7682]_  | ~\new_[10084]_ );
  assign \new_[6082]_  = (~\new_[7106]_  | ~\new_[11453]_ ) & (~\new_[7682]_  | ~\new_[9616]_ );
  assign \new_[6083]_  = (~\new_[7361]_  | ~\new_[11453]_ ) & (~\new_[7682]_  | ~\new_[9589]_ );
  assign \new_[6084]_  = (~\new_[7362]_  | ~\new_[11453]_ ) & (~\new_[7995]_  | ~\new_[11515]_ );
  assign \new_[6085]_  = (~\new_[7360]_  | ~\new_[11453]_ ) & (~\new_[7682]_  | ~\new_[9844]_ );
  assign \new_[6086]_  = ~\new_[6343]_ ;
  assign \new_[6087]_  = ~\new_[6344]_ ;
  assign \new_[6088]_  = ~\new_[6345]_ ;
  assign \new_[6089]_  = ~\new_[6343]_ ;
  assign \new_[6090]_  = ~\new_[6343]_ ;
  assign \new_[6091]_  = ~\new_[10291]_  | ~\new_[12695]_  | ~\new_[11814]_ ;
  assign \new_[6092]_  = ~\new_[7247]_  | ~\new_[6683]_ ;
  assign \new_[6093]_  = ~\new_[7249]_  | ~\new_[6683]_ ;
  assign \new_[6094]_  = ~\new_[7095]_  | ~\new_[6683]_ ;
  assign \new_[6095]_  = ~\new_[6359]_ ;
  assign \new_[6096]_  = ~\new_[7256]_  | ~\new_[6683]_ ;
  assign \new_[6097]_  = ~\new_[7999]_  | ~\new_[7296]_  | ~\new_[7180]_ ;
  assign \new_[6098]_  = ~\new_[12109]_  | ~\new_[12170]_  | ~\new_[6283]_ ;
  assign \new_[6099]_  = ~\new_[7258]_  | ~\new_[6683]_ ;
  assign \new_[6100]_  = ~\new_[7259]_  | ~\new_[6683]_ ;
  assign \new_[6101]_  = ~\new_[8001]_  | ~\new_[12236]_  | ~\new_[6735]_  | ~\new_[11449]_ ;
  assign \new_[6102]_  = ~\new_[9308]_  & (~\new_[7370]_  | ~\new_[7479]_ );
  assign \new_[6103]_  = ~\new_[7168]_  & (~\new_[7017]_  | ~\new_[7498]_ );
  assign \new_[6104]_  = ~\new_[7294]_  & (~\new_[7017]_  | ~\new_[7504]_ );
  assign \new_[6105]_  = (~\new_[7293]_  | ~\new_[7289]_ ) & (~\new_[7059]_  | ~\new_[10265]_ );
  assign \new_[6106]_  = (~\new_[12455]_  | ~\new_[10265]_ ) & (~\new_[12786]_  | ~\new_[10102]_ );
  assign \new_[6107]_  = ~\new_[3042]_  | ~\new_[3138]_  | ~\new_[6718]_  | ~\new_[10931]_ ;
  assign \new_[6108]_  = \new_[7759]_  | \new_[12687]_ ;
  assign \new_[6109]_  = ~\new_[11306]_  | ~\new_[7496]_ ;
  assign \new_[6110]_  = ~\new_[11306]_  | ~\new_[7501]_ ;
  assign \new_[6111]_  = ~\new_[11306]_  | ~\new_[7505]_ ;
  assign \new_[6112]_  = ~\new_[6735]_  & (~\new_[10268]_  | ~\new_[12274]_ );
  assign \new_[6113]_  = \new_[7301]_  | \new_[6722]_ ;
  assign \new_[6114]_  = ~\new_[12735]_  & ~\new_[6722]_ ;
  assign \new_[6115]_  = ~\new_[11894]_  | ~\new_[9109]_ ;
  assign \new_[6116]_  = ~\new_[11439]_ ;
  assign \new_[6117]_  = ~\new_[11894]_  | ~\new_[10111]_ ;
  assign \new_[6118]_  = ~\new_[11894]_  | ~\new_[11860]_ ;
  assign \new_[6119]_  = ~\new_[11894]_  | (~\new_[11776]_  & ~\new_[10955]_ );
  assign \new_[6120]_  = u5_dv_r_reg;
  assign \new_[6121]_  = ~\new_[7419]_  & ~\new_[6723]_ ;
  assign \new_[6122]_  = ~\new_[7305]_  | ~\new_[12384]_ ;
  assign \new_[6123]_  = \new_[6733]_  & \new_[12384]_ ;
  assign \new_[6124]_  = (~\new_[9241]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[9979]_ );
  assign \new_[6125]_  = (~\new_[8890]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9401]_ );
  assign \new_[6126]_  = (~\new_[9279]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[10099]_ );
  assign \new_[6127]_  = (~\new_[9281]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[9661]_ );
  assign \new_[6128]_  = (~\new_[8710]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9963]_ );
  assign \new_[6129]_  = (~\new_[9275]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[10104]_ );
  assign \new_[6130]_  = (~\new_[9277]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[10128]_ );
  assign \new_[6131]_  = (~\new_[8802]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[8805]_ );
  assign \new_[6132]_  = (~\new_[8882]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[10011]_ );
  assign \new_[6133]_  = (~\new_[9141]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[9388]_ );
  assign \new_[6134]_  = (~\new_[8921]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9680]_ );
  assign \new_[6135]_  = (~\new_[9065]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[10263]_ );
  assign \new_[6136]_  = (~\new_[9188]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9995]_ );
  assign \new_[6137]_  = (~\new_[8884]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[9845]_ );
  assign \new_[6138]_  = (~\new_[9068]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[10237]_ );
  assign \new_[6139]_  = (~\new_[9071]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9660]_ );
  assign \new_[6140]_  = (~\new_[8883]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9641]_ );
  assign \new_[6141]_  = (~\new_[8926]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[10052]_ );
  assign \new_[6142]_  = (~\new_[9032]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[10019]_ );
  assign \new_[6143]_  = (~\new_[9073]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[9391]_ );
  assign \new_[6144]_  = (~\new_[9047]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[9595]_ );
  assign \new_[6145]_  = (~\new_[8892]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9978]_ );
  assign \new_[6146]_  = (~\new_[9573]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[10083]_ );
  assign \new_[6147]_  = (~\new_[8930]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9619]_ );
  assign \new_[6148]_  = (~\new_[8887]_  | ~\new_[7109]_ ) & (~\new_[7216]_  | ~\new_[9599]_ );
  assign \new_[6149]_  = (~\new_[9278]_  | ~\new_[7109]_ ) & (~\new_[7061]_  | ~\new_[9604]_ );
  assign \new_[6150]_  = (~\new_[9169]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[9407]_ );
  assign \new_[6151]_  = (~\new_[9069]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[10037]_ );
  assign \new_[6152]_  = (~\new_[9328]_  | ~\new_[7109]_ ) & (~\new_[7060]_  | ~\new_[10136]_ );
  assign \new_[6153]_  = ~\new_[7586]_  | (~\new_[11774]_  & ~\new_[10208]_ );
  assign \new_[6154]_  = (~\new_[9284]_  | ~\new_[12790]_ ) & (~\new_[7077]_  | ~\new_[10011]_ );
  assign \new_[6155]_  = ~\new_[7556]_  | (~\new_[7020]_  & ~\new_[9177]_ );
  assign \new_[6156]_  = ~\new_[7475]_  | (~\new_[7075]_  & ~\new_[10150]_ );
  assign \new_[6157]_  = ~\new_[7569]_  | (~\new_[7020]_  & ~\new_[9305]_ );
  assign \new_[6158]_  = ~\new_[7555]_  | (~\new_[11774]_  & ~\new_[9715]_ );
  assign \new_[6159]_  = ~\new_[6540]_ ;
  assign \new_[6160]_  = ~\new_[7053]_  & (~\new_[7067]_  | ~\new_[10039]_ );
  assign \new_[6161]_  = ~\new_[6778]_  & (~\new_[7329]_  | ~\new_[10099]_ );
  assign \new_[6162]_  = (~\new_[12780]_  | ~\new_[9938]_ ) & (~\new_[11864]_  | ~\new_[10031]_ );
  assign \new_[6163]_  = (~\new_[12385]_  | ~\new_[9937]_ ) & (~\new_[7060]_  | ~\new_[9936]_ );
  assign \new_[6164]_  = ~\new_[7161]_  | ~\new_[7323]_  | ~\new_[7370]_  | ~\new_[7111]_ ;
  assign \new_[6165]_  = (~\new_[11997]_  | ~\new_[9591]_ ) & (~\new_[6826]_  | ~\new_[9979]_ );
  assign \new_[6166]_  = (~\new_[11997]_  | ~\new_[10102]_ ) & (~\new_[6826]_  | ~\new_[10039]_ );
  assign \new_[6167]_  = (~\new_[11997]_  | ~\new_[9584]_ ) & (~\new_[12002]_  | ~\new_[9401]_ );
  assign \new_[6168]_  = (~\new_[11997]_  | ~\new_[9588]_ ) & (~\new_[12002]_  | ~\new_[9661]_ );
  assign \new_[6169]_  = (~\new_[11997]_  | ~\new_[9933]_ ) & (~\new_[12002]_  | ~\new_[9963]_ );
  assign \new_[6170]_  = (~\new_[11997]_  | ~\new_[9592]_ ) & (~\new_[12002]_  | ~\new_[10104]_ );
  assign \new_[6171]_  = (~\new_[11997]_  | ~\new_[12293]_ ) & (~\new_[6828]_  | ~\new_[10128]_ );
  assign \new_[6172]_  = (~\new_[11997]_  | ~\new_[9960]_ ) & (~\new_[6828]_  | ~\new_[10011]_ );
  assign \new_[6173]_  = (~\new_[11997]_  | ~\new_[9612]_ ) & (~\new_[6828]_  | ~\new_[9680]_ );
  assign \new_[6174]_  = (~\new_[11997]_  | ~\new_[9603]_ ) & (~\new_[6828]_  | ~\new_[10263]_ );
  assign \new_[6175]_  = (~\new_[11997]_  | ~\new_[9842]_ ) & (~\new_[12002]_  | ~\new_[9995]_ );
  assign \new_[6176]_  = (~\new_[7059]_  | ~\new_[9848]_ ) & (~\new_[11553]_  | ~\new_[9577]_ );
  assign \new_[6177]_  = (~\new_[11997]_  | ~\new_[9678]_ ) & (~\new_[12002]_  | ~\new_[9845]_ );
  assign \new_[6178]_  = (~\new_[11997]_  | ~\new_[9489]_ ) & (~\new_[6828]_  | ~\new_[10237]_ );
  assign \new_[6179]_  = (~\new_[11997]_  | ~\new_[9593]_ ) & (~\new_[6828]_  | ~\new_[9660]_ );
  assign \new_[6180]_  = (~\new_[11997]_  | ~\new_[9601]_ ) & (~\new_[12002]_  | ~\new_[9641]_ );
  assign \new_[6181]_  = (~\new_[11997]_  | ~\new_[10064]_ ) & (~\new_[6826]_  | ~\new_[10111]_ );
  assign \new_[6182]_  = (~\new_[7059]_  | ~\new_[11504]_ ) & (~\new_[11553]_  | ~\new_[9640]_ );
  assign \new_[6183]_  = (~\new_[11997]_  | ~\new_[9585]_ ) & (~\new_[6828]_  | ~\new_[10052]_ );
  assign \new_[6184]_  = (~\new_[11997]_  | ~\new_[9863]_ ) & (~\new_[6828]_  | ~\new_[10037]_ );
  assign \new_[6185]_  = (~\new_[11997]_  | ~\new_[9864]_ ) & (~\new_[6826]_  | ~\new_[11860]_ );
  assign \new_[6186]_  = (~\new_[7059]_  | ~\new_[10045]_ ) & (~\new_[11553]_  | ~\new_[9285]_ );
  assign \new_[6187]_  = ~\new_[7204]_  & (~\new_[7008]_  | ~\new_[9694]_ );
  assign \new_[6188]_  = (~\new_[11997]_  | ~\new_[9602]_ ) & (~\new_[6826]_  | ~\new_[9987]_ );
  assign \new_[6189]_  = (~\new_[11997]_  | ~\new_[9614]_ ) & (~\new_[6828]_  | ~\new_[10019]_ );
  assign \new_[6190]_  = (~\new_[11997]_  | ~\new_[9613]_ ) & (~\new_[12002]_  | ~\new_[9978]_ );
  assign \new_[6191]_  = (~\new_[11997]_  | ~\new_[9408]_ ) & (~\new_[6828]_  | ~\new_[9599]_ );
  assign \new_[6192]_  = (~\new_[11997]_  | ~\new_[9824]_ ) & (~\new_[6826]_  | ~\new_[9980]_ );
  assign \new_[6193]_  = (~\new_[11997]_  | ~\new_[9609]_ ) & (~\new_[6828]_  | ~\new_[10083]_ );
  assign \new_[6194]_  = (~\new_[7059]_  | ~\new_[10127]_ ) & (~\new_[11553]_  | ~\new_[9575]_ );
  assign \new_[6195]_  = (~\new_[11997]_  | ~\new_[11962]_ ) & (~\new_[6826]_  | ~\new_[9684]_ );
  assign \new_[6196]_  = (~\new_[11997]_  | ~\new_[11521]_ ) & (~\new_[6828]_  | ~\new_[9604]_ );
  assign \new_[6197]_  = (~\new_[11997]_  | ~\new_[9850]_ ) & (~\new_[6826]_  | ~\new_[10137]_ );
  assign \new_[6198]_  = (~\new_[11997]_  | ~\new_[10047]_ ) & (~\new_[6826]_  | ~\new_[12110]_ );
  assign \new_[6199]_  = (~\new_[11997]_  | ~\new_[11928]_ ) & (~\new_[6826]_  | ~\new_[9665]_ );
  assign \new_[6200]_  = (~\new_[11997]_  | ~\new_[9874]_ ) & (~\new_[6826]_  | ~\new_[9990]_ );
  assign \new_[6201]_  = (~\new_[11997]_  | ~\new_[9596]_ ) & (~\new_[6826]_  | ~\new_[10136]_ );
  assign \new_[6202]_  = ~\new_[6804]_  | ~\wb_addr_i[22] ;
  assign \new_[6203]_  = ~\new_[6806]_  | ~\wb_addr_i[23] ;
  assign \new_[6204]_  = ~\new_[11716]_  | ~\wb_addr_i[24] ;
  assign \new_[6205]_  = ~\new_[7238]_  | ~\new_[10097]_ ;
  assign \new_[6206]_  = ~\new_[6809]_  | ~\new_[10039]_ ;
  assign \new_[6207]_  = ~\new_[12749]_  | ~\new_[10054]_ ;
  assign \new_[6208]_  = ~\new_[6663]_  & ~\new_[7069]_ ;
  assign \new_[6209]_  = ~\new_[12747]_  | ~\new_[9912]_ ;
  assign \new_[6210]_  = ~\new_[12751]_  | ~\new_[10065]_ ;
  assign \new_[6211]_  = ~\new_[12751]_  | ~\new_[10053]_ ;
  assign \new_[6212]_  = ~\new_[6808]_  | ~\new_[10104]_ ;
  assign \new_[6213]_  = ~\new_[12747]_  | ~\new_[10046]_ ;
  assign \new_[6214]_  = ~\new_[12747]_  | ~\new_[10078]_ ;
  assign \new_[6215]_  = ~\new_[10177]_  | ~\new_[7825]_  | ~\new_[7116]_ ;
  assign \new_[6216]_  = ~\new_[12750]_  | ~\new_[9849]_ ;
  assign \new_[6217]_  = ~\new_[12747]_  | ~\new_[10140]_ ;
  assign \new_[6218]_  = ~\new_[12751]_  | ~\new_[10081]_ ;
  assign \new_[6219]_  = ~\new_[12751]_  | ~\new_[10130]_ ;
  assign \new_[6220]_  = ~\new_[12751]_  | ~\new_[9985]_ ;
  assign \new_[6221]_  = ~\new_[12751]_  | ~\new_[10082]_ ;
  assign \new_[6222]_  = ~\new_[11320]_  | ~\new_[7776]_  | ~\new_[7116]_ ;
  assign \new_[6223]_  = ~\new_[11773]_  | ~\new_[9418]_ ;
  assign \new_[6224]_  = ~\new_[6809]_  | ~\new_[10126]_ ;
  assign \new_[6225]_  = ~\new_[12747]_  | ~\new_[9668]_ ;
  assign \new_[6226]_  = ~\new_[12751]_  | ~\new_[9807]_ ;
  assign \new_[6227]_  = ~\new_[12751]_  | ~\new_[9970]_ ;
  assign \new_[6228]_  = ~\new_[12749]_  | ~\new_[10071]_ ;
  assign \new_[6229]_  = ~\new_[12751]_  | ~\new_[9839]_ ;
  assign \new_[6230]_  = ~\new_[11313]_  | ~\new_[7776]_  | ~\new_[7116]_ ;
  assign \new_[6231]_  = ~\new_[12751]_  | ~\new_[9847]_ ;
  assign \new_[6232]_  = ~\new_[6809]_  | ~\new_[9987]_ ;
  assign \new_[6233]_  = ~\new_[12747]_  | ~\new_[9649]_ ;
  assign \new_[6234]_  = ~\new_[12747]_  | ~\new_[9965]_ ;
  assign \new_[6235]_  = ~\new_[12751]_  | ~\new_[9856]_ ;
  assign \new_[6236]_  = ~\new_[12093]_  | ~\new_[7776]_  | ~\new_[7116]_ ;
  assign \new_[6237]_  = ~\new_[6808]_  | ~\new_[10083]_ ;
  assign \new_[6238]_  = ~\new_[12747]_  | ~\new_[10049]_ ;
  assign \new_[6239]_  = ~\new_[12747]_  | ~\new_[10087]_ ;
  assign \new_[6240]_  = ~\new_[12747]_  | ~\new_[10127]_ ;
  assign \new_[6241]_  = ~\new_[12751]_  | ~\new_[9606]_ ;
  assign \new_[6242]_  = ~\new_[12751]_  | ~\new_[11452]_ ;
  assign \new_[6243]_  = ~\new_[11773]_  | ~\new_[9618]_ ;
  assign \new_[6244]_  = ~\new_[6808]_  | ~\new_[9657]_ ;
  assign \new_[6245]_  = ~\new_[11773]_  | ~\new_[9682]_ ;
  assign \new_[6246]_  = ~\new_[12751]_  | ~\new_[9846]_ ;
  assign \new_[6247]_  = ~\new_[11353]_  | ~\new_[7776]_  | ~\new_[7116]_ ;
  assign \new_[6248]_  = ~\new_[12751]_  | ~\new_[9967]_ ;
  assign \new_[6249]_  = ~\new_[12750]_  | ~\new_[9871]_ ;
  assign \new_[6250]_  = ~\new_[6807]_  | ~\new_[9675]_ ;
  assign \new_[6251]_  = ~\new_[7238]_  | ~\new_[9709]_ ;
  assign \new_[6252]_  = ~\new_[12751]_  | ~\new_[10044]_ ;
  assign \new_[6253]_  = ~\new_[11367]_  | ~\new_[7776]_  | ~\new_[7116]_ ;
  assign \new_[6254]_  = ~\new_[7238]_  | ~\new_[9619]_ ;
  assign \new_[6255]_  = ~\new_[12747]_  | ~\new_[10050]_ ;
  assign \new_[6256]_  = ~\new_[12769]_  & ~\new_[12385]_ ;
  assign \new_[6257]_  = ~\new_[6807]_  | ~\new_[9567]_ ;
  assign \new_[6258]_  = ~\new_[6807]_  | ~\new_[9707]_ ;
  assign \new_[6259]_  = ~\new_[12751]_  | ~\new_[10056]_ ;
  assign \new_[6260]_  = ~\new_[11361]_  | ~\new_[7776]_  | ~\new_[7116]_ ;
  assign \new_[6261]_  = ~\new_[12747]_  | ~\new_[10089]_ ;
  assign \new_[6262]_  = ~\new_[12751]_  | ~\new_[10107]_ ;
  assign \new_[6263]_  = ~\new_[12751]_  | ~\new_[10118]_ ;
  assign \new_[6264]_  = ~\new_[12751]_  | ~\new_[10063]_ ;
  assign \new_[6265]_  = ~\new_[12751]_  | ~\new_[9608]_ ;
  assign \new_[6266]_  = ~\new_[6808]_  | ~\new_[9990]_ ;
  assign \new_[6267]_  = ~\new_[6268]_ ;
  assign \new_[6268]_  = ~\new_[7180]_ ;
  assign \new_[6269]_  = ~\new_[12273]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6270]_  = ~\new_[11735]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6271]_  = ~\new_[11298]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6272]_  = ~\new_[12089]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6273]_  = ~\new_[10108]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6274]_  = ~n5021 | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6275]_  = ~\new_[10164]_  | ~\new_[12655]_  | ~\new_[8748]_ ;
  assign \new_[6276]_  = ~\new_[7059]_  | ~\new_[9967]_ ;
  assign \new_[6277]_  = ~\new_[12785]_  | ~\new_[7865]_  | ~\new_[12388]_ ;
  assign \new_[6278]_  = ~\new_[7059]_  | ~\new_[9871]_ ;
  assign \new_[6279]_  = ~\new_[7059]_  | ~\new_[10089]_ ;
  assign \new_[6280]_  = ~\new_[12044]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6281]_  = ~\new_[10509]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6282]_  = ~\new_[6639]_ ;
  assign \new_[6283]_  = ~\new_[7185]_ ;
  assign \new_[6284]_  = ~\new_[7185]_ ;
  assign \new_[6285]_  = ~\new_[6668]_  | ~\wb_addr_i[21] ;
  assign \new_[6286]_  = ~\new_[6668]_  | ~\wb_addr_i[22] ;
  assign \new_[6287]_  = ~\new_[6665]_  | ~\new_[9388]_ ;
  assign \new_[6288]_  = ~\new_[6665]_  | ~\new_[11772]_ ;
  assign \new_[6289]_  = ~\new_[7366]_  & ~\new_[6064]_ ;
  assign \new_[6290]_  = ~\new_[6669]_  & ~\new_[7714]_ ;
  assign \new_[6291]_  = ~\new_[6667]_  & ~\new_[11718]_ ;
  assign \new_[6292]_  = ~\new_[12783]_  | (~\new_[10148]_  & ~\new_[9648]_ );
  assign \new_[6293]_  = (~\new_[11264]_  | ~\wb_addr_i[7] ) & (~\new_[6836]_  | ~\wb_addr_i[6] );
  assign \new_[6294]_  = (~\new_[11264]_  | ~\wb_addr_i[5] ) & (~\new_[7373]_  | ~\wb_addr_i[4] );
  assign \new_[6295]_  = (~\new_[11264]_  | ~\wb_addr_i[12] ) & (~\new_[6836]_  | ~\wb_addr_i[11] );
  assign \new_[6296]_  = (~\new_[11264]_  | ~\wb_addr_i[18] ) & (~\new_[7373]_  | ~\wb_addr_i[17] );
  assign \new_[6297]_  = (~\new_[11264]_  | ~\wb_addr_i[21] ) & (~\new_[6836]_  | ~\wb_addr_i[20] );
  assign \new_[6298]_  = (~\new_[11264]_  | ~\wb_addr_i[13] ) & (~\new_[7373]_  | ~\wb_addr_i[12] );
  assign \new_[6299]_  = (~\new_[11264]_  | ~\wb_addr_i[14] ) & (~\new_[7373]_  | ~\wb_addr_i[13] );
  assign \new_[6300]_  = (~\new_[11264]_  | ~\wb_addr_i[16] ) & (~\new_[7373]_  | ~\wb_addr_i[15] );
  assign \new_[6301]_  = (~\new_[11264]_  | ~\wb_addr_i[17] ) & (~\new_[7373]_  | ~\wb_addr_i[16] );
  assign \new_[6302]_  = (~\new_[11264]_  | ~\wb_addr_i[19] ) & (~\new_[7373]_  | ~\wb_addr_i[18] );
  assign \new_[6303]_  = (~\new_[11264]_  | ~\wb_addr_i[20] ) & (~\new_[7373]_  | ~\wb_addr_i[19] );
  assign \new_[6304]_  = (~\new_[11264]_  | ~\wb_addr_i[22] ) & (~\new_[6836]_  | ~\wb_addr_i[21] );
  assign \new_[6305]_  = ~\new_[6661]_ ;
  assign \new_[6306]_  = (~\new_[11264]_  | ~\wb_addr_i[24] ) & (~\new_[6836]_  | ~\wb_addr_i[23] );
  assign \new_[6307]_  = (~\new_[11264]_  | ~\wb_addr_i[25] ) & (~\new_[6836]_  | ~\wb_addr_i[24] );
  assign \new_[6308]_  = (~\new_[11264]_  | ~\wb_addr_i[6] ) & (~\new_[6836]_  | ~\wb_addr_i[5] );
  assign \new_[6309]_  = (~\new_[11264]_  | ~\wb_addr_i[8] ) & (~\new_[6836]_  | ~\wb_addr_i[7] );
  assign \new_[6310]_  = (~\new_[11264]_  | ~\wb_addr_i[9] ) & (~\new_[6836]_  | ~\wb_addr_i[8] );
  assign \new_[6311]_  = (~\new_[11264]_  | ~\wb_addr_i[4] ) & (~\new_[7373]_  | ~\wb_addr_i[3] );
  assign \new_[6312]_  = (~\new_[11264]_  | ~\wb_addr_i[11] ) & (~\new_[7373]_  | ~\wb_addr_i[10] );
  assign \new_[6313]_  = (~\new_[11264]_  | ~\wb_addr_i[10] ) & (~\new_[7373]_  | ~\wb_addr_i[9] );
  assign \new_[6314]_  = (~\new_[11264]_  | ~\wb_addr_i[15] ) & (~\new_[7373]_  | ~\wb_addr_i[14] );
  assign \new_[6315]_  = ~\new_[6836]_  | ~\new_[10164]_ ;
  assign \new_[6316]_  = ~\new_[6663]_ ;
  assign \new_[6317]_  = ~\new_[12238]_ ;
  assign \new_[6318]_  = \\u2_u0_b0_last_row_reg[6] ;
  assign \new_[6319]_  = ~\new_[6836]_  | ~\wb_addr_i[2] ;
  assign \new_[6320]_  = ~\new_[6664]_ ;
  assign \new_[6321]_  = ~\new_[6720]_ ;
  assign \new_[6322]_  = ~\new_[6666]_ ;
  assign \new_[6323]_  = \\u2_u0_b3_last_row_reg[8] ;
  assign \new_[6324]_  = \\u2_u1_b2_last_row_reg[0] ;
  assign \new_[6325]_  = ~\new_[12534]_  | ~\new_[9839]_ ;
  assign \new_[6326]_  = \\u2_u1_b2_last_row_reg[8] ;
  assign \new_[6327]_  = \new_[10068]_  & \new_[12566]_ ;
  assign \new_[6328]_  = ~\new_[12564]_  | ~\new_[12566]_  | ~\new_[10839]_ ;
  assign \new_[6329]_  = \\u2_u1_b3_last_row_reg[10] ;
  assign \new_[6330]_  = \\u2_u1_b3_last_row_reg[1] ;
  assign \new_[6331]_  = \\u2_u0_b0_last_row_reg[4] ;
  assign \new_[6332]_  = ~\\u2_u0_b0_last_row_reg[12] ;
  assign \new_[6333]_  = \\u2_u1_b3_last_row_reg[0] ;
  assign \new_[6334]_  = \\u2_u1_b2_last_row_reg[7] ;
  assign \new_[6335]_  = \\u2_u1_b2_last_row_reg[9] ;
  assign \new_[6336]_  = ~\new_[6838]_  | ~\new_[7125]_ ;
  assign \new_[6337]_  = ~\new_[6839]_  | ~\new_[7126]_ ;
  assign \new_[6338]_  = ~\new_[11160]_  | ~\new_[12622]_ ;
  assign \new_[6339]_  = ~\new_[11143]_  | ~\new_[12622]_ ;
  assign \new_[6340]_  = ~\new_[11261]_  | ~\new_[12622]_ ;
  assign \new_[6341]_  = \\u2_u1_b2_last_row_reg[3] ;
  assign \new_[6342]_  = (~\new_[7157]_  | ~\new_[10127]_ ) & (~\new_[7571]_  | ~\new_[9109]_ );
  assign \new_[6343]_  = ~\new_[12593]_ ;
  assign \new_[6344]_  = ~\new_[12593]_ ;
  assign \new_[6345]_  = ~\new_[12593]_ ;
  assign \new_[6346]_  = \new_[12593]_ ;
  assign \new_[6347]_  = \new_[7351]_  & \new_[11453]_ ;
  assign \new_[6348]_  = ~\new_[7352]_  | ~\new_[11453]_ ;
  assign \new_[6349]_  = ~\new_[7308]_  | ~\new_[7830]_  | ~\new_[8050]_  | ~\new_[7711]_ ;
  assign \new_[6350]_  = ~\new_[6948]_  | ~\new_[10463]_ ;
  assign \new_[6351]_  = ~\new_[6948]_  | ~\new_[10508]_ ;
  assign \new_[6352]_  = ~\new_[6948]_  | ~\new_[10502]_ ;
  assign \new_[6353]_  = ~\new_[10463]_  | ~\new_[6949]_ ;
  assign \new_[6354]_  = ~\new_[10508]_  | ~\new_[6949]_ ;
  assign \new_[6355]_  = ~\new_[10502]_  | ~\new_[6949]_ ;
  assign \new_[6356]_  = ~\new_[7357]_  | ~\new_[11453]_ ;
  assign \new_[6357]_  = ~\new_[7358]_  | ~\new_[11453]_ ;
  assign \new_[6358]_  = ~\new_[7359]_  | ~\new_[11453]_ ;
  assign \new_[6359]_  = ~\new_[3176]_  | ~\new_[10941]_  | ~\new_[7163]_ ;
  assign \new_[6360]_  = ~\new_[7101]_  | ~\new_[11453]_ ;
  assign \new_[6361]_  = ~\new_[7356]_  | ~\new_[11453]_ ;
  assign \new_[6362]_  = \\u2_u1_b2_last_row_reg[1] ;
  assign \new_[6363]_  = \new_[6997]_  | \new_[12075]_ ;
  assign \new_[6364]_  = ~\new_[6676]_ ;
  assign \new_[6365]_  = ~\new_[11774]_  & ~\new_[11505]_ ;
  assign \new_[6366]_  = ~\\u2_u1_b2_last_row_reg[12] ;
  assign \new_[6367]_  = ~\new_[6972]_  & ~\new_[7172]_ ;
  assign \new_[6368]_  = \\u2_u1_b2_last_row_reg[11] ;
  assign \new_[6369]_  = ~\new_[6814]_  | ~\new_[11453]_ ;
  assign \new_[6370]_  = \\u2_u1_b1_last_row_reg[8] ;
  assign \new_[6371]_  = ~\new_[7107]_  | ~\new_[11453]_ ;
  assign \new_[6372]_  = ~\new_[6815]_  | ~\new_[11453]_ ;
  assign \new_[6373]_  = ~\new_[7261]_  | ~\new_[11453]_ ;
  assign \new_[6374]_  = (~\new_[11248]_  | ~\new_[12618]_ ) & (~\new_[10994]_  | ~\new_[12622]_ );
  assign \new_[6375]_  = ~\new_[7262]_  | ~\new_[11453]_ ;
  assign \new_[6376]_  = ~\new_[6677]_ ;
  assign \new_[6377]_  = ~\new_[11573]_  | ~\new_[11881]_  | ~\new_[6998]_  | ~\new_[11572]_ ;
  assign \new_[6378]_  = ~\\u2_u1_b1_last_row_reg[12] ;
  assign \new_[6379]_  = ~\new_[10126]_  & (~\new_[7164]_  | ~\new_[10367]_ );
  assign \new_[6380]_  = ~\new_[9987]_  & (~\new_[7166]_  | ~\new_[10367]_ );
  assign \new_[6381]_  = ~\new_[7438]_  & (~\new_[7171]_  | ~\new_[7317]_ );
  assign \new_[6382]_  = \\u2_u0_b3_last_row_reg[9] ;
  assign \new_[6383]_  = ~\new_[7432]_  & (~\new_[7171]_  | ~\new_[7660]_ );
  assign \new_[6384]_  = ~\new_[7176]_  | ~\new_[7183]_ ;
  assign \new_[6385]_  = \\u2_u1_b1_last_row_reg[4] ;
  assign \new_[6386]_  = \\u2_u1_b1_last_row_reg[7] ;
  assign \new_[6387]_  = \\u2_u1_b1_last_row_reg[6] ;
  assign \new_[6388]_  = \\u2_u1_b1_last_row_reg[5] ;
  assign \new_[6389]_  = \\u2_u1_b1_last_row_reg[2] ;
  assign \new_[6390]_  = \\u2_u1_b0_last_row_reg[0] ;
  assign \new_[6391]_  = ~\new_[12070]_  & ~\new_[1433]_ ;
  assign \new_[6392]_  = \\u2_u1_b1_last_row_reg[10] ;
  assign \new_[6393]_  = ~\new_[6681]_ ;
  assign \new_[6394]_  = ~\new_[7021]_  & ~\new_[7065]_ ;
  assign \new_[6395]_  = ~\new_[10838]_  | ~\new_[10367]_  | ~\new_[7523]_ ;
  assign \new_[6396]_  = ~\new_[8740]_  & ~\new_[7292]_ ;
  assign \new_[6397]_  = \new_[7021]_  | \new_[7577]_ ;
  assign \new_[6398]_  = ~\new_[7163]_  | ~\new_[10961]_  | ~\new_[10931]_ ;
  assign \new_[6399]_  = ~\new_[10818]_  | ~\new_[11776]_  | ~\new_[7523]_ ;
  assign \new_[6400]_  = ~\new_[10938]_  | ~\new_[11776]_  | ~\new_[7191]_ ;
  assign \new_[6401]_  = \\u2_u1_b0_last_row_reg[7] ;
  assign \new_[6402]_  = ~\new_[9785]_  | ~\new_[11776]_  | ~\new_[7523]_ ;
  assign \new_[6403]_  = \\u2_u1_b0_last_row_reg[9] ;
  assign \new_[6404]_  = \\u2_u1_b0_last_row_reg[5] ;
  assign \new_[6405]_  = \\u2_u1_b0_last_row_reg[2] ;
  assign \new_[6406]_  = ~\new_[10933]_  | ~\new_[10367]_  | ~\new_[7191]_ ;
  assign \new_[6407]_  = \\u2_u0_b0_last_row_reg[0] ;
  assign \new_[6408]_  = \\u2_u0_b0_last_row_reg[10] ;
  assign \new_[6409]_  = \\u2_u0_b0_last_row_reg[11] ;
  assign \new_[6410]_  = \\u2_u0_b0_last_row_reg[1] ;
  assign \new_[6411]_  = \\u2_u0_b0_last_row_reg[2] ;
  assign \new_[6412]_  = \\u2_u0_b0_last_row_reg[3] ;
  assign \new_[6413]_  = \\u2_u0_b0_last_row_reg[5] ;
  assign \new_[6414]_  = \\u2_u0_b0_last_row_reg[9] ;
  assign \new_[6415]_  = \\u2_u0_b1_last_row_reg[10] ;
  assign \new_[6416]_  = ~\\u2_u0_b1_last_row_reg[12] ;
  assign \new_[6417]_  = \\u2_u0_b1_last_row_reg[4] ;
  assign \new_[6418]_  = \\u2_u0_b1_last_row_reg[6] ;
  assign \new_[6419]_  = \\u2_u0_b1_last_row_reg[9] ;
  assign \new_[6420]_  = \\u2_u0_b2_last_row_reg[10] ;
  assign \new_[6421]_  = ~\\u2_u0_b2_last_row_reg[12] ;
  assign \new_[6422]_  = \\u2_u0_b2_last_row_reg[2] ;
  assign \new_[6423]_  = \\u2_u0_b2_last_row_reg[4] ;
  assign \new_[6424]_  = \\u2_u0_b2_last_row_reg[5] ;
  assign \new_[6425]_  = \\u2_u0_b2_last_row_reg[8] ;
  assign \new_[6426]_  = \\u2_u0_b2_last_row_reg[9] ;
  assign \new_[6427]_  = \\u2_u0_b2_last_row_reg[3] ;
  assign \new_[6428]_  = \\u2_u0_b3_last_row_reg[11] ;
  assign \new_[6429]_  = \\u2_u0_b3_last_row_reg[5] ;
  assign \new_[6430]_  = \\u2_u1_b0_last_row_reg[11] ;
  assign \new_[6431]_  = ~\\u2_u1_b0_last_row_reg[12] ;
  assign \new_[6432]_  = ~\new_[11313]_  | ~\new_[10367]_  | ~\new_[7191]_ ;
  assign \new_[6433]_  = \\u2_u1_b0_last_row_reg[3] ;
  assign \new_[6434]_  = \\u2_u1_b0_last_row_reg[4] ;
  assign \new_[6435]_  = \\u2_u1_b0_last_row_reg[6] ;
  assign \new_[6436]_  = \\u2_u1_b0_last_row_reg[8] ;
  assign \new_[6437]_  = \\u2_u1_b1_last_row_reg[0] ;
  assign \new_[6438]_  = \\u2_u1_b1_last_row_reg[11] ;
  assign \new_[6439]_  = \\u2_u1_b1_last_row_reg[1] ;
  assign \new_[6440]_  = \\u2_u1_b1_last_row_reg[3] ;
  assign \new_[6441]_  = \\u2_u1_b1_last_row_reg[9] ;
  assign \new_[6442]_  = \\u2_u1_b2_last_row_reg[10] ;
  assign \new_[6443]_  = \\u2_u1_b2_last_row_reg[2] ;
  assign \new_[6444]_  = \\u2_u1_b2_last_row_reg[4] ;
  assign \new_[6445]_  = \\u2_u1_b2_last_row_reg[5] ;
  assign \new_[6446]_  = \\u2_u1_b2_last_row_reg[6] ;
  assign \new_[6447]_  = \\u2_u1_b3_last_row_reg[11] ;
  assign \new_[6448]_  = ~\\u2_u1_b3_last_row_reg[12] ;
  assign \new_[6449]_  = ~\new_[9903]_  | ~\new_[10367]_  | ~\new_[7191]_ ;
  assign \new_[6450]_  = \\u2_u1_b3_last_row_reg[3] ;
  assign \new_[6451]_  = \\u2_u1_b3_last_row_reg[5] ;
  assign \new_[6452]_  = \\u2_u1_b3_last_row_reg[7] ;
  assign \new_[6453]_  = \\u2_u1_b3_last_row_reg[6] ;
  assign \new_[6454]_  = \\u2_u1_b3_last_row_reg[8] ;
  assign \new_[6455]_  = \\u2_u0_b3_last_row_reg[0] ;
  assign \new_[6456]_  = ~\new_[12054]_  | ~\new_[10367]_  | ~\new_[7191]_ ;
  assign \new_[6457]_  = ~\new_[7019]_  & ~\new_[11987]_ ;
  assign \new_[6458]_  = \\u2_u1_b0_last_row_reg[10] ;
  assign \new_[6459]_  = ~\new_[7363]_  | ~\new_[11846]_ ;
  assign \new_[6460]_  = ~\new_[6688]_ ;
  assign \new_[6461]_  = \new_[7014]_  | \new_[7573]_ ;
  assign \new_[6462]_  = ~\new_[12598]_  | ~\new_[10367]_  | ~\new_[7523]_ ;
  assign \new_[6463]_  = ~\new_[7298]_  | ~\new_[7911]_ ;
  assign \new_[6464]_  = ~\new_[7197]_  | ~\new_[7671]_  | ~\new_[7219]_ ;
  assign \new_[6465]_  = ~\new_[7016]_  & ~\new_[12794]_ ;
  assign \new_[6466]_  = ~\new_[7864]_  & ~\new_[7012]_ ;
  assign \new_[6467]_  = \\u2_u1_b0_last_row_reg[1] ;
  assign \new_[6468]_  = ~\new_[11310]_  | ~\new_[10367]_  | ~\new_[7191]_ ;
  assign \new_[6469]_  = ~\new_[10960]_  | ~\new_[10367]_  | ~\new_[7191]_ ;
  assign \new_[6470]_  = ~\new_[10634]_  | ~\new_[10367]_  | ~\new_[7523]_ ;
  assign \new_[6471]_  = \\u2_u0_b0_last_row_reg[7] ;
  assign \new_[6472]_  = \new_[7025]_  | \new_[7600]_ ;
  assign \new_[6473]_  = \new_[7033]_  | \new_[7600]_ ;
  assign \new_[6474]_  = \new_[7038]_  | \new_[7600]_ ;
  assign \new_[6475]_  = ~\new_[7042]_  & ~\new_[7600]_ ;
  assign \new_[6476]_  = ~\new_[7040]_  & ~\new_[7600]_ ;
  assign \new_[6477]_  = ~\new_[7027]_  & ~\new_[7600]_ ;
  assign \new_[6478]_  = ~\new_[7028]_  & ~\new_[7600]_ ;
  assign \new_[6479]_  = \new_[7044]_  | \new_[7600]_ ;
  assign \new_[6480]_  = ~\new_[7032]_  & ~\new_[7600]_ ;
  assign \new_[6481]_  = ~\new_[7029]_  & ~\new_[7600]_ ;
  assign \new_[6482]_  = ~\new_[7034]_  & ~\new_[7600]_ ;
  assign \new_[6483]_  = ~\new_[7030]_  & ~\new_[7600]_ ;
  assign \new_[6484]_  = \new_[7036]_  | \new_[7600]_ ;
  assign \new_[6485]_  = \new_[7026]_  | \new_[7600]_ ;
  assign \new_[6486]_  = \new_[7041]_  | \new_[7600]_ ;
  assign \new_[6487]_  = \new_[7035]_  | \new_[7600]_ ;
  assign \new_[6488]_  = \new_[7031]_  | \new_[7600]_ ;
  assign \new_[6489]_  = \new_[7043]_  | \new_[7600]_ ;
  assign \new_[6490]_  = \\u2_u0_b3_last_row_reg[3] ;
  assign \new_[6491]_  = \new_[7037]_  | \new_[7600]_ ;
  assign \new_[6492]_  = ~\new_[7024]_  & ~\new_[7600]_ ;
  assign \new_[6493]_  = \new_[7045]_  | \new_[7600]_ ;
  assign \new_[6494]_  = \new_[7039]_  | \new_[7600]_ ;
  assign \new_[6495]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7647]_ ;
  assign \new_[6496]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7648]_ ;
  assign \new_[6497]_  = ~n3951 | ~\new_[7054]_  | ~\new_[12672]_ ;
  assign \new_[6498]_  = ~\new_[11491]_  | ~\new_[7001]_  | ~\new_[7766]_ ;
  assign \new_[6499]_  = ~\new_[12398]_  | ~\new_[6823]_  | ~\new_[7482]_ ;
  assign \new_[6500]_  = ~\new_[11491]_  | ~\new_[7001]_  | ~\new_[7483]_ ;
  assign \new_[6501]_  = ~\new_[12398]_  | ~\new_[6823]_  | ~\new_[7484]_ ;
  assign \new_[6502]_  = ~\new_[12398]_  | ~\new_[6822]_  | ~\new_[7486]_ ;
  assign \new_[6503]_  = ~\new_[12398]_  | ~\new_[6824]_  | ~\new_[7312]_ ;
  assign \new_[6504]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7500]_ ;
  assign \new_[6505]_  = ~\new_[12398]_  | ~\new_[6822]_  | ~\new_[7313]_ ;
  assign \new_[6506]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7504]_ ;
  assign \new_[6507]_  = ~\new_[12398]_  | ~\new_[6822]_  | ~\new_[7314]_ ;
  assign \new_[6508]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7767]_ ;
  assign \new_[6509]_  = ~\new_[12398]_  | ~\new_[6822]_  | ~\new_[7489]_ ;
  assign \new_[6510]_  = ~\new_[11491]_  | ~\new_[7001]_  | ~\new_[7491]_ ;
  assign \new_[6511]_  = ~\new_[12398]_  | ~\new_[6824]_  | ~\new_[7492]_ ;
  assign \new_[6512]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7493]_ ;
  assign \new_[6513]_  = \\u2_u0_b1_last_row_reg[5] ;
  assign \new_[6514]_  = ~\new_[12398]_  | ~\new_[6823]_  | ~\new_[7495]_ ;
  assign \new_[6515]_  = ~\new_[11491]_  | ~\new_[7001]_  | ~\new_[7497]_ ;
  assign \new_[6516]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7653]_ ;
  assign \new_[6517]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7488]_ ;
  assign \new_[6518]_  = \\u2_u0_b3_last_row_reg[7] ;
  assign \new_[6519]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7509]_ ;
  assign \new_[6520]_  = ~\new_[11491]_  | ~\new_[6824]_  | ~\new_[7517]_ ;
  assign \new_[6521]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7511]_ ;
  assign \new_[6522]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7499]_ ;
  assign \new_[6523]_  = \\u2_u1_b3_last_row_reg[4] ;
  assign \new_[6524]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7652]_ ;
  assign \new_[6525]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7315]_ ;
  assign \new_[6526]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7519]_ ;
  assign \new_[6527]_  = \new_[3176]_  ^ \new_[7163]_ ;
  assign \new_[6528]_  = ~\new_[12398]_  | ~\new_[6823]_  | ~\new_[7318]_ ;
  assign \new_[6529]_  = \\u2_u0_b3_last_row_reg[4] ;
  assign \new_[6530]_  = ~\new_[11491]_  | ~\new_[6825]_  | ~\new_[7320]_ ;
  assign \new_[6531]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7516]_ ;
  assign \new_[6532]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7660]_ ;
  assign \new_[6533]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7505]_ ;
  assign \new_[6534]_  = ~\new_[12398]_  | ~\new_[6824]_  | ~\new_[7321]_ ;
  assign \new_[6535]_  = ~\new_[11307]_  & (~\new_[1643]_  | ~\new_[7593]_ );
  assign \new_[6536]_  = ~\new_[11491]_  | ~\new_[6821]_  | ~\new_[7322]_ ;
  assign \new_[6537]_  = \\u2_u0_b3_last_row_reg[6] ;
  assign \new_[6538]_  = ~\new_[7673]_  | (~\new_[7182]_  & ~\new_[10101]_ );
  assign \new_[6539]_  = ~\new_[7670]_  | (~\new_[7182]_  & ~\new_[9927]_ );
  assign \new_[6540]_  = ~\new_[7004]_  & (~\new_[12665]_  | ~\new_[12002]_ );
  assign \new_[6541]_  = ~\new_[10057]_  & (~\new_[7112]_  | ~\new_[7136]_ );
  assign \new_[6542]_  = \\u2_u0_b3_last_row_reg[1] ;
  assign \new_[6543]_  = ~u0_wp_err_reg;
  assign \new_[6544]_  = \\u2_u0_b3_last_row_reg[2] ;
  assign \new_[6545]_  = (~\new_[10223]_  | ~\new_[12664]_ ) & (~\new_[7682]_  | ~\new_[9584]_ );
  assign \new_[6546]_  = (~\new_[10512]_  | ~\new_[12664]_ ) & (~\new_[7682]_  | ~\new_[9588]_ );
  assign \new_[6547]_  = (~\new_[9620]_  | ~\new_[7537]_ ) & (~\new_[7239]_  | ~\new_[9388]_ );
  assign \new_[6548]_  = ~\\u2_u0_b3_last_row_reg[12] ;
  assign \new_[6549]_  = (~\new_[7588]_  | ~\new_[10265]_ ) & (~\new_[7239]_  | ~\new_[10039]_ );
  assign \new_[6550]_  = \\u2_u0_b3_last_row_reg[10] ;
  assign \new_[6551]_  = (~\new_[11997]_  | ~\new_[9615]_ ) & (~\new_[6828]_  | ~\new_[10126]_ );
  assign \new_[6552]_  = \\u2_u0_b2_last_row_reg[7] ;
  assign \new_[6553]_  = (~\new_[11997]_  | ~\new_[9855]_ ) & (~\new_[7287]_  | ~\new_[9958]_ );
  assign \new_[6554]_  = (~\new_[11997]_  | ~\new_[9598]_ ) & (~\new_[7113]_  | ~\new_[9326]_ );
  assign \new_[6555]_  = (~\new_[11997]_  | ~\new_[10210]_ ) & (~\new_[7113]_  | ~\new_[9611]_ );
  assign \new_[6556]_  = (~\new_[11997]_  | ~\new_[9865]_ ) & (~\new_[7113]_  | ~\new_[9853]_ );
  assign \new_[6557]_  = (~\new_[11997]_  | ~\new_[9969]_ ) & (~\new_[7287]_  | ~\new_[9644]_ );
  assign \new_[6558]_  = (~\new_[11997]_  | ~\new_[9906]_ ) & (~\new_[7287]_  | ~\new_[9582]_ );
  assign \new_[6559]_  = (~\new_[11997]_  | ~\new_[9837]_ ) & (~\new_[7287]_  | ~\new_[9104]_ );
  assign \new_[6560]_  = (~\new_[11997]_  | ~\new_[9857]_ ) & (~\new_[7113]_  | ~\new_[9682]_ );
  assign \new_[6561]_  = (~\new_[11997]_  | ~\new_[9663]_ ) & (~\new_[7113]_  | ~\new_[9374]_ );
  assign \new_[6562]_  = \\u2_u0_b2_last_row_reg[1] ;
  assign \new_[6563]_  = (~\new_[11997]_  | ~\new_[9581]_ ) & (~\new_[7287]_  | ~\new_[10097]_ );
  assign \new_[6564]_  = (~\new_[11997]_  | ~\new_[9862]_ ) & (~\new_[7287]_  | ~\new_[9675]_ );
  assign \new_[6565]_  = (~\new_[11997]_  | ~\new_[9840]_ ) & (~\new_[7113]_  | ~\new_[9709]_ );
  assign \new_[6566]_  = (~\new_[11997]_  | ~\new_[11973]_ ) & (~\new_[7113]_  | ~\new_[10115]_ );
  assign \new_[6567]_  = (~\new_[11997]_  | ~\new_[9818]_ ) & (~\new_[7287]_  | ~\new_[9567]_ );
  assign \new_[6568]_  = (~\new_[11997]_  | ~\new_[9659]_ ) & (~\new_[7113]_  | ~\new_[9707]_ );
  assign \new_[6569]_  = (~\new_[11997]_  | ~\new_[9746]_ ) & (~\new_[7287]_  | ~\new_[9389]_ );
  assign \new_[6570]_  = \\u2_u0_b2_last_row_reg[0] ;
  assign \new_[6571]_  = ~\new_[7061]_  | ~\new_[10039]_ ;
  assign \new_[6572]_  = ~\new_[12273]_  | ~\new_[7777]_  | ~\new_[7117]_ ;
  assign \new_[6573]_  = ~\new_[7022]_  | ~\new_[9401]_ ;
  assign \new_[6574]_  = ~\new_[7076]_  | ~\new_[9479]_ ;
  assign \new_[6575]_  = \\u2_u0_b1_last_row_reg[7] ;
  assign \new_[6576]_  = ~\new_[7060]_  | (~\new_[11776]_  & ~\new_[10922]_ );
  assign \new_[6577]_  = ~\new_[10743]_  | ~\new_[7825]_  | ~\new_[7267]_ ;
  assign \new_[6578]_  = \new_[7069]_  | \new_[8840]_ ;
  assign \new_[6579]_  = ~\new_[7022]_  | ~\new_[10099]_ ;
  assign \new_[6580]_  = ~\new_[7022]_  | ~\new_[9661]_ ;
  assign \new_[6581]_  = ~\new_[7022]_  | ~\new_[9963]_ ;
  assign \new_[6582]_  = \\u2_u0_b2_last_row_reg[11] ;
  assign \new_[6583]_  = ~\new_[7067]_  | ~\new_[10097]_ ;
  assign \new_[6584]_  = ~\new_[7022]_  | ~\new_[9680]_ ;
  assign \new_[6585]_  = ~\new_[7022]_  | ~\new_[9995]_ ;
  assign \new_[6586]_  = ~\new_[7022]_  | ~\new_[9845]_ ;
  assign \new_[6587]_  = ~\new_[7022]_  | ~\new_[10237]_ ;
  assign \new_[6588]_  = \\u2_u0_b2_last_row_reg[6] ;
  assign \new_[6589]_  = ~\new_[10243]_  | ~\new_[7825]_  | ~\new_[7286]_ ;
  assign \new_[6590]_  = ~\new_[7022]_  | ~\new_[9660]_ ;
  assign \new_[6591]_  = ~\new_[7061]_  | ~\new_[10126]_ ;
  assign \new_[6592]_  = ~\new_[7022]_  | ~\new_[9641]_ ;
  assign \new_[6593]_  = ~\new_[7076]_  | ~\new_[10137]_ ;
  assign \new_[6594]_  = ~\new_[11298]_  | ~\new_[7823]_  | ~\new_[7117]_ ;
  assign \new_[6595]_  = ~\new_[7022]_  | ~\new_[10287]_ ;
  assign \new_[6596]_  = ~\new_[11316]_  | ~\new_[7825]_  | ~\new_[7286]_ ;
  assign \new_[6597]_  = ~\new_[12089]_  | ~\new_[7823]_  | ~\new_[7117]_ ;
  assign \new_[6598]_  = ~\new_[7067]_  | ~\new_[9936]_ ;
  assign \new_[6599]_  = ~\new_[7061]_  | ~\new_[9987]_ ;
  assign \new_[6600]_  = ~\new_[7076]_  | ~\new_[9958]_ ;
  assign \new_[6601]_  = ~\new_[7067]_  | ~\new_[9958]_ ;
  assign \new_[6602]_  = ~\new_[7076]_  | ~\new_[9389]_ ;
  assign \new_[6603]_  = ~\new_[7067]_  | ~\new_[9665]_ ;
  assign \new_[6604]_  = ~\new_[10802]_  | ~\new_[7825]_  | ~\new_[7267]_ ;
  assign \new_[6605]_  = ~\new_[7076]_  | ~\new_[9326]_ ;
  assign \new_[6606]_  = \\u2_u1_b3_last_row_reg[9] ;
  assign \new_[6607]_  = ~\new_[7067]_  | ~\new_[9326]_ ;
  assign \new_[6608]_  = ~\new_[7076]_  | ~\new_[9611]_ ;
  assign \new_[6609]_  = ~\new_[7067]_  | ~\new_[9611]_ ;
  assign \new_[6610]_  = ~\new_[7076]_  | ~\new_[9644]_ ;
  assign \new_[6611]_  = ~\new_[7067]_  | ~\new_[9644]_ ;
  assign \new_[6612]_  = ~\new_[10164]_  | ~\new_[7825]_  | ~\new_[7267]_ ;
  assign \new_[6613]_  = ~\new_[7067]_  | ~\new_[9104]_ ;
  assign \new_[6614]_  = \\u2_u0_b1_last_row_reg[8] ;
  assign \new_[6615]_  = ~\new_[12748]_  | ~\new_[10153]_ ;
  assign \new_[6616]_  = ~\new_[7022]_  | ~\new_[10019]_ ;
  assign \new_[6617]_  = ~\new_[7079]_  | ~\new_[8002]_ ;
  assign \new_[6618]_  = ~\new_[12044]_  | ~\new_[7823]_  | ~\new_[7117]_ ;
  assign \new_[6619]_  = ~\new_[7022]_  | ~\new_[9407]_ ;
  assign \new_[6620]_  = ~\new_[7263]_  | ~\new_[7523]_ ;
  assign \new_[6621]_  = ~\new_[11864]_  | ~\new_[11776]_ ;
  assign \new_[6622]_  = ~\new_[7067]_  | ~\new_[9675]_ ;
  assign \new_[6623]_  = ~\new_[7067]_  | ~\new_[9709]_ ;
  assign \new_[6624]_  = ~\new_[7008]_  | ~\new_[9870]_ ;
  assign \new_[6625]_  = ~\new_[7067]_  | ~\new_[9619]_ ;
  assign \new_[6626]_  = ~\new_[7022]_  | ~\new_[9599]_ ;
  assign \new_[6627]_  = ~\new_[7067]_  | ~\new_[9567]_ ;
  assign \new_[6628]_  = ~\new_[7022]_  | ~\new_[9604]_ ;
  assign \new_[6629]_  = ~\new_[7067]_  | ~\new_[9389]_ ;
  assign \new_[6630]_  = ~\new_[7067]_  | ~\new_[10137]_ ;
  assign \new_[6631]_  = ~\new_[7022]_  | ~\new_[10037]_ ;
  assign \new_[6632]_  = ~\new_[12171]_  | ~\new_[12235]_  | ~\new_[12234]_ ;
  assign \new_[6633]_  = \\u2_u0_b0_last_row_reg[8] ;
  assign \new_[6634]_  = ~\new_[7008]_  | (~\new_[10511]_  & ~\new_[11355]_ );
  assign \new_[6635]_  = \new_[9064]_  | \new_[7264]_ ;
  assign \new_[6636]_  = \new_[6840]_  | \new_[10772]_ ;
  assign \new_[6637]_  = ~\new_[9785]_  | ~\new_[7109]_  | ~\new_[10572]_ ;
  assign \new_[6638]_  = ~\new_[7059]_  | (~\new_[10511]_  & ~\new_[12044]_ );
  assign \new_[6639]_  = ~\new_[6736]_ ;
  assign \new_[6640]_  = ~\new_[7185]_ ;
  assign \new_[6641]_  = ~\new_[7185]_ ;
  assign \new_[6642]_  = ~\new_[6738]_ ;
  assign \new_[6643]_  = \\u2_u1_b3_last_row_reg[2] ;
  assign \new_[6644]_  = \\u2_u0_b1_last_row_reg[11] ;
  assign \new_[6645]_  = \\u2_u0_b1_last_row_reg[3] ;
  assign n2931 = u5_wb_wait_r2_reg;
  assign \new_[6647]_  = \\u2_u0_b1_last_row_reg[2] ;
  assign \new_[6648]_  = \new_[3178]_  | \new_[7266]_ ;
  assign \new_[6649]_  = \new_[11050]_  | \new_[7266]_ ;
  assign \new_[6650]_  = \new_[3113]_  | \new_[6999]_ ;
  assign \new_[6651]_  = \\u2_u0_b1_last_row_reg[1] ;
  assign \new_[6652]_  = \new_[11864]_ ;
  assign \new_[6653]_  = \\u2_u0_b1_last_row_reg[0] ;
  assign \new_[6654]_  = ~\new_[11719]_ ;
  assign \new_[6655]_  = ~\new_[9855]_  & (~\new_[7288]_  | ~\new_[10148]_ );
  assign \new_[6656]_  = ~\new_[6729]_ ;
  assign \new_[6657]_  = ~\new_[6729]_ ;
  assign \new_[6658]_  = ~\new_[6729]_ ;
  assign \new_[6659]_  = ~\new_[6729]_ ;
  assign \new_[6660]_  = ~\new_[6729]_ ;
  assign \new_[6661]_  = (~\new_[11264]_  | ~\wb_addr_i[23] ) & (~\new_[6836]_  | ~\wb_addr_i[22] );
  assign \new_[6662]_  = ~\new_[7288]_  & ~\new_[12577]_ ;
  assign \new_[6663]_  = ~\new_[6317]_ ;
  assign \new_[6664]_  = \new_[11553]_ ;
  assign \new_[6665]_  = ~\new_[6827]_ ;
  assign \new_[6666]_  = \new_[11726]_  & \new_[7288]_ ;
  assign \new_[6667]_  = ~\new_[7827]_  | ~\new_[7288]_ ;
  assign \new_[6668]_  = ~\new_[6834]_ ;
  assign \new_[6669]_  = ~\new_[7717]_  | ~\new_[7288]_ ;
  assign \new_[6670]_  = ~\new_[6835]_ ;
  assign \new_[6671]_  = ~\new_[7131]_  & ~\new_[10036]_ ;
  assign \new_[6672]_  = ~\new_[7372]_ ;
  assign \new_[6673]_  = ~\new_[11038]_  | ~\new_[12621]_ ;
  assign \new_[6674]_  = \new_[12779]_  | \new_[7420]_ ;
  assign \new_[6675]_  = ~\new_[7155]_  | (~\new_[10190]_  & ~\new_[10743]_ );
  assign \new_[6676]_  = \new_[7537]_  | \new_[7141]_ ;
  assign \new_[6677]_  = ~\new_[11510]_  | ~\new_[7135]_ ;
  assign \new_[6678]_  = ~\new_[7154]_  & ~\new_[7573]_ ;
  assign \new_[6679]_  = \new_[11864]_ ;
  assign \new_[6680]_  = (~\new_[11500]_  | ~\new_[10043]_ ) & (~\new_[7682]_  | ~\new_[9850]_ );
  assign \new_[6681]_  = ~\new_[11453]_ ;
  assign \new_[6682]_  = \new_[11453]_ ;
  assign \new_[6683]_  = \new_[11453]_ ;
  assign \new_[6684]_  = \new_[11453]_ ;
  assign \new_[6685]_  = \new_[7186]_  | \new_[12384]_ ;
  assign \new_[6686]_  = ~\new_[6972]_ ;
  assign \new_[6687]_  = ~\new_[11505]_ ;
  assign \new_[6688]_  = ~\new_[12071]_  | ~\new_[7183]_ ;
  assign \new_[6689]_  = ~\new_[7370]_  | ~\new_[7176]_ ;
  assign \new_[6690]_  = \new_[7634]_  & \new_[7183]_ ;
  assign \new_[6691]_  = ~\new_[7184]_  & ~\new_[7190]_ ;
  assign \new_[6692]_  = \new_[9631]_  | \new_[7183]_ ;
  assign \new_[6693]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7481]_ ;
  assign \new_[6694]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7650]_ ;
  assign \new_[6695]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7510]_ ;
  assign \new_[6696]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7311]_ ;
  assign \new_[6697]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7487]_ ;
  assign \new_[6698]_  = ~\new_[11491]_  | ~\new_[7110]_  | ~\new_[7769]_ ;
  assign \new_[6699]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7490]_ ;
  assign \new_[6700]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7494]_ ;
  assign \new_[6701]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7502]_ ;
  assign \new_[6702]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7659]_ ;
  assign \new_[6703]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7310]_ ;
  assign \new_[6704]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7503]_ ;
  assign \new_[6705]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7514]_ ;
  assign \new_[6706]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7506]_ ;
  assign \new_[6707]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7507]_ ;
  assign \new_[6708]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7485]_ ;
  assign \new_[6709]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7508]_ ;
  assign \new_[6710]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7656]_ ;
  assign \new_[6711]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7658]_ ;
  assign \new_[6712]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7498]_ ;
  assign \new_[6713]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7515]_ ;
  assign \new_[6714]_  = ~\new_[7111]_  & (~\new_[7316]_  | ~\new_[11491]_ );
  assign \new_[6715]_  = ~\new_[11491]_  | ~\new_[7110]_  | ~\new_[7518]_ ;
  assign \new_[6716]_  = ~\new_[11491]_  | ~\new_[7110]_  | ~\new_[7768]_ ;
  assign \new_[6717]_  = ~\new_[12398]_  | ~\new_[7110]_  | ~\new_[7512]_ ;
  assign \new_[6718]_  = \new_[10961]_  & \new_[7163]_ ;
  assign \new_[6719]_  = ~\new_[12234]_  | ~\new_[11419]_  | ~\new_[8001]_  | ~\new_[12235]_ ;
  assign \new_[6720]_  = ~\new_[11553]_ ;
  assign \new_[6721]_  = ~\new_[12664]_  | ~\new_[3438]_ ;
  assign \new_[6722]_  = ~\new_[12665]_  | ~\new_[7197]_ ;
  assign \new_[6723]_  = ~\new_[7564]_  | ~\new_[7219]_ ;
  assign \new_[6724]_  = ~\new_[11773]_  | ~\new_[9930]_ ;
  assign \new_[6725]_  = ~\new_[7216]_  | ~\new_[10111]_ ;
  assign \new_[6726]_  = ~\new_[7216]_  | ~\new_[11860]_ ;
  assign \new_[6727]_  = ~\new_[7329]_  | ~\new_[9853]_ ;
  assign \new_[6728]_  = ~\new_[7329]_  | ~\new_[9582]_ ;
  assign \new_[6729]_  = ~\new_[7008]_ ;
  assign \new_[6730]_  = ~\new_[7190]_  & (~\new_[8145]_  | ~\new_[7708]_ );
  assign \new_[6731]_  = ~\new_[7216]_  | ~\new_[12110]_ ;
  assign \new_[6732]_  = ~\new_[7216]_  | ~\new_[9990]_ ;
  assign \new_[6733]_  = ~\new_[7018]_ ;
  assign \new_[6734]_  = ~\new_[7019]_ ;
  assign \new_[6735]_  = ~\new_[7021]_ ;
  assign \new_[6736]_  = ~\new_[7187]_  & (~\new_[7370]_  | ~\new_[11993]_ );
  assign \new_[6737]_  = ~\new_[12602]_  & (~n3451 | ~\new_[10148]_ );
  assign \new_[6738]_  = ~\new_[7186]_ ;
  assign \new_[6739]_  = (~\new_[7369]_  | ~\new_[9342]_ ) & (~\new_[7597]_  | ~\wb_addr_i[15] );
  assign \new_[6740]_  = (~\new_[7369]_  | ~\new_[9351]_ ) & (~\new_[7597]_  | ~\wb_addr_i[16] );
  assign \new_[6741]_  = \new_[7116]_  & \new_[10291]_ ;
  assign \new_[6742]_  = \new_[7116]_  & \new_[10250]_ ;
  assign \new_[6743]_  = \new_[7116]_  & \new_[10827]_ ;
  assign \new_[6744]_  = \new_[7267]_  & \new_[10959]_ ;
  assign \new_[6745]_  = \new_[7267]_  & \new_[10955]_ ;
  assign \new_[6746]_  = \new_[7286]_  & \new_[11355]_ ;
  assign \new_[6747]_  = \new_[7116]_  & \new_[11348]_ ;
  assign \new_[6748]_  = \new_[7286]_  & \new_[10928]_ ;
  assign \new_[6749]_  = \new_[7117]_  & \new_[10963]_ ;
  assign \new_[6750]_  = \new_[7117]_  & \new_[11576]_ ;
  assign \new_[6751]_  = \new_[7286]_  & \new_[10962]_ ;
  assign \new_[6752]_  = \new_[7286]_  & \new_[11331]_ ;
  assign \new_[6753]_  = \new_[7117]_  & \new_[11343]_ ;
  assign \new_[6754]_  = \new_[7117]_  & \new_[10818]_ ;
  assign \new_[6755]_  = \new_[7116]_  & \new_[10922]_ ;
  assign \new_[6756]_  = \new_[7286]_  & \new_[11340]_ ;
  assign \new_[6757]_  = \new_[7116]_  & \new_[11492]_ ;
  assign \new_[6758]_  = \new_[7286]_  & \new_[10938]_ ;
  assign \new_[6759]_  = \new_[7286]_  & \new_[11735]_ ;
  assign \new_[6760]_  = \new_[7286]_  & \new_[10526]_ ;
  assign \new_[6761]_  = \new_[7117]_  & \new_[10919]_ ;
  assign \new_[6762]_  = \new_[7116]_  & \new_[10496]_ ;
  assign \new_[6763]_  = \new_[7286]_  & \new_[10217]_ ;
  assign \new_[6764]_  = \new_[7267]_  & n5021;
  assign \new_[6765]_  = \new_[7267]_  & \new_[12567]_ ;
  assign \new_[6766]_  = \new_[7267]_  & \new_[11363]_ ;
  assign \new_[6767]_  = \new_[7116]_  & \new_[12453]_ ;
  assign \new_[6768]_  = \new_[7267]_  & \new_[9903]_ ;
  assign \new_[6769]_  = \new_[7117]_  & \new_[11356]_ ;
  assign \new_[6770]_  = \new_[7116]_  & \new_[9968]_ ;
  assign \new_[6771]_  = \new_[7116]_  & \new_[12755]_ ;
  assign \new_[6772]_  = \new_[7286]_  & \new_[12610]_ ;
  assign \new_[6773]_  = \new_[7286]_  & \new_[10419]_ ;
  assign \new_[6774]_  = \new_[7286]_  & \new_[11526]_ ;
  assign \new_[6775]_  = \new_[7286]_  & \new_[10509]_ ;
  assign \new_[6776]_  = ~\new_[7421]_  & ~\new_[8891]_ ;
  assign \new_[6777]_  = ~\new_[7421]_  & ~\new_[9051]_ ;
  assign \new_[6778]_  = ~\new_[7421]_  & ~\new_[9042]_ ;
  assign \new_[6779]_  = ~\new_[7421]_  & ~\new_[9137]_ ;
  assign \new_[6780]_  = ~\new_[7421]_  & ~\new_[9125]_ ;
  assign \new_[6781]_  = ~\new_[7421]_  & ~\new_[9034]_ ;
  assign \new_[6782]_  = ~\new_[7421]_  & ~\new_[9286]_ ;
  assign \new_[6783]_  = ~\new_[7421]_  & ~\new_[9365]_ ;
  assign \new_[6784]_  = ~\new_[7421]_  & ~\new_[9120]_ ;
  assign \new_[6785]_  = ~\new_[7421]_  & ~\new_[9074]_ ;
  assign \new_[6786]_  = ~\new_[6827]_  | ~\new_[7111]_ ;
  assign \new_[6787]_  = ~\new_[7421]_  & ~\new_[9122]_ ;
  assign \new_[6788]_  = ~\new_[7421]_  & ~\new_[9132]_ ;
  assign \new_[6789]_  = ~\new_[7421]_  & ~\new_[9159]_ ;
  assign \new_[6790]_  = ~\new_[7421]_  & ~\new_[9079]_ ;
  assign \new_[6791]_  = ~\new_[7421]_  & ~\new_[9095]_ ;
  assign \new_[6792]_  = ~\new_[7421]_  & ~\new_[9046]_ ;
  assign \new_[6793]_  = ~\new_[7421]_  & ~\new_[9091]_ ;
  assign \new_[6794]_  = ~\new_[7421]_  & ~\new_[9112]_ ;
  assign \new_[6795]_  = ~\new_[7421]_  & ~\new_[9325]_ ;
  assign \new_[6796]_  = ~\new_[7421]_  & ~\new_[8899]_ ;
  assign \new_[6797]_  = ~\new_[7421]_  & ~\new_[9049]_ ;
  assign \new_[6798]_  = ~\new_[7421]_  & ~\new_[9097]_ ;
  assign \new_[6799]_  = ~\new_[7421]_  & ~\new_[9084]_ ;
  assign \new_[6800]_  = ~\new_[7421]_  & ~\new_[9124]_ ;
  assign \new_[6801]_  = ~\new_[7421]_  & ~\new_[9098]_ ;
  assign \new_[6802]_  = ~\new_[7421]_  & ~\new_[9088]_ ;
  assign \new_[6803]_  = ~\new_[7421]_  & ~\new_[9149]_ ;
  assign \new_[6804]_  = ~\new_[6837]_ ;
  assign \new_[6805]_  = ~\new_[12736]_  | ~\new_[7363]_ ;
  assign \new_[6806]_  = ~\new_[7074]_ ;
  assign \new_[6807]_  = ~\new_[7075]_ ;
  assign \new_[6808]_  = ~\new_[7078]_ ;
  assign \new_[6809]_  = ~\new_[7020]_ ;
  assign \new_[6810]_  = \new_[7008]_ ;
  assign \new_[6811]_  = (~\new_[9713]_  | ~\new_[7807]_ ) & (~\new_[7763]_  | ~\new_[10767]_ );
  assign \new_[6812]_  = ~\new_[7707]_  & (~\new_[11731]_  | ~\new_[11726]_ );
  assign \new_[6813]_  = \new_[9709]_  ? \new_[7763]_  : \new_[11328]_ ;
  assign \new_[6814]_  = \new_[10115]_  ? \new_[7763]_  : \new_[11367]_ ;
  assign \new_[6815]_  = \new_[9684]_  ? \new_[7763]_  : \new_[11361]_ ;
  assign \new_[6816]_  = \new_[9599]_  ? \new_[7763]_  : \new_[10419]_ ;
  assign \new_[6817]_  = \new_[9990]_  ? \new_[7763]_  : \new_[10509]_ ;
  assign \new_[6818]_  = \new_[9407]_  ? \new_[7763]_  : \new_[10526]_ ;
  assign \new_[6819]_  = \new_[10037]_  ? \new_[7763]_  : \new_[10919]_ ;
  assign \new_[6820]_  = ~\new_[9896]_  | ~\new_[7291]_ ;
  assign \new_[6821]_  = ~\new_[7111]_ ;
  assign \new_[6822]_  = ~\new_[7111]_ ;
  assign \new_[6823]_  = ~\new_[7111]_ ;
  assign \new_[6824]_  = ~\new_[7111]_ ;
  assign \new_[6825]_  = ~\new_[7111]_ ;
  assign \new_[6826]_  = ~\new_[7112]_ ;
  assign \new_[6827]_  = ~\new_[12002]_ ;
  assign \new_[6828]_  = \new_[12002]_ ;
  assign \new_[6829]_  = ~\new_[6828]_ ;
  assign \new_[6830]_  = ~\new_[7266]_ ;
  assign \new_[6831]_  = ~\new_[7266]_ ;
  assign \new_[6832]_  = \new_[7115]_ ;
  assign \new_[6833]_  = \new_[7373]_  | \new_[7288]_ ;
  assign \new_[6834]_  = ~\new_[7701]_  | ~\new_[11726]_ ;
  assign \new_[6835]_  = ~\new_[7286]_ ;
  assign \new_[6836]_  = ~\new_[11727]_ ;
  assign \new_[6837]_  = ~\new_[7701]_  | ~\new_[11718]_  | ~\new_[7717]_ ;
  assign \new_[6838]_  = ~\new_[11014]_  | ~\new_[12619]_ ;
  assign \new_[6839]_  = ~\new_[11206]_  | ~\new_[12622]_ ;
  assign \new_[6840]_  = ~\new_[7386]_  & (~\new_[7385]_  | ~\new_[11333]_ );
  assign \new_[6841]_  = ~\new_[12737]_  | (~\new_[7866]_  & ~\new_[7479]_ );
  assign n3316 = \new_[2833]_  ? \new_[7433]_  : \new_[6455]_ ;
  assign n3191 = \new_[2721]_  ? \new_[7433]_  : \new_[6428]_ ;
  assign n3381 = \new_[2769]_  ? \new_[7433]_  : \new_[11063]_ ;
  assign n3366 = \new_[2839]_  ? \new_[7433]_  : \new_[6542]_ ;
  assign n3376 = \new_[2840]_  ? \new_[7433]_  : \new_[6544]_ ;
  assign n3336 = \new_[2829]_  ? \new_[7433]_  : \new_[6490]_ ;
  assign n3356 = \new_[2841]_  ? \new_[7433]_  : \new_[6529]_ ;
  assign n3196 = \new_[2842]_  ? \new_[7433]_  : \new_[6429]_ ;
  assign n3346 = \new_[2830]_  ? \new_[7433]_  : \new_[6518]_ ;
  assign n3361 = \new_[2843]_  ? \new_[7433]_  : \new_[6537]_ ;
  assign n2946 = \new_[2845]_  ? \new_[7433]_  : \new_[6323]_ ;
  assign n3026 = \new_[2768]_  ? \new_[7433]_  : \new_[6382]_ ;
  assign n2981 = \new_[2833]_  ? \new_[7430]_  : \new_[6333]_ ;
  assign n2961 = \new_[2720]_  ? \new_[7430]_  : \new_[6329]_ ;
  assign n3281 = \new_[2721]_  ? \new_[7430]_  : \new_[6447]_ ;
  assign n3286 = \new_[2769]_  ? \new_[7430]_  : \new_[11147]_ ;
  assign n2966 = \new_[2839]_  ? \new_[7430]_  : \new_[6330]_ ;
  assign n3436 = \new_[2840]_  ? \new_[7430]_  : \new_[6643]_ ;
  assign n3291 = \new_[2829]_  ? \new_[7430]_  : \new_[6450]_ ;
  assign n3351 = \new_[2841]_  ? \new_[7430]_  : \new_[6523]_ ;
  assign n3296 = \new_[2842]_  ? \new_[7430]_  : \new_[6451]_ ;
  assign n3306 = \new_[2843]_  ? \new_[7430]_  : \new_[6453]_ ;
  assign n3301 = \new_[2830]_  ? \new_[7430]_  : \new_[6452]_ ;
  assign n3311 = \new_[2845]_  ? \new_[7430]_  : \new_[6454]_ ;
  assign \new_[6866]_  = \\u0_cs_reg[0] ;
  assign n3421 = \new_[2768]_  ? \new_[7430]_  : \new_[6606]_ ;
  assign n3386 = \new_[2720]_  ? \new_[7433]_  : \new_[6550]_ ;
  assign n3426 = \new_[2845]_  ? \new_[7431]_  : \new_[6614]_ ;
  assign n3186 = \new_[2829]_  ? \new_[7439]_  : \new_[6427]_ ;
  assign n3086 = \new_[2833]_  ? \new_[12201]_  : \new_[6407]_ ;
  assign n3091 = \new_[2720]_  ? \new_[12201]_  : \new_[6408]_ ;
  assign n3096 = \new_[2721]_  ? \new_[12201]_  : \new_[6409]_ ;
  assign n2976 = \new_[2769]_  ? \new_[12201]_  : \new_[11180]_ ;
  assign n3101 = \new_[2839]_  ? \new_[12201]_  : \new_[6410]_ ;
  assign n3106 = \new_[2840]_  ? \new_[12201]_  : \new_[6411]_ ;
  assign n3111 = \new_[2829]_  ? \new_[12201]_  : \new_[6412]_ ;
  assign n2971 = \new_[2841]_  ? \new_[12201]_  : \new_[6331]_ ;
  assign n3116 = \new_[2842]_  ? \new_[12201]_  : \new_[6413]_ ;
  assign n2941 = \new_[2843]_  ? \new_[12201]_  : \new_[6318]_ ;
  assign n3331 = \new_[2830]_  ? \new_[12201]_  : \new_[6471]_ ;
  assign n3431 = \new_[2845]_  ? \new_[12201]_  : \new_[6633]_ ;
  assign n3121 = \new_[2768]_  ? \new_[12201]_  : \new_[6414]_ ;
  assign n3466 = \new_[2833]_  ? \new_[7431]_  : \new_[6653]_ ;
  assign n3166 = \new_[2841]_  ? \new_[7439]_  : \new_[6423]_ ;
  assign n3441 = \new_[2721]_  ? \new_[7431]_  : \new_[6644]_ ;
  assign n3131 = \new_[2769]_  ? \new_[7431]_  : \new_[11025]_ ;
  assign n3461 = \new_[2839]_  ? \new_[7431]_  : \new_[6651]_ ;
  assign n3456 = \new_[2840]_  ? \new_[7431]_  : \new_[6647]_ ;
  assign n3446 = \new_[2829]_  ? \new_[7431]_  : \new_[6645]_ ;
  assign n3136 = \new_[2841]_  ? \new_[7431]_  : \new_[6417]_ ;
  assign n3341 = \new_[2842]_  ? \new_[7431]_  : \new_[6513]_ ;
  assign n3141 = \new_[2843]_  ? \new_[7431]_  : \new_[6418]_ ;
  assign \new_[6894]_  = ~\new_[12567]_  | ~\new_[11776]_  | ~\new_[7418]_ ;
  assign n3406 = \new_[2830]_  ? \new_[7431]_  : \new_[6575]_ ;
  assign n3146 = \new_[2768]_  ? \new_[7431]_  : \new_[6419]_ ;
  assign n3401 = \new_[2833]_  ? \new_[7439]_  : \new_[6570]_ ;
  assign n3151 = \new_[2720]_  ? \new_[7439]_  : \new_[6420]_ ;
  assign n3411 = \new_[2721]_  ? \new_[7439]_  : \new_[6582]_ ;
  assign n3156 = \new_[2769]_  ? \new_[7439]_  : \new_[11139]_ ;
  assign n3171 = \new_[2842]_  ? \new_[7439]_  : \new_[6424]_ ;
  assign n3416 = \new_[2843]_  ? \new_[7439]_  : \new_[6588]_ ;
  assign n3391 = \new_[2830]_  ? \new_[7439]_  : \new_[6552]_ ;
  assign n3176 = \new_[2845]_  ? \new_[7439]_  : \new_[6425]_ ;
  assign n3181 = \new_[2768]_  ? \new_[7439]_  : \new_[6426]_ ;
  assign n3056 = \new_[2833]_  ? \new_[12208]_  : \new_[6390]_ ;
  assign n3321 = \new_[2720]_  ? \new_[12208]_  : \new_[6458]_ ;
  assign n3201 = \new_[2721]_  ? \new_[12208]_  : \new_[6430]_ ;
  assign n3206 = \new_[2769]_  ? \new_[12208]_  : \new_[11183]_ ;
  assign n3326 = \new_[2839]_  ? \new_[12208]_  : \new_[6467]_ ;
  assign n3081 = \new_[2840]_  ? \new_[12208]_  : \new_[6405]_ ;
  assign n3211 = \new_[2829]_  ? \new_[12208]_  : \new_[6433]_ ;
  assign n3216 = \new_[2841]_  ? \new_[12208]_  : \new_[6434]_ ;
  assign n3076 = \new_[2842]_  ? \new_[12208]_  : \new_[6404]_ ;
  assign n3221 = \new_[2843]_  ? \new_[12208]_  : \new_[6435]_ ;
  assign n3066 = \new_[2830]_  ? \new_[12208]_  : \new_[6401]_ ;
  assign n3226 = \new_[2845]_  ? \new_[12208]_  : \new_[6436]_ ;
  assign n3071 = \new_[2768]_  ? \new_[12208]_  : \new_[6403]_ ;
  assign n3231 = \new_[2833]_  ? \new_[7427]_  : \new_[6437]_ ;
  assign n3061 = \new_[2720]_  ? \new_[7427]_  : \new_[6392]_ ;
  assign n3236 = \new_[2721]_  ? \new_[7427]_  : \new_[6438]_ ;
  assign n3021 = \new_[2769]_  ? \new_[7427]_  : \new_[11004]_ ;
  assign n3241 = \new_[2839]_  ? \new_[7427]_  : \new_[6439]_ ;
  assign n3051 = \new_[2840]_  ? \new_[7427]_  : \new_[6389]_ ;
  assign n3246 = \new_[2829]_  ? \new_[7427]_  : \new_[6440]_ ;
  assign n3031 = \new_[2841]_  ? \new_[7427]_  : \new_[6385]_ ;
  assign n3046 = \new_[2842]_  ? \new_[7427]_  : \new_[6388]_ ;
  assign n3041 = \new_[2843]_  ? \new_[7427]_  : \new_[6387]_ ;
  assign n3036 = \new_[2830]_  ? \new_[7427]_  : \new_[6386]_ ;
  assign n3016 = \new_[2845]_  ? \new_[7427]_  : \new_[6370]_ ;
  assign n2951 = \new_[2833]_  ? \new_[7429]_  : \new_[6324]_ ;
  assign n3251 = \new_[2768]_  ? \new_[7427]_  : \new_[6441]_ ;
  assign n3256 = \new_[2720]_  ? \new_[7429]_  : \new_[6442]_ ;
  assign n3011 = \new_[2721]_  ? \new_[7429]_  : \new_[6368]_ ;
  assign n3006 = \new_[2769]_  ? \new_[7429]_  : \new_[11123]_ ;
  assign n3001 = \new_[2839]_  ? \new_[7429]_  : \new_[6362]_ ;
  assign n3261 = \new_[2840]_  ? \new_[7429]_  : \new_[6443]_ ;
  assign n2996 = \new_[2829]_  ? \new_[7429]_  : \new_[6341]_ ;
  assign n3266 = \new_[2841]_  ? \new_[7429]_  : \new_[6444]_ ;
  assign n3271 = \new_[2842]_  ? \new_[7429]_  : \new_[6445]_ ;
  assign n3276 = \new_[2843]_  ? \new_[7429]_  : \new_[6446]_ ;
  assign n2986 = \new_[2830]_  ? \new_[7429]_  : \new_[6334]_ ;
  assign n2956 = \new_[2845]_  ? \new_[7429]_  : \new_[6326]_ ;
  assign n2991 = \new_[2768]_  ? \new_[7429]_  : \new_[6335]_ ;
  assign n3161 = \new_[2840]_  ? \new_[7439]_  : \new_[6422]_ ;
  assign n3396 = \new_[2839]_  ? \new_[7439]_  : \new_[6562]_ ;
  assign n3126 = \new_[2720]_  ? \new_[7431]_  : \new_[6415]_ ;
  assign \new_[6948]_  = ~\new_[7307]_  & ~\new_[11404]_ ;
  assign \new_[6949]_  = ~\new_[7307]_  & ~\new_[11403]_ ;
  assign \new_[6950]_  = ~\new_[10291]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[6951]_  = ~\new_[12273]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6952]_  = ~\new_[10922]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6953]_  = ~\new_[10743]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[6954]_  = ~\new_[11355]_  | ~\new_[10367]_  | ~\new_[7417]_ ;
  assign \new_[6955]_  = ~\new_[11363]_  | ~\new_[11776]_  | ~\new_[7418]_ ;
  assign \new_[6956]_  = ~\new_[10963]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6957]_  = ~\new_[11576]_  | ~\new_[11776]_  | ~\new_[7418]_ ;
  assign \new_[6958]_  = ~\new_[9647]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6959]_  = ~\new_[11332]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6960]_  = ~\new_[10177]_  | ~\new_[10367]_  | ~\new_[7417]_ ;
  assign \new_[6961]_  = ~\new_[11343]_  | ~\new_[10367]_  | ~\new_[7772]_ ;
  assign \new_[6962]_  = ~\new_[11356]_  | ~\new_[10367]_  | ~\new_[7772]_ ;
  assign \new_[6963]_  = ~\new_[11340]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6964]_  = ~\new_[11492]_  | ~\new_[11776]_  | ~\new_[7417]_ ;
  assign \new_[6965]_  = ~\new_[11320]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6966]_  = ~\new_[11298]_  | ~\new_[11776]_  | ~\new_[7417]_ ;
  assign \new_[6967]_  = ~\new_[12089]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6968]_  = ~\new_[11500]_  | ~\new_[10045]_ ;
  assign \new_[6969]_  = ~\new_[11500]_  | ~\new_[9856]_ ;
  assign \new_[6970]_  = ~\new_[12554]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[6971]_  = ~\new_[11500]_  | ~\new_[9594]_ ;
  assign \new_[6972]_  = ~\new_[7363]_  | ~\new_[7296]_  | ~\new_[7999]_ ;
  assign \new_[6973]_  = ~\new_[10250]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6974]_  = ~\new_[12755]_  | ~\new_[11776]_  | ~\new_[7417]_ ;
  assign \new_[6975]_  = \new_[7291]_  & \new_[9772]_ ;
  assign \new_[6976]_  = ~\new_[11500]_  | ~\new_[10059]_ ;
  assign \new_[6977]_  = ~\new_[11353]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6978]_  = ~\new_[7294]_  & ~\new_[7432]_ ;
  assign \new_[6979]_  = ~\new_[10164]_  | ~\new_[11776]_  | ~\new_[7418]_ ;
  assign \new_[6980]_  = ~\new_[11328]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6981]_  = ~\new_[11366]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[6982]_  = ~\new_[11500]_  | ~\new_[9870]_ ;
  assign \new_[6983]_  = ~\new_[10419]_  | ~\new_[10367]_  | ~\new_[7417]_ ;
  assign \new_[6984]_  = ~\new_[7156]_ ;
  assign \new_[6985]_  = ~\new_[7156]_ ;
  assign \new_[6986]_  = ~\new_[7156]_ ;
  assign \new_[6987]_  = ~\new_[11500]_  | ~\new_[10056]_ ;
  assign \new_[6988]_  = ~\new_[11526]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6989]_  = ~\new_[12044]_  | ~\new_[11776]_  | ~\new_[7417]_ ;
  assign \new_[6990]_  = ~\new_[10509]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[6991]_  = ~\new_[10526]_  | ~\new_[10367]_  | ~\new_[7417]_ ;
  assign \new_[6992]_  = ~\new_[10919]_  | ~\new_[10367]_  | ~\new_[7521]_ ;
  assign \new_[6993]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7480]_ ;
  assign \new_[6994]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7651]_ ;
  assign \new_[6995]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7496]_ ;
  assign \new_[6996]_  = ~\new_[11491]_  | ~\new_[7289]_  | ~\new_[7501]_ ;
  assign \new_[6997]_  = ~\new_[7865]_  | ~\new_[12388]_  | ~\new_[7365]_ ;
  assign \new_[6998]_  = ~\new_[7160]_ ;
  assign \new_[6999]_  = ~\new_[7115]_ ;
  assign \new_[7000]_  = ~\new_[7541]_  | (~\new_[7422]_  & ~\new_[10827]_ );
  assign \new_[7001]_  = ~\new_[7111]_ ;
  assign \new_[7002]_  = \new_[3225]_  ^ \new_[7587]_ ;
  assign \new_[7003]_  = ~\new_[12512]_ ;
  assign \new_[7004]_  = ~\new_[11263]_  & ~\new_[12665]_ ;
  assign \new_[7005]_  = ~\new_[7168]_ ;
  assign \new_[7006]_  = ~\new_[7329]_  | (~\new_[11776]_  & ~\new_[10963]_ );
  assign \new_[7007]_  = ~\new_[7169]_ ;
  assign \new_[7008]_  = \new_[12472]_ ;
  assign \new_[7009]_  = ~\new_[7226]_  | ~\new_[10083]_ ;
  assign \new_[7010]_  = ~\new_[7326]_  | ~\new_[12069]_ ;
  assign \new_[7011]_  = ~\new_[11434]_ ;
  assign \new_[7012]_  = ~\new_[11774]_  | ~\new_[12382]_ ;
  assign \new_[7013]_  = \new_[12787]_  | \new_[7572]_ ;
  assign \new_[7014]_  = ~\new_[12477]_  | ~\new_[7774]_ ;
  assign \new_[7015]_  = ~\new_[7226]_  | ~\new_[9978]_ ;
  assign \new_[7016]_  = ~\new_[12584]_  | ~\new_[12382]_ ;
  assign \new_[7017]_  = ~\new_[7633]_  | ~\new_[12697]_  | ~\new_[11263]_ ;
  assign \new_[7018]_  = ~\new_[12665]_  & ~\new_[12697]_ ;
  assign \new_[7019]_  = ~\new_[7924]_  & ~\new_[7328]_ ;
  assign \new_[7020]_  = ~\new_[11773]_ ;
  assign \new_[7021]_  = ~\new_[11450]_ ;
  assign \new_[7022]_  = \new_[7238]_ ;
  assign \new_[7023]_  = (~\new_[7708]_  | ~\new_[11058]_ ) & (~\new_[2927]_  | ~\new_[1711]_ );
  assign \new_[7024]_  = (~\new_[7369]_  | ~\new_[9350]_ ) & (~\new_[7597]_  | ~\wb_addr_i[17] );
  assign \new_[7025]_  = (~\new_[7369]_  | ~\new_[9334]_ ) & (~\new_[7597]_  | ~\wb_addr_i[2] );
  assign \new_[7026]_  = (~\new_[7369]_  | ~\new_[9339]_ ) & (~\new_[7597]_  | ~\wb_addr_i[5] );
  assign \new_[7027]_  = (~\new_[7369]_  | ~\new_[9184]_ ) & (~\new_[7597]_  | ~\wb_addr_i[20] );
  assign \new_[7028]_  = (~\new_[7369]_  | ~\new_[9366]_ ) & (~\new_[7597]_  | ~\wb_addr_i[21] );
  assign \new_[7029]_  = (~\new_[7369]_  | ~\new_[9257]_ ) & (~\new_[7597]_  | ~\wb_addr_i[23] );
  assign \new_[7030]_  = (~\new_[7369]_  | ~\new_[9306]_ ) & (~\new_[7597]_  | ~\wb_addr_i[25] );
  assign \new_[7031]_  = (~\new_[7369]_  | ~\new_[9179]_ ) & (~\new_[7597]_  | ~\wb_addr_i[8] );
  assign \new_[7032]_  = (~\new_[7369]_  | ~\new_[9207]_ ) & (~\new_[7597]_  | ~\wb_addr_i[22] );
  assign \new_[7033]_  = (~\new_[7369]_  | ~\new_[9333]_ ) & (~\new_[7597]_  | ~\wb_addr_i[12] );
  assign \new_[7034]_  = (~\new_[7369]_  | ~\new_[9369]_ ) & (~\new_[7597]_  | ~\wb_addr_i[24] );
  assign \new_[7035]_  = (~\new_[7369]_  | ~\new_[9176]_ ) & (~\new_[7597]_  | ~\wb_addr_i[7] );
  assign \new_[7036]_  = (~\new_[7369]_  | ~\new_[9332]_ ) & (~\new_[7597]_  | ~\wb_addr_i[4] );
  assign \new_[7037]_  = (~\new_[7369]_  | ~\new_[9380]_ ) & (~\new_[7597]_  | ~\wb_addr_i[11] );
  assign \new_[7038]_  = (~\new_[7369]_  | ~\new_[9362]_ ) & (~\new_[7597]_  | ~\wb_addr_i[14] );
  assign \new_[7039]_  = (~\new_[7369]_  | ~\new_[9347]_ ) & (~\new_[7597]_  | ~\wb_addr_i[9] );
  assign \new_[7040]_  = (~\new_[7369]_  | ~\new_[9373]_ ) & (~\new_[7597]_  | ~\wb_addr_i[19] );
  assign \new_[7041]_  = (~\new_[7369]_  | ~\new_[9364]_ ) & (~\new_[7597]_  | ~\wb_addr_i[6] );
  assign \new_[7042]_  = (~\new_[7369]_  | ~\new_[9335]_ ) & (~\new_[7597]_  | ~\wb_addr_i[18] );
  assign \new_[7043]_  = (~\new_[7369]_  | ~\new_[9331]_ ) & (~\new_[7597]_  | ~\wb_addr_i[13] );
  assign \new_[7044]_  = (~\new_[7369]_  | ~\new_[9354]_ ) & (~\new_[7597]_  | ~\wb_addr_i[3] );
  assign \new_[7045]_  = (~\new_[7369]_  | ~\new_[9337]_ ) & (~\new_[7597]_  | ~\wb_addr_i[10] );
  assign \new_[7046]_  = ~\new_[12453]_  | ~\new_[10367]_  | ~\new_[7772]_ ;
  assign \new_[7047]_  = \new_[7267]_  & \new_[12598]_ ;
  assign \new_[7048]_  = \new_[7267]_  & \new_[10808]_ ;
  assign \new_[7049]_  = \new_[7286]_  & \new_[10838]_ ;
  assign \new_[7050]_  = \new_[7286]_  & \new_[9785]_ ;
  assign \new_[7051]_  = \new_[7267]_  & \new_[10634]_ ;
  assign \new_[7052]_  = ~\new_[7421]_  & ~\new_[8905]_ ;
  assign \new_[7053]_  = ~\new_[7421]_  & ~\new_[9642]_ ;
  assign \new_[7054]_  = ~\new_[7190]_ ;
  assign \new_[7055]_  = ~\new_[7421]_  & ~\new_[9288]_ ;
  assign \new_[7056]_  = ~\new_[7421]_  & ~\new_[9081]_ ;
  assign \new_[7057]_  = ~\new_[7421]_  & ~\new_[9090]_ ;
  assign \new_[7058]_  = ~\new_[7421]_  & ~\new_[9664]_ ;
  assign \new_[7059]_  = ~\new_[7213]_ ;
  assign \new_[7060]_  = ~\new_[7136]_ ;
  assign \new_[7061]_  = ~\new_[7134]_ ;
  assign n3371 = ~\new_[9806]_  | ~\new_[7268]_ ;
  assign \new_[7063]_  = ~\new_[7365]_  | ~\new_[12736]_ ;
  assign \new_[7064]_  = ~\new_[7421]_  & ~\new_[8903]_ ;
  assign \new_[7065]_  = ~\new_[7219]_ ;
  assign \new_[7066]_  = ~\new_[12780]_  & ~n3451;
  assign \new_[7067]_  = ~\new_[7227]_ ;
  assign \new_[7068]_  = ~\new_[7421]_  & ~\new_[9080]_ ;
  assign \new_[7069]_  = ~\new_[12234]_  | ~\new_[12736]_ ;
  assign \new_[7070]_  = ~\new_[7421]_  & ~\new_[8929]_ ;
  assign \new_[7071]_  = ~\new_[10496]_  | ~\new_[11776]_  | ~\new_[7772]_ ;
  assign \new_[7072]_  = ~\new_[7235]_ ;
  assign \new_[7073]_  = ~\new_[10846]_  | ~\new_[7592]_  | ~\new_[11973]_ ;
  assign \new_[7074]_  = ~\new_[7274]_  | ~\new_[7714]_ ;
  assign \new_[7075]_  = ~\new_[7238]_ ;
  assign \new_[7076]_  = \new_[7238]_ ;
  assign \new_[7077]_  = ~\new_[7182]_ ;
  assign \new_[7078]_  = ~\new_[11773]_ ;
  assign \new_[7079]_  = ~\new_[12472]_ ;
  assign \new_[7080]_  = \new_[9383]_  ? \new_[7763]_  : \new_[10291]_ ;
  assign \new_[7081]_  = \new_[10099]_  ? \new_[7763]_  : \new_[11355]_ ;
  assign \new_[7082]_  = \new_[9963]_  ? \new_[7763]_  : \new_[10928]_ ;
  assign \new_[7083]_  = \new_[10104]_  ? \new_[7763]_  : \new_[9997]_ ;
  assign \new_[7084]_  = \new_[10128]_  ? \new_[7763]_  : \new_[11576]_ ;
  assign \new_[7085]_  = \new_[9607]_  ? \new_[7763]_  : \new_[10962]_ ;
  assign \new_[7086]_  = \new_[9604]_  ? \new_[7763]_  : \new_[11526]_ ;
  assign \new_[7087]_  = \new_[10097]_  ? \new_[7763]_  : \new_[11353]_ ;
  assign \new_[7088]_  = \new_[10011]_  ? \new_[7763]_  : \new_[11332]_ ;
  assign \new_[7089]_  = \new_[9680]_  ? \new_[7763]_  : \new_[10177]_ ;
  assign \new_[7090]_  = \new_[10263]_  ? \new_[7763]_  : \new_[11343]_ ;
  assign \new_[7091]_  = \new_[9619]_  ? \new_[7763]_  : \new_[11356]_ ;
  assign \new_[7092]_  = \new_[9845]_  ? \new_[7763]_  : \new_[11340]_ ;
  assign \new_[7093]_  = \new_[10237]_  ? \new_[7763]_  : \new_[10243]_ ;
  assign \new_[7094]_  = \new_[9660]_  ? \new_[7763]_  : \new_[11320]_ ;
  assign \new_[7095]_  = \new_[9418]_  ? \new_[7763]_  : \new_[10938]_ ;
  assign \new_[7096]_  = \new_[10126]_  ? \new_[7763]_  : \new_[11735]_ ;
  assign \new_[7097]_  = \new_[9641]_  ? \new_[7763]_  : \new_[9913]_ ;
  assign \new_[7098]_  = \new_[10287]_  ? \new_[7763]_  : \new_[11316]_ ;
  assign \new_[7099]_  = \new_[9567]_  ? \new_[7763]_  : \new_[11310]_ ;
  assign \new_[7100]_  = \new_[9958]_  ? \new_[7763]_  : \new_[10802]_ ;
  assign \new_[7101]_  = \new_[9326]_  ? \new_[7763]_  : \new_[12093]_ ;
  assign \new_[7102]_  = \new_[9388]_  ? \new_[7763]_  : \new_[10743]_ ;
  assign \new_[7103]_  = \new_[9644]_  ? \new_[7763]_  : \new_[10164]_ ;
  assign \new_[7104]_  = \new_[9655]_  ? \new_[7763]_  : \new_[12453]_ ;
  assign \new_[7105]_  = \new_[10019]_  ? \new_[7763]_  : \new_[10902]_ ;
  assign \new_[7106]_  = \new_[8977]_  ? \new_[7763]_  : \new_[10496]_ ;
  assign \new_[7107]_  = \new_[9707]_  ? \new_[7763]_  : \new_[11313]_ ;
  assign \new_[7108]_  = \new_[9675]_  ? \new_[7763]_  : \new_[10955]_ ;
  assign \new_[7109]_  = ~\new_[7264]_ ;
  assign \new_[7110]_  = \new_[7289]_ ;
  assign \new_[7111]_  = ~\new_[7289]_ ;
  assign \new_[7112]_  = ~\new_[7287]_ ;
  assign \new_[7113]_  = \new_[12002]_ ;
  assign \new_[7114]_  = \new_[3138]_  ^ \new_[7604]_ ;
  assign \new_[7115]_  = ~\new_[7266]_ ;
  assign \new_[7116]_  = ~\new_[7367]_ ;
  assign \new_[7117]_  = ~\new_[7367]_ ;
  assign \new_[7118]_  = ~\new_[7717]_  | ~\new_[7373]_ ;
  assign \new_[7119]_  = \\u3_u0_rd_adr_reg[3] ;
  assign \new_[7120]_  = \new_[11101]_  ? \new_[12622]_  : \new_[11244]_ ;
  assign \new_[7121]_  = \new_[11225]_  ? \new_[12622]_  : \new_[11044]_ ;
  assign \new_[7122]_  = ~\new_[10955]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7123]_  = \new_[11024]_  ? \new_[12622]_  : \new_[11002]_ ;
  assign \new_[7124]_  = \new_[11169]_  ? \new_[12622]_  : \new_[11216]_ ;
  assign \new_[7125]_  = ~\new_[11037]_  | ~\new_[12621]_ ;
  assign \new_[7126]_  = ~\new_[11155]_  | ~\new_[12621]_ ;
  assign \new_[7127]_  = ~\new_[7271]_ ;
  assign \new_[7128]_  = ~\new_[7272]_ ;
  assign \new_[7129]_  = ~\new_[7273]_ ;
  assign \new_[7130]_  = \new_[7731]_  | \new_[7689]_ ;
  assign \new_[7131]_  = ~\new_[11572]_  | ~\new_[7385]_  | ~\new_[10516]_ ;
  assign \new_[7132]_  = ~\new_[7728]_  & ~\new_[7689]_ ;
  assign \new_[7133]_  = ~\new_[10411]_  | ~\new_[11776]_  | ~\new_[7744]_ ;
  assign \new_[7134]_  = ~\new_[7327]_ ;
  assign \new_[7135]_  = u2_bank_open_reg;
  assign \new_[7136]_  = ~\new_[11813]_ ;
  assign \new_[7137]_  = ~\new_[10827]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7138]_  = ~\new_[11348]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7139]_  = ~\new_[10928]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7140]_  = ~\new_[11361]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7141]_  = ~\new_[7479]_  | ~\new_[12573]_ ;
  assign \new_[7142]_  = ~\new_[10808]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7143]_  = \new_[12070]_  | \new_[9774]_ ;
  assign \new_[7144]_  = ~\new_[10243]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7145]_  = ~\new_[9913]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7146]_  = ~\new_[11316]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7147]_  = ~\new_[10802]_  | ~\new_[11776]_  | ~\new_[7744]_ ;
  assign \new_[7148]_  = ~\new_[12093]_  | ~\new_[11776]_  | ~\new_[7744]_ ;
  assign \new_[7149]_  = ~n5021 | ~\new_[11776]_  | ~\new_[7744]_ ;
  assign \new_[7150]_  = \\u3_u0_rd_adr_reg[0] ;
  assign \new_[7151]_  = \\u3_u0_rd_adr_reg[2] ;
  assign \new_[7152]_  = \\u3_u0_rd_adr_reg[1] ;
  assign \new_[7153]_  = ~\new_[12610]_  | ~\new_[11776]_  | ~\new_[7744]_ ;
  assign \new_[7154]_  = ~\new_[7689]_  | ~\new_[12605]_ ;
  assign \new_[7155]_  = ~\new_[7283]_ ;
  assign \new_[7156]_  = ~\new_[7428]_  | ~\new_[10001]_ ;
  assign \new_[7157]_  = ~\new_[12536]_ ;
  assign \new_[7158]_  = ~\new_[9946]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7159]_  = ~\new_[7438]_  & (~\new_[7806]_  | ~\new_[12696]_ );
  assign \new_[7160]_  = ~\new_[9055]_  | ~\new_[7770]_  | ~\new_[10240]_  | ~\new_[10516]_ ;
  assign \new_[7161]_  = ~\new_[12075]_ ;
  assign \new_[7162]_  = ~\new_[10902]_  | ~\new_[10367]_  | ~\new_[7744]_ ;
  assign \new_[7163]_  = \new_[7587]_  & \new_[3225]_ ;
  assign \new_[7164]_  = ~\new_[7664]_  & ~\new_[11881]_ ;
  assign \new_[7165]_  = ~\new_[12673]_  | ~\new_[9785]_ ;
  assign \new_[7166]_  = ~\new_[7664]_  & ~\new_[10160]_ ;
  assign \new_[7167]_  = ~\new_[7292]_ ;
  assign \new_[7168]_  = \new_[7662]_  & \new_[12696]_ ;
  assign \new_[7169]_  = ~\new_[7191]_  | ~\new_[7366]_ ;
  assign \new_[7170]_  = ~\new_[11297]_  | ~\new_[9849]_ ;
  assign \new_[7171]_  = ~\new_[7633]_  | ~\new_[11263]_  | ~\new_[12697]_ ;
  assign \new_[7172]_  = ~\new_[11846]_ ;
  assign \new_[7173]_  = ~\new_[7925]_  & ~\new_[7368]_ ;
  assign \new_[7174]_  = ~\new_[7298]_ ;
  assign \new_[7175]_  = ~\new_[7226]_  & ~\new_[7560]_ ;
  assign \new_[7176]_  = ~\new_[11894]_ ;
  assign \new_[7177]_  = ~\new_[7538]_  & ~\new_[8016]_ ;
  assign \new_[7178]_  = ~\new_[7301]_ ;
  assign \new_[7179]_  = ~\new_[7545]_  & ~\new_[7690]_ ;
  assign \new_[7180]_  = ~\new_[10799]_  | ~\new_[10933]_  | ~\new_[7525]_  | ~\new_[10471]_ ;
  assign \new_[7181]_  = u2_row_same_reg;
  assign \new_[7182]_  = \new_[11774]_ ;
  assign \new_[7183]_  = ~\new_[10964]_  | ~\new_[11140]_  | ~\new_[7532]_  | ~\new_[12040]_ ;
  assign \new_[7184]_  = ~\new_[7662]_  & (~\new_[7805]_  | ~\new_[11337]_ );
  assign \new_[7185]_  = ~\new_[11808]_ ;
  assign \new_[7186]_  = ~\new_[7305]_ ;
  assign \new_[7187]_  = ~\new_[7309]_ ;
  assign \new_[7188]_  = ~\new_[7421]_  & ~\new_[9096]_ ;
  assign \new_[7189]_  = ~\new_[7995]_  | ~\new_[10062]_ ;
  assign \new_[7190]_  = ~\new_[12238]_  | ~\new_[11776]_ ;
  assign \new_[7191]_  = ~\new_[7664]_ ;
  assign \new_[7192]_  = ~\new_[7421]_  & ~\new_[9083]_ ;
  assign \new_[7193]_  = ~\new_[7421]_  & ~\new_[9192]_ ;
  assign \new_[7194]_  = ~\new_[7421]_  & ~\new_[9030]_ ;
  assign \new_[7195]_  = ~\new_[7421]_  & ~\new_[9289]_ ;
  assign \new_[7196]_  = ~\new_[7421]_  & ~\new_[9568]_ ;
  assign \new_[7197]_  = ~\new_[12238]_  & ~\new_[7419]_ ;
  assign \new_[7198]_  = ~\new_[7995]_  | ~\new_[9659]_ ;
  assign \new_[7199]_  = ~\new_[7421]_  & ~\new_[9287]_ ;
  assign \new_[7200]_  = ~\new_[7682]_  | ~\new_[9621]_ ;
  assign \new_[7201]_  = ~\new_[7421]_  & ~\new_[8987]_ ;
  assign \new_[7202]_  = ~\new_[7421]_  & ~\new_[9296]_ ;
  assign \new_[7203]_  = ~\new_[7421]_  & ~\new_[9291]_ ;
  assign \new_[7204]_  = ~\new_[7421]_  & ~\new_[9290]_ ;
  assign \new_[7205]_  = ~\new_[7421]_  & ~\new_[9078]_ ;
  assign \new_[7206]_  = ~\new_[7421]_  & ~\new_[9037]_ ;
  assign \new_[7207]_  = ~\new_[7421]_  & ~\new_[9578]_ ;
  assign \new_[7208]_  = ~\new_[7421]_  & ~\new_[9115]_ ;
  assign \new_[7209]_  = ~\new_[7995]_  | ~\new_[9598]_ ;
  assign \new_[7210]_  = ~\new_[7421]_  & ~\new_[9133]_ ;
  assign \new_[7211]_  = ~\new_[7421]_  & ~\new_[9322]_ ;
  assign \new_[7212]_  = ~\new_[7421]_  & ~\new_[9101]_ ;
  assign \new_[7213]_  = \new_[7326]_ ;
  assign \new_[7214]_  = ~\new_[7682]_  | ~\new_[9586]_ ;
  assign \new_[7215]_  = \new_[7327]_ ;
  assign \new_[7216]_  = \new_[7327]_ ;
  assign \new_[7217]_  = ~\new_[7995]_  | ~\new_[11962]_ ;
  assign \new_[7218]_  = ~\new_[7421]_  & ~\new_[9239]_ ;
  assign \new_[7219]_  = \new_[11420]_ ;
  assign \new_[7220]_  = ~\new_[12388]_  | ~\new_[7681]_ ;
  assign \new_[7221]_  = ~\new_[7421]_  & ~\new_[8910]_ ;
  assign \new_[7222]_  = \new_[7863]_  & \new_[7421]_ ;
  assign \new_[7223]_  = ~\new_[7421]_  & ~\new_[9113]_ ;
  assign \new_[7224]_  = ~\new_[7421]_  & ~\new_[9094]_ ;
  assign \new_[7225]_  = ~\new_[7995]_  | ~\new_[11973]_ ;
  assign \new_[7226]_  = ~\new_[12236]_ ;
  assign \new_[7227]_  = ~\new_[7329]_ ;
  assign \new_[7228]_  = ~\new_[7421]_  & ~\new_[9087]_ ;
  assign \new_[7229]_  = ~\new_[7421]_  & ~\new_[8896]_ ;
  assign \new_[7230]_  = ~\new_[7421]_  & ~\new_[9040]_ ;
  assign \new_[7231]_  = ~\new_[7421]_  & ~\new_[9139]_ ;
  assign \new_[7232]_  = ~\new_[7421]_  & ~\new_[8900]_ ;
  assign \new_[7233]_  = ~\new_[7421]_  & ~\new_[9298]_ ;
  assign \new_[7234]_  = ~\new_[7995]_  | ~\new_[9581]_ ;
  assign \new_[7235]_  = ~\new_[7564]_ ;
  assign \new_[7236]_  = ~\new_[11298]_  | ~\new_[12792]_  | ~\new_[10393]_ ;
  assign \new_[7237]_  = ~\new_[12089]_  | ~\new_[12792]_  | ~\new_[10393]_ ;
  assign \new_[7238]_  = ~\new_[11774]_ ;
  assign \new_[7239]_  = ~\new_[7343]_ ;
  assign \new_[7240]_  = ~\new_[12598]_  | ~\new_[12793]_  | ~\new_[10657]_ ;
  assign \new_[7241]_  = ~\new_[11337]_  | ~\new_[12792]_  | ~\new_[10657]_ ;
  assign \new_[7242]_  = ~\new_[12386]_  | ~\new_[8003]_ ;
  assign \new_[7243]_  = ~\new_[9785]_  | ~\new_[12790]_  | ~\new_[10393]_ ;
  assign \new_[7244]_  = ~\new_[12044]_  | ~\new_[12792]_  | ~\new_[10393]_ ;
  assign \new_[7245]_  = (~\new_[10155]_  | ~\new_[7807]_ ) & (~\new_[7909]_  | ~\new_[10920]_ );
  assign \new_[7246]_  = ~\new_[7421]_  & (~\new_[9307]_  | ~\new_[10846]_ );
  assign \new_[7247]_  = \new_[9401]_  ? \new_[7763]_  : \new_[10827]_ ;
  assign \new_[7248]_  = \new_[9665]_  ? \new_[7763]_  : \new_[10960]_ ;
  assign \new_[7249]_  = \new_[9661]_  ? \new_[7763]_  : \new_[11348]_ ;
  assign \new_[7250]_  = \new_[9374]_  ? \new_[7763]_  : \new_[12610]_ ;
  assign \new_[7251]_  = \new_[9987]_  ? \new_[7763]_  : \new_[10108]_ ;
  assign \new_[7252]_  = \new_[9611]_  ? \new_[7763]_  : n5021;
  assign \new_[7253]_  = \new_[9853]_  ? \new_[7763]_  : \new_[12567]_ ;
  assign \new_[7254]_  = \new_[9582]_  ? \new_[7763]_  : \new_[11363]_ ;
  assign \new_[7255]_  = \new_[9104]_  ? \new_[7763]_  : \new_[10411]_ ;
  assign \new_[7256]_  = \new_[9618]_  ? \new_[7763]_  : \new_[9903]_ ;
  assign \new_[7257]_  = \new_[9682]_  ? \new_[7763]_  : \new_[9674]_ ;
  assign \new_[7258]_  = \new_[9978]_  ? \new_[7763]_  : \new_[11337]_ ;
  assign \new_[7259]_  = \new_[9710]_  ? \new_[7763]_  : \new_[11323]_ ;
  assign \new_[7260]_  = \new_[9389]_  ? \new_[7763]_  : \new_[10933]_ ;
  assign \new_[7261]_  = \new_[12110]_  ? \new_[7763]_  : \new_[12044]_ ;
  assign \new_[7262]_  = \new_[10136]_  ? \new_[7909]_  : \new_[10634]_ ;
  assign \new_[7263]_  = ~\new_[7363]_ ;
  assign \new_[7264]_  = ~\new_[7560]_ ;
  assign \new_[7265]_  = \\u4_rfr_cnt_reg[3] ;
  assign \new_[7266]_  = ~\new_[7366]_ ;
  assign \new_[7267]_  = ~\new_[7367]_ ;
  assign \new_[7268]_  = ~\new_[7610]_  | ~wb_we_i;
  assign \new_[7269]_  = \new_[11103]_  ? \new_[12622]_  : \new_[11035]_ ;
  assign \new_[7270]_  = (~\new_[8084]_  | ~\new_[7612]_ ) & (~\new_[7727]_  | ~\new_[11166]_ );
  assign \new_[7271]_  = (~\new_[8084]_  | ~\new_[7618]_ ) & (~\new_[7727]_  | ~\new_[7813]_ );
  assign \new_[7272]_  = (~\new_[8084]_  | ~\new_[7616]_ ) & (~\new_[7727]_  | ~\new_[7828]_ );
  assign \new_[7273]_  = (~\new_[8084]_  | ~\new_[7732]_ ) & (~\new_[7727]_  | ~\new_[7851]_ );
  assign \new_[7274]_  = \new_[7827]_  & \new_[7701]_ ;
  assign \new_[7275]_  = \\u4_rfr_cnt_reg[5] ;
  assign n3471 = \new_[6866]_  ? n5766 : \new_[7765]_ ;
  assign \new_[7277]_  = ~\new_[12049]_  & ~\new_[10286]_ ;
  assign \new_[7278]_  = \\u4_rfr_cnt_reg[6] ;
  assign \new_[7279]_  = \\u4_rfr_cnt_reg[4] ;
  assign \new_[7280]_  = u0_u0_init_req_reg;
  assign \new_[7281]_  = \\u4_rfr_cnt_reg[7] ;
  assign \new_[7282]_  = ~\new_[11374]_ ;
  assign \new_[7283]_  = ~\new_[7635]_  | ~\new_[7990]_ ;
  assign \new_[7284]_  = \\u4_rfr_cnt_reg[2] ;
  assign \new_[7285]_  = \\u4_rfr_cnt_reg[1] ;
  assign \new_[7286]_  = ~\new_[7367]_ ;
  assign \new_[7287]_  = ~\new_[12234]_ ;
  assign \new_[7288]_  = ~\new_[7372]_ ;
  assign \new_[7289]_  = ~\new_[7365]_ ;
  assign \new_[7290]_  = ~\new_[11507]_  | ~\new_[11058]_ ;
  assign \new_[7291]_  = \new_[12664]_  & \new_[10553]_ ;
  assign \new_[7292]_  = \new_[7662]_  | \new_[8957]_ ;
  assign \new_[7293]_  = \new_[7649]_  & \new_[12398]_ ;
  assign \new_[7294]_  = ~\new_[7664]_  & ~\new_[12697]_ ;
  assign \new_[7295]_  = ~\new_[7428]_ ;
  assign \new_[7296]_  = \new_[11502]_  & \new_[7669]_ ;
  assign \new_[7297]_  = ~\new_[12672]_  & ~\new_[10818]_ ;
  assign \new_[7298]_  = ~\new_[11472]_ ;
  assign \new_[7299]_  = ~\new_[7438]_ ;
  assign \new_[7300]_  = ~\new_[7443]_ ;
  assign \new_[7301]_  = \new_[8740]_  | \new_[7662]_ ;
  assign \new_[7302]_  = \new_[7665]_  | \new_[10549]_ ;
  assign \new_[7303]_  = ~\new_[7826]_  | ~\new_[7615]_  | ~\new_[12169]_ ;
  assign \new_[7304]_  = ~\new_[12491]_  & (~\new_[7873]_  | ~\new_[9906]_ );
  assign \new_[7305]_  = ~\new_[7668]_  & (~\new_[12385]_  | ~\new_[10517]_ );
  assign \new_[7306]_  = (~\new_[9375]_  | ~\new_[7683]_ ) & (~\new_[7873]_  | ~\new_[9864]_ );
  assign \new_[7307]_  = ~\new_[7478]_ ;
  assign \new_[7308]_  = ~\new_[10918]_  | ~\new_[8399]_  | ~\new_[10915]_  | ~\new_[7712]_ ;
  assign \new_[7309]_  = ~\new_[7599]_  | ~\new_[10378]_ ;
  assign \new_[7310]_  = ~\new_[7805]_  & ~\new_[10799]_ ;
  assign \new_[7311]_  = ~\new_[7806]_  & ~\new_[10722]_ ;
  assign \new_[7312]_  = ~\new_[7806]_  & ~\new_[10809]_ ;
  assign \new_[7313]_  = ~\new_[7806]_  & ~\new_[11334]_ ;
  assign \new_[7314]_  = ~\new_[7806]_  & ~\new_[11344]_ ;
  assign \new_[7315]_  = ~\new_[7805]_  & ~\new_[11324]_ ;
  assign \new_[7316]_  = ~\new_[7513]_ ;
  assign \new_[7317]_  = ~\new_[7805]_  & ~\new_[12052]_ ;
  assign \new_[7318]_  = ~\new_[7806]_  & ~\new_[10771]_ ;
  assign \new_[7319]_  = ~\new_[7516]_ ;
  assign \new_[7320]_  = ~\new_[7806]_  & ~\new_[11529]_ ;
  assign \new_[7321]_  = ~\new_[7806]_  & ~\new_[10715]_ ;
  assign \new_[7322]_  = ~\new_[7806]_  & ~\new_[10783]_ ;
  assign \new_[7323]_  = ~\new_[7588]_  | ~\new_[10378]_ ;
  assign \new_[7324]_  = ~\new_[7591]_  | ~\new_[12000]_ ;
  assign \new_[7325]_  = ~\new_[12307]_  | ~\new_[9603]_ ;
  assign \new_[7326]_  = \new_[9565]_  | \new_[7596]_ ;
  assign \new_[7327]_  = \new_[11813]_ ;
  assign \new_[7328]_  = ~\new_[11320]_  | ~\new_[11573]_  | ~\new_[7700]_ ;
  assign \new_[7329]_  = \new_[7543]_ ;
  assign \new_[7330]_  = ~\new_[12307]_  | ~\new_[9596]_ ;
  assign \new_[7331]_  = ~\new_[12273]_  | ~\new_[12792]_  | ~\new_[10393]_ ;
  assign \new_[7332]_  = ~\new_[11343]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7333]_  = ~\new_[9913]_  | ~\new_[12790]_  | ~\new_[10314]_ ;
  assign \new_[7334]_  = ~\new_[11316]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7335]_  = ~\new_[10108]_  | ~\new_[12789]_  | ~\new_[10393]_ ;
  assign \new_[7336]_  = ~\new_[10802]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7337]_  = ~\new_[12093]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7338]_  = ~n5021 | ~\new_[12792]_  | ~\new_[10657]_ ;
  assign \new_[7339]_  = ~\new_[10164]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7340]_  = ~\new_[10411]_  | ~\new_[12789]_  | ~\new_[10314]_ ;
  assign \new_[7341]_  = \new_[3177]_  ^ \new_[7725]_ ;
  assign \new_[7342]_  = ~\new_[10902]_  | ~\new_[12790]_  | ~\new_[10314]_ ;
  assign \new_[7343]_  = ~\new_[7571]_ ;
  assign \new_[7344]_  = \new_[7571]_ ;
  assign \new_[7345]_  = ~\new_[12780]_  | (~\new_[10148]_  & ~\new_[12755]_ );
  assign \new_[7346]_  = ~\new_[10933]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7347]_  = ~\new_[11735]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7348]_  = ~\new_[9946]_  | ~\new_[12792]_  | ~\new_[10657]_ ;
  assign \new_[7349]_  = ~\new_[10919]_  | ~\new_[12790]_  | ~\new_[10314]_ ;
  assign \new_[7350]_  = ~\new_[10509]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7351]_  = \new_[9627]_  ? \new_[7763]_  : \new_[10818]_ ;
  assign \new_[7352]_  = \new_[9979]_  ? \new_[7909]_  : \new_[9998]_ ;
  assign \new_[7353]_  = \new_[10039]_  ? \new_[7763]_  : \new_[12273]_ ;
  assign \new_[7354]_  = \new_[10031]_  ? \new_[7909]_  : \new_[10922]_ ;
  assign \new_[7355]_  = \new_[9930]_  ? \new_[7909]_  : \new_[11492]_ ;
  assign \new_[7356]_  = \new_[9980]_  ? \new_[7909]_  : \new_[12598]_ ;
  assign \new_[7357]_  = \new_[10111]_  ? \new_[7763]_  : \new_[11298]_ ;
  assign \new_[7358]_  = \new_[11860]_  ? \new_[7763]_  : \new_[12089]_ ;
  assign \new_[7359]_  = \new_[9936]_  ? \new_[7909]_  : \new_[9785]_ ;
  assign \new_[7360]_  = \new_[9391]_  ? \new_[7909]_  : \new_[12755]_ ;
  assign \new_[7361]_  = \new_[9950]_  ? \new_[7909]_  : \new_[12554]_ ;
  assign \new_[7362]_  = \new_[9107]_  ? \new_[7909]_  : \new_[10250]_ ;
  assign \new_[7363]_  = ~\new_[8705]_  | ~\new_[10022]_  | ~\new_[7698]_  | ~\new_[12543]_ ;
  assign \new_[7364]_  = ~\new_[11264]_  | ~\wb_addr_i[2] ;
  assign \new_[7365]_  = ~\new_[11720]_ ;
  assign \new_[7366]_  = ~\new_[7633]_ ;
  assign \new_[7367]_  = ~\new_[7593]_ ;
  assign \new_[7368]_  = ~\new_[12667]_  | ~\new_[7700]_  | ~\new_[11362]_ ;
  assign \new_[7369]_  = ~\new_[7597]_ ;
  assign \new_[7370]_  = ~\new_[7599]_ ;
  assign n3501 = \new_[7742]_  | \new_[7713]_ ;
  assign \new_[7372]_  = \new_[11731]_  | \new_[7707]_ ;
  assign \new_[7373]_  = ~\new_[11727]_ ;
  assign \new_[7374]_  = \new_[3179]_  ^ \new_[7837]_ ;
  assign \new_[7375]_  = (~\new_[2074]_  & ~\new_[12622]_ ) | (~\new_[2090]_  & ~\new_[12621]_ );
  assign \new_[7376]_  = (~\new_[2133]_  & ~\new_[12620]_ ) | (~\new_[2111]_  & ~\new_[12621]_ );
  assign \new_[7377]_  = \new_[9010]_  ^ \new_[7854]_ ;
  assign \new_[7378]_  = \new_[9023]_  ^ \new_[7856]_ ;
  assign \new_[7379]_  = \new_[9017]_  ^ \new_[7857]_ ;
  assign \new_[7380]_  = \new_[9015]_  ^ \new_[7858]_ ;
  assign \new_[7381]_  = \\u0_cs_reg[1] ;
  assign \new_[7382]_  = \\u0_u0_csc_reg[0] ;
  assign \new_[7383]_  = ~\new_[7765]_  | ~\new_[8023]_ ;
  assign \new_[7384]_  = ~\new_[8084]_  | ~\new_[8051]_ ;
  assign \new_[7385]_  = ~\new_[12309]_  & ~\new_[10912]_ ;
  assign \new_[7386]_  = ~\new_[12309]_  & ~\new_[10493]_ ;
  assign \new_[7387]_  = ~\new_[8084]_  | ~\new_[11028]_ ;
  assign \new_[7388]_  = ~\new_[8084]_  | ~\new_[11223]_ ;
  assign \new_[7389]_  = ~\new_[7682]_  | ~\new_[9937]_ ;
  assign \new_[7390]_  = u0_u1_lmr_req_reg;
  assign \new_[7391]_  = \new_[8401]_  | \new_[12171]_ ;
  assign \new_[7392]_  = ~\new_[7765]_  | ~\new_[11188]_ ;
  assign \new_[7393]_  = ~\new_[7765]_  | ~\new_[8063]_ ;
  assign \new_[7394]_  = ~\new_[7765]_  | ~\new_[8072]_ ;
  assign \new_[7395]_  = ~\new_[8084]_  | ~\new_[11243]_ ;
  assign \new_[7396]_  = ~\new_[8084]_  | ~\new_[11066]_ ;
  assign \new_[7397]_  = ~\new_[7765]_  | ~\new_[11093]_ ;
  assign \new_[7398]_  = ~\new_[8084]_  | ~\new_[11240]_ ;
  assign \new_[7399]_  = ~\new_[8084]_  | ~\new_[11082]_ ;
  assign \new_[7400]_  = ~\new_[7765]_  | ~\new_[11220]_ ;
  assign \new_[7401]_  = ~\new_[8084]_  | ~\new_[11245]_ ;
  assign \new_[7402]_  = ~\new_[7765]_  | ~\new_[8061]_ ;
  assign \new_[7403]_  = ~\new_[8084]_  | ~\new_[11043]_ ;
  assign \new_[7404]_  = ~\new_[8084]_  | ~\new_[11250]_ ;
  assign \new_[7405]_  = ~\new_[7765]_  | ~\new_[11022]_ ;
  assign \new_[7406]_  = ~\new_[8084]_  | ~\new_[11249]_ ;
  assign \new_[7407]_  = ~\new_[7765]_  | ~\new_[11241]_ ;
  assign \new_[7408]_  = ~\new_[7765]_  | ~\new_[11013]_ ;
  assign \new_[7409]_  = ~\new_[7765]_  | ~\new_[11234]_ ;
  assign \new_[7410]_  = ~\new_[7765]_  | ~\new_[8078]_ ;
  assign \new_[7411]_  = ~\new_[7765]_  | ~\new_[8067]_ ;
  assign \new_[7412]_  = ~\new_[8084]_  | ~\new_[8048]_ ;
  assign \new_[7413]_  = ~\new_[7765]_  | ~\new_[8052]_ ;
  assign \new_[7414]_  = ~\new_[7765]_  | ~\new_[8068]_ ;
  assign \new_[7415]_  = ~\new_[7765]_  | ~\new_[8043]_ ;
  assign \new_[7416]_  = \\u4_rfr_cnt_reg[0] ;
  assign \new_[7417]_  = ~\new_[7663]_ ;
  assign \new_[7418]_  = ~\new_[7631]_ ;
  assign \new_[7419]_  = ~\new_[12234]_ ;
  assign \new_[7420]_  = ~\new_[7689]_  | ~\new_[7747]_ ;
  assign \new_[7421]_  = ~\new_[7592]_ ;
  assign \new_[7422]_  = ~\new_[7675]_ ;
  assign \new_[7423]_  = ~\new_[12673]_  | ~\new_[12089]_ ;
  assign \new_[7424]_  = ~\new_[12673]_  | ~\new_[12567]_ ;
  assign \new_[7425]_  = ~\new_[12673]_  | ~\new_[11363]_ ;
  assign \new_[7426]_  = \new_[12384]_  & \new_[12555]_ ;
  assign \new_[7427]_  = ~\new_[10463]_  | ~\new_[7773]_ ;
  assign \new_[7428]_  = ~\new_[11554]_  & ~\new_[3438]_ ;
  assign \new_[7429]_  = ~\new_[10508]_  | ~\new_[7773]_ ;
  assign \new_[7430]_  = ~\new_[7773]_  | ~\new_[10502]_ ;
  assign \new_[7431]_  = ~\new_[7771]_  | ~\new_[10463]_ ;
  assign \new_[7432]_  = ~\new_[11263]_  & ~\new_[7992]_ ;
  assign \new_[7433]_  = ~\new_[7771]_  | ~\new_[10502]_ ;
  assign n3486 = ~\new_[7676]_  | ~\new_[9986]_ ;
  assign n3496 = ~\new_[12507]_  & (~\new_[7783]_  | ~\new_[7779]_ );
  assign n3491 = ~\new_[12507]_  & (~\new_[7784]_  | ~\new_[7780]_ );
  assign n3476 = ~\new_[12507]_  & (~\new_[7785]_  | ~\new_[7781]_ );
  assign \new_[7438]_  = ~\new_[11263]_  & ~\new_[7861]_ ;
  assign \new_[7439]_  = ~\new_[7771]_  | ~\new_[10508]_ ;
  assign \new_[7440]_  = \new_[8001]_  & \new_[11419]_ ;
  assign n3481 = \new_[7778]_  | \new_[7775]_ ;
  assign \new_[7442]_  = \new_[8742]_  | \new_[12171]_ ;
  assign \new_[7443]_  = \new_[12384]_  & \new_[12554]_ ;
  assign \new_[7444]_  = ~\new_[9634]_  | ~\new_[12384]_ ;
  assign \new_[7445]_  = ~\new_[10291]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7446]_  = ~\new_[9998]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7447]_  = ~\new_[10922]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7448]_  = ~\new_[10164]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7449]_  = ~\new_[10933]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7450]_  = ~\new_[10250]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7451]_  = ~\new_[11363]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7452]_  = ~\new_[10962]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7453]_  = ~\new_[9946]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7454]_  = ~\new_[10411]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7455]_  = ~\new_[11343]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7456]_  = ~n5021 | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7457]_  = ~\new_[10818]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7458]_  = ~\new_[12755]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7459]_  = ~\new_[9785]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7460]_  = ~\new_[10802]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7461]_  = ~\new_[12093]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7462]_  = ~\new_[12567]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7463]_  = ~\new_[11367]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7464]_  = ~\new_[12453]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7465]_  = ~\new_[10496]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7466]_  = ~\new_[11353]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7467]_  = ~\new_[10634]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[7468]_  = ~\new_[10955]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7469]_  = ~\new_[11328]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7470]_  = ~\new_[11313]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7471]_  = ~\new_[11356]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7472]_  = ~\new_[11310]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7473]_  = ~\new_[11361]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7474]_  = ~\new_[10960]_  | ~\new_[11485]_  | ~\new_[12398]_ ;
  assign \new_[7475]_  = ~\new_[12453]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7476]_  = (~\new_[9316]_  | ~\new_[7873]_ ) & (~\new_[12492]_  | ~\new_[10210]_ );
  assign \new_[7477]_  = (~\new_[9315]_  | ~\new_[12492]_ ) & (~\new_[7873]_  | ~\new_[9969]_ );
  assign \new_[7478]_  = (~\new_[4242]_  & ~\new_[9998]_  & ~\new_[10724]_ ) | (~\new_[7782]_  & ~\new_[10747]_  & ~\new_[10902]_ );
  assign \new_[7479]_  = ~\new_[12455]_ ;
  assign \new_[7480]_  = ~\new_[7691]_  & ~\new_[12400]_ ;
  assign \new_[7481]_  = ~\new_[7806]_  & ~\new_[10402]_ ;
  assign \new_[7482]_  = ~\new_[7691]_  & ~\new_[12184]_ ;
  assign \new_[7483]_  = ~\new_[7806]_  & ~\new_[11349]_ ;
  assign \new_[7484]_  = ~\new_[7691]_  & ~\new_[11737]_ ;
  assign \new_[7485]_  = ~\new_[7708]_  & ~\new_[11364]_ ;
  assign \new_[7486]_  = ~\new_[7691]_  & ~\new_[11575]_ ;
  assign \new_[7487]_  = ~\new_[7708]_  & ~\new_[10752]_ ;
  assign \new_[7488]_  = \new_[7692]_  & n5021;
  assign \new_[7489]_  = ~\new_[7691]_  & ~\new_[11341]_ ;
  assign \new_[7490]_  = ~\new_[7806]_  & ~\new_[11493]_ ;
  assign \new_[7491]_  = ~\new_[7691]_  & ~\new_[10673]_ ;
  assign \new_[7492]_  = ~\new_[7708]_  & ~\new_[11321]_ ;
  assign \new_[7493]_  = ~\new_[7708]_  & ~\new_[11012]_ ;
  assign \new_[7494]_  = ~\new_[7708]_  & ~\new_[11881]_ ;
  assign \new_[7495]_  = ~\new_[7708]_  & ~\new_[10872]_ ;
  assign \new_[7496]_  = ~\new_[7806]_  & ~\new_[11299]_ ;
  assign \new_[7497]_  = ~\new_[7708]_  & ~\new_[11317]_ ;
  assign \new_[7498]_  = ~\new_[7708]_  & ~\new_[11329]_ ;
  assign \new_[7499]_  = ~\new_[7806]_  & ~\new_[12555]_ ;
  assign \new_[7500]_  = ~\new_[7708]_  & ~\new_[12611]_ ;
  assign \new_[7501]_  = \new_[7907]_  & \new_[12089]_ ;
  assign \new_[7502]_  = ~\new_[7708]_  & ~\new_[10160]_ ;
  assign \new_[7503]_  = ~\new_[7708]_  & ~\new_[10897]_ ;
  assign \new_[7504]_  = ~\new_[7708]_  & ~\new_[11311]_ ;
  assign \new_[7505]_  = ~\new_[7806]_  & ~\new_[12045]_ ;
  assign \new_[7506]_  = ~\new_[7708]_  & ~\new_[12564]_ ;
  assign \new_[7507]_  = \new_[7692]_  & \new_[10164]_ ;
  assign \new_[7508]_  = ~\new_[7708]_  & ~\new_[10676]_ ;
  assign \new_[7509]_  = ~\new_[7654]_ ;
  assign \new_[7510]_  = ~\new_[7655]_ ;
  assign \new_[7511]_  = ~\new_[7708]_  & ~\new_[10704]_ ;
  assign \new_[7512]_  = ~\new_[7657]_ ;
  assign \new_[7513]_  = ~\new_[7708]_  & ~\new_[11338]_ ;
  assign \new_[7514]_  = ~\new_[7708]_  & ~\new_[12094]_ ;
  assign \new_[7515]_  = ~\new_[7708]_  & ~\new_[11368]_ ;
  assign \new_[7516]_  = ~\new_[7708]_  & ~\new_[10767]_ ;
  assign \new_[7517]_  = ~\new_[7806]_  & ~\new_[10724]_ ;
  assign \new_[7518]_  = ~\new_[7708]_  & ~\new_[12401]_ ;
  assign \new_[7519]_  = ~\new_[7708]_  & ~\new_[10579]_ ;
  assign \new_[7520]_  = \new_[12553]_  & \new_[10551]_ ;
  assign \new_[7521]_  = ~\new_[7629]_ ;
  assign \new_[7522]_  = \new_[7628]_ ;
  assign \new_[7523]_  = ~\new_[7628]_ ;
  assign \new_[7524]_  = ~\new_[7685]_  | ~\new_[12293]_ ;
  assign \new_[7525]_  = ~\new_[7687]_  & ~\new_[11919]_ ;
  assign \new_[7526]_  = ~\new_[7685]_  | ~\new_[9929]_ ;
  assign \new_[7527]_  = ~\new_[7685]_  | ~\new_[9960]_ ;
  assign \new_[7528]_  = \new_[7682]_  & \new_[9975]_ ;
  assign \new_[7529]_  = ~\new_[7682]_  | ~\new_[9824]_ ;
  assign \new_[7530]_  = ~\new_[7995]_  | ~\new_[9489]_ ;
  assign \new_[7531]_  = \new_[7680]_  & \new_[8714]_ ;
  assign \new_[7532]_  = ~\new_[10578]_  & ~\new_[7687]_ ;
  assign \new_[7533]_  = ~\new_[7682]_  | ~\new_[10064]_ ;
  assign \new_[7534]_  = \new_[12791]_  | \new_[10529]_ ;
  assign \new_[7535]_  = ~\new_[7682]_  | ~\new_[9864]_ ;
  assign \new_[7536]_  = \new_[7682]_  & \new_[9613]_ ;
  assign \new_[7537]_  = ~\new_[12537]_  | ~\new_[7681]_ ;
  assign \new_[7538]_  = ~\new_[11577]_ ;
  assign \new_[7539]_  = ~\new_[11502]_ ;
  assign \new_[7540]_  = ~\new_[7615]_ ;
  assign \new_[7541]_  = ~\new_[7693]_  | ~\new_[10086]_ ;
  assign \new_[7542]_  = \new_[7682]_  & \new_[9609]_ ;
  assign \new_[7543]_  = ~\new_[12438]_  & ~\new_[8359]_ ;
  assign \new_[7544]_  = ~\new_[7682]_  | ~\new_[10047]_ ;
  assign \new_[7545]_  = ~\new_[7688]_  | ~\new_[7822]_ ;
  assign \new_[7546]_  = ~\new_[7682]_  | ~\new_[9596]_ ;
  assign \new_[7547]_  = ~\new_[7666]_ ;
  assign \new_[7548]_  = ~\new_[10291]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7549]_  = ~\new_[12492]_  | ~\new_[9591]_ ;
  assign \new_[7550]_  = ~\new_[10827]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7551]_  = ~\new_[11355]_  | ~\new_[12789]_  | ~\new_[10657]_ ;
  assign \new_[7552]_  = ~\new_[11348]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7553]_  = ~\new_[11323]_  | ~\new_[12790]_  | ~\new_[10393]_ ;
  assign \new_[7554]_  = ~\new_[10928]_  | ~\new_[12793]_  | ~\new_[10657]_ ;
  assign \new_[7555]_  = ~\new_[12755]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7556]_  = ~\new_[10496]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7557]_  = ~\new_[11353]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7558]_  = ~\new_[10963]_  | ~\new_[12789]_  | ~\new_[10393]_ ;
  assign \new_[7559]_  = ~\new_[9647]_  | ~\new_[12792]_  | ~\new_[10657]_ ;
  assign \new_[7560]_  = ~\new_[7671]_ ;
  assign \new_[7561]_  = ~\new_[10808]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7562]_  = ~\new_[11340]_  | ~\new_[12790]_  | ~\new_[10314]_ ;
  assign \new_[7563]_  = ~\new_[11492]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7564]_  = ~\new_[7672]_ ;
  assign \new_[7565]_  = ~\new_[10243]_  | ~\new_[12790]_  | ~\new_[10314]_ ;
  assign \new_[7566]_  = ~\new_[11320]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7567]_  = ~\new_[12054]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7568]_  = ~\new_[10526]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7569]_  = ~\new_[10250]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7570]_  = ~\new_[10955]_  | ~\new_[12793]_  | ~\new_[10657]_ ;
  assign \new_[7571]_  = ~\new_[7674]_ ;
  assign \new_[7572]_  = ~\new_[7674]_ ;
  assign \new_[7573]_  = ~\new_[12781]_  | ~\new_[7679]_ ;
  assign \new_[7574]_  = ~\new_[9903]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7575]_  = ~\new_[12554]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7576]_  = ~\new_[10419]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7577]_  = ~\new_[11419]_ ;
  assign \new_[7578]_  = ~\new_[10177]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7579]_  = ~\new_[12610]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7580]_  = ~\new_[10938]_  | ~\new_[12793]_  | ~\new_[10393]_ ;
  assign \new_[7581]_  = ~\new_[11328]_  | ~\new_[12793]_  | ~\new_[10314]_ ;
  assign \new_[7582]_  = ~\new_[11356]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7583]_  = ~\new_[11310]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7584]_  = ~\new_[11313]_  | ~\new_[12790]_  | ~\new_[10657]_ ;
  assign \new_[7585]_  = ~\new_[11526]_  | ~\new_[12789]_  | ~\new_[10657]_ ;
  assign \new_[7586]_  = ~\new_[10922]_  | ~\new_[12792]_  | ~\new_[10314]_ ;
  assign \new_[7587]_  = \new_[7725]_  & \new_[3177]_ ;
  assign \new_[7588]_  = ~\new_[7681]_ ;
  assign \new_[7589]_  = ~\new_[8488]_  & ~\new_[11723]_ ;
  assign \new_[7590]_  = ~\new_[10493]_  & ~\new_[7809]_ ;
  assign \new_[7591]_  = ~\new_[12383]_ ;
  assign \new_[7592]_  = ~\new_[7747]_ ;
  assign \new_[7593]_  = ~\new_[8172]_  & ~\new_[7811]_ ;
  assign \new_[7594]_  = \\u0_u0_csc_reg[4] ;
  assign \new_[7595]_  = \\u0_u0_csc_reg[7] ;
  assign \new_[7596]_  = ~\new_[10715]_  | ~\new_[11921]_  | ~\new_[11319]_  | ~\new_[9405]_ ;
  assign \new_[7597]_  = ~\new_[8028]_  | ~\new_[8810]_  | ~\new_[11835]_  | ~\new_[8188]_ ;
  assign \new_[7598]_  = \\u0_u0_csc_reg[16] ;
  assign \new_[7599]_  = ~\new_[12537]_ ;
  assign \new_[7600]_  = ~\new_[7811]_ ;
  assign \new_[7601]_  = \\u0_u0_csc_reg[18] ;
  assign \new_[7602]_  = \new_[11001]_  ? \new_[12622]_  : \new_[11137]_ ;
  assign \new_[7603]_  = \new_[10985]_  ? \new_[12622]_  : \new_[11027]_ ;
  assign \new_[7604]_  = ~\new_[10877]_  | ~\new_[7837]_  | ~\new_[10941]_ ;
  assign \new_[7605]_  = \new_[11047]_  ? \new_[12622]_  : \new_[11076]_ ;
  assign \new_[7606]_  = \\u0_u0_csc_reg[13] ;
  assign \new_[7607]_  = \\u0_u0_csc_reg[14] ;
  assign \new_[7608]_  = ~\new_[7838]_  & ~\new_[8399]_ ;
  assign n3521 = ~\new_[7821]_  & ~\new_[10124]_ ;
  assign \new_[7610]_  = ~\new_[7852]_  & ~\new_[10151]_ ;
  assign n3506 = ~\new_[7820]_  & ~\new_[10091]_ ;
  assign \new_[7612]_  = \\u0_u0_csc_reg[11] ;
  assign \new_[7613]_  = \\u0_u0_csc_reg[15] ;
  assign \new_[7614]_  = \new_[3169]_  ^ \new_[7989]_ ;
  assign \new_[7615]_  = ~\new_[12308]_  & ~\new_[12492]_ ;
  assign \new_[7616]_  = \\u0_u0_csc_reg[2] ;
  assign \new_[7617]_  = ~u0_u1_init_req_reg;
  assign \new_[7618]_  = \\u0_u0_csc_reg[1] ;
  assign \new_[7619]_  = \\u0_u0_csc_reg[5] ;
  assign \new_[7620]_  = \\u0_u0_csc_reg[17] ;
  assign \new_[7621]_  = \\u0_u0_csc_reg[22] ;
  assign \new_[7622]_  = \\u0_u0_csc_reg[12] ;
  assign \new_[7623]_  = \\u0_u0_csc_reg[8] ;
  assign \new_[7624]_  = \\u0_u0_csc_reg[9] ;
  assign \new_[7625]_  = \\u0_u0_csc_reg[6] ;
  assign \new_[7626]_  = u0_u0_lmr_req_reg;
  assign \new_[7627]_  = ~\new_[8016]_  & (~\new_[12673]_  | ~\new_[10838]_ );
  assign \new_[7628]_  = ~\new_[7772]_ ;
  assign \new_[7629]_  = ~\new_[7744]_ ;
  assign \new_[7630]_  = ~\new_[7744]_ ;
  assign \new_[7631]_  = ~\new_[7744]_ ;
  assign \new_[7632]_  = ~\new_[10203]_  | ~\new_[12398]_  | ~\new_[12672]_  | ~\new_[10481]_ ;
  assign \new_[7633]_  = ~\new_[7690]_ ;
  assign \new_[7634]_  = \new_[12388]_  & \new_[7865]_ ;
  assign \new_[7635]_  = ~\new_[7689]_ ;
  assign \new_[7636]_  = ~\new_[11976]_  | ~\new_[9938]_ ;
  assign \new_[7637]_  = ~\new_[11976]_  | ~\new_[9937]_ ;
  assign n3541 = ~\new_[10124]_  & (~\new_[8035]_  | ~\new_[7931]_ );
  assign \new_[7639]_  = ~\new_[11976]_  | ~\new_[11515]_ ;
  assign \new_[7640]_  = ~\new_[11976]_  | ~\new_[10084]_ ;
  assign \new_[7641]_  = ~\new_[11976]_  | ~\new_[9616]_ ;
  assign \new_[7642]_  = ~\new_[11976]_  | ~\new_[9844]_ ;
  assign n3536 = ~\new_[7819]_  & ~\new_[10091]_ ;
  assign n3511 = ~\new_[7816]_  & ~\new_[10124]_ ;
  assign n3516 = ~\new_[7817]_  & ~\new_[10124]_ ;
  assign n3531 = ~\new_[7818]_  & ~\new_[10091]_ ;
  assign \new_[7647]_  = ~\new_[7806]_  & ~\new_[11889]_ ;
  assign \new_[7648]_  = ~\new_[7806]_  & ~\new_[10747]_ ;
  assign \new_[7649]_  = ~\new_[7805]_  & ~\new_[12274]_ ;
  assign \new_[7650]_  = n3451 & \new_[10922]_ ;
  assign \new_[7651]_  = ~\new_[7805]_  & ~\new_[10551]_ ;
  assign \new_[7652]_  = ~\new_[7806]_  & ~\new_[12599]_ ;
  assign \new_[7653]_  = \new_[7907]_  & \new_[10892]_ ;
  assign \new_[7654]_  = ~\new_[7804]_  | ~\new_[12453]_ ;
  assign \new_[7655]_  = ~n3451 | ~\new_[10743]_ ;
  assign \new_[7656]_  = n3451 & \new_[10496]_ ;
  assign \new_[7657]_  = ~n3451 | ~\new_[10509]_ ;
  assign \new_[7658]_  = n3451 & \new_[10250]_ ;
  assign \new_[7659]_  = n3451 & \new_[12756]_ ;
  assign \new_[7660]_  = ~\new_[7805]_  & ~\new_[11393]_ ;
  assign \new_[7661]_  = ~\new_[7769]_ ;
  assign \new_[7662]_  = ~\new_[7861]_ ;
  assign \new_[7663]_  = ~\new_[7744]_ ;
  assign \new_[7664]_  = ~\new_[7772]_ ;
  assign \new_[7665]_  = \new_[12697]_  | \new_[10369]_ ;
  assign \new_[7666]_  = ~\new_[2606]_  | ~\new_[8030]_  | ~\new_[8413]_ ;
  assign n3526 = ~\new_[8486]_  | ~\new_[7789]_ ;
  assign \new_[7668]_  = ~\new_[12385]_  & ~\new_[8003]_ ;
  assign \new_[7669]_  = ~\new_[9561]_  | ~\new_[10404]_  | ~\new_[7788]_  | ~\new_[8714]_ ;
  assign \new_[7670]_  = ~\new_[11363]_  | ~\new_[12792]_  | ~\new_[10657]_ ;
  assign \new_[7671]_  = ~\new_[10345]_  | ~\new_[9561]_  | ~\new_[12649]_  | ~\new_[8175]_ ;
  assign \new_[7672]_  = ~\new_[10030]_  & ~\new_[12211]_ ;
  assign \new_[7673]_  = ~\new_[12567]_  | ~\new_[12794]_  | ~\new_[10657]_ ;
  assign \new_[7674]_  = ~\new_[8877]_  | ~\new_[10204]_  | ~\new_[12649]_  | ~\new_[8175]_ ;
  assign \new_[7675]_  = ~\new_[7814]_  & (~\new_[10207]_  | ~\new_[10275]_ );
  assign \new_[7676]_  = (~\new_[8148]_  | ~\new_[11794]_ ) & (~\new_[8017]_  | ~\new_[7150]_ );
  assign \new_[7677]_  = ~\new_[2577]_  | ~\new_[7911]_ ;
  assign \new_[7678]_  = ~\new_[12169]_ ;
  assign \new_[7679]_  = ~\new_[10152]_  | ~\new_[9142]_  | ~\new_[12463]_  | ~\new_[12543]_ ;
  assign \new_[7680]_  = \new_[8795]_  & \new_[12091]_ ;
  assign \new_[7681]_  = ~\new_[12456]_ ;
  assign \new_[7682]_  = ~\new_[7863]_ ;
  assign \new_[7683]_  = ~\new_[7786]_ ;
  assign \new_[7684]_  = ~\new_[7786]_ ;
  assign \new_[7685]_  = \new_[12308]_ ;
  assign \new_[7686]_  = ~\new_[7911]_  & ~\new_[8014]_ ;
  assign \new_[7687]_  = \new_[9565]_  | \new_[12213]_ ;
  assign \new_[7688]_  = ~\new_[7913]_  | ~\new_[11835]_ ;
  assign \new_[7689]_  = ~\new_[9559]_  | ~\new_[10579]_  | ~\new_[12156]_  | ~\new_[10892]_ ;
  assign \new_[7690]_  = \new_[8172]_  & \new_[7986]_ ;
  assign \new_[7691]_  = ~\new_[7804]_ ;
  assign \new_[7692]_  = ~\new_[7805]_ ;
  assign \new_[7693]_  = ~\new_[7814]_ ;
  assign \new_[7694]_  = \\u0_u1_csc_reg[16] ;
  assign \new_[7695]_  = ~\new_[10029]_  | ~\new_[9318]_  | ~\new_[8169]_  | ~\new_[8025]_ ;
  assign \new_[7696]_  = ~\new_[8173]_  | ~\new_[8186]_  | ~\new_[8026]_  | ~\new_[8187]_ ;
  assign \new_[7697]_  = \\u0_u0_csc_reg[21] ;
  assign \new_[7698]_  = ~\new_[11723]_ ;
  assign \new_[7699]_  = ~\new_[7920]_  | ~\new_[10811]_ ;
  assign \new_[7700]_  = ~\new_[7809]_ ;
  assign \new_[7701]_  = \new_[7707]_  & \new_[11732]_ ;
  assign \new_[7702]_  = \\u0_u1_csc_reg[17] ;
  assign \new_[7703]_  = \\u0_u1_csc_reg[19] ;
  assign \new_[7704]_  = \\u0_u0_csc_reg[19] ;
  assign \new_[7705]_  = ~\new_[8202]_  | ~\new_[10946]_  | ~\new_[10454]_  | ~\new_[10762]_ ;
  assign \new_[7706]_  = \\u0_u0_csc_reg[20] ;
  assign \new_[7707]_  = ~\new_[11728]_ ;
  assign \new_[7708]_  = ~n3451;
  assign \new_[7709]_  = ~\\u0_u1_csc_reg[13] ;
  assign \new_[7710]_  = ~\\u0_u1_csc_reg[15] ;
  assign \new_[7711]_  = ~\new_[10708]_  | ~\new_[8399]_  | ~\new_[7957]_  | ~\new_[10929]_ ;
  assign \new_[7712]_  = ~\new_[7976]_  & ~\new_[10975]_ ;
  assign \new_[7713]_  = ~\new_[11404]_  & (~\new_[8398]_  | ~\new_[8731]_ );
  assign \new_[7714]_  = ~\new_[11718]_ ;
  assign \new_[7715]_  = \\u0_u0_csc_reg[10] ;
  assign \new_[7716]_  = \\u0_u1_csc_reg[10] ;
  assign \new_[7717]_  = ~\new_[7827]_ ;
  assign \new_[7718]_  = ~\\u0_u1_csc_reg[12] ;
  assign n3561 = ~\new_[7930]_  & ~\new_[10091]_ ;
  assign \new_[7720]_  = \\u0_u0_csc_reg[27] ;
  assign \new_[7721]_  = ~\new_[8399]_  | ~\new_[7978]_  | ~\new_[10793]_ ;
  assign \new_[7722]_  = \\u0_u1_csc_reg[5] ;
  assign \new_[7723]_  = \\u0_u1_csc_reg[7] ;
  assign \new_[7724]_  = \\u0_u1_csc_reg[9] ;
  assign \new_[7725]_  = \new_[7989]_  & \new_[3169]_ ;
  assign n3546 = \new_[7381]_  ? n5766 : \new_[8085]_ ;
  assign \new_[7727]_  = \new_[7991]_  & \new_[8085]_ ;
  assign \new_[7728]_  = ~\new_[7990]_  | ~\new_[3036]_ ;
  assign \new_[7729]_  = \\u0_u0_csc_reg[28] ;
  assign \new_[7730]_  = \\u0_u1_csc_reg[21] ;
  assign \new_[7731]_  = \new_[7990]_  | \new_[10485]_ ;
  assign \new_[7732]_  = \\u0_u0_csc_reg[3] ;
  assign \new_[7733]_  = \\u0_u1_csc_reg[4] ;
  assign \new_[7734]_  = \\u0_u0_csc_reg[23] ;
  assign \new_[7735]_  = \\u0_u0_csc_reg[25] ;
  assign \new_[7736]_  = ~\\u0_u1_csc_reg[14] ;
  assign \new_[7737]_  = \\u0_u1_csc_reg[20] ;
  assign \new_[7738]_  = \\u0_u1_csc_reg[22] ;
  assign \new_[7739]_  = ~\\u0_u1_csc_reg[26] ;
  assign \new_[7740]_  = ~\\u0_u1_csc_reg[27] ;
  assign \new_[7741]_  = \\u0_u0_csc_reg[30] ;
  assign \new_[7742]_  = ~\new_[8395]_  & ~\new_[11403]_ ;
  assign \new_[7743]_  = \\u0_u0_csc_reg[31] ;
  assign \new_[7744]_  = ~\new_[7992]_ ;
  assign \new_[7745]_  = \\u0_u0_csc_reg[29] ;
  assign \new_[7746]_  = ~\\u0_u1_csc_reg[30] ;
  assign \new_[7747]_  = ~\new_[7787]_ ;
  assign \new_[7748]_  = ~\\u0_u1_csc_reg[24] ;
  assign \new_[7749]_  = \\u0_u0_csc_reg[26] ;
  assign \new_[7750]_  = ~\new_[7786]_ ;
  assign \new_[7751]_  = ~\\u0_u1_csc_reg[31] ;
  assign \new_[7752]_  = ~\new_[12673]_  | ~\new_[10922]_ ;
  assign \new_[7753]_  = ~\new_[12673]_  | ~\new_[12755]_ ;
  assign \new_[7754]_  = ~\new_[12673]_  | ~n5021;
  assign \new_[7755]_  = ~\new_[12673]_  | ~\new_[10164]_ ;
  assign \new_[7756]_  = ~\new_[12673]_  | ~\new_[12453]_ ;
  assign \new_[7757]_  = ~\new_[12673]_  | ~\new_[10496]_ ;
  assign \new_[7758]_  = ~\new_[12673]_  | ~\new_[10250]_ ;
  assign \new_[7759]_  = \new_[1645]_  | \new_[7992]_ ;
  assign \new_[7760]_  = ~\new_[7994]_  | ~\new_[10960]_ ;
  assign \new_[7761]_  = \\u0_u0_csc_reg[24] ;
  assign n3551 = ~\new_[10120]_  | ~\new_[10012]_  | ~\new_[8038]_ ;
  assign \new_[7763]_  = ~\new_[7807]_ ;
  assign n3556 = ~\new_[7997]_  | ~\new_[7996]_ ;
  assign \new_[7765]_  = ~\new_[7991]_ ;
  assign \new_[7766]_  = ~\new_[7921]_  & ~\new_[10698]_ ;
  assign \new_[7767]_  = ~\new_[7921]_  & ~\new_[10920]_ ;
  assign \new_[7768]_  = ~\new_[7921]_  & ~\new_[10348]_ ;
  assign \new_[7769]_  = ~\new_[7921]_  & ~\new_[11314]_ ;
  assign \new_[7770]_  = ~\new_[7885]_  & ~\new_[9297]_ ;
  assign \new_[7771]_  = ~\new_[11404]_  & ~\new_[8015]_ ;
  assign \new_[7772]_  = ~\new_[7992]_ ;
  assign \new_[7773]_  = ~\new_[11403]_  & ~\new_[8015]_ ;
  assign \new_[7774]_  = ~\new_[12478]_ ;
  assign \new_[7775]_  = ~\new_[11403]_  & (~\new_[9248]_  | ~\new_[10198]_ );
  assign \new_[7776]_  = ~\new_[7824]_ ;
  assign \new_[7777]_  = ~\new_[7824]_ ;
  assign \new_[7778]_  = ~\new_[11404]_  & (~\new_[10026]_  | ~\new_[10138]_ );
  assign \new_[7779]_  = ~\new_[8148]_  | ~\new_[7150]_ ;
  assign \new_[7780]_  = ~\new_[8148]_  | ~\new_[7152]_ ;
  assign \new_[7781]_  = ~\new_[8148]_  | ~\new_[7151]_ ;
  assign \new_[7782]_  = ~\new_[11456]_  | ~\new_[8014]_ ;
  assign \new_[7783]_  = ~\new_[8017]_  | ~\new_[7152]_ ;
  assign \new_[7784]_  = ~\new_[8017]_  | ~\new_[7151]_ ;
  assign \new_[7785]_  = ~\new_[8017]_  | ~\new_[11794]_ ;
  assign \new_[7786]_  = ~\new_[12308]_ ;
  assign \new_[7787]_  = ~\new_[12464]_  & ~\new_[8698]_ ;
  assign \new_[7788]_  = ~\new_[12440]_  & ~\new_[9376]_ ;
  assign \new_[7789]_  = ~\new_[10370]_  | ~\new_[7382]_  | ~\new_[8024]_  | ~\new_[8177]_ ;
  assign n3596 = ~\new_[10299]_  & (~\new_[8155]_  | ~\new_[8304]_ );
  assign n3636 = ~\new_[10299]_  & (~\new_[8156]_  | ~\new_[8388]_ );
  assign n3586 = ~\new_[10299]_  & (~\new_[8157]_  | ~\new_[8306]_ );
  assign n3591 = ~\new_[10299]_  & (~\new_[8158]_  | ~\new_[8307]_ );
  assign n3576 = ~\new_[10299]_  & (~\new_[8160]_  | ~\new_[8309]_ );
  assign n3626 = ~\new_[10299]_  & (~\new_[8161]_  | ~\new_[8308]_ );
  assign n3631 = ~\new_[10299]_  & (~\new_[8288]_  | ~\new_[8167]_ );
  assign n3601 = ~\new_[10299]_  & (~\new_[8159]_  | ~\new_[8220]_ );
  assign \new_[7798]_  = \\u1_u0_out_r_reg[11] ;
  assign n3571 = ~\new_[10299]_  & (~\new_[8300]_  | ~\new_[8166]_ );
  assign n3641 = ~\new_[10299]_  & (~\new_[8163]_  | ~\new_[8348]_ );
  assign n3581 = ~\new_[10299]_  & (~\new_[8286]_  | ~\new_[8165]_ );
  assign n3651 = ~\new_[10299]_  & (~\new_[8164]_  | ~\new_[8346]_ );
  assign n3646 = ~\new_[10299]_  & (~\new_[8162]_  | ~\new_[8338]_ );
  assign \new_[7804]_  = ~\new_[7921]_ ;
  assign \new_[7805]_  = \new_[7921]_ ;
  assign \new_[7806]_  = ~\new_[7907]_ ;
  assign \new_[7807]_  = ~\new_[7909]_ ;
  assign \new_[7808]_  = ~\new_[8029]_  | ~\new_[10811]_ ;
  assign \new_[7809]_  = ~\new_[12091]_ ;
  assign \new_[7810]_  = ~\new_[8027]_  | ~\new_[10811]_ ;
  assign \new_[7811]_  = ~\new_[7986]_ ;
  assign \new_[7812]_  = \\u0_u1_csc_reg[18] ;
  assign \new_[7813]_  = \\u0_u1_csc_reg[1] ;
  assign \new_[7814]_  = ~\new_[10240]_  | ~\new_[11572]_  | ~\new_[8020]_  | ~\new_[9957]_ ;
  assign n3451 = ~\new_[7921]_ ;
  assign \new_[7816]_  = ~\new_[8040]_  & (~\new_[7275]_  | ~\new_[8369]_ );
  assign \new_[7817]_  = ~\new_[8041]_  & (~\new_[7278]_  | ~\new_[8369]_ );
  assign \new_[7818]_  = ~\new_[8042]_  & (~\new_[8369]_  | ~\new_[7281]_ );
  assign \new_[7819]_  = ~\new_[8036]_  & (~\new_[7284]_  | ~\new_[8369]_ );
  assign \new_[7820]_  = ~\new_[8037]_  & (~\new_[7265]_  | ~\new_[8369]_ );
  assign \new_[7821]_  = ~\new_[8039]_  & (~\new_[7279]_  | ~\new_[8369]_ );
  assign \new_[7822]_  = ~\new_[8172]_  | ~\new_[11835]_  | ~\new_[8188]_ ;
  assign \new_[7823]_  = \new_[7994]_ ;
  assign \new_[7824]_  = ~\new_[7994]_ ;
  assign \new_[7825]_  = \new_[7994]_ ;
  assign \new_[7826]_  = ~\new_[12491]_ ;
  assign \new_[7827]_  = \new_[11201]_  ? \new_[12623]_  : \new_[11099]_ ;
  assign \new_[7828]_  = \\u0_u1_csc_reg[2] ;
  assign n3566 = \new_[8152]_  ? \new_[10299]_  : \poc_o[0] ;
  assign \new_[7830]_  = ~\new_[7285]_  | ~\new_[11256]_  | ~\new_[10762]_  | ~\new_[8202]_ ;
  assign \wb_data_o[10]  = \\u6_wb_data_o_reg[10] ;
  assign \wb_data_o[2]  = \\u6_wb_data_o_reg[2] ;
  assign \new_[7833]_  = \\u0_u1_csc_reg[8] ;
  assign \wb_data_o[7]  = \\u6_wb_data_o_reg[7] ;
  assign \wb_data_o[3]  = \\u6_wb_data_o_reg[3] ;
  assign \wb_data_o[0]  = \\u6_wb_data_o_reg[0] ;
  assign \new_[7837]_  = ~\new_[10498]_  & ~\new_[8031]_ ;
  assign \new_[7838]_  = ~\new_[7957]_ ;
  assign \new_[7839]_  = ~\\u0_u1_csc_reg[25] ;
  assign \wb_data_o[11]  = \\u6_wb_data_o_reg[11] ;
  assign \wb_data_o[14]  = \\u6_wb_data_o_reg[14] ;
  assign \wb_data_o[1]  = \\u6_wb_data_o_reg[1] ;
  assign \wb_data_o[5]  = \\u6_wb_data_o_reg[5] ;
  assign \wb_data_o[9]  = \\u6_wb_data_o_reg[9] ;
  assign \wb_data_o[6]  = \\u6_wb_data_o_reg[6] ;
  assign \wb_data_o[4]  = \\u6_wb_data_o_reg[4] ;
  assign \wb_data_o[12]  = \\u6_wb_data_o_reg[12] ;
  assign \wb_data_o[15]  = \\u6_wb_data_o_reg[15] ;
  assign \wb_data_o[8]  = \\u6_wb_data_o_reg[8] ;
  assign \new_[7850]_  = \\u0_u1_csc_reg[0] ;
  assign \new_[7851]_  = \\u0_u1_csc_reg[3] ;
  assign \new_[7852]_  = (~\new_[8216]_  | ~\new_[7833]_ ) & (~\new_[8217]_  | ~\new_[7623]_ );
  assign \wb_data_o[13]  = \\u6_wb_data_o_reg[13] ;
  assign \new_[7854]_  = \new_[8105]_  ^ \new_[8104]_ ;
  assign \new_[7855]_  = ~\new_[8046]_  | ~\new_[10811]_ ;
  assign \new_[7856]_  = \new_[8111]_  ^ \new_[8106]_ ;
  assign \new_[7857]_  = \new_[8110]_  ^ \new_[8107]_ ;
  assign \new_[7858]_  = \new_[8108]_  ^ \new_[8109]_ ;
  assign \new_[7859]_  = ~\new_[12173]_ ;
  assign n3656 = ~\new_[8112]_  | ~\new_[8102]_ ;
  assign \new_[7861]_  = ~\new_[8030]_  | ~\new_[11779]_ ;
  assign \new_[7862]_  = \new_[8016]_  | \new_[8748]_ ;
  assign \new_[7863]_  = ~\new_[7995]_ ;
  assign \new_[7864]_  = ~\new_[12383]_  | ~\new_[8003]_ ;
  assign \new_[7865]_  = \new_[8013]_  & \new_[8005]_ ;
  assign \new_[7866]_  = ~\new_[8030]_  | ~\new_[11062]_ ;
  assign n3611 = ~\new_[8000]_  | (~\new_[7617]_  & ~\new_[8772]_ );
  assign n3616 = ~\new_[10120]_  | (~\new_[8151]_  & ~\new_[10299]_ );
  assign n3606 = ~\new_[10012]_  | (~\new_[8153]_  & ~\new_[10299]_ );
  assign n3621 = \new_[8154]_  ? \new_[10299]_  : \poc_o[1] ;
  assign \new_[7871]_  = ~\new_[11987]_ ;
  assign \new_[7872]_  = \new_[8362]_  ^ \new_[3180]_ ;
  assign \new_[7873]_  = ~\new_[12170]_ ;
  assign \new_[7874]_  = ~\new_[8003]_ ;
  assign \new_[7875]_  = ~\new_[8004]_ ;
  assign n3686 = ~\new_[10299]_  & (~\new_[8299]_  | ~\new_[8317]_ );
  assign n3666 = ~\new_[10299]_  & (~\new_[8295]_  | ~\new_[8312]_ );
  assign n3826 = ~\new_[10299]_  & (~\new_[8298]_  | ~\new_[8336]_ );
  assign n3816 = ~\new_[10299]_  & (~\new_[8303]_  | ~\new_[8313]_ );
  assign n3716 = ~\new_[10299]_  & (~\new_[8297]_  | ~\new_[8318]_ );
  assign n3736 = ~\new_[10299]_  & (~\new_[8291]_  | ~\new_[8314]_ );
  assign n3791 = ~\new_[10299]_  & (~\new_[8293]_  | ~\new_[8315]_ );
  assign n3746 = ~\new_[10299]_  & (~\new_[8294]_  | ~\new_[8340]_ );
  assign n3761 = ~\new_[10299]_  & (~\new_[8290]_  | ~\new_[8345]_ );
  assign \new_[7885]_  = ~\new_[9991]_  | ~\new_[10211]_  | ~\new_[10157]_  | ~\new_[8347]_ ;
  assign \new_[7886]_  = ~\new_[8189]_  & ~\new_[11833]_ ;
  assign n3706 = ~\new_[10282]_  & (~\new_[8440]_  | ~\new_[8321]_ );
  assign n3711 = ~\new_[10282]_  & (~\new_[8591]_  | ~\new_[8322]_ );
  assign n3696 = ~\new_[10282]_  & (~\new_[8442]_  | ~\new_[8325]_ );
  assign n3676 = ~\new_[10282]_  & (~\new_[8628]_  | ~\new_[8328]_ );
  assign n3801 = ~\new_[10299]_  & (~\new_[8292]_  | ~\new_[8305]_ );
  assign n3776 = ~\new_[10282]_  & (~\new_[8447]_  | ~\new_[8342]_ );
  assign n3741 = ~\new_[10282]_  & (~\new_[8626]_  | ~\new_[8344]_ );
  assign n3811 = ~\new_[10282]_  & (~\new_[8448]_  | ~\new_[8329]_ );
  assign n3781 = ~\new_[10282]_  & (~\new_[8452]_  | ~\new_[8330]_ );
  assign n3786 = ~\new_[10282]_  & (~\new_[8592]_  | ~\new_[8331]_ );
  assign n3806 = ~\new_[10282]_  & (~\new_[8597]_  | ~\new_[8332]_ );
  assign n3821 = ~\new_[10282]_  & (~\new_[8594]_  | ~\new_[8333]_ );
  assign n3751 = ~\new_[10282]_  & (~\new_[8595]_  | ~\new_[8320]_ );
  assign n3721 = ~\new_[10282]_  & (~\new_[8596]_  | ~\new_[8319]_ );
  assign n3726 = ~\new_[10282]_  & (~\new_[8450]_  | ~\new_[8341]_ );
  assign n3756 = ~\new_[10299]_  & (~\new_[8289]_  | ~\new_[8337]_ );
  assign n3701 = ~\new_[10299]_  & (~\new_[8301]_  | ~\new_[8339]_ );
  assign n3661 = ~\new_[10282]_  & (~\new_[8630]_  | ~\new_[8326]_ );
  assign n3796 = ~\new_[10299]_  & (~\new_[8302]_  | ~\new_[8316]_ );
  assign n3681 = ~\new_[10299]_  & (~\new_[8287]_  | ~\new_[8310]_ );
  assign \new_[7907]_  = ~\new_[8030]_ ;
  assign \new_[7908]_  = ~u5_wb_write_go_r_reg;
  assign \new_[7909]_  = ~\new_[8014]_ ;
  assign \new_[7910]_  = ~\new_[8170]_  | ~\new_[10811]_ ;
  assign \new_[7911]_  = ~\new_[11456]_ ;
  assign \new_[7912]_  = ~\new_[8171]_  | ~\new_[10811]_ ;
  assign \new_[7913]_  = \new_[8188]_  & \new_[8353]_ ;
  assign \new_[7914]_  = ~\\u0_u1_tms_reg[30] ;
  assign \new_[7915]_  = ~\new_[10872]_  | ~\new_[10920]_  | ~\new_[10658]_  | ~\new_[8356]_ ;
  assign \wb_data_o[31]  = \\u6_wb_data_o_reg[31] ;
  assign \new_[7917]_  = ~\\u0_u1_tms_reg[13] ;
  assign \new_[7918]_  = ~\new_[11256]_  | ~\new_[8202]_  | ~\new_[10929]_ ;
  assign \new_[7919]_  = \\u0_u1_tms_reg[27] ;
  assign \new_[7920]_  = ~\new_[8026]_ ;
  assign \new_[7921]_  = \new_[8030]_ ;
  assign \new_[7922]_  = ~\\u0_u1_tms_reg[15] ;
  assign \wb_data_o[24]  = \\u6_wb_data_o_reg[24] ;
  assign \new_[7924]_  = ~\new_[8175]_  | ~\new_[8795]_ ;
  assign \new_[7925]_  = ~\new_[9681]_  | ~\new_[8175]_  | ~\new_[10276]_ ;
  assign \new_[7926]_  = \\u0_u1_tms_reg[8] ;
  assign \new_[7927]_  = \\u0_u1_tms_reg[7] ;
  assign \wb_data_o[26]  = \\u6_wb_data_o_reg[26] ;
  assign \new_[7929]_  = ~\\u0_u1_csc_reg[29] ;
  assign \new_[7930]_  = \new_[7416]_  ^ \new_[8369]_ ;
  assign \new_[7931]_  = ~\new_[10537]_  | ~\new_[8191]_ ;
  assign \new_[7932]_  = ~\\u0_u1_tms_reg[28] ;
  assign \new_[7933]_  = ~\\u0_u1_csc_reg[11] ;
  assign \new_[7934]_  = \\u0_u1_tms_reg[0] ;
  assign \new_[7935]_  = ~\\u0_u1_tms_reg[29] ;
  assign \new_[7936]_  = ~\\u0_u1_tms_reg[16] ;
  assign \new_[7937]_  = \\u0_u1_tms_reg[3] ;
  assign \new_[7938]_  = \\u0_u1_tms_reg[10] ;
  assign \new_[7939]_  = ~\\u0_u1_tms_reg[23] ;
  assign n3731 = ~\new_[10282]_  & (~\new_[8522]_  | ~\new_[8334]_ );
  assign \new_[7941]_  = ~\\u0_u1_tms_reg[17] ;
  assign \new_[7942]_  = \\u0_u1_tms_reg[24] ;
  assign \new_[7943]_  = ~\\u0_u1_tms_reg[12] ;
  assign \new_[7944]_  = \\u0_u1_tms_reg[25] ;
  assign \new_[7945]_  = \\u0_u1_tms_reg[5] ;
  assign \wb_data_o[17]  = \\u6_wb_data_o_reg[17] ;
  assign n3771 = ~\new_[10282]_  & (~\new_[8446]_  | ~\new_[8343]_ );
  assign n3671 = ~\new_[10282]_  & (~\new_[8443]_  | ~\new_[8327]_ );
  assign \wb_data_o[18]  = \\u6_wb_data_o_reg[18] ;
  assign \new_[7950]_  = ~\\u0_u1_tms_reg[18] ;
  assign \new_[7951]_  = \\u0_u1_csc_reg[6] ;
  assign \wb_data_o[20]  = \\u6_wb_data_o_reg[20] ;
  assign \wb_data_o[23]  = \\u6_wb_data_o_reg[23] ;
  assign n3691 = ~\new_[10282]_  & (~\new_[8454]_  | ~\new_[8323]_ );
  assign n3766 = ~\new_[10282]_  & (~\new_[8441]_  | ~\new_[8324]_ );
  assign \new_[7956]_  = ~\new_[8190]_  & ~\new_[11833]_ ;
  assign \new_[7957]_  = \new_[8202]_  & \new_[10930]_ ;
  assign \wb_data_o[19]  = \\u6_wb_data_o_reg[19] ;
  assign \wb_data_o[29]  = \\u6_wb_data_o_reg[29] ;
  assign \new_[7960]_  = \\u0_u1_csc_reg[23] ;
  assign \wb_data_o[21]  = \\u6_wb_data_o_reg[21] ;
  assign \wb_data_o[25]  = \\u6_wb_data_o_reg[25] ;
  assign \wb_data_o[16]  = \\u6_wb_data_o_reg[16] ;
  assign \wb_data_o[27]  = \\u6_wb_data_o_reg[27] ;
  assign \wb_data_o[30]  = \\u6_wb_data_o_reg[30] ;
  assign \new_[7966]_  = \\u4_ps_cnt_reg[7] ;
  assign \wb_data_o[28]  = \\u6_wb_data_o_reg[28] ;
  assign \new_[7968]_  = ~\\u0_u1_tms_reg[11] ;
  assign \new_[7969]_  = ~\\u0_u1_tms_reg[14] ;
  assign \new_[7970]_  = ~\\u0_u1_tms_reg[20] ;
  assign \new_[7971]_  = \\u0_u1_tms_reg[26] ;
  assign \new_[7972]_  = \\u0_u1_tms_reg[2] ;
  assign \new_[7973]_  = ~\\u0_u1_tms_reg[31] ;
  assign \new_[7974]_  = \\u0_u1_tms_reg[4] ;
  assign \new_[7975]_  = \\u0_u1_tms_reg[6] ;
  assign \new_[7976]_  = ~\new_[7265]_  | ~\new_[7281]_  | ~\new_[8204]_  | ~\new_[7416]_ ;
  assign \new_[7977]_  = \\u4_ps_cnt_reg[4] ;
  assign \new_[7978]_  = ~\new_[8203]_  & ~\new_[10353]_ ;
  assign \new_[7979]_  = ~\\u0_u1_csc_reg[28] ;
  assign \wb_data_o[22]  = \\u6_wb_data_o_reg[22] ;
  assign \new_[7981]_  = ~\\u0_u1_tms_reg[19] ;
  assign \new_[7982]_  = \\u0_u1_tms_reg[9] ;
  assign \new_[7983]_  = \\u0_u1_tms_reg[1] ;
  assign \new_[7984]_  = ~\\u0_u1_tms_reg[22] ;
  assign \new_[7985]_  = ~\\u0_u1_tms_reg[21] ;
  assign \new_[7986]_  = ~\new_[11835]_  & ~\new_[11947]_ ;
  assign \new_[7987]_  = \new_[8489]_  | \new_[9043]_  | \new_[8259]_  | \new_[8791]_ ;
  assign \new_[7988]_  = ~\new_[8015]_ ;
  assign \new_[7989]_  = ~\new_[8031]_ ;
  assign \new_[7990]_  = ~\new_[12577]_  & (~\new_[12282]_  | ~\new_[10679]_ );
  assign \new_[7991]_  = ~\new_[8084]_ ;
  assign \new_[7992]_  = ~\new_[8143]_  | ~\new_[11778]_ ;
  assign \new_[7993]_  = ~\new_[8094]_ ;
  assign \new_[7994]_  = ~\new_[8143]_  | ~\new_[8813]_ ;
  assign \new_[7995]_  = ~\new_[7999]_ ;
  assign \new_[7996]_  = ~\new_[7390]_  | ~\new_[9803]_  | ~\new_[8263]_ ;
  assign \new_[7997]_  = \new_[8168]_  | \new_[8263]_ ;
  assign \new_[7998]_  = \new_[8850]_  | \new_[12633]_ ;
  assign \new_[7999]_  = \new_[12633]_  | \new_[8697]_ ;
  assign \new_[8000]_  = ~\new_[10523]_  | ~\new_[7850]_  | ~\new_[8285]_  | ~\new_[8168]_ ;
  assign \new_[8001]_  = \new_[8857]_  | \new_[12633]_ ;
  assign \new_[8002]_  = \new_[9028]_  | \new_[12633]_ ;
  assign \new_[8003]_  = \new_[12633]_  | \new_[8853]_ ;
  assign \new_[8004]_  = ~\new_[12090]_  | ~\new_[8456]_  | ~\new_[12392]_ ;
  assign \new_[8005]_  = \new_[12633]_  | \new_[8854]_ ;
  assign n3936 = ~\new_[10282]_  & (~\new_[8455]_  | ~\new_[8640]_ );
  assign n3836 = ~\new_[10282]_  & (~\new_[8444]_  | ~\new_[8642]_ );
  assign n3841 = ~\new_[10282]_  & (~\new_[8445]_  | ~\new_[8668]_ );
  assign n3881 = ~\new_[10282]_  & (~\new_[8453]_  | ~\new_[8644]_ );
  assign n3846 = ~\new_[10282]_  & (~\new_[8449]_  | ~\new_[8645]_ );
  assign n3941 = ~\new_[10282]_  & (~\new_[8439]_  | ~\new_[8639]_ );
  assign n3861 = ~\new_[10282]_  & (~\new_[8451]_  | ~\new_[8647]_ );
  assign \new_[8013]_  = ~\new_[10113]_  | ~\new_[9262]_  | ~\new_[8358]_  | ~\new_[11753]_ ;
  assign \new_[8014]_  = ~\new_[11510]_  & ~\new_[8862]_ ;
  assign \new_[8015]_  = ~\new_[11510]_  | ~\new_[10959]_ ;
  assign \new_[8016]_  = ~\new_[11510]_  & ~\new_[2055]_ ;
  assign \new_[8017]_  = ~\new_[8148]_ ;
  assign \new_[8018]_  = ~\new_[10481]_  | ~\new_[8311]_ ;
  assign \new_[8019]_  = ~\new_[8150]_ ;
  assign \new_[8020]_  = ~\new_[8349]_  & ~\new_[8773]_ ;
  assign \new_[8021]_  = ~\new_[9648]_  & (~\new_[8485]_  | ~\new_[9566]_ );
  assign \new_[8022]_  = ~\new_[8368]_  & ~\new_[12469]_ ;
  assign \new_[8023]_  = \\u0_u0_tms_reg[8] ;
  assign \new_[8024]_  = u0_u0_init_req_we_reg;
  assign \new_[8025]_  = ~\new_[8791]_  & ~\new_[8360]_ ;
  assign \new_[8026]_  = (~\new_[10324]_  | ~\new_[12763]_ ) & (~\new_[10289]_  | ~\new_[11309]_ );
  assign \new_[8027]_  = ~\new_[8187]_ ;
  assign \new_[8028]_  = ~\new_[8172]_ ;
  assign \new_[8029]_  = ~\new_[8173]_ ;
  assign \new_[8030]_  = \new_[8143]_ ;
  assign \new_[8031]_  = ~\new_[8362]_  | ~\new_[3180]_ ;
  assign \new_[8032]_  = ~\\u0_u0_tms_reg[14] ;
  assign n3831 = ~\new_[8367]_  | (~\new_[8723]_  & ~\new_[11235]_ );
  assign \new_[8034]_  = ~\\u0_u0_tms_reg[12] ;
  assign \new_[8035]_  = ~\new_[7285]_  | ~\new_[8369]_ ;
  assign \new_[8036]_  = ~\new_[9747]_  & ~\new_[8369]_ ;
  assign \new_[8037]_  = ~\new_[8978]_  & ~\new_[8369]_ ;
  assign \new_[8038]_  = \new_[8284]_  | \new_[10299]_ ;
  assign \new_[8039]_  = ~\new_[9145]_  & ~\new_[8369]_ ;
  assign \new_[8040]_  = ~\new_[9417]_  & ~\new_[8369]_ ;
  assign \new_[8041]_  = ~\new_[9186]_  & ~\new_[8369]_ ;
  assign \new_[8042]_  = ~\new_[8972]_  & ~\new_[8369]_ ;
  assign \new_[8043]_  = \\u0_u0_tms_reg[9] ;
  assign \new_[8044]_  = ~\new_[8393]_  & ~\new_[12469]_ ;
  assign \new_[8045]_  = ~\\u0_u0_tms_reg[31] ;
  assign \new_[8046]_  = ~\new_[8186]_ ;
  assign \new_[8047]_  = ~\\u0_u0_tms_reg[11] ;
  assign \new_[8048]_  = \\u0_u0_tms_reg[4] ;
  assign \new_[8049]_  = \\u4_ps_cnt_reg[3] ;
  assign \new_[8050]_  = ~\new_[9726]_  | ~\new_[11256]_  | ~\new_[10915]_  | ~\new_[8492]_ ;
  assign \new_[8051]_  = \\u0_u0_tms_reg[6] ;
  assign \new_[8052]_  = \\u0_u0_tms_reg[5] ;
  assign \new_[8053]_  = ~\\u0_u0_tms_reg[30] ;
  assign \new_[8054]_  = ~\\u0_u0_tms_reg[23] ;
  assign \new_[8055]_  = ~\\u0_u0_tms_reg[24] ;
  assign \new_[8056]_  = ~\\u0_u0_tms_reg[17] ;
  assign \new_[8057]_  = ~\\u0_u0_tms_reg[18] ;
  assign \new_[8058]_  = ~\\u0_u0_tms_reg[20] ;
  assign \new_[8059]_  = ~\\u0_u0_tms_reg[19] ;
  assign \new_[8060]_  = ~\\u0_u0_tms_reg[13] ;
  assign \new_[8061]_  = \\u0_u0_tms_reg[1] ;
  assign n3931 = \new_[8540]_  ? \new_[10300]_  : \new_[8427]_ ;
  assign \new_[8063]_  = \\u0_u0_tms_reg[0] ;
  assign \new_[8064]_  = ~\\u0_u0_tms_reg[15] ;
  assign \new_[8065]_  = ~\\u0_u0_tms_reg[21] ;
  assign \new_[8066]_  = ~\\u0_u0_tms_reg[29] ;
  assign \new_[8067]_  = \\u0_u0_tms_reg[3] ;
  assign \new_[8068]_  = \\u0_u0_tms_reg[7] ;
  assign n3856 = \new_[8539]_  ? \new_[10300]_  : \new_[8433]_ ;
  assign \new_[8070]_  = ~\new_[8403]_  | ~\new_[10320]_ ;
  assign \new_[8071]_  = \\u4_ps_cnt_reg[0] ;
  assign \new_[8072]_  = \\u0_u0_tms_reg[10] ;
  assign \new_[8073]_  = ~\\u0_u0_tms_reg[16] ;
  assign \new_[8074]_  = ~\\u0_u0_tms_reg[25] ;
  assign \new_[8075]_  = \\u4_ps_cnt_reg[6] ;
  assign \new_[8076]_  = ~\\u0_u0_tms_reg[26] ;
  assign \new_[8077]_  = \\u4_ps_cnt_reg[1] ;
  assign \new_[8078]_  = \\u0_u0_tms_reg[2] ;
  assign \new_[8079]_  = \\u4_ps_cnt_reg[2] ;
  assign \new_[8080]_  = ~\\u0_u0_tms_reg[27] ;
  assign \new_[8081]_  = \\u4_ps_cnt_reg[5] ;
  assign \new_[8082]_  = ~\\u0_u0_tms_reg[28] ;
  assign \new_[8083]_  = ~\\u0_u0_tms_reg[22] ;
  assign \new_[8084]_  = ~\new_[8406]_  & (~\new_[7623]_  | ~wb_we_i);
  assign \new_[8085]_  = ~\new_[8405]_  & (~\new_[7833]_  | ~wb_we_i);
  assign n3896 = \new_[8751]_  ? \new_[10300]_  : \new_[8424]_ ;
  assign n3871 = \new_[8757]_  ? \new_[10300]_  : \new_[8428]_ ;
  assign n3901 = \new_[8750]_  ? \new_[10300]_  : \new_[8436]_ ;
  assign n3906 = \new_[8747]_  ? \new_[10300]_  : \new_[8434]_ ;
  assign n3911 = \new_[8755]_  ? \new_[10300]_  : \new_[8432]_ ;
  assign n3916 = \new_[8756]_  ? \new_[10300]_  : \new_[8435]_ ;
  assign \new_[8092]_  = ~\new_[8404]_  & (~\new_[8821]_  | ~\new_[2056]_ );
  assign \new_[8093]_  = (~\new_[9745]_  | ~\new_[8407]_ ) & (~\new_[8821]_  | ~\new_[2070]_ );
  assign \new_[8094]_  = ~\new_[3036]_  | ~\new_[11776]_  | ~\new_[8413]_ ;
  assign n3886 = \new_[8956]_  ? \new_[10300]_  : \new_[8425]_ ;
  assign n3921 = \new_[8838]_  ? \new_[10300]_  : \new_[8438]_ ;
  assign n3891 = \new_[8958]_  ? \new_[10300]_  : \new_[8429]_ ;
  assign n3926 = \new_[8833]_  ? \new_[10300]_  : \new_[8426]_ ;
  assign n3946 = \new_[8832]_  ? \new_[10300]_  : \new_[8431]_ ;
  assign n3876 = \new_[8538]_  ? \new_[10300]_  : \new_[8437]_ ;
  assign n3851 = \new_[8542]_  ? \new_[10300]_  : \new_[8423]_ ;
  assign \new_[8102]_  = ~\new_[7626]_  | ~\new_[9915]_  | ~\new_[8415]_ ;
  assign n3866 = \new_[8541]_  ? \new_[10300]_  : \new_[8430]_ ;
  assign \new_[8104]_  = \new_[8575]_  ^ \new_[8574]_ ;
  assign \new_[8105]_  = \new_[8576]_  ^ \new_[8588]_ ;
  assign \new_[8106]_  = \new_[8578]_  ^ \new_[8577]_ ;
  assign \new_[8107]_  = \new_[8581]_  ^ \new_[8711]_ ;
  assign \new_[8108]_  = \new_[8583]_  ^ \new_[8587]_ ;
  assign \new_[8109]_  = \new_[8582]_  ^ \new_[8585]_ ;
  assign \new_[8110]_  = \new_[8584]_  ^ \new_[8580]_ ;
  assign \new_[8111]_  = \new_[8579]_  ^ \new_[8586]_ ;
  assign \new_[8112]_  = \new_[8177]_  | \new_[8415]_ ;
  assign n4206 = ~\new_[10282]_  & (~\new_[8605]_  | ~\new_[8670]_ );
  assign n4041 = ~\new_[10282]_  & (~\new_[8609]_  | ~\new_[8732]_ );
  assign n4046 = ~\new_[10282]_  & (~\new_[8603]_  | ~\new_[8650]_ );
  assign n4141 = ~\new_[8479]_  & ~n4566;
  assign n4026 = ~\new_[10282]_  & (~\new_[8702]_  | ~\new_[8633]_ );
  assign n4221 = ~\new_[10282]_  & (~\new_[8608]_  | ~\new_[8653]_ );
  assign n4111 = ~\new_[10282]_  & (~\new_[8624]_  | ~\new_[8643]_ );
  assign n4001 = ~\new_[10282]_  & (~\new_[8593]_  | ~\new_[8651]_ );
  assign n4016 = ~\new_[10282]_  & (~\new_[8521]_  | ~\new_[8648]_ );
  assign n3956 = ~\new_[10282]_  & (~\new_[8614]_  | ~\new_[8636]_ );
  assign n4151 = ~\new_[10282]_  & (~\new_[8600]_  | ~\new_[8735]_ );
  assign n4056 = ~\new_[10282]_  & (~\new_[8601]_  | ~\new_[8649]_ );
  assign n3966 = ~\new_[10282]_  & (~\new_[8623]_  | ~\new_[8654]_ );
  assign n4081 = ~\new_[10282]_  & (~\new_[8604]_  | ~\new_[8635]_ );
  assign n4161 = ~\new_[10282]_  & (~\new_[8606]_  | ~\new_[8652]_ );
  assign n4226 = ~\new_[10282]_  & (~\new_[8607]_  | ~\new_[8665]_ );
  assign n4051 = ~\new_[10282]_  & (~\new_[8610]_  | ~\new_[8655]_ );
  assign n4061 = ~\new_[10282]_  & (~\new_[8627]_  | ~\new_[8667]_ );
  assign n4171 = ~\new_[10282]_  & (~\new_[8613]_  | ~\new_[8672]_ );
  assign n4176 = ~\new_[10282]_  & (~\new_[8615]_  | ~\new_[8657]_ );
  assign n4031 = ~\new_[10282]_  & (~\new_[8616]_  | ~\new_[8669]_ );
  assign n4066 = ~\new_[10282]_  & (~\new_[8618]_  | ~\new_[8659]_ );
  assign n3986 = ~\new_[10282]_  & (~\new_[8621]_  | ~\new_[8673]_ );
  assign n4211 = ~\new_[10282]_  & (~\new_[8622]_  | ~\new_[8662]_ );
  assign n4216 = ~\new_[10282]_  & (~\new_[8625]_  | ~\new_[8675]_ );
  assign n4186 = ~\new_[10282]_  & (~\new_[8619]_  | ~\new_[8660]_ );
  assign n4021 = ~\new_[10282]_  & (~\new_[8612]_  | ~\new_[8664]_ );
  assign n4006 = ~\new_[10282]_  & (~\new_[8629]_  | ~\new_[8656]_ );
  assign n4166 = ~\new_[10282]_  & (~\new_[8611]_  | ~\new_[8676]_ );
  assign n3991 = ~\new_[10282]_  & (~\new_[8620]_  | ~\new_[8661]_ );
  assign \new_[8143]_  = ~\new_[12282]_ ;
  assign \new_[8144]_  = ~\new_[8957]_  & ~\new_[9902]_ ;
  assign \new_[8145]_  = ~n3951 | ~\new_[11323]_ ;
  assign \new_[8146]_  = ~\new_[8957]_  & ~\new_[11299]_ ;
  assign \new_[8147]_  = ~\new_[8957]_  & ~\new_[12045]_ ;
  assign \new_[8148]_  = ~\new_[1646]_  & ~\new_[8957]_ ;
  assign \new_[8149]_  = \\u0_csc_mask_r_reg[0] ;
  assign \new_[8150]_  = ~\new_[12585]_  | ~\new_[9706]_  | ~\new_[11753]_  | ~\new_[8714]_ ;
  assign \new_[8151]_  = (~n4236 | ~\wb_data_i[1] ) & (~\new_[8856]_  | ~\new_[7618]_ );
  assign \new_[8152]_  = \wb_data_i[4]  ? \new_[8856]_  : \new_[7594]_ ;
  assign \new_[8153]_  = (~n4236 | ~\wb_data_i[2] ) & (~\new_[8856]_  | ~\new_[7616]_ );
  assign \new_[8154]_  = \wb_data_i[5]  ? \new_[8856]_  : \new_[7619]_ ;
  assign \new_[8155]_  = ~\new_[8856]_  | ~\new_[7612]_ ;
  assign \new_[8156]_  = ~\new_[8856]_  | ~\new_[7622]_ ;
  assign \new_[8157]_  = ~\new_[8856]_  | ~\new_[7606]_ ;
  assign \new_[8158]_  = ~\new_[8856]_  | ~\new_[7607]_ ;
  assign \new_[8159]_  = ~\new_[8856]_  | ~\new_[7613]_ ;
  assign \new_[8160]_  = ~\new_[8856]_  | ~\new_[7598]_ ;
  assign \new_[8161]_  = ~\new_[8856]_  | ~\new_[7620]_ ;
  assign \new_[8162]_  = ~\new_[8856]_  | ~\new_[7624]_ ;
  assign \new_[8163]_  = ~\new_[8856]_  | ~\new_[7623]_ ;
  assign \new_[8164]_  = ~\new_[8856]_  | ~\new_[7625]_ ;
  assign \new_[8165]_  = ~n4236 | ~\wb_data_i[18] ;
  assign \new_[8166]_  = ~n4236 | ~\wb_data_i[7] ;
  assign \new_[8167]_  = ~n4236 | ~\wb_data_i[22] ;
  assign \new_[8168]_  = ~u0_u1_inited_reg;
  assign \new_[8169]_  = ~\new_[8475]_  & ~\new_[8970]_ ;
  assign \new_[8170]_  = \new_[10330]_  ? \new_[12764]_  : \new_[10351]_ ;
  assign \new_[8171]_  = \new_[10347]_  ? \new_[12764]_  : \new_[10368]_ ;
  assign \new_[8172]_  = ~\new_[8353]_ ;
  assign \new_[8173]_  = (~\new_[12625]_  | ~\new_[10279]_ ) & (~\new_[10333]_  | ~\new_[12764]_ );
  assign \new_[8174]_  = ~\new_[9681]_  | ~\new_[8714]_  | ~\new_[10452]_ ;
  assign \new_[8175]_  = \new_[8714]_ ;
  assign n4181 = ~\new_[10282]_  & (~\new_[8617]_  | ~\new_[8663]_ );
  assign \new_[8177]_  = ~u0_u0_inited_reg;
  assign n3971 = ~\new_[10282]_  & (~\new_[8631]_  | ~\new_[8674]_ );
  assign \new_[8179]_  = \\u0_csc_mask_r_reg[1] ;
  assign n4196 = ~\new_[10282]_  & (~\new_[8744]_  | ~\new_[8658]_ );
  assign n3976 = ~\new_[10282]_  & (~\new_[8590]_  | ~\new_[8638]_ );
  assign n4156 = ~\new_[10282]_  & (~\new_[8602]_  | ~\new_[8666]_ );
  assign n4036 = ~\new_[10282]_  & (~\new_[8599]_  | ~\new_[8741]_ );
  assign n4086 = ~\new_[10282]_  & (~\new_[8598]_  | ~\new_[8646]_ );
  assign \new_[8185]_  = u0_sreq_cs_le_reg;
  assign \new_[8186]_  = (~\new_[10360]_  | ~\new_[12624]_ ) & (~\new_[10277]_  | ~\new_[12626]_ );
  assign \new_[8187]_  = (~\new_[10311]_  | ~\new_[12763]_ ) & (~\new_[10327]_  | ~\new_[12626]_ );
  assign \new_[8188]_  = ~\new_[11947]_ ;
  assign \new_[8189]_  = ~\new_[8482]_  & (~\new_[8821]_  | ~\new_[2137]_ );
  assign \new_[8190]_  = ~\new_[8493]_  & (~\new_[8821]_  | ~\new_[2138]_ );
  assign \new_[8191]_  = ~\new_[8369]_ ;
  assign \new_[8192]_  = \new_[8487]_  & \new_[10160]_ ;
  assign n4011 = ~\new_[10282]_  & (~\new_[8632]_  | ~\new_[8641]_ );
  assign \new_[8194]_  = \\u0_csc_mask_r_reg[9] ;
  assign \new_[8195]_  = \\u0_csc_mask_r_reg[10] ;
  assign \new_[8196]_  = \\u0_csc_mask_r_reg[2] ;
  assign \new_[8197]_  = ~u5_cmd_asserted2_reg;
  assign \new_[8198]_  = \\u0_csc_mask_r_reg[4] ;
  assign \new_[8199]_  = \\u0_csc_mask_r_reg[5] ;
  assign \new_[8200]_  = \\u0_csc_mask_r_reg[6] ;
  assign \new_[8201]_  = \\u0_csc_mask_r_reg[7] ;
  assign \new_[8202]_  = \new_[8492]_  & \new_[7416]_ ;
  assign \new_[8203]_  = ~\new_[10946]_  | ~\new_[8492]_  | ~\new_[10930]_ ;
  assign \new_[8204]_  = \new_[8492]_  & \new_[10930]_ ;
  assign \new_[8205]_  = \\u0_csc_mask_r_reg[8] ;
  assign n3996 = \new_[8758]_  ? \new_[10300]_  : \new_[8527]_ ;
  assign n4131 = \new_[8753]_  ? \new_[10300]_  : \new_[8526]_ ;
  assign n4146 = \new_[8745]_  ? \new_[10300]_  : \new_[8528]_ ;
  assign n4106 = \new_[8759]_  ? \new_[10300]_  : \new_[8525]_ ;
  assign n3961 = \new_[8746]_  ? \new_[10300]_  : \new_[8730]_ ;
  assign n4191 = ~\new_[8476]_  & ~n4566;
  assign n4136 = \new_[8752]_  ? \new_[10300]_  : \new_[8728]_ ;
  assign n3981 = \new_[8754]_  ? \new_[10300]_  : \new_[8530]_ ;
  assign n4121 = \new_[8760]_  ? \new_[10300]_  : \new_[8537]_ ;
  assign \new_[8215]_  = ~\new_[8408]_  & ~\new_[10747]_ ;
  assign \new_[8216]_  = ~\new_[8405]_ ;
  assign \new_[8217]_  = ~\new_[8406]_ ;
  assign \new_[8218]_  = ~\new_[8408]_  & ~\new_[11364]_ ;
  assign \new_[8219]_  = ~\new_[12283]_  & ~\new_[1643]_ ;
  assign \new_[8220]_  = ~n4236 | ~\wb_data_i[15] ;
  assign n4126 = \new_[8959]_  ? \new_[10300]_  : \new_[8531]_ ;
  assign n4071 = \new_[8837]_  ? \new_[10300]_  : \new_[8534]_ ;
  assign n4076 = \new_[8828]_  ? \new_[10300]_  : \new_[8532]_ ;
  assign n4101 = \new_[8835]_  ? \new_[10300]_  : \new_[8533]_ ;
  assign n4091 = \new_[8834]_  ? \new_[10300]_  : \new_[8529]_ ;
  assign n4201 = \new_[8955]_  ? \new_[10300]_  : \new_[8536]_ ;
  assign n4096 = \new_[8836]_  ? \new_[10300]_  : \new_[8535]_ ;
  assign n4116 = \new_[8829]_  ? \new_[10300]_  : \new_[8726]_ ;
  assign \new_[8229]_  = \\u0_csc_mask_r_reg[3] ;
  assign \new_[8230]_  = u5_no_wb_cycle_reg;
  assign \new_[8231]_  = ~n4501 | ~\new_[11735]_ ;
  assign \new_[8232]_  = \\u0_csr_r2_reg[6] ;
  assign n4331 = \new_[8543]_  | \new_[10299]_ ;
  assign n4246 = \new_[8546]_  | \new_[10299]_ ;
  assign n4241 = \new_[8548]_  | \new_[10299]_ ;
  assign n4321 = \new_[8547]_  | \new_[10299]_ ;
  assign n4336 = \new_[8549]_  | \new_[10299]_ ;
  assign n4371 = \new_[8550]_  | \new_[10299]_ ;
  assign n4301 = \new_[8551]_  | \new_[10299]_ ;
  assign n4306 = \new_[8552]_  | \new_[10299]_ ;
  assign n4316 = \new_[8553]_  | \new_[10299]_ ;
  assign n4341 = \new_[8572]_  | \new_[10299]_ ;
  assign n4421 = \new_[8555]_  | \new_[10299]_ ;
  assign n4291 = \new_[8556]_  | \new_[10299]_ ;
  assign n4296 = \new_[8557]_  | \new_[10299]_ ;
  assign n4376 = \new_[8558]_  | \new_[10299]_ ;
  assign n4406 = \new_[8559]_  | \new_[10299]_ ;
  assign n4416 = \new_[8560]_  | \new_[10299]_ ;
  assign n4396 = \new_[8562]_  | \new_[10299]_ ;
  assign n4351 = \new_[8565]_  | \new_[10299]_ ;
  assign n4266 = \new_[8566]_  | \new_[10299]_ ;
  assign n4281 = \new_[8567]_  | \new_[10299]_ ;
  assign n4276 = \new_[8568]_  | \new_[10299]_ ;
  assign n4231 = \new_[8571]_  | \new_[10299]_ ;
  assign n4251 = \new_[8570]_  | \new_[10299]_ ;
  assign n4311 = \new_[8554]_  | \new_[10299]_ ;
  assign n4256 = \new_[8564]_  | \new_[10299]_ ;
  assign \new_[8258]_  = ~\new_[1643]_  & (~n4626 | ~\new_[10851]_ );
  assign \new_[8259]_  = ~\new_[12274]_  | ~\new_[11889]_  | ~\new_[9406]_  | ~\new_[8776]_ ;
  assign \new_[8260]_  = \\u0_csr_r2_reg[4] ;
  assign \new_[8261]_  = \\u1_u0_out_r_reg[9] ;
  assign \new_[8262]_  = ~\new_[8840]_  & ~\new_[12597]_ ;
  assign \new_[8263]_  = ~\new_[10523]_  | ~\new_[8589]_ ;
  assign \new_[8264]_  = ~\new_[8957]_  & ~\new_[10722]_ ;
  assign \new_[8265]_  = ~\new_[8957]_  & ~\new_[11575]_ ;
  assign \new_[8266]_  = ~\new_[8957]_  & ~\new_[11334]_ ;
  assign \new_[8267]_  = ~\new_[8957]_  & ~\new_[10752]_ ;
  assign \new_[8268]_  = ~\new_[8957]_  & ~\new_[10920]_ ;
  assign \new_[8269]_  = ~\new_[8957]_  & ~\new_[11341]_ ;
  assign \new_[8270]_  = ~\new_[8957]_  & ~\new_[10673]_ ;
  assign \new_[8271]_  = ~\new_[8957]_  & ~\new_[11321]_ ;
  assign \new_[8272]_  = ~\new_[8957]_  & ~\new_[10872]_ ;
  assign \new_[8273]_  = ~\new_[8957]_  & ~\new_[11317]_ ;
  assign \new_[8274]_  = \new_[12398]_  & \new_[12089]_ ;
  assign \new_[8275]_  = ~\new_[8840]_  & ~\new_[10783]_ ;
  assign \new_[8276]_  = ~\new_[8957]_  & ~\new_[11012]_ ;
  assign \new_[8277]_  = ~\new_[8957]_  & ~\new_[11324]_ ;
  assign \new_[8278]_  = ~\new_[8840]_  & ~\new_[10715]_ ;
  assign \new_[8279]_  = ~\new_[8957]_  & ~\new_[10724]_ ;
  assign \new_[8280]_  = ~\new_[8957]_  & ~\new_[10704]_ ;
  assign \new_[8281]_  = ~\new_[8957]_  & ~\new_[10771]_ ;
  assign \new_[8282]_  = ~\new_[8957]_  & ~\new_[10698]_ ;
  assign \new_[8283]_  = ~\new_[8957]_  & ~\new_[11529]_ ;
  assign \new_[8284]_  = (~n4236 | ~\wb_data_i[0] ) & (~\new_[8856]_  | ~\new_[7382]_ );
  assign \new_[8285]_  = u0_u1_init_req_we_reg;
  assign \new_[8286]_  = ~\new_[8856]_  | ~\new_[7601]_ ;
  assign \new_[8287]_  = ~\new_[8856]_  | ~\new_[7704]_ ;
  assign \new_[8288]_  = ~\new_[8856]_  | ~\new_[7621]_ ;
  assign \new_[8289]_  = ~\new_[8856]_  | ~\new_[7734]_ ;
  assign \new_[8290]_  = ~\new_[8856]_  | ~\new_[7735]_ ;
  assign \new_[8291]_  = ~\new_[8856]_  | ~\new_[7729]_ ;
  assign \new_[8292]_  = ~\new_[8856]_  | ~\new_[7745]_ ;
  assign \new_[8293]_  = ~\new_[8856]_  | ~\new_[7741]_ ;
  assign \new_[8294]_  = ~\new_[8856]_  | ~\new_[7732]_ ;
  assign \new_[8295]_  = ~\new_[8856]_  | ~\new_[7697]_ ;
  assign \new_[8296]_  = \\u0_csr_r2_reg[0] ;
  assign \new_[8297]_  = ~\new_[8856]_  | ~\new_[7720]_ ;
  assign \new_[8298]_  = ~\new_[8856]_  | ~\new_[7761]_ ;
  assign \new_[8299]_  = ~\new_[8856]_  | ~\new_[7706]_ ;
  assign \new_[8300]_  = ~\new_[8856]_  | ~\new_[7595]_ ;
  assign \new_[8301]_  = ~\new_[8856]_  | ~\new_[7715]_ ;
  assign \new_[8302]_  = ~\new_[8856]_  | ~\new_[7743]_ ;
  assign \new_[8303]_  = ~\new_[8856]_  | ~\new_[7749]_ ;
  assign \new_[8304]_  = ~n4236 | ~\wb_data_i[11] ;
  assign \new_[8305]_  = ~n4236 | ~\wb_data_i[29] ;
  assign \new_[8306]_  = ~n4236 | ~\wb_data_i[13] ;
  assign \new_[8307]_  = ~n4236 | ~\wb_data_i[14] ;
  assign \new_[8308]_  = ~n4236 | ~\wb_data_i[17] ;
  assign \new_[8309]_  = ~n4236 | ~\wb_data_i[16] ;
  assign \new_[8310]_  = ~n4236 | ~\wb_data_i[19] ;
  assign \new_[8311]_  = ~n3951;
  assign \new_[8312]_  = ~n4236 | ~\wb_data_i[21] ;
  assign \new_[8313]_  = ~n4236 | ~\wb_data_i[26] ;
  assign \new_[8314]_  = ~n4236 | ~\wb_data_i[28] ;
  assign \new_[8315]_  = ~n4236 | ~\wb_data_i[30] ;
  assign \new_[8316]_  = ~n4236 | ~\wb_data_i[31] ;
  assign \new_[8317]_  = ~n4236 | ~\wb_data_i[20] ;
  assign \new_[8318]_  = ~n4236 | ~\wb_data_i[27] ;
  assign \new_[8319]_  = ~n4521 | ~\wb_data_i[5] ;
  assign \new_[8320]_  = ~n4521 | ~\wb_data_i[4] ;
  assign \new_[8321]_  = ~n4521 | ~\wb_data_i[10] ;
  assign \new_[8322]_  = ~n4521 | ~\wb_data_i[12] ;
  assign \new_[8323]_  = ~n4521 | ~\wb_data_i[13] ;
  assign \new_[8324]_  = ~n4521 | ~\wb_data_i[14] ;
  assign \new_[8325]_  = ~n4521 | ~\wb_data_i[15] ;
  assign \new_[8326]_  = ~n4521 | ~\wb_data_i[16] ;
  assign \new_[8327]_  = ~n4521 | ~\wb_data_i[17] ;
  assign \new_[8328]_  = ~n4521 | ~\wb_data_i[19] ;
  assign \new_[8329]_  = ~n4521 | ~\wb_data_i[24] ;
  assign \new_[8330]_  = ~n4521 | ~\wb_data_i[26] ;
  assign \new_[8331]_  = ~n4521 | ~\wb_data_i[27] ;
  assign \new_[8332]_  = ~n4521 | ~\wb_data_i[30] ;
  assign \new_[8333]_  = ~n4521 | ~\wb_data_i[31] ;
  assign \new_[8334]_  = ~n4521 | ~\wb_data_i[9] ;
  assign \new_[8335]_  = ~\new_[8456]_ ;
  assign \new_[8336]_  = ~n4236 | ~\wb_data_i[24] ;
  assign \new_[8337]_  = ~n4236 | ~\wb_data_i[23] ;
  assign \new_[8338]_  = ~n4236 | ~\wb_data_i[9] ;
  assign \new_[8339]_  = ~n4236 | ~\wb_data_i[10] ;
  assign \new_[8340]_  = ~n4236 | ~\wb_data_i[3] ;
  assign \new_[8341]_  = ~n4521 | ~\wb_data_i[7] ;
  assign \new_[8342]_  = ~n4521 | ~\wb_data_i[22] ;
  assign \new_[8343]_  = ~n4521 | ~\wb_data_i[20] ;
  assign \new_[8344]_  = ~n4521 | ~\wb_data_i[21] ;
  assign \new_[8345]_  = ~n4236 | ~\wb_data_i[25] ;
  assign \new_[8346]_  = ~n4236 | ~\wb_data_i[6] ;
  assign \new_[8347]_  = ~\new_[8701]_  & ~\new_[12319]_ ;
  assign \new_[8348]_  = ~n4236 | ~\wb_data_i[8] ;
  assign \new_[8349]_  = ~\new_[11573]_  | ~\new_[11317]_  | ~\new_[8694]_  | ~\new_[10469]_ ;
  assign \new_[8350]_  = ~\\u0_csr_r_reg[7] ;
  assign \new_[8351]_  = (~\new_[6866]_  | ~\new_[11308]_ ) & (~\new_[9569]_  | ~\new_[12764]_ );
  assign \new_[8352]_  = \\u0_csr_r2_reg[1] ;
  assign \new_[8353]_  = (~\new_[2494]_  | ~\new_[11308]_ ) & (~\new_[2369]_  | ~\new_[12617]_ );
  assign \new_[8354]_  = \new_[7381]_  ? \new_[12626]_  : \new_[9136]_ ;
  assign \new_[8355]_  = \\u0_csr_r2_reg[2] ;
  assign \new_[8356]_  = ~\new_[8703]_  & ~n5001;
  assign \new_[8357]_  = ~\new_[9658]_  | ~\new_[10553]_  | ~\new_[10549]_ ;
  assign \new_[8358]_  = \new_[10253]_  & \new_[8714]_ ;
  assign \new_[8359]_  = ~\new_[10928]_  | ~\new_[12667]_  | ~\new_[8714]_  | ~\new_[11354]_ ;
  assign \new_[8360]_  = ~\new_[10802]_  | ~\new_[10771]_  | ~\new_[8706]_  | ~\new_[10157]_ ;
  assign \new_[8361]_  = ~\new_[8720]_  & ~\new_[9997]_ ;
  assign \new_[8362]_  = \\u1_u0_out_r_reg[12] ;
  assign n4271 = ~\new_[8724]_  & ~n4566;
  assign \new_[8364]_  = ~\\u0_csr_r_reg[6] ;
  assign \new_[8365]_  = \\u0_csr_r_reg[9] ;
  assign \new_[8366]_  = \\u1_u0_out_r_reg[7] ;
  assign \new_[8367]_  = ~\new_[8723]_  | ~\new_[11235]_ ;
  assign \new_[8368]_  = (~\new_[8818]_  | ~\new_[8820]_ ) & (~\new_[9170]_  | ~\new_[1843]_ );
  assign \new_[8369]_  = ~u4_rfr_ce_reg;
  assign n4401 = ~\new_[8762]_  & ~n4566;
  assign n4411 = ~\new_[8764]_  & ~n4566;
  assign n4381 = ~\new_[8743]_  & ~n4566;
  assign n4361 = ~\new_[8845]_  & ~n4566;
  assign n4346 = \new_[8561]_  | \new_[10299]_ ;
  assign n4356 = \new_[8569]_  | \new_[10299]_ ;
  assign n4286 = \new_[8563]_  | \new_[10299]_ ;
  assign n4386 = \new_[8573]_  | \new_[10299]_ ;
  assign \new_[8378]_  = \\u0_csr_r2_reg[3] ;
  assign mc_vpen_pad_o = \\u0_csr_r_reg[1] ;
  assign \new_[8380]_  = ~\\u0_csr_r_reg[3] ;
  assign n4326 = \new_[8737]_  | \new_[10299]_ ;
  assign \new_[8382]_  = \\u0_csr_r_reg[8] ;
  assign n4261 = \new_[8545]_  | \new_[10299]_ ;
  assign n4366 = \new_[8544]_  | \new_[10299]_ ;
  assign \new_[8385]_  = \new_[8733]_  | \new_[12469]_ ;
  assign n4391 = ~n4566 & (~\new_[9161]_  | ~\new_[8851]_ );
  assign \new_[8387]_  = \\u0_csr_r_reg[2] ;
  assign \new_[8388]_  = ~n4236 | ~\wb_data_i[12] ;
  assign \new_[8389]_  = ~\\u0_csr_r_reg[4] ;
  assign \new_[8390]_  = \\u0_csr_r2_reg[7] ;
  assign \new_[8391]_  = \new_[1796]_  ? \new_[8820]_  : \new_[9409]_ ;
  assign \new_[8392]_  = \new_[1955]_  ? \new_[8820]_  : \new_[8765]_ ;
  assign \new_[8393]_  = (~\new_[8761]_  | ~\new_[8820]_ ) & (~\new_[9170]_  | ~\new_[1842]_ );
  assign \new_[8394]_  = \new_[8740]_  | \new_[8840]_ ;
  assign \new_[8395]_  = ~\new_[8495]_  & ~\new_[8497]_ ;
  assign \new_[8396]_  = ~\\u0_csr_r_reg[5] ;
  assign \new_[8397]_  = ~\new_[8957]_  & ~\new_[11349]_ ;
  assign \new_[8398]_  = ~\new_[8496]_  & (~\new_[8763]_  | ~\new_[10435]_ );
  assign \new_[8399]_  = \\u0_csr_r_reg[10] ;
  assign \new_[8400]_  = \\u0_csr_r2_reg[5] ;
  assign \new_[8401]_  = ~\new_[8740]_  & (~\new_[8749]_  | ~\new_[11337]_ );
  assign \new_[8402]_  = ~\new_[8738]_  & (~\new_[8821]_  | ~\new_[1454]_ );
  assign \new_[8403]_  = ~\new_[8739]_  & (~\new_[8821]_  | ~\new_[1519]_ );
  assign \new_[8404]_  = ~\new_[9204]_  & ~\new_[8821]_ ;
  assign \new_[8405]_  = ~\new_[8844]_  | ~\new_[8990]_  | ~\new_[9749]_  | ~\new_[9733]_ ;
  assign \new_[8406]_  = ~\new_[8843]_  | ~\new_[8841]_  | ~\new_[9382]_  | ~\new_[9788]_ ;
  assign \new_[8407]_  = ~\new_[8821]_ ;
  assign \new_[8408]_  = ~\new_[8748]_ ;
  assign \new_[8409]_  = \\u1_u0_out_r_reg[4] ;
  assign \new_[8410]_  = u6_wb_first_r_reg;
  assign n4431 = \new_[8772]_  | \new_[11221]_ ;
  assign n4436 = ~\new_[8786]_  | ~\new_[8177]_ ;
  assign \new_[8413]_  = ~\new_[1645]_  & ~\new_[11779]_ ;
  assign \new_[8414]_  = ~\new_[8840]_  & ~\new_[12274]_ ;
  assign \new_[8415]_  = ~\new_[10370]_  | ~\new_[8804]_ ;
  assign \new_[8416]_  = ~\new_[8840]_  & ~\new_[12184]_ ;
  assign \new_[8417]_  = ~\new_[8840]_  & ~\new_[10754]_ ;
  assign \new_[8418]_  = ~\new_[8840]_  & ~\new_[9889]_ ;
  assign \new_[8419]_  = ~\new_[8840]_  & ~\new_[10160]_ ;
  assign \new_[8420]_  = ~\new_[8840]_  & ~\new_[12555]_ ;
  assign \new_[8421]_  = ~\new_[8840]_  & ~\new_[11881]_ ;
  assign n4446 = ~\new_[8947]_  | ~\new_[10163]_  | ~\new_[10863]_ ;
  assign \new_[8423]_  = ~\new_[8779]_  | (~\new_[9795]_  & ~\new_[10201]_ );
  assign \new_[8424]_  = ~\new_[8769]_  | (~\new_[9793]_  & ~\new_[10201]_ );
  assign \new_[8425]_  = ~\new_[8784]_  | (~\new_[9801]_  & ~\new_[10201]_ );
  assign \new_[8426]_  = ~\new_[8768]_  | (~\new_[9723]_  & ~\new_[10201]_ );
  assign \new_[8427]_  = ~\new_[8777]_  | (~\new_[9792]_  & ~\new_[10201]_ );
  assign \new_[8428]_  = ~\new_[8781]_  | (~\new_[9966]_  & ~\new_[10201]_ );
  assign \new_[8429]_  = ~\new_[8770]_  | (~\new_[9735]_  & ~\new_[10201]_ );
  assign \new_[8430]_  = ~\new_[8778]_  | (~\new_[9798]_  & ~\new_[10201]_ );
  assign \new_[8431]_  = ~\new_[8771]_  | (~\new_[9796]_  & ~\new_[10201]_ );
  assign \new_[8432]_  = ~\new_[8775]_  | (~\new_[9799]_  & ~\new_[10201]_ );
  assign \new_[8433]_  = ~\new_[8780]_  | (~\new_[9797]_  & ~\new_[10201]_ );
  assign \new_[8434]_  = ~\new_[8785]_  | (~\new_[9873]_  & ~\new_[10201]_ );
  assign \new_[8435]_  = ~\new_[8774]_  | (~\new_[9794]_  & ~\new_[10201]_ );
  assign \new_[8436]_  = ~\new_[8782]_  | (~\new_[9741]_  & ~\new_[10201]_ );
  assign \new_[8437]_  = ~\new_[8783]_  | (~\new_[9800]_  & ~\new_[10201]_ );
  assign \new_[8438]_  = ~\new_[8767]_  | (~\new_[9935]_  & ~\new_[10201]_ );
  assign \new_[8439]_  = ~\new_[9026]_  | ~\new_[7851]_ ;
  assign \new_[8440]_  = ~\new_[9026]_  | ~\new_[7716]_ ;
  assign \new_[8441]_  = ~\new_[9026]_  | ~\new_[11156]_ ;
  assign \new_[8442]_  = ~\new_[9026]_  | ~\new_[11175]_ ;
  assign \new_[8443]_  = ~\new_[9026]_  | ~\new_[7702]_ ;
  assign \new_[8444]_  = ~\new_[9026]_  | ~\new_[7812]_ ;
  assign \new_[8445]_  = ~\new_[9026]_  | ~\new_[7813]_ ;
  assign \new_[8446]_  = ~\new_[9026]_  | ~\new_[7737]_ ;
  assign \new_[8447]_  = ~\new_[9026]_  | ~\new_[7738]_ ;
  assign \new_[8448]_  = ~\new_[9026]_  | ~\new_[11036]_ ;
  assign \new_[8449]_  = ~\new_[9026]_  | ~\new_[7828]_ ;
  assign \new_[8450]_  = ~\new_[9026]_  | ~\new_[7723]_ ;
  assign \new_[8451]_  = ~\new_[9026]_  | ~\new_[7833]_ ;
  assign \new_[8452]_  = ~\new_[9026]_  | ~\new_[11092]_ ;
  assign \new_[8453]_  = ~\new_[9026]_  | ~\new_[11186]_ ;
  assign \new_[8454]_  = ~\new_[9026]_  | ~\new_[11089]_ ;
  assign \new_[8455]_  = ~\new_[9026]_  | ~\new_[7850]_ ;
  assign \new_[8456]_  = ~\new_[8864]_  & ~\new_[12099]_ ;
  assign \new_[8457]_  = ~\new_[11390]_ ;
  assign n4491 = \wb_data_i[8]  ? \new_[8870]_  : \new_[8205]_ ;
  assign n4451 = \wb_data_i[9]  ? \new_[8870]_  : \new_[8194]_ ;
  assign n4496 = \wb_data_i[3]  ? \new_[8870]_  : \new_[8229]_ ;
  assign n4456 = \wb_data_i[10]  ? \new_[8870]_  : \new_[8195]_ ;
  assign n4461 = \wb_data_i[2]  ? \new_[8870]_  : \new_[8196]_ ;
  assign n4441 = \wb_data_i[1]  ? \new_[8870]_  : \new_[8179]_ ;
  assign n4476 = \wb_data_i[5]  ? \new_[8870]_  : \new_[8199]_ ;
  assign n4481 = \wb_data_i[6]  ? \new_[8870]_  : \new_[8200]_ ;
  assign n4486 = \wb_data_i[7]  ? \new_[8870]_  : \new_[8201]_ ;
  assign n4471 = \wb_data_i[4]  ? \new_[8870]_  : \new_[8198]_ ;
  assign n4426 = \wb_data_i[0]  ? \new_[8870]_  : \new_[8149]_ ;
  assign \new_[8469]_  = ~\new_[2094]_  | ~\new_[11309]_ ;
  assign \new_[8470]_  = ~\new_[2108]_  | ~\new_[12764]_ ;
  assign \new_[8471]_  = ~\new_[2103]_  | ~\new_[11309]_ ;
  assign \new_[8472]_  = ~\new_[2116]_  | ~\new_[11876]_ ;
  assign \new_[8473]_  = ~\new_[2131]_  | ~\new_[12766]_ ;
  assign \new_[8474]_  = ~\new_[2081]_  | ~\new_[12767]_ ;
  assign \new_[8475]_  = ~\new_[9957]_  | ~\new_[11572]_  | ~\new_[8880]_  | ~\new_[8912]_ ;
  assign \new_[8476]_  = ~\new_[8799]_  & (~\new_[9493]_  | ~\new_[7977]_ );
  assign \new_[8477]_  = ~\new_[8714]_ ;
  assign n4466 = (~\new_[8197]_  & ~n5306) | (~\new_[10072]_  & ~\new_[1433]_ );
  assign \new_[8479]_  = ~\new_[8798]_  & (~\new_[9493]_  | ~\new_[7966]_ );
  assign \new_[8480]_  = ~\new_[10072]_  | ~\new_[11776]_ ;
  assign \new_[8481]_  = \\u1_u0_out_r_reg[10] ;
  assign \new_[8482]_  = ~\new_[9163]_  & ~\new_[8821]_ ;
  assign \new_[8483]_  = \\u1_u0_out_r_reg[8] ;
  assign \new_[8484]_  = (~\new_[9725]_  | ~\new_[8820]_ ) & (~\new_[9170]_  | ~\new_[1657]_ );
  assign \new_[8485]_  = \new_[1841]_  ^ \new_[9170]_ ;
  assign \new_[8486]_  = ~\new_[7280]_  | ~\new_[8786]_ ;
  assign \new_[8487]_  = ~\new_[8820]_  & ~\new_[12469]_ ;
  assign \new_[8488]_  = ~\new_[11337]_  | ~\new_[12731]_  | ~\new_[9570]_  | ~\new_[10196]_ ;
  assign \new_[8489]_  = ~\new_[10246]_  | ~\new_[10348]_  | ~\new_[8789]_  | ~\new_[10029]_ ;
  assign \new_[8490]_  = \new_[9724]_  ? \new_[8821]_  : \new_[1611]_ ;
  assign \new_[8491]_  = \new_[1453]_  ^ \new_[8821]_ ;
  assign \new_[8492]_  = u4_rfr_early_reg;
  assign \new_[8493]_  = ~\new_[9400]_  & ~\new_[8821]_ ;
  assign mc_rp_pad_o_ = u7_mc_rp_reg;
  assign \new_[8495]_  = (~\new_[9198]_  & ~\new_[10007]_  & ~\new_[10482]_ ) | (~\new_[10459]_  & ~\new_[9195]_  & ~\new_[10109]_ );
  assign \new_[8496]_  = (~\new_[9194]_  & ~\new_[10074]_  & ~\new_[10413]_ ) | (~\new_[10408]_  & ~\new_[9353]_  & ~\new_[10085]_ );
  assign \new_[8497]_  = (~\new_[9196]_  & ~\new_[9983]_  & ~\new_[10484]_ ) | (~\new_[10457]_  & ~\new_[9193]_  & ~\new_[10008]_ );
  assign \new_[8498]_  = \new_[11777]_  & \new_[10933]_ ;
  assign \new_[8499]_  = ~\new_[11528]_ ;
  assign \new_[8500]_  = \new_[11777]_  & \new_[11356]_ ;
  assign \new_[8501]_  = \new_[11777]_  & \new_[11363]_ ;
  assign \new_[8502]_  = \new_[11777]_  & \new_[11576]_ ;
  assign \new_[8503]_  = \new_[11777]_  & \new_[12273]_ ;
  assign \new_[8504]_  = \new_[11777]_  & \new_[9785]_ ;
  assign \new_[8505]_  = \new_[11777]_  & \new_[10802]_ ;
  assign \new_[8506]_  = \new_[11777]_  & \new_[12093]_ ;
  assign \new_[8507]_  = \new_[11777]_  & n5021;
  assign \new_[8508]_  = \new_[11777]_  & \new_[12567]_ ;
  assign \new_[8509]_  = \new_[11777]_  & \new_[10164]_ ;
  assign \new_[8510]_  = \new_[11777]_  & \new_[10411]_ ;
  assign \new_[8511]_  = \new_[11777]_  & \new_[9674]_ ;
  assign \new_[8512]_  = \new_[11777]_  & \new_[12610]_ ;
  assign \new_[8513]_  = \new_[11777]_  & \new_[10955]_ ;
  assign \new_[8514]_  = \new_[11777]_  & \new_[11353]_ ;
  assign \new_[8515]_  = \new_[11777]_  & \new_[10496]_ ;
  assign \new_[8516]_  = \new_[11777]_  & \new_[11328]_ ;
  assign \new_[8517]_  = \new_[11777]_  & \new_[11367]_ ;
  assign \new_[8518]_  = \new_[11777]_  & \new_[11310]_ ;
  assign \new_[8519]_  = \new_[11777]_  & \new_[11313]_ ;
  assign \new_[8520]_  = \new_[11777]_  & \new_[10960]_ ;
  assign \new_[8521]_  = n4651 | \new_[11217]_ ;
  assign \new_[8522]_  = ~\new_[9026]_  | ~\new_[7724]_ ;
  assign n4501 = ~\new_[11435]_ ;
  assign \new_[8524]_  = ~\new_[8957]_  & ~\new_[12052]_ ;
  assign \new_[8525]_  = \new_[9242]_  ? \new_[10201]_  : \new_[9016]_ ;
  assign \new_[8526]_  = \new_[9243]_  ? \new_[10201]_  : \new_[9025]_ ;
  assign \new_[8527]_  = \new_[9246]_  ? \new_[10201]_  : \new_[9019]_ ;
  assign \new_[8528]_  = \new_[9199]_  ? \new_[10201]_  : \new_[8998]_ ;
  assign \new_[8529]_  = \new_[9270]_  ? \new_[10201]_  : \new_[9157]_ ;
  assign \new_[8530]_  = \new_[9497]_  ? \new_[10201]_  : \new_[9009]_ ;
  assign \new_[8531]_  = \new_[9495]_  ? \new_[10201]_  : \new_[9013]_ ;
  assign \new_[8532]_  = \new_[9496]_  ? \new_[10201]_  : \new_[8993]_ ;
  assign \new_[8533]_  = \new_[9498]_  ? \new_[10201]_  : \new_[8996]_ ;
  assign \new_[8534]_  = \new_[9416]_  ? \new_[10201]_  : \new_[8994]_ ;
  assign \new_[8535]_  = \new_[9244]_  ? \new_[10201]_  : \new_[9014]_ ;
  assign \new_[8536]_  = \new_[9415]_  ? \new_[10201]_  : \new_[8995]_ ;
  assign \new_[8537]_  = \new_[9397]_  ? \new_[10201]_  : \new_[9005]_ ;
  assign \new_[8538]_  = ~\new_[9215]_  | ~\new_[9909]_  | ~\new_[9429]_  | ~\new_[9470]_ ;
  assign \new_[8539]_  = ~\new_[9218]_  | ~\new_[9778]_  | ~\new_[9474]_  | ~\new_[9471]_ ;
  assign \new_[8540]_  = ~\new_[9213]_  | ~\new_[9758]_  | ~\new_[9452]_  | ~\new_[9466]_ ;
  assign \new_[8541]_  = ~\new_[9219]_  | ~\new_[9907]_  | ~\new_[9450]_  | ~\new_[9469]_ ;
  assign \new_[8542]_  = ~\new_[9209]_  | ~\new_[9754]_  | ~\new_[9455]_  | ~\new_[9431]_ ;
  assign \new_[8543]_  = \new_[8063]_  ? n4691 : \wb_data_i[0] ;
  assign \new_[8544]_  = \new_[8072]_  ? n4691 : \wb_data_i[10] ;
  assign \new_[8545]_  = \new_[11243]_  ? n4691 : \wb_data_i[11] ;
  assign \new_[8546]_  = \new_[11066]_  ? n4691 : \wb_data_i[12] ;
  assign \new_[8547]_  = \new_[11093]_  ? n4691 : \wb_data_i[13] ;
  assign \new_[8548]_  = \new_[11188]_  ? n4691 : \wb_data_i[14] ;
  assign \new_[8549]_  = \new_[11240]_  ? n4691 : \wb_data_i[15] ;
  assign \new_[8550]_  = \new_[11082]_  ? n4691 : \wb_data_i[16] ;
  assign \new_[8551]_  = \new_[11220]_  ? n4691 : \wb_data_i[17] ;
  assign \new_[8552]_  = \new_[11245]_  ? n4691 : \wb_data_i[18] ;
  assign \new_[8553]_  = \new_[11223]_  ? n4691 : \wb_data_i[19] ;
  assign \new_[8554]_  = \new_[11043]_  ? n4691 : \wb_data_i[20] ;
  assign \new_[8555]_  = \new_[11250]_  ? n4691 : \wb_data_i[22] ;
  assign \new_[8556]_  = \new_[11249]_  ? n4691 : \wb_data_i[23] ;
  assign \new_[8557]_  = \new_[11028]_  ? n4691 : \wb_data_i[24] ;
  assign \new_[8558]_  = \new_[11241]_  ? n4691 : \wb_data_i[25] ;
  assign \new_[8559]_  = \new_[11234]_  ? n4691 : \wb_data_i[27] ;
  assign \new_[8560]_  = \new_[10986]_  ? n4691 : \wb_data_i[28] ;
  assign \new_[8561]_  = \new_[10991]_  ? n4691 : \wb_data_i[29] ;
  assign \new_[8562]_  = \new_[8078]_  ? n4691 : \wb_data_i[2] ;
  assign \new_[8563]_  = \new_[11226]_  ? n4691 : \wb_data_i[30] ;
  assign \new_[8564]_  = \new_[11074]_  ? n4691 : \wb_data_i[31] ;
  assign \new_[8565]_  = \new_[8067]_  ? n4691 : \wb_data_i[3] ;
  assign \new_[8566]_  = \new_[8048]_  ? n4691 : \wb_data_i[4] ;
  assign \new_[8567]_  = \new_[8052]_  ? n4691 : \wb_data_i[5] ;
  assign \new_[8568]_  = \new_[8051]_  ? n4691 : \wb_data_i[6] ;
  assign \new_[8569]_  = \new_[8068]_  ? n4691 : \wb_data_i[7] ;
  assign \new_[8570]_  = \new_[8043]_  ? n4691 : \wb_data_i[9] ;
  assign \new_[8571]_  = \new_[8023]_  ? n4691 : \wb_data_i[8] ;
  assign \new_[8572]_  = \new_[11022]_  ? n4691 : \wb_data_i[21] ;
  assign \new_[8573]_  = \new_[11013]_  ? n4691 : \wb_data_i[26] ;
  assign \new_[8574]_  = \new_[8993]_  ^ \new_[9157]_ ;
  assign \new_[8575]_  = \new_[9014]_  ^ \new_[9013]_ ;
  assign \new_[8576]_  = \new_[8996]_  ^ \new_[11797]_ ;
  assign \new_[8577]_  = \new_[8992]_  ^ \new_[9022]_ ;
  assign \new_[8578]_  = \new_[9158]_  ^ \new_[9024]_ ;
  assign \new_[8579]_  = \new_[8997]_  ^ \new_[9011]_ ;
  assign \new_[8580]_  = \new_[9016]_  ^ \new_[9025]_ ;
  assign \new_[8581]_  = \new_[8999]_  ^ \new_[9009]_ ;
  assign \new_[8582]_  = \new_[9012]_  ^ \new_[9000]_ ;
  assign \new_[8583]_  = \new_[9002]_  ^ \new_[9008]_ ;
  assign \new_[8584]_  = \new_[9005]_  ^ \new_[9131]_ ;
  assign \new_[8585]_  = \new_[9162]_  ^ \new_[9003]_ ;
  assign \new_[8586]_  = \new_[9018]_  ^ \new_[9021]_ ;
  assign \new_[8587]_  = \new_[9001]_  ^ \new_[9020]_ ;
  assign \new_[8588]_  = \new_[8994]_  ^ \new_[8995]_ ;
  assign \new_[8589]_  = u0_u1_lmr_req_we_reg;
  assign \new_[8590]_  = n4651 | \new_[7922]_ ;
  assign \new_[8591]_  = ~\new_[9026]_  | ~\new_[11247]_ ;
  assign \new_[8592]_  = ~\new_[9026]_  | ~\new_[11088]_ ;
  assign \new_[8593]_  = ~\new_[9026]_  | ~\new_[11008]_ ;
  assign \new_[8594]_  = ~\new_[9026]_  | ~\new_[11190]_ ;
  assign \new_[8595]_  = ~\new_[9026]_  | ~\new_[7733]_ ;
  assign \new_[8596]_  = ~\new_[9026]_  | ~\new_[7722]_ ;
  assign \new_[8597]_  = ~\new_[9026]_  | ~\new_[10978]_ ;
  assign \new_[8598]_  = ~\new_[9026]_  | ~\new_[7951]_ ;
  assign \new_[8599]_  = n4651 | \new_[10982]_ ;
  assign \new_[8600]_  = n4651 | \new_[7968]_ ;
  assign \new_[8601]_  = n4651 | \new_[7943]_ ;
  assign \new_[8602]_  = n4651 | \new_[7969]_ ;
  assign \new_[8603]_  = n4651 | \new_[7941]_ ;
  assign \new_[8604]_  = n4651 | \new_[7950]_ ;
  assign \new_[8605]_  = n4651 | \new_[7981]_ ;
  assign \new_[8606]_  = n4651 | \new_[7970]_ ;
  assign \new_[8607]_  = n4651 | \new_[7985]_ ;
  assign \new_[8608]_  = n4651 | \new_[7984]_ ;
  assign \new_[8609]_  = n4651 | \new_[7939]_ ;
  assign \new_[8610]_  = n4651 | \new_[11023]_ ;
  assign \new_[8611]_  = n4651 | \new_[11054]_ ;
  assign \new_[8612]_  = n4651 | \new_[7935]_ ;
  assign \new_[8613]_  = n4651 | \new_[10981]_ ;
  assign \new_[8614]_  = n4651 | \new_[7914]_ ;
  assign \new_[8615]_  = n4651 | \new_[7973]_ ;
  assign \new_[8616]_  = n4651 | \new_[11032]_ ;
  assign \new_[8617]_  = n4651 | \new_[10999]_ ;
  assign \new_[8618]_  = n4651 | \new_[11149]_ ;
  assign \new_[8619]_  = n4651 | \new_[11172]_ ;
  assign \new_[8620]_  = n4651 | \new_[11157]_ ;
  assign \new_[8621]_  = n4651 | \new_[11163]_ ;
  assign \new_[8622]_  = n4651 | \new_[11077]_ ;
  assign \new_[8623]_  = n4651 | \new_[7917]_ ;
  assign \new_[8624]_  = ~\new_[9026]_  | ~\new_[7960]_ ;
  assign \new_[8625]_  = n4651 | \new_[11152]_ ;
  assign \new_[8626]_  = ~\new_[9026]_  | ~\new_[7730]_ ;
  assign \new_[8627]_  = n4651 | \new_[11118]_ ;
  assign \new_[8628]_  = ~\new_[9026]_  | ~\new_[7703]_ ;
  assign \new_[8629]_  = n4651 | \new_[7932]_ ;
  assign \new_[8630]_  = ~\new_[9026]_  | ~\new_[7694]_ ;
  assign \new_[8631]_  = n4651 | \new_[11096]_ ;
  assign \new_[8632]_  = ~\new_[9026]_  | ~\new_[11166]_ ;
  assign \new_[8633]_  = ~n4651 | ~\wb_data_i[16] ;
  assign n3951 = ~\new_[11779]_ ;
  assign \new_[8635]_  = ~n4651 | ~\wb_data_i[18] ;
  assign \new_[8636]_  = ~n4651 | ~\wb_data_i[30] ;
  assign \new_[8637]_  = ~\new_[8773]_ ;
  assign \new_[8638]_  = ~n4651 | ~\wb_data_i[15] ;
  assign \new_[8639]_  = ~n4521 | ~\wb_data_i[3] ;
  assign \new_[8640]_  = ~n4521 | ~\wb_data_i[0] ;
  assign \new_[8641]_  = ~n4521 | ~\wb_data_i[11] ;
  assign \new_[8642]_  = ~n4521 | ~\wb_data_i[18] ;
  assign \new_[8643]_  = ~n4521 | ~\wb_data_i[23] ;
  assign \new_[8644]_  = ~n4521 | ~\wb_data_i[25] ;
  assign \new_[8645]_  = ~n4521 | ~\wb_data_i[2] ;
  assign \new_[8646]_  = ~n4521 | ~\wb_data_i[6] ;
  assign \new_[8647]_  = ~n4521 | ~\wb_data_i[8] ;
  assign \new_[8648]_  = ~n4651 | ~\wb_data_i[0] ;
  assign \new_[8649]_  = ~n4651 | ~\wb_data_i[12] ;
  assign \new_[8650]_  = ~n4651 | ~\wb_data_i[17] ;
  assign \new_[8651]_  = ~n4521 | ~\wb_data_i[29] ;
  assign \new_[8652]_  = ~n4651 | ~\wb_data_i[20] ;
  assign \new_[8653]_  = ~n4651 | ~\wb_data_i[22] ;
  assign \new_[8654]_  = ~n4651 | ~\wb_data_i[13] ;
  assign \new_[8655]_  = ~n4651 | ~\wb_data_i[24] ;
  assign \new_[8656]_  = ~n4651 | ~\wb_data_i[28] ;
  assign \new_[8657]_  = ~n4651 | ~\wb_data_i[31] ;
  assign \new_[8658]_  = ~n4521 | ~\wb_data_i[28] ;
  assign \new_[8659]_  = ~n4651 | ~\wb_data_i[5] ;
  assign \new_[8660]_  = ~n4651 | ~\wb_data_i[6] ;
  assign \new_[8661]_  = ~n4651 | ~\wb_data_i[7] ;
  assign \new_[8662]_  = ~n4651 | ~\wb_data_i[9] ;
  assign \new_[8663]_  = ~n4651 | ~\wb_data_i[4] ;
  assign \new_[8664]_  = ~n4651 | ~\wb_data_i[29] ;
  assign \new_[8665]_  = ~n4651 | ~\wb_data_i[21] ;
  assign \new_[8666]_  = ~n4651 | ~\wb_data_i[14] ;
  assign \new_[8667]_  = ~n4651 | ~\wb_data_i[25] ;
  assign \new_[8668]_  = ~n4521 | ~\wb_data_i[1] ;
  assign \new_[8669]_  = ~n4651 | ~\wb_data_i[3] ;
  assign \new_[8670]_  = ~n4651 | ~\wb_data_i[19] ;
  assign \new_[8671]_  = ~\new_[8858]_  & ~\new_[10316]_ ;
  assign \new_[8672]_  = ~n4651 | ~\wb_data_i[2] ;
  assign \new_[8673]_  = ~n4651 | ~\wb_data_i[8] ;
  assign \new_[8674]_  = ~n4651 | ~\wb_data_i[27] ;
  assign \new_[8675]_  = ~n4651 | ~\wb_data_i[1] ;
  assign \new_[8676]_  = ~n4651 | ~\wb_data_i[26] ;
  assign n4516 = ~\new_[8855]_  | (~\new_[9236]_  & ~\new_[11051]_ );
  assign n4526 = \new_[8296]_  ? \new_[9045]_  : \wb_data_i[24] ;
  assign n4571 = \new_[8378]_  ? \new_[9045]_  : \wb_data_i[27] ;
  assign n4506 = \new_[8232]_  ? \new_[9045]_  : \wb_data_i[30] ;
  assign n4601 = \new_[8390]_  ? \new_[9045]_  : \wb_data_i[31] ;
  assign n4576 = mc_vpen_pad_o ? \new_[9045]_  : \wb_data_i[1] ;
  assign n4591 = \new_[8387]_  ? \new_[9045]_  : \wb_data_i[2] ;
  assign n4596 = \new_[11203]_  ? \new_[9045]_  : \wb_data_i[4] ;
  assign n4606 = \new_[11253]_  ? \new_[9045]_  : \wb_data_i[5] ;
  assign n4551 = \new_[11042]_  ? \new_[9045]_  : \wb_data_i[6] ;
  assign n4531 = \new_[11126]_  ? \new_[9045]_  : \wb_data_i[7] ;
  assign \new_[8688]_  = u6_read_go_r1_reg;
  assign n4536 = \new_[8352]_  ? \new_[9045]_  : \wb_data_i[25] ;
  assign n4511 = \new_[8260]_  ? \new_[9045]_  : \wb_data_i[28] ;
  assign n4611 = \new_[8399]_  ? \new_[9045]_  : \wb_data_i[10] ;
  assign n4541 = \new_[8355]_  ? \new_[9045]_  : \wb_data_i[26] ;
  assign n4556 = \new_[8365]_  ? \new_[9045]_  : \wb_data_i[9] ;
  assign \new_[8694]_  = ~\new_[9265]_  & ~\new_[8872]_ ;
  assign \new_[8695]_  = ~\new_[11359]_  | ~\new_[12401]_  | ~\new_[12543]_  | ~\new_[9054]_ ;
  assign \new_[8696]_  = ~\new_[10466]_  | ~\new_[12555]_  | ~\new_[12459]_  | ~\new_[9057]_ ;
  assign \new_[8697]_  = ~\new_[11298]_  | ~\new_[11881]_  | ~\new_[8945]_  | ~\new_[9916]_ ;
  assign \new_[8698]_  = ~\new_[11310]_  | ~\new_[11314]_  | ~\new_[12543]_  | ~\new_[9146]_ ;
  assign \new_[8699]_  = ~\new_[10450]_  | ~\new_[12756]_  | ~\new_[9570]_  | ~\new_[9056]_ ;
  assign \new_[8700]_  = ~\new_[11311]_  | ~\new_[11313]_  | ~\new_[12543]_  | ~\new_[9146]_ ;
  assign \new_[8701]_  = ~\new_[10017]_  | ~\new_[9730]_  | ~\new_[8867]_  | ~\new_[10209]_ ;
  assign \new_[8702]_  = n4651 | \new_[7936]_ ;
  assign \new_[8703]_  = ~\new_[9357]_  | ~\new_[11335]_  | ~\new_[10301]_  | ~\new_[10143]_ ;
  assign \new_[8704]_  = ~\\u3_mc_dp_o_reg[3] ;
  assign \new_[8705]_  = ~\new_[12730]_  & ~\new_[11353]_ ;
  assign \new_[8706]_  = \new_[8881]_  & \new_[9730]_ ;
  assign \new_[8707]_  = ~\new_[12337]_  | ~\new_[8881]_  | ~\new_[9318]_ ;
  assign \new_[8708]_  = ~\new_[10959]_  | ~\new_[12040]_  | ~\new_[11168]_ ;
  assign \new_[8709]_  = ~\new_[10265]_  & (~\new_[10461]_  | ~\new_[10511]_ );
  assign \new_[8710]_  = \new_[10572]_  & \new_[10928]_ ;
  assign \new_[8711]_  = \new_[9019]_  ^ \new_[8998]_ ;
  assign \new_[8712]_  = ~\new_[9902]_  | ~\new_[10195]_ ;
  assign \new_[8713]_  = ~\new_[12755]_  | ~\new_[9902]_ ;
  assign \new_[8714]_  = ~\new_[12447]_ ;
  assign n4616 = \new_[8400]_  ? \new_[9045]_  : \wb_data_i[29] ;
  assign n4586 = \new_[8382]_  ? \new_[9045]_  : \wb_data_i[8] ;
  assign \new_[8717]_  = ~\\u3_mc_dp_o_reg[2] ;
  assign \new_[8718]_  = ~\\u3_mc_dp_o_reg[0] ;
  assign n4581 = \new_[11213]_  ? \new_[9045]_  : \wb_data_i[3] ;
  assign \new_[8720]_  = ~\new_[9396]_  | ~\new_[8880]_ ;
  assign \new_[8721]_  = ~\\u3_mc_dp_o_reg[1] ;
  assign n4546 = ~\new_[8812]_ ;
  assign \new_[8723]_  = ~\new_[11131]_  | ~\new_[8967]_  | ~\new_[11026]_ ;
  assign \new_[8724]_  = ~\new_[8961]_  & (~\new_[9493]_  | ~\new_[8049]_ );
  assign \new_[8725]_  = ~\new_[10089]_  & (~\new_[10805]_  | ~\new_[10511]_ );
  assign \new_[8726]_  = \new_[9499]_  ? \new_[10201]_  : \new_[11797]_ ;
  assign \new_[8727]_  = \new_[11777]_  & \new_[9946]_ ;
  assign \new_[8728]_  = \new_[9247]_  ? \new_[10201]_  : \new_[9131]_ ;
  assign n4561 = ~\new_[8950]_  | (~\new_[9238]_  & ~\new_[11131]_ );
  assign \new_[8730]_  = \new_[9240]_  ? \new_[10201]_  : \new_[8999]_ ;
  assign \new_[8731]_  = ~\new_[10293]_  | ~\new_[10386]_  | ~\new_[8842]_  | ~\new_[10427]_ ;
  assign \new_[8732]_  = ~n4651 | ~\wb_data_i[23] ;
  assign \new_[8733]_  = \new_[9343]_  | \new_[9170]_ ;
  assign \new_[8734]_  = u6_write_go_r1_reg;
  assign \new_[8735]_  = ~n4651 | ~\wb_data_i[11] ;
  assign n4566 = ~\new_[8824]_  & (~\new_[10521]_  | ~\new_[10449]_ );
  assign \new_[8737]_  = \new_[8061]_  ? n4691 : \wb_data_i[1] ;
  assign \new_[8738]_  = ~\new_[10518]_  & ~\new_[8821]_ ;
  assign \new_[8739]_  = ~\new_[10002]_  & ~\new_[8821]_ ;
  assign \new_[8740]_  = ~\new_[11490]_  & ~\new_[12398]_ ;
  assign \new_[8741]_  = ~n4651 | ~\wb_data_i[10] ;
  assign \new_[8742]_  = ~\new_[11490]_  & (~\new_[11491]_  | ~\new_[12610]_ );
  assign \new_[8743]_  = ~\new_[8822]_  & (~\new_[9493]_  | ~\new_[8075]_ );
  assign \new_[8744]_  = ~\new_[9026]_  | ~\new_[11198]_ ;
  assign \new_[8745]_  = ~\new_[9449]_  | ~\new_[9919]_  | ~\new_[9650]_  | ~\new_[9893]_ ;
  assign \new_[8746]_  = ~\new_[9656]_  | ~\new_[9900]_  | ~\new_[9464]_  | ~\new_[9767]_ ;
  assign \new_[8747]_  = ~\new_[9458]_  | ~\new_[9427]_  | ~\new_[9208]_  | ~\new_[9766]_ ;
  assign \new_[8748]_  = ~\new_[11525]_ ;
  assign \new_[8749]_  = ~\new_[11490]_ ;
  assign \new_[8750]_  = ~\new_[9398]_  | ~\new_[9435]_  | ~\new_[9210]_  | ~\new_[9777]_ ;
  assign \new_[8751]_  = ~\new_[9434]_  | ~\new_[9423]_  | ~\new_[9206]_  | ~\new_[9771]_ ;
  assign \new_[8752]_  = ~\new_[9465]_  | ~\new_[9920]_  | ~\new_[9637]_  | ~\new_[9898]_ ;
  assign \new_[8753]_  = ~\new_[9440]_  | ~\new_[9757]_  | ~\new_[9438]_  | ~\new_[9769]_ ;
  assign \new_[8754]_  = ~\new_[9402]_  | ~\new_[9759]_  | ~\new_[9425]_  | ~\new_[9770]_ ;
  assign \new_[8755]_  = ~\new_[9445]_  | ~\new_[9432]_  | ~\new_[9217]_  | ~\new_[9780]_ ;
  assign \new_[8756]_  = ~\new_[9436]_  | ~\new_[9459]_  | ~\new_[9212]_  | ~\new_[9891]_ ;
  assign \new_[8757]_  = ~\new_[9428]_  | ~\new_[9451]_  | ~\new_[9214]_  | ~\new_[9901]_ ;
  assign \new_[8758]_  = ~\new_[9463]_  | ~\new_[9910]_  | ~\new_[9433]_  | ~\new_[9875]_ ;
  assign \new_[8759]_  = ~\new_[9467]_  | ~\new_[9761]_  | ~\new_[9468]_  | ~\new_[9881]_ ;
  assign \new_[8760]_  = ~\new_[9475]_  | ~\new_[9760]_  | ~\new_[9426]_  | ~\new_[9869]_ ;
  assign \new_[8761]_  = ~\new_[8981]_  | (~\new_[9669]_  & ~\new_[1842]_ );
  assign \new_[8762]_  = ~\new_[8980]_  & (~\new_[9493]_  | ~\new_[8079]_ );
  assign \new_[8763]_  = ~\new_[8991]_  & ~\new_[10006]_ ;
  assign \new_[8764]_  = ~\new_[8988]_  & (~\new_[9493]_  | ~\new_[8081]_ );
  assign \new_[8765]_  = ~\new_[8989]_  | (~\new_[9695]_  & ~\new_[1955]_ );
  assign \new_[8766]_  = \\u1_u0_out_r_reg[5] ;
  assign \new_[8767]_  = ~\new_[9003]_  | ~\new_[10201]_ ;
  assign \new_[8768]_  = ~\new_[9012]_  | ~\new_[10201]_ ;
  assign \new_[8769]_  = ~\new_[8992]_  | ~\new_[10201]_ ;
  assign \new_[8770]_  = ~\new_[9020]_  | ~\new_[10201]_ ;
  assign \new_[8771]_  = ~\new_[9008]_  | ~\new_[10201]_ ;
  assign \new_[8772]_  = \new_[9007]_  & \new_[9136]_ ;
  assign \new_[8773]_  = ~\new_[12400]_  | ~\new_[10322]_  | ~\new_[9044]_  | ~\new_[11338]_ ;
  assign \new_[8774]_  = ~\new_[9021]_  | ~\new_[10201]_ ;
  assign \new_[8775]_  = ~\new_[9022]_  | ~\new_[10201]_ ;
  assign \new_[8776]_  = ~\new_[9140]_  & ~\new_[10213]_ ;
  assign \new_[8777]_  = ~\new_[9000]_  | ~\new_[10201]_ ;
  assign \new_[8778]_  = ~\new_[8997]_  | ~\new_[10201]_ ;
  assign \new_[8779]_  = ~\new_[9162]_  | ~\new_[10201]_ ;
  assign \new_[8780]_  = ~\new_[9018]_  | ~\new_[10201]_ ;
  assign \new_[8781]_  = ~\new_[9158]_  | ~\new_[10201]_ ;
  assign \new_[8782]_  = ~\new_[9024]_  | ~\new_[10201]_ ;
  assign \new_[8783]_  = ~\new_[9011]_  | ~\new_[10201]_ ;
  assign \new_[8784]_  = ~\new_[9002]_  | ~\new_[10201]_ ;
  assign \new_[8785]_  = ~\new_[9001]_  | ~\new_[10201]_ ;
  assign \new_[8786]_  = ~\new_[9007]_  | ~\new_[10949]_ ;
  assign n4626 = ~\new_[10499]_  | ~\new_[9031]_ ;
  assign n4236 = ~\new_[8856]_ ;
  assign \new_[8789]_  = ~\new_[9035]_  & ~\new_[9819]_ ;
  assign \new_[8790]_  = ~\new_[10123]_  | ~\new_[12090]_  | ~\new_[9693]_ ;
  assign \new_[8791]_  = ~\new_[9991]_  | ~\new_[11351]_  | ~\new_[9267]_  | ~\new_[10209]_ ;
  assign \new_[8792]_  = \new_[10572]_  & \new_[9648]_ ;
  assign n4646 = ~\new_[8387]_  & ~n4706;
  assign \new_[8794]_  = ~\new_[11892]_  | ~\new_[11889]_  | ~\new_[1480]_ ;
  assign \new_[8795]_  = \new_[9058]_  & \new_[12444]_ ;
  assign \new_[8796]_  = \new_[12731]_  & \new_[11353]_ ;
  assign \new_[8797]_  = \new_[10432]_  & \new_[12731]_ ;
  assign \new_[8798]_  = ~\new_[9126]_  & ~\new_[9493]_ ;
  assign \new_[8799]_  = ~\new_[9151]_  & ~\new_[9493]_ ;
  assign \new_[8800]_  = ~\new_[9103]_  | ~\new_[10598]_ ;
  assign \new_[8801]_  = \new_[10572]_  & \new_[10164]_ ;
  assign \new_[8802]_  = \new_[10572]_  & \new_[9379]_ ;
  assign \new_[8803]_  = \new_[10572]_  & \new_[10496]_ ;
  assign \new_[8804]_  = u0_u0_lmr_req_we_reg;
  assign \new_[8805]_  = ~\new_[9894]_ ;
  assign \new_[8806]_  = ~\new_[10268]_  | ~\new_[10920]_ ;
  assign \new_[8807]_  = ~\new_[8197]_  & ~\new_[10658]_ ;
  assign n4636 = \new_[11205]_  ^ \new_[9367]_ ;
  assign \new_[8809]_  = u0_rf_we_reg;
  assign \new_[8810]_  = u6_wr_hold_reg;
  assign mc_zz_pad_o = u7_mc_zz_o_reg;
  assign \new_[8812]_  = ~\new_[11026]_  | ~\new_[11235]_  | ~\new_[9156]_  | ~\new_[10361]_ ;
  assign \new_[8813]_  = u5_lookup_ready2_reg;
  assign n4641 = ~\new_[8824]_ ;
  assign n4621 = \new_[10836]_  ^ \new_[9959]_ ;
  assign \new_[8816]_  = \\u1_u0_out_r_reg[6] ;
  assign \new_[8817]_  = \new_[9781]_  | \new_[9170]_ ;
  assign \new_[8818]_  = \new_[1843]_  ^ \new_[9175]_ ;
  assign n4631 = \new_[11026]_  ^ \new_[9173]_ ;
  assign \new_[8820]_  = ~\new_[9170]_ ;
  assign \new_[8821]_  = n4741 | \new_[10072]_ ;
  assign \new_[8822]_  = ~\new_[9187]_  & ~\new_[9493]_ ;
  assign \poc_o[0]  = \\u0_poc_reg[0] ;
  assign \new_[8824]_  = \new_[9943]_  | \new_[10684]_  | \new_[10653]_  | \new_[10648]_ ;
  assign n4671 = \new_[9411]_  ? \new_[10221]_  : n5646;
  assign n4676 = \new_[9410]_  ? \new_[10221]_  : n5671;
  assign n4666 = \new_[9414]_  ? \new_[10221]_  : n5481;
  assign \new_[8828]_  = ~\new_[9437]_  | ~\new_[9387]_  | ~\new_[9787]_ ;
  assign \new_[8829]_  = ~\new_[9444]_  | ~\new_[9430]_  | ~\new_[9887]_ ;
  assign \new_[8830]_  = ~\new_[9211]_  & ~\new_[10268]_ ;
  assign \new_[8831]_  = \new_[9211]_  & \new_[10511]_ ;
  assign \new_[8832]_  = ~\new_[9421]_  | ~\new_[9597]_  | ~\new_[9784]_ ;
  assign \new_[8833]_  = ~\new_[9654]_  | ~\new_[9447]_  | ~\new_[9802]_ ;
  assign \new_[8834]_  = ~\new_[9645]_  | ~\new_[9456]_  | ~\new_[9858]_ ;
  assign \new_[8835]_  = ~\new_[9461]_  | ~\new_[9457]_  | ~\new_[9775]_ ;
  assign \new_[8836]_  = ~\new_[9442]_  | ~\new_[9462]_  | ~\new_[9876]_ ;
  assign \new_[8837]_  = ~\new_[9472]_  | ~\new_[9605]_  | ~\new_[9773]_ ;
  assign \new_[8838]_  = ~\new_[9473]_  | ~\new_[9453]_  | ~\new_[9786]_ ;
  assign n4656 = ~\new_[9403]_  & (~\new_[9638]_  | ~\new_[10445]_ );
  assign \new_[8840]_  = ~\new_[11491]_ ;
  assign \new_[8841]_  = ~\new_[9370]_  & (~\new_[10337]_  | ~\new_[10434]_ );
  assign \new_[8842]_  = ~\new_[9384]_  & ~\new_[10080]_ ;
  assign \new_[8843]_  = ~\new_[9227]_  & (~\new_[10094]_  | ~\new_[10429]_ );
  assign \new_[8844]_  = ~\new_[9235]_  & (~\new_[10093]_  | ~\new_[10480]_ );
  assign \new_[8845]_  = \new_[8071]_  ^ \new_[9493]_ ;
  assign n4681 = \new_[9336]_  & wb_cyc_i;
  assign \new_[8847]_  = ~\new_[12595]_  & ~\new_[12097]_  & ~\new_[12545]_ ;
  assign \new_[8848]_  = ~\new_[3036]_  | ~wb_cyc_i | ~\new_[9557]_ ;
  assign n4651 = \new_[9255]_  & \new_[10042]_ ;
  assign \new_[8850]_  = ~\new_[10906]_  | ~\new_[10897]_  | ~\new_[9262]_  | ~\new_[9805]_ ;
  assign \new_[8851]_  = ~\new_[10535]_  | ~\new_[9237]_ ;
  assign \poc_o[22]  = \\u0_poc_reg[22] ;
  assign \new_[8853]_  = ~\new_[12454]_  | ~\new_[10514]_  | ~\new_[12585]_  | ~\new_[9413]_ ;
  assign \new_[8854]_  = ~\new_[10253]_  | ~\new_[11316]_  | ~\new_[9262]_  | ~\new_[10021]_ ;
  assign \new_[8855]_  = ~\new_[9236]_  | ~\new_[11051]_ ;
  assign \new_[8856]_  = ~\new_[9245]_  | ~\new_[10041]_ ;
  assign \new_[8857]_  = ~\new_[12089]_  | ~\new_[10252]_  | ~\new_[9262]_  | ~\new_[9562]_ ;
  assign \new_[8858]_  = ~\new_[9263]_  & (~\new_[11396]_  | ~\new_[11328]_ );
  assign \poc_o[25]  = \\u0_poc_reg[25] ;
  assign n5871 = \\u7_mc_dqm_r_reg[0] ;
  assign \new_[8861]_  = \new_[1463]_  ^ \new_[9460]_ ;
  assign \new_[8862]_  = ~u5_tmr_done_reg;
  assign \new_[8863]_  = ~\new_[9034]_ ;
  assign \new_[8864]_  = ~\new_[9268]_  | ~\new_[12544]_ ;
  assign \poc_o[23]  = \\u0_poc_reg[23] ;
  assign \new_[8866]_  = ~\new_[11914]_  | ~\new_[11259]_ ;
  assign \new_[8867]_  = \new_[9267]_  & \new_[12559]_ ;
  assign \new_[8868]_  = ~\new_[9095]_ ;
  assign \new_[8869]_  = ~\new_[10827]_  | ~\new_[12667]_  | ~\new_[11357]_  | ~\new_[11349]_ ;
  assign \new_[8870]_  = ~\new_[10205]_  | ~\new_[9269]_  | ~\new_[10519]_ ;
  assign \new_[8871]_  = ~\new_[9042]_ ;
  assign \new_[8872]_  = ~\new_[12312]_  | ~\new_[10531]_  | ~\new_[12316]_  | ~\new_[12318]_ ;
  assign \new_[8873]_  = ~\new_[9051]_ ;
  assign \new_[8874]_  = \new_[10698]_  & \new_[12667]_ ;
  assign \new_[8875]_  = ~\new_[9341]_  & ~\new_[9249]_ ;
  assign \new_[8876]_  = \new_[10722]_  & \new_[12667]_ ;
  assign \new_[8877]_  = \new_[12667]_  & \new_[11346]_ ;
  assign \poc_o[24]  = \\u0_poc_reg[24] ;
  assign \poc_o[26]  = \\u0_poc_reg[26] ;
  assign \new_[8880]_  = \new_[9355]_  & \new_[11357]_ ;
  assign \new_[8881]_  = \new_[9314]_  & \new_[11920]_ ;
  assign \new_[8882]_  = \new_[10572]_  & \new_[11332]_ ;
  assign \new_[8883]_  = \new_[10572]_  & \new_[9913]_ ;
  assign \new_[8884]_  = \new_[10572]_  & \new_[11340]_ ;
  assign \new_[8885]_  = \new_[10572]_  & \new_[9903]_ ;
  assign \poc_o[21]  = \\u0_poc_reg[21] ;
  assign \new_[8887]_  = \new_[10572]_  & \new_[10419]_ ;
  assign \new_[8888]_  = \new_[10572]_  & \new_[10411]_ ;
  assign \new_[8889]_  = \new_[10572]_  & \new_[10250]_ ;
  assign \new_[8890]_  = \new_[10572]_  & \new_[10827]_ ;
  assign \new_[8891]_  = ~\new_[9092]_ ;
  assign \new_[8892]_  = \new_[10572]_  & \new_[11337]_ ;
  assign \new_[8893]_  = \\u1_col_adr_reg[0] ;
  assign \new_[8894]_  = \new_[10572]_  & \new_[12093]_ ;
  assign \new_[8895]_  = ~\new_[9079]_ ;
  assign \new_[8896]_  = ~\new_[10846]_  | (~\new_[10148]_  & ~\new_[11361]_ );
  assign \new_[8897]_  = ~\new_[9137]_ ;
  assign \new_[8898]_  = ~\new_[9120]_ ;
  assign \new_[8899]_  = ~\new_[9123]_ ;
  assign \new_[8900]_  = ~\new_[9117]_ ;
  assign \new_[8901]_  = ~\new_[9090]_ ;
  assign \new_[8902]_  = ~\new_[9074]_ ;
  assign \new_[8903]_  = ~\new_[9093]_ ;
  assign \new_[8904]_  = ~\new_[9046]_ ;
  assign \new_[8905]_  = ~\new_[9089]_ ;
  assign \new_[8906]_  = ~\new_[9037]_ ;
  assign \new_[8907]_  = ~\new_[9098]_ ;
  assign \new_[8908]_  = ~\new_[9149]_ ;
  assign \new_[8909]_  = ~\new_[8987]_ ;
  assign \new_[8910]_  = ~\new_[9102]_ ;
  assign \poc_o[17]  = \\u0_poc_reg[17] ;
  assign \new_[8912]_  = ~\new_[11343]_  & ~\new_[10177]_ ;
  assign \new_[8913]_  = ~\new_[8197]_  & ~\new_[11338]_ ;
  assign \new_[8914]_  = ~\new_[10268]_  | ~\new_[11575]_ ;
  assign \poc_o[13]  = \\u0_poc_reg[13] ;
  assign n5786 = \\u7_mc_dqm_r_reg[2] ;
  assign \new_[8917]_  = ~\new_[12052]_  | ~\new_[9902]_ ;
  assign \new_[8918]_  = ~\new_[8197]_  & ~\new_[12094]_ ;
  assign \new_[8919]_  = ~\new_[10268]_  | ~\new_[10485]_ ;
  assign \new_[8920]_  = ~\new_[10268]_  & ~\new_[12274]_ ;
  assign \new_[8921]_  = \new_[10572]_  & \new_[10177]_ ;
  assign \new_[8922]_  = ~\new_[9091]_ ;
  assign \new_[8923]_  = ~\new_[9112]_ ;
  assign \poc_o[1]  = \\u0_poc_reg[1] ;
  assign \poc_o[28]  = \\u0_poc_reg[28] ;
  assign \new_[8926]_  = \new_[10572]_  & \new_[11316]_ ;
  assign \poc_o[11]  = \\u0_poc_reg[11] ;
  assign \poc_o[16]  = \\u0_poc_reg[16] ;
  assign \new_[8929]_  = ~\new_[9118]_ ;
  assign \new_[8930]_  = \new_[10572]_  & \new_[11356]_ ;
  assign \new_[8931]_  = ~\new_[9124]_ ;
  assign \poc_o[19]  = \\u0_poc_reg[19] ;
  assign \poc_o[10]  = \\u0_poc_reg[10] ;
  assign \poc_o[15]  = \\u0_poc_reg[15] ;
  assign \poc_o[18]  = \\u0_poc_reg[18] ;
  assign \poc_o[20]  = \\u0_poc_reg[20] ;
  assign \poc_o[9]  = \\u0_poc_reg[9] ;
  assign \poc_o[31]  = \\u0_poc_reg[31] ;
  assign \new_[8939]_  = \\u1_col_adr_reg[7] ;
  assign \new_[8940]_  = \\u1_col_adr_reg[5] ;
  assign n5711 = \\u7_mc_dqm_r_reg[3] ;
  assign n5891 = \\u7_mc_dqm_r_reg[1] ;
  assign \new_[8943]_  = ~\new_[9132]_ ;
  assign \poc_o[14]  = \\u0_poc_reg[14] ;
  assign \new_[8945]_  = ~\new_[9961]_  & ~\new_[9752]_ ;
  assign \poc_o[5]  = \\u0_poc_reg[5] ;
  assign \new_[8947]_  = ~\new_[9007]_ ;
  assign \poc_o[29]  = \\u0_poc_reg[29] ;
  assign \poc_o[27]  = \\u0_poc_reg[27] ;
  assign \new_[8950]_  = ~\new_[9238]_  | ~\new_[11131]_ ;
  assign \new_[8951]_  = \\u1_col_adr_reg[6] ;
  assign n4661 = \new_[9412]_  ? \new_[10221]_  : n5476;
  assign \new_[8953]_  = ~\new_[11363]_  | ~\new_[10575]_  | ~\new_[12585]_  | ~\new_[9882]_ ;
  assign n4521 = ~\new_[9026]_ ;
  assign \new_[8955]_  = ~\new_[9424]_  | ~\new_[9443]_  | ~\new_[9783]_ ;
  assign \new_[8956]_  = ~\new_[9454]_  | ~\new_[9439]_  | ~\new_[9779]_ ;
  assign \new_[8957]_  = ~\new_[12398]_ ;
  assign \new_[8958]_  = ~\new_[9441]_  | ~\new_[9448]_  | ~\new_[9782]_ ;
  assign \new_[8959]_  = ~\new_[9446]_  | ~\new_[9422]_  | ~\new_[9768]_ ;
  assign \poc_o[12]  = \\u0_poc_reg[12] ;
  assign \new_[8961]_  = ~\new_[9344]_  & ~\new_[9493]_ ;
  assign \poc_o[3]  = \\u0_poc_reg[3] ;
  assign \poc_o[2]  = \\u0_poc_reg[2] ;
  assign \poc_o[7]  = \\u0_poc_reg[7] ;
  assign \poc_o[8]  = \\u0_poc_reg[8] ;
  assign \new_[8966]_  = \\u1_col_adr_reg[2] ;
  assign \new_[8967]_  = ~\new_[9238]_  & ~\new_[10671]_ ;
  assign \poc_o[6]  = \\u0_poc_reg[6] ;
  assign \new_[8969]_  = \\u1_col_adr_reg[4] ;
  assign \new_[8970]_  = \new_[10213]_  | \new_[9205]_ ;
  assign \new_[8971]_  = \\u1_col_adr_reg[3] ;
  assign \new_[8972]_  = \new_[7281]_  ^ \new_[9399]_ ;
  assign \new_[8973]_  = \\u1_col_adr_reg[1] ;
  assign \poc_o[30]  = \\u0_poc_reg[30] ;
  assign \poc_o[4]  = \\u0_poc_reg[4] ;
  assign \new_[8976]_  = ~u0_init_ack_r_reg;
  assign \new_[8977]_  = ~\new_[9177]_ ;
  assign \new_[8978]_  = \new_[7265]_  ^ \new_[10176]_ ;
  assign \new_[8979]_  = ~\\u3_mc_data_o_reg[7] ;
  assign \new_[8980]_  = ~\new_[9835]_  & ~\new_[9493]_ ;
  assign \new_[8981]_  = ~\new_[9669]_  | ~\new_[1842]_ ;
  assign \new_[8982]_  = \new_[1464]_  ^ \new_[9949]_ ;
  assign \new_[8983]_  = ~\new_[9622]_  | ~\new_[10846]_ ;
  assign \new_[8984]_  = ~\\u3_mc_data_o_reg[24] ;
  assign \new_[8985]_  = ~\\u3_mc_data_o_reg[25] ;
  assign \new_[8986]_  = ~\\u3_mc_data_o_reg[9] ;
  assign \new_[8987]_  = ~\new_[9615]_  | ~\new_[10846]_ ;
  assign \new_[8988]_  = ~\new_[10105]_  & ~\new_[9493]_ ;
  assign \new_[8989]_  = ~\new_[9695]_  | ~\new_[1955]_ ;
  assign \new_[8990]_  = ~\new_[9583]_  & (~\new_[10103]_  | ~\new_[10415]_ );
  assign \new_[8991]_  = ~\new_[10141]_  | ~\new_[10365]_  | ~\new_[9762]_  | ~\new_[10357]_ ;
  assign \new_[8992]_  = ~\new_[9552]_  | ~\new_[9501]_ ;
  assign \new_[8993]_  = ~\new_[9520]_  | ~\new_[9545]_ ;
  assign \new_[8994]_  = ~\new_[9531]_  | ~\new_[9513]_ ;
  assign \new_[8995]_  = ~\new_[9550]_  | ~\new_[9544]_ ;
  assign \new_[8996]_  = ~\new_[9543]_  | ~\new_[9523]_ ;
  assign \new_[8997]_  = ~\new_[9539]_  | ~\new_[9540]_ ;
  assign \new_[8998]_  = ~\new_[9392]_  | ~\new_[9533]_ ;
  assign \new_[8999]_  = ~\new_[9511]_  | ~\new_[9506]_ ;
  assign \new_[9000]_  = ~\new_[9687]_  | ~\new_[9507]_ ;
  assign \new_[9001]_  = ~\new_[9529]_  | ~\new_[9527]_ ;
  assign \new_[9002]_  = ~\new_[9549]_  | ~\new_[9510]_ ;
  assign \new_[9003]_  = ~\new_[9532]_  | ~\new_[9512]_ ;
  assign \new_[9004]_  = ~\\u3_mc_data_o_reg[0] ;
  assign \new_[9005]_  = ~\new_[9515]_  | ~\new_[9667]_ ;
  assign n4691 = ~\new_[9624]_  & ~\new_[10041]_ ;
  assign \new_[9007]_  = ~n4946 & ~\new_[8976]_ ;
  assign \new_[9008]_  = ~\new_[9394]_  | ~\new_[9509]_ ;
  assign \new_[9009]_  = ~\new_[9522]_  | ~\new_[9505]_ ;
  assign \new_[9010]_  = ~\new_[9600]_  | ~\new_[9546]_ ;
  assign \new_[9011]_  = ~\new_[9636]_  | ~\new_[9541]_ ;
  assign \new_[9012]_  = ~\new_[9508]_  | ~\new_[9673]_ ;
  assign \new_[9013]_  = ~\new_[9677]_  | ~\new_[9547]_ ;
  assign \new_[9014]_  = ~\new_[9526]_  | ~\new_[9517]_ ;
  assign \new_[9015]_  = ~\new_[9553]_  | ~\new_[9521]_ ;
  assign \new_[9016]_  = ~\new_[9551]_  | ~\new_[11789]_ ;
  assign \new_[9017]_  = ~\new_[9514]_  | ~\new_[9555]_ ;
  assign \new_[9018]_  = ~\new_[9530]_  | ~\new_[9518]_ ;
  assign \new_[9019]_  = ~\new_[9504]_  | ~\new_[9537]_ ;
  assign \new_[9020]_  = ~\new_[9534]_  | ~\new_[9528]_ ;
  assign \new_[9021]_  = ~\new_[9542]_  | ~\new_[9538]_ ;
  assign \new_[9022]_  = ~\new_[9503]_  | ~\new_[9652]_ ;
  assign \new_[9023]_  = ~\new_[9524]_  | ~\new_[9500]_ ;
  assign \new_[9024]_  = ~\new_[9502]_  | ~\new_[9688]_ ;
  assign \new_[9025]_  = ~\new_[9535]_  | ~\new_[9536]_ ;
  assign \new_[9026]_  = \new_[9690]_  | \new_[10042]_ ;
  assign \new_[9027]_  = ~\\u3_mc_data_o_reg[20] ;
  assign \new_[9028]_  = ~\new_[11364]_  | ~\new_[10496]_  | ~\new_[12585]_  | ~\new_[9882]_ ;
  assign \new_[9029]_  = ~\\u3_mc_data_o_reg[3] ;
  assign \new_[9030]_  = ~\new_[11515]_  | ~\new_[10846]_ ;
  assign \new_[9031]_  = ~\new_[10009]_  | ~\new_[10488]_  | ~\new_[10300]_  | ~\new_[10445]_ ;
  assign \new_[9032]_  = \new_[10572]_  & \new_[10902]_ ;
  assign n4686 = \new_[11100]_  ^ \new_[9947]_ ;
  assign \new_[9034]_  = ~\new_[9592]_  | ~\new_[10846]_ ;
  assign \new_[9035]_  = ~\new_[10396]_  | ~\new_[10228]_  | ~\new_[9730]_ ;
  assign \new_[9036]_  = ~\\u3_mc_data_o_reg[26] ;
  assign \new_[9037]_  = ~\new_[9598]_  | ~\new_[10846]_ ;
  assign n4696 = \new_[9563]_  & \new_[10400]_ ;
  assign n4711 = \new_[9556]_  & \new_[10488]_ ;
  assign \new_[9040]_  = ~\new_[9294]_ ;
  assign \new_[9041]_  = ~\new_[10488]_  | ~\new_[11016]_  | ~\new_[10412]_  | ~\new_[10400]_ ;
  assign \new_[9042]_  = ~\new_[9587]_  | ~\new_[10846]_ ;
  assign \new_[9043]_  = ~\new_[11573]_  | ~\new_[11321]_  | ~\new_[10143]_  | ~\new_[10469]_ ;
  assign \new_[9044]_  = ~\new_[9216]_ ;
  assign \new_[9045]_  = ~\new_[10112]_  & ~\new_[9639]_ ;
  assign \new_[9046]_  = ~\new_[9585]_  | ~\new_[10846]_ ;
  assign \new_[9047]_  = \new_[10572]_  & \new_[12598]_ ;
  assign \new_[9048]_  = \new_[10572]_  & \new_[10291]_ ;
  assign \new_[9049]_  = ~\new_[9613]_  | ~\new_[10846]_ ;
  assign \new_[9050]_  = ~\\u3_mc_data_o_reg[16] ;
  assign \new_[9051]_  = ~\new_[9584]_  | ~\new_[10846]_ ;
  assign \new_[9052]_  = ~\\u3_mc_data_o_reg[1] ;
  assign n4706 = u5_suspended_reg;
  assign \new_[9054]_  = \new_[11356]_  & \new_[11351]_ ;
  assign \new_[9055]_  = \new_[10029]_  & \new_[10771]_ ;
  assign \new_[9056]_  = \new_[11338]_  & \new_[12731]_ ;
  assign \new_[9057]_  = \new_[10250]_  & \new_[12731]_ ;
  assign \new_[9058]_  = ~\new_[9376]_ ;
  assign \new_[9059]_  = ~\new_[10902]_  & ~\new_[11919]_ ;
  assign \new_[9060]_  = ~\new_[10018]_  | ~\new_[12337]_ ;
  assign \new_[9061]_  = ~\\u3_mc_data_o_reg[19] ;
  assign \new_[9062]_  = \new_[10572]_  & n5021;
  assign \new_[9063]_  = ~\new_[10529]_  & ~\new_[10747]_ ;
  assign \new_[9064]_  = \new_[10572]_  & \new_[11493]_ ;
  assign \new_[9065]_  = \new_[10572]_  & \new_[11343]_ ;
  assign \new_[9066]_  = \new_[10572]_  & \new_[12610]_ ;
  assign \new_[9067]_  = \new_[10572]_  & \new_[11363]_ ;
  assign \new_[9068]_  = \new_[10572]_  & \new_[10243]_ ;
  assign \new_[9069]_  = \new_[10572]_  & \new_[10919]_ ;
  assign \new_[9070]_  = \new_[10572]_  & \new_[11310]_ ;
  assign \new_[9071]_  = \new_[10572]_  & \new_[11320]_ ;
  assign \new_[9072]_  = \new_[10572]_  & \new_[12453]_ ;
  assign \new_[9073]_  = \new_[10572]_  & \new_[12755]_ ;
  assign \new_[9074]_  = ~\new_[9603]_  | ~\new_[10846]_ ;
  assign \new_[9075]_  = \new_[10572]_  & \new_[9946]_ ;
  assign \new_[9076]_  = ~\\u3_mc_data_o_reg[13] ;
  assign \new_[9077]_  = ~\new_[9365]_ ;
  assign \new_[9078]_  = ~\new_[9358]_ ;
  assign \new_[9079]_  = ~\new_[9489]_  | ~\new_[10846]_ ;
  assign \new_[9080]_  = ~\new_[9349]_ ;
  assign \new_[9081]_  = ~\new_[9285]_ ;
  assign \new_[9082]_  = ~\new_[9286]_ ;
  assign \new_[9083]_  = ~\new_[9329]_ ;
  assign \new_[9084]_  = ~\new_[9609]_  | ~\new_[10846]_ ;
  assign \new_[9085]_  = ~\new_[9287]_ ;
  assign \new_[9086]_  = \new_[10572]_  & \new_[11328]_ ;
  assign \new_[9087]_  = ~\new_[9378]_ ;
  assign \new_[9088]_  = ~\new_[9323]_ ;
  assign \new_[9089]_  = \new_[9591]_  & \new_[10846]_ ;
  assign \new_[9090]_  = ~\new_[9602]_  | ~\new_[10846]_ ;
  assign \new_[9091]_  = ~\new_[9601]_  | ~\new_[10846]_ ;
  assign \new_[9092]_  = \new_[9621]_  & \new_[10846]_ ;
  assign \new_[9093]_  = \new_[9589]_  & \new_[10846]_ ;
  assign \new_[9094]_  = ~\new_[9293]_ ;
  assign \new_[9095]_  = ~\new_[9593]_  | ~\new_[10846]_ ;
  assign \new_[9096]_  = ~\new_[12000]_  | ~\new_[10846]_ ;
  assign \new_[9097]_  = ~\new_[9295]_ ;
  assign \new_[9098]_  = ~\new_[9614]_  | ~\new_[10846]_ ;
  assign \new_[9099]_  = ~\new_[9192]_ ;
  assign \new_[9100]_  = ~\\u3_mc_data_o_reg[18] ;
  assign \new_[9101]_  = ~\new_[9616]_  | ~\new_[10846]_ ;
  assign \new_[9102]_  = \new_[9663]_  & \new_[10846]_ ;
  assign \new_[9103]_  = u5_pack_le1_reg;
  assign \new_[9104]_  = ~\new_[9954]_ ;
  assign n4701 = ~\new_[9685]_  | ~\new_[9988]_ ;
  assign \new_[9106]_  = ~\\u3_mc_data_o_reg[29] ;
  assign \new_[9107]_  = ~\new_[9305]_ ;
  assign \new_[9108]_  = ~\new_[9924]_ ;
  assign \new_[9109]_  = ~\new_[9714]_ ;
  assign \new_[9110]_  = ~\new_[8197]_  & ~\new_[10676]_ ;
  assign \new_[9111]_  = ~\new_[1433]_  | ~\new_[11341]_ ;
  assign \new_[9112]_  = ~\new_[11521]_  | ~\new_[10846]_ ;
  assign \new_[9113]_  = ~\new_[9292]_ ;
  assign \new_[9114]_  = ~\new_[9290]_ ;
  assign \new_[9115]_  = ~\new_[9321]_ ;
  assign \new_[9116]_  = ~\\u3_mc_data_o_reg[15] ;
  assign \new_[9117]_  = \new_[9581]_  & \new_[10846]_ ;
  assign \new_[9118]_  = \new_[9596]_  & \new_[10846]_ ;
  assign \new_[9119]_  = ~\\u3_mc_data_o_reg[10] ;
  assign \new_[9120]_  = ~\new_[9612]_  | ~\new_[10846]_ ;
  assign \new_[9121]_  = u5_burst_act_rd_reg;
  assign \new_[9122]_  = ~\new_[9324]_ ;
  assign \new_[9123]_  = \new_[9586]_  & \new_[10846]_ ;
  assign \new_[9124]_  = ~\new_[9408]_  | ~\new_[10846]_ ;
  assign \new_[9125]_  = ~\new_[9330]_ ;
  assign \new_[9126]_  = \new_[7966]_  ^ \new_[9722]_ ;
  assign \new_[9127]_  = ~\\u3_mc_data_o_reg[11] ;
  assign \new_[9128]_  = ~\\u3_mc_data_o_reg[21] ;
  assign \new_[9129]_  = ~\\u3_mc_data_o_reg[27] ;
  assign \new_[9130]_  = ~\\u3_mc_data_o_reg[31] ;
  assign \new_[9131]_  = ~\new_[9666]_  | ~\new_[9525]_ ;
  assign \new_[9132]_  = ~\new_[9678]_  | ~\new_[10846]_ ;
  assign \new_[9133]_  = ~\new_[9338]_ ;
  assign \new_[9134]_  = ~\new_[10488]_  | (~\new_[11258]_  & ~\new_[11361]_ );
  assign \new_[9135]_  = ~\\u3_mc_data_o_reg[28] ;
  assign \new_[9136]_  = \\u0_spec_req_cs_reg[1] ;
  assign \new_[9137]_  = ~\new_[9588]_  | ~\new_[10846]_ ;
  assign \new_[9138]_  = ~\\u3_mc_data_o_reg[22] ;
  assign \new_[9139]_  = ~\new_[9346]_ ;
  assign \new_[9140]_  = ~\new_[10516]_  | ~\new_[12441]_  | ~\new_[10016]_  | ~\new_[10240]_ ;
  assign \new_[9141]_  = \new_[10572]_  & \new_[10743]_ ;
  assign \new_[9142]_  = \new_[12400]_  & \new_[11351]_ ;
  assign \new_[9143]_  = ~\\u3_mc_data_o_reg[5] ;
  assign \new_[9144]_  = ~\new_[8197]_  & ~\new_[10872]_ ;
  assign \new_[9145]_  = \new_[10975]_  ^ \new_[9726]_ ;
  assign \new_[9146]_  = \new_[12399]_  & \new_[11351]_ ;
  assign \new_[9147]_  = ~\\u3_mc_data_o_reg[17] ;
  assign \new_[9148]_  = ~\\u3_mc_data_o_reg[30] ;
  assign \new_[9149]_  = ~\new_[9393]_  | ~\new_[10846]_ ;
  assign \new_[9150]_  = ~\\u3_mc_data_o_reg[14] ;
  assign \new_[9151]_  = \new_[7977]_  ^ \new_[9727]_ ;
  assign \new_[9152]_  = ~\\u3_mc_data_o_reg[6] ;
  assign \new_[9153]_  = \\u1_u0_out_r_reg[3] ;
  assign \new_[9154]_  = ~\\u3_mc_data_o_reg[8] ;
  assign \new_[9155]_  = ~\\u3_mc_data_o_reg[23] ;
  assign \new_[9156]_  = ~\new_[10671]_  & ~\new_[9494]_ ;
  assign \new_[9157]_  = ~\new_[9516]_  | ~\new_[9698]_ ;
  assign \new_[9158]_  = ~\new_[9548]_  | ~\new_[9708]_ ;
  assign \new_[9159]_  = ~\new_[12306]_  | ~\new_[10846]_ ;
  assign \new_[9160]_  = \new_[10572]_  & \new_[10802]_ ;
  assign \new_[9161]_  = ~\new_[9493]_  | ~\new_[8077]_ ;
  assign \new_[9162]_  = ~\new_[9554]_  | ~\new_[9519]_ ;
  assign \new_[9163]_  = \new_[2137]_  ^ \new_[9711]_ ;
  assign \new_[9164]_  = \new_[11209]_  ^ \new_[9721]_ ;
  assign \new_[9165]_  = \new_[10572]_  & \new_[12054]_ ;
  assign \new_[9166]_  = ~\\u3_mc_data_o_reg[12] ;
  assign \new_[9167]_  = ~\\u3_mc_data_o_reg[4] ;
  assign \new_[9168]_  = ~\new_[9742]_ ;
  assign \new_[9169]_  = \new_[10572]_  & \new_[10526]_ ;
  assign \new_[9170]_  = \new_[9404]_  & \new_[10940]_ ;
  assign \new_[9171]_  = ~\\u3_mc_data_o_reg[2] ;
  assign n4716 = \new_[10820]_  ^ \new_[9890]_ ;
  assign \new_[9173]_  = \new_[10303]_  & \new_[9890]_ ;
  assign n4901 = \new_[10833]_  ? \new_[10132]_  : \poc_o[7] ;
  assign \new_[9175]_  = \new_[9934]_  & \new_[10381]_ ;
  assign \new_[9176]_  = \\u1_sram_addr_reg[5] ;
  assign \new_[9177]_  = ~\new_[10154]_  | ~\new_[10496]_ ;
  assign \new_[9178]_  = ~\new_[9608]_ ;
  assign \new_[9179]_  = \\u1_sram_addr_reg[6] ;
  assign n4726 = \new_[10843]_  ? \new_[10132]_  : \poc_o[22] ;
  assign n4836 = \new_[10935]_  ? \new_[10132]_  : \poc_o[31] ;
  assign n4866 = \new_[10852]_  ? \new_[10132]_  : \poc_o[5] ;
  assign n4896 = \new_[10968]_  ? \new_[10132]_  : \poc_o[2] ;
  assign \new_[9184]_  = \\u1_sram_addr_reg[18] ;
  assign n4791 = \new_[10835]_  ? \new_[10132]_  : \poc_o[28] ;
  assign \new_[9186]_  = \new_[7278]_  ^ \new_[10095]_ ;
  assign \new_[9187]_  = \new_[8075]_  ^ \new_[10066]_ ;
  assign \new_[9188]_  = \new_[10572]_  & \new_[10808]_ ;
  assign n4771 = \new_[10860]_  ? \new_[10132]_  : \poc_o[17] ;
  assign \new_[9190]_  = ~\new_[9620]_ ;
  assign \new_[9191]_  = ~\new_[11779]_ ;
  assign \new_[9192]_  = ~\new_[9929]_  | ~\new_[10846]_ ;
  assign \new_[9193]_  = ~\new_[10363]_  | ~\new_[10379]_  | ~\new_[9755]_  | ~\new_[10377]_ ;
  assign \new_[9194]_  = ~\new_[10366]_  | ~\new_[10384]_  | ~\new_[9765]_  | ~\new_[10362]_ ;
  assign \new_[9195]_  = ~\new_[10382]_  | ~\new_[10385]_  | ~\new_[9763]_  | ~\new_[10380]_ ;
  assign \new_[9196]_  = ~\new_[10295]_  | ~\new_[10375]_  | ~\new_[9764]_  | ~\new_[10372]_ ;
  assign n4746 = \new_[10814]_  ? \new_[10132]_  : \poc_o[23] ;
  assign \new_[9198]_  = ~\new_[10376]_  | ~\new_[10387]_  | ~\new_[9776]_  | ~\new_[10315]_ ;
  assign \new_[9199]_  = ~\new_[10069]_  | ~\new_[9811]_ ;
  assign n4816 = \new_[10896]_  ? \new_[10132]_  : \poc_o[15] ;
  assign \new_[9201]_  = ~\new_[12094]_  & ~\new_[9752]_ ;
  assign \new_[9202]_  = \new_[9951]_  & \new_[12094]_ ;
  assign n4811 = \new_[10885]_  ? \new_[10132]_  : \poc_o[10] ;
  assign \new_[9204]_  = ~\new_[9716]_  & (~\new_[10162]_  | ~\new_[2056]_ );
  assign \new_[9205]_  = ~\new_[12337]_ ;
  assign \new_[9206]_  = (~\new_[10116]_  | ~\new_[8179]_ ) & (~\new_[10236]_  | ~\poc_o[1] );
  assign \new_[9207]_  = \\u1_sram_addr_reg[20] ;
  assign \new_[9208]_  = (~\new_[10116]_  | ~\new_[8194]_ ) & (~\new_[10236]_  | ~\poc_o[9] );
  assign \new_[9209]_  = (~\new_[10116]_  | ~\new_[8195]_ ) & (~\new_[8399]_  | ~\new_[10249]_ );
  assign \new_[9210]_  = (~\new_[10116]_  | ~\new_[8199]_ ) & (~\new_[10236]_  | ~\poc_o[5] );
  assign \new_[9211]_  = u5_ir_cnt_done_reg;
  assign \new_[9212]_  = (~\new_[10116]_  | ~\new_[8198]_ ) & (~\new_[10236]_  | ~\poc_o[4] );
  assign \new_[9213]_  = (~\new_[10116]_  | ~\new_[8205]_ ) & (~\new_[8382]_  | ~\new_[10249]_ );
  assign \new_[9214]_  = (~\new_[10116]_  | ~\new_[8229]_ ) & (~\new_[10236]_  | ~\poc_o[3] );
  assign \new_[9215]_  = (~\new_[10116]_  | ~\new_[8149]_ ) & (~\new_[10439]_  | ~\new_[10249]_ );
  assign \new_[9216]_  = ~\new_[11311]_  | ~\new_[10211]_  | ~\new_[10346]_  | ~\new_[12611]_ ;
  assign \new_[9217]_  = (~\new_[10116]_  | ~\new_[8200]_ ) & (~\new_[10236]_  | ~\poc_o[6] );
  assign \new_[9218]_  = (~\new_[10116]_  | ~\new_[8196]_ ) & (~\new_[10236]_  | ~\poc_o[2] );
  assign \new_[9219]_  = (~\new_[10116]_  | ~\new_[8201]_ ) & (~\new_[11126]_  | ~\new_[10249]_ );
  assign n4731 = \new_[10923]_  ? \new_[10132]_  : \poc_o[25] ;
  assign n4936 = \new_[10947]_  ? \new_[10132]_  : \poc_o[30] ;
  assign n4876 = \new_[10879]_  ? \new_[10132]_  : \poc_o[27] ;
  assign n4786 = \new_[10844]_  ? \new_[10132]_  : \poc_o[1] ;
  assign n4806 = \new_[10847]_  ? \new_[10132]_  : \poc_o[19] ;
  assign n4721 = \new_[10845]_  ? \new_[10132]_  : \poc_o[0] ;
  assign n4831 = \new_[10908]_  ? \new_[10132]_  : \poc_o[9] ;
  assign \new_[9227]_  = ~\new_[9728]_  | (~\new_[10227]_  & ~\new_[10447]_ );
  assign n4861 = \new_[10828]_  ? \new_[10132]_  : \poc_o[14] ;
  assign n4941 = \new_[10869]_  ? \new_[10132]_  : \poc_o[4] ;
  assign n4776 = \new_[10825]_  ? \new_[10132]_  : \poc_o[13] ;
  assign n4821 = \new_[10868]_  ? \new_[10132]_  : \poc_o[18] ;
  assign n4796 = \new_[10878]_  ? \new_[10132]_  : \poc_o[11] ;
  assign n4891 = \new_[10916]_  ? \new_[10132]_  : \poc_o[3] ;
  assign n4916 = \new_[10819]_  ? \new_[10132]_  : \poc_o[6] ;
  assign \new_[9235]_  = ~\new_[9790]_  | (~\new_[10269]_  & ~\new_[10447]_ );
  assign \new_[9236]_  = ~\new_[11131]_  | ~\new_[10683]_  | ~\new_[9852]_  | ~\new_[10820]_ ;
  assign \new_[9237]_  = ~\new_[9493]_ ;
  assign \new_[9238]_  = ~\new_[11100]_  | ~\new_[11202]_  | ~\new_[9959]_  | ~\new_[10836]_ ;
  assign \new_[9239]_  = ~\new_[9575]_ ;
  assign \new_[9240]_  = ~\new_[9971]_  | ~\new_[9962]_ ;
  assign \new_[9241]_  = \new_[10572]_  & \new_[10838]_ ;
  assign \new_[9242]_  = ~\new_[10134]_  | ~\new_[9886]_ ;
  assign \new_[9243]_  = ~\new_[10027]_  | ~\new_[9884]_ ;
  assign \new_[9244]_  = ~\new_[10149]_  | ~\new_[9812]_ ;
  assign \new_[9245]_  = ~\new_[9624]_ ;
  assign \new_[9246]_  = ~\new_[9982]_  | ~\new_[9751]_ ;
  assign \new_[9247]_  = ~\new_[10025]_  | ~\new_[9809]_ ;
  assign \new_[9248]_  = ~\new_[9810]_  & (~\new_[11178]_  | ~\new_[10502]_ );
  assign \new_[9249]_  = ~\new_[10767]_  | ~\new_[10157]_  | ~\new_[10724]_ ;
  assign n4926 = \wb_addr_i[5]  ? \new_[10125]_  : \new_[8971]_ ;
  assign n4921 = \wb_addr_i[6]  ? \new_[10125]_  : \new_[8969]_ ;
  assign n4841 = \wb_addr_i[9]  ? \new_[10125]_  : \new_[8939]_ ;
  assign n4881 = \wb_addr_i[8]  ? \new_[10125]_  : \new_[8951]_ ;
  assign n4911 = \wb_addr_i[4]  ? \new_[10125]_  : \new_[8966]_ ;
  assign \new_[9255]_  = ~\new_[9690]_ ;
  assign n4766 = \wb_addr_i[2]  ? \new_[10125]_  : \new_[8893]_ ;
  assign \new_[9257]_  = \\u1_sram_addr_reg[21] ;
  assign n4931 = \wb_addr_i[3]  ? \new_[10125]_  : \new_[8973]_ ;
  assign n4761 = \new_[10832]_  ? \new_[10132]_  : \poc_o[21] ;
  assign \new_[9260]_  = ~\new_[11833]_  & ~\new_[9942]_ ;
  assign \new_[9261]_  = ~\new_[11252]_  & ~\new_[11919]_ ;
  assign \new_[9262]_  = ~\new_[12719]_  & ~\new_[9752]_ ;
  assign \new_[9263]_  = ~\new_[10503]_  & ~\new_[12732]_ ;
  assign n4736 = n5871 ? \new_[10488]_  : \wb_sel_i[0] ;
  assign \new_[9265]_  = ~\new_[9951]_  | ~\new_[10301]_ ;
  assign \new_[9266]_  = ~\new_[10692]_  & ~\new_[12730]_ ;
  assign \new_[9267]_  = ~\new_[9883]_  & ~\new_[10286]_ ;
  assign \new_[9268]_  = ~\new_[12594]_ ;
  assign \new_[9269]_  = ~\new_[9639]_ ;
  assign \new_[9270]_  = ~\new_[10144]_  | ~\new_[9808]_ ;
  assign n4856 = n5891 ? \new_[10488]_  : \wb_sel_i[1] ;
  assign \new_[9272]_  = \new_[1581]_  ^ \new_[9981]_ ;
  assign \new_[9273]_  = \new_[10572]_  & \new_[10955]_ ;
  assign \new_[9274]_  = \new_[10572]_  & \new_[11367]_ ;
  assign \new_[9275]_  = \new_[10572]_  & \new_[9997]_ ;
  assign \new_[9276]_  = \new_[10572]_  & \new_[10960]_ ;
  assign \new_[9277]_  = \new_[10572]_  & \new_[11576]_ ;
  assign \new_[9278]_  = \new_[10572]_  & \new_[11526]_ ;
  assign \new_[9279]_  = \new_[10572]_  & \new_[11355]_ ;
  assign \new_[9280]_  = \new_[10572]_  & \new_[12567]_ ;
  assign \new_[9281]_  = \new_[10572]_  & \new_[11348]_ ;
  assign \new_[9282]_  = \new_[10572]_  & \new_[10933]_ ;
  assign n4906 = \new_[10817]_  ? \new_[10132]_  : \poc_o[8] ;
  assign \new_[9284]_  = ~\new_[10529]_  & ~\new_[11334]_ ;
  assign \new_[9285]_  = \new_[9864]_  & \new_[10846]_ ;
  assign \new_[9286]_  = ~\new_[12293]_  | ~\new_[10846]_ ;
  assign \new_[9287]_  = ~\new_[9857]_  | ~\new_[10846]_ ;
  assign \new_[9288]_  = ~\new_[9640]_ ;
  assign \new_[9289]_  = ~\new_[9577]_ ;
  assign \new_[9290]_  = ~\new_[9937]_  | ~\new_[10846]_ ;
  assign \new_[9291]_  = ~\new_[9746]_  | ~\new_[10846]_ ;
  assign \new_[9292]_  = \new_[9862]_  & \new_[10846]_ ;
  assign \new_[9293]_  = \new_[9840]_  & \new_[10846]_ ;
  assign \new_[9294]_  = \new_[9850]_  & \new_[10846]_ ;
  assign \new_[9295]_  = \new_[9824]_  & \new_[10846]_ ;
  assign \new_[9296]_  = ~\new_[9844]_  | ~\new_[10846]_ ;
  assign \new_[9297]_  = \new_[11012]_  ^ \new_[11320]_ ;
  assign \new_[9298]_  = ~\new_[9579]_ ;
  assign \new_[9299]_  = \new_[9914]_  & \new_[10724]_ ;
  assign \new_[9300]_  = \new_[10572]_  & \new_[10818]_ ;
  assign n4781 = n5786 ? \new_[10488]_  : \wb_sel_i[2] ;
  assign \new_[9302]_  = ~\new_[9591]_ ;
  assign \new_[9303]_  = ~\new_[9668]_ ;
  assign \new_[9304]_  = ~\new_[9657]_ ;
  assign \new_[9305]_  = ~\new_[10517]_  | ~\new_[10250]_ ;
  assign \new_[9306]_  = \\u1_sram_addr_reg[23] ;
  assign \new_[9307]_  = ~\new_[9659]_ ;
  assign \new_[9308]_  = ~\new_[9848]_ ;
  assign \new_[9309]_  = ~\new_[11045]_  | ~\new_[11321]_ ;
  assign n4851 = n5711 ? \new_[10488]_  : \wb_sel_i[3] ;
  assign \new_[9311]_  = \new_[12667]_  & \new_[11343]_ ;
  assign \new_[9312]_  = ~\new_[8197]_  & ~\new_[11329]_ ;
  assign n4756 = \new_[10939]_  ? \new_[10132]_  : \poc_o[26] ;
  assign \new_[9314]_  = ~\new_[12044]_  & ~\new_[10509]_ ;
  assign \new_[9315]_  = ~\new_[12577]_  | ~\new_[10658]_ ;
  assign \new_[9316]_  = ~\new_[12577]_  | ~\new_[10749]_ ;
  assign \new_[9317]_  = ~\new_[8197]_  & ~\new_[12052]_ ;
  assign \new_[9318]_  = ~\new_[9946]_  & ~\new_[10960]_ ;
  assign \new_[9319]_  = ~\new_[8197]_  & ~\new_[12401]_ ;
  assign \new_[9320]_  = ~\new_[8197]_  & ~\new_[10897]_ ;
  assign \new_[9321]_  = \new_[9865]_  & \new_[10846]_ ;
  assign \new_[9322]_  = ~\new_[9938]_  | ~\new_[10846]_ ;
  assign \new_[9323]_  = \new_[9863]_  & \new_[10846]_ ;
  assign \new_[9324]_  = \new_[9842]_  & \new_[10846]_ ;
  assign \new_[9325]_  = ~\new_[9646]_ ;
  assign \new_[9326]_  = ~\new_[9691]_ ;
  assign \new_[9327]_  = ~\new_[9649]_ ;
  assign \new_[9328]_  = \new_[10572]_  & \new_[10634]_ ;
  assign \new_[9329]_  = \new_[9906]_  & \new_[10846]_ ;
  assign \new_[9330]_  = \new_[9933]_  & \new_[10846]_ ;
  assign \new_[9331]_  = \\u1_sram_addr_reg[11] ;
  assign \new_[9332]_  = \\u1_sram_addr_reg[2] ;
  assign \new_[9333]_  = \\u1_sram_addr_reg[10] ;
  assign \new_[9334]_  = \\u1_sram_addr_reg[0] ;
  assign \new_[9335]_  = \\u1_sram_addr_reg[16] ;
  assign \new_[9336]_  = ~\new_[10009]_  | (~\new_[10412]_  & ~\new_[10481]_ );
  assign \new_[9337]_  = \\u1_sram_addr_reg[8] ;
  assign \new_[9338]_  = \new_[9837]_  & \new_[10846]_ ;
  assign \new_[9339]_  = \\u1_sram_addr_reg[3] ;
  assign \new_[9340]_  = ~\new_[9590]_ ;
  assign \new_[9341]_  = ~\new_[10551]_  | ~\new_[10383]_  | ~\new_[10397]_ ;
  assign \new_[9342]_  = \\u1_sram_addr_reg[13] ;
  assign \new_[9343]_  = ~\new_[9940]_  & (~\new_[10280]_  | ~\new_[1712]_ );
  assign \new_[9344]_  = \new_[8049]_  ^ \new_[9999]_ ;
  assign \new_[9345]_  = ~\new_[9958]_ ;
  assign \new_[9346]_  = \new_[11928]_  & \new_[10846]_ ;
  assign \new_[9347]_  = \\u1_sram_addr_reg[7] ;
  assign \new_[9348]_  = \new_[10572]_  & \new_[11361]_ ;
  assign \new_[9349]_  = \new_[10846]_  & \new_[9874]_ ;
  assign \new_[9350]_  = \\u1_sram_addr_reg[15] ;
  assign \new_[9351]_  = \\u1_sram_addr_reg[14] ;
  assign n4751 = \new_[10942]_  ? \new_[10132]_  : \poc_o[24] ;
  assign \new_[9353]_  = ~\new_[10321]_  | ~\new_[10272]_  | ~\new_[9756]_  | ~\new_[10281]_ ;
  assign \new_[9354]_  = \\u1_sram_addr_reg[1] ;
  assign \new_[9355]_  = ~\new_[10827]_  & ~\new_[12273]_ ;
  assign n4846 = \wb_addr_i[7]  ? \new_[10125]_  : \new_[8940]_ ;
  assign \new_[9357]_  = ~\new_[10108]_  & ~\new_[11298]_ ;
  assign \new_[9358]_  = \new_[9855]_  & \new_[10846]_ ;
  assign n4741 = \new_[9716]_  & \new_[10926]_ ;
  assign n4801 = \new_[10943]_  ? \new_[10132]_  : \poc_o[16] ;
  assign \new_[9361]_  = ~\new_[12523]_ ;
  assign \new_[9362]_  = \\u1_sram_addr_reg[12] ;
  assign \new_[9363]_  = \new_[1579]_  ^ \new_[10090]_ ;
  assign \new_[9364]_  = \\u1_sram_addr_reg[4] ;
  assign \new_[9365]_  = ~\new_[9960]_  | ~\new_[10846]_ ;
  assign \new_[9366]_  = \\u1_sram_addr_reg[19] ;
  assign \new_[9367]_  = \new_[9959]_  & \new_[10361]_ ;
  assign n4871 = \new_[10867]_  ? \new_[10132]_  : \poc_o[29] ;
  assign \new_[9369]_  = \\u1_sram_addr_reg[22] ;
  assign \new_[9370]_  = ~\new_[9791]_  | ~\new_[7382]_ ;
  assign \new_[9371]_  = ~\new_[8197]_  & ~\new_[11311]_ ;
  assign \new_[9372]_  = ~\new_[9391]_ ;
  assign \new_[9373]_  = \\u1_sram_addr_reg[17] ;
  assign \new_[9374]_  = ~\new_[9717]_ ;
  assign \new_[9375]_  = ~\new_[12577]_  | ~\new_[12177]_ ;
  assign \new_[9376]_  = \new_[9701]_ ;
  assign n4826 = \new_[10972]_  ? \new_[10132]_  : \poc_o[20] ;
  assign \new_[9378]_  = \new_[9818]_  & \new_[10846]_ ;
  assign \new_[9379]_  = ~\new_[10809]_ ;
  assign \new_[9380]_  = \\u1_sram_addr_reg[9] ;
  assign n4886 = \new_[10901]_  ? \new_[10132]_  : \poc_o[12] ;
  assign \new_[9382]_  = ~\new_[9789]_  & (~\new_[10273]_  | ~\new_[10448]_ );
  assign \new_[9383]_  = ~\new_[12003]_ ;
  assign \new_[9384]_  = ~\new_[10294]_  | ~\new_[10373]_  | ~\new_[10147]_ ;
  assign \new_[9385]_  = \new_[1580]_  ^ \new_[10260]_ ;
  assign n5046 = \wb_data_i[11]  ? \new_[10221]_  : n5556;
  assign \new_[9387]_  = (~\new_[10995]_  | ~\new_[10186]_ ) & (~\new_[7812]_  | ~\new_[10245]_ );
  assign \new_[9388]_  = ~\new_[9861]_ ;
  assign \new_[9389]_  = ~\new_[9739]_ ;
  assign \new_[9390]_  = \new_[10572]_  & \new_[11313]_ ;
  assign \new_[9391]_  = ~\new_[9715]_ ;
  assign \new_[9392]_  = (~\new_[11792]_  | ~\new_[4382]_ ) & (~\new_[12670]_  | ~\new_[4355]_ );
  assign \new_[9393]_  = ~\new_[10088]_  & ~\new_[10715]_ ;
  assign \new_[9394]_  = (~\new_[11792]_  | ~\new_[4370]_ ) & (~\new_[12670]_  | ~\new_[4345]_ );
  assign n5106 = \new_[10710]_  ^ \new_[10175]_ ;
  assign \new_[9396]_  = ~\new_[10036]_  & ~\new_[10213]_ ;
  assign \new_[9397]_  = ~\new_[10033]_  | ~\new_[10076]_ ;
  assign \new_[9398]_  = (~\new_[8052]_  | ~\new_[10242]_ ) & (~\new_[7619]_  | ~\new_[10188]_ );
  assign \new_[9399]_  = ~\new_[10918]_  | ~\new_[10028]_  | ~\new_[10708]_ ;
  assign \new_[9400]_  = \new_[2138]_  ^ \new_[10170]_ ;
  assign \new_[9401]_  = ~\new_[9718]_ ;
  assign \new_[9402]_  = (~\new_[7761]_  | ~\new_[10188]_ ) & (~\new_[8296]_  | ~\new_[10249]_ );
  assign \new_[9403]_  = ~\new_[11946]_  | ~wb_cyc_i;
  assign \new_[9404]_  = ~\new_[10114]_  & ~\new_[1955]_ ;
  assign \new_[9405]_  = \new_[10079]_  & \new_[11526]_ ;
  assign \new_[9406]_  = \new_[10786]_  & \new_[9992]_ ;
  assign \new_[9407]_  = ~\new_[9732]_ ;
  assign \new_[9408]_  = ~\new_[10088]_  & ~\new_[10771]_ ;
  assign \new_[9409]_  = \new_[1796]_  ^ \new_[10225]_ ;
  assign \new_[9410]_  = \new_[10182]_  ^ \new_[10178]_ ;
  assign \new_[9411]_  = \new_[10179]_  ^ \new_[10184]_ ;
  assign \new_[9412]_  = \new_[10181]_  ^ \new_[10183]_ ;
  assign \new_[9413]_  = \new_[10253]_  & \new_[10411]_ ;
  assign \new_[9414]_  = \new_[10180]_  ^ \new_[10185]_ ;
  assign \new_[9415]_  = ~\new_[9993]_  | ~\new_[10077]_ ;
  assign \new_[9416]_  = ~\new_[10032]_  | ~\new_[10038]_ ;
  assign \new_[9417]_  = \new_[7275]_  ^ \new_[10266]_ ;
  assign \new_[9418]_  = ~\new_[9924]_ ;
  assign \new_[9419]_  = \new_[1582]_  ^ \new_[10193]_ ;
  assign n5071 = ~\new_[10058]_  | (~\new_[8185]_  & ~\new_[11141]_ );
  assign \new_[9421]_  = (~\new_[7606]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[13] );
  assign \new_[9422]_  = (~\new_[11007]_  | ~\new_[10186]_ ) & (~\new_[7694]_  | ~\new_[10245]_ );
  assign \new_[9423]_  = (~\new_[8061]_  | ~\new_[10242]_ ) & (~\new_[10188]_  | ~\new_[7618]_ );
  assign \new_[9424]_  = (~\new_[7621]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[22] );
  assign \new_[9425]_  = (~\new_[7942]_  | ~\new_[10186]_ ) & (~\new_[11036]_  | ~\new_[10245]_ );
  assign \new_[9426]_  = (~\new_[7944]_  | ~\new_[10186]_ ) & (~\new_[11186]_  | ~\new_[10245]_ );
  assign \new_[9427]_  = (~\new_[10242]_  | ~\new_[8043]_ ) & (~\new_[10188]_  | ~\new_[7624]_ );
  assign \new_[9428]_  = (~\new_[8067]_  | ~\new_[10242]_ ) & (~\new_[10188]_  | ~\new_[7732]_ );
  assign \new_[9429]_  = (~\new_[8063]_  | ~\new_[10242]_ ) & (~\new_[10188]_  | ~\new_[7382]_ );
  assign \new_[9430]_  = (~\new_[11046]_  | ~\new_[10186]_ ) & (~\new_[7730]_  | ~\new_[10245]_ );
  assign \new_[9431]_  = (~\new_[7938]_  | ~\new_[10186]_ ) & (~\new_[7716]_  | ~\new_[10245]_ );
  assign \new_[9432]_  = (~\new_[8051]_  | ~\new_[10242]_ ) & (~\new_[7625]_  | ~\new_[10188]_ );
  assign \new_[9433]_  = (~\new_[7971]_  | ~\new_[10186]_ ) & (~\new_[11092]_  | ~\new_[10245]_ );
  assign \new_[9434]_  = (~\new_[7983]_  | ~\new_[10186]_ ) & (~\new_[10245]_  | ~\new_[7813]_ );
  assign \new_[9435]_  = (~\new_[7945]_  | ~\new_[10186]_ ) & (~\new_[7722]_  | ~\new_[10245]_ );
  assign \new_[9436]_  = (~\new_[7974]_  | ~\new_[10186]_ ) & (~\new_[7733]_  | ~\new_[10245]_ );
  assign \new_[9437]_  = (~\new_[7601]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[18] );
  assign \new_[9438]_  = (~\new_[7919]_  | ~\new_[10186]_ ) & (~\new_[11088]_  | ~\new_[10245]_ );
  assign \new_[9439]_  = (~\new_[11018]_  | ~\new_[10186]_ ) & (~\new_[11166]_  | ~\new_[10245]_ );
  assign \new_[9440]_  = (~\new_[7720]_  | ~\new_[10188]_ ) & (~\new_[8378]_  | ~\new_[10249]_ );
  assign \new_[9441]_  = (~\new_[7607]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[14] );
  assign \new_[9442]_  = (~\new_[7734]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[23] );
  assign \new_[9443]_  = (~\new_[10980]_  | ~\new_[10186]_ ) & (~\new_[7738]_  | ~\new_[10245]_ );
  assign \new_[9444]_  = (~\new_[7697]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[21] );
  assign \new_[9445]_  = (~\new_[7975]_  | ~\new_[10186]_ ) & (~\new_[7951]_  | ~\new_[10245]_ );
  assign \new_[9446]_  = (~\new_[7598]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[16] );
  assign \new_[9447]_  = (~\new_[11134]_  | ~\new_[10186]_ ) & (~\new_[11175]_  | ~\new_[10245]_ );
  assign \new_[9448]_  = (~\new_[11127]_  | ~\new_[10186]_ ) & (~\new_[11156]_  | ~\new_[10245]_ );
  assign \new_[9449]_  = (~\new_[7729]_  | ~\new_[10188]_ ) & (~\new_[8260]_  | ~\new_[10249]_ );
  assign \new_[9450]_  = (~\new_[8068]_  | ~\new_[10242]_ ) & (~\new_[7595]_  | ~\new_[10188]_ );
  assign \new_[9451]_  = (~\new_[7937]_  | ~\new_[10186]_ ) & (~\new_[10245]_  | ~\new_[7851]_ );
  assign \new_[9452]_  = (~\new_[8023]_  | ~\new_[10242]_ ) & (~\new_[7623]_  | ~\new_[10188]_ );
  assign \new_[9453]_  = (~\new_[11056]_  | ~\new_[10186]_ ) & (~\new_[11247]_  | ~\new_[10245]_ );
  assign \new_[9454]_  = (~\new_[7612]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[11] );
  assign \new_[9455]_  = (~\new_[8072]_  | ~\new_[10242]_ ) & (~\new_[7715]_  | ~\new_[10188]_ );
  assign \new_[9456]_  = (~\new_[11010]_  | ~\new_[10186]_ ) & (~\new_[7737]_  | ~\new_[10245]_ );
  assign \new_[9457]_  = (~\new_[10983]_  | ~\new_[10186]_ ) & (~\new_[7703]_  | ~\new_[10245]_ );
  assign \new_[9458]_  = (~\new_[10186]_  | ~\new_[7982]_ ) & (~\new_[10245]_  | ~\new_[7724]_ );
  assign \new_[9459]_  = (~\new_[8048]_  | ~\new_[10242]_ ) & (~\new_[7594]_  | ~\new_[10188]_ );
  assign \new_[9460]_  = ~\new_[10505]_  | ~\new_[10932]_  | ~\new_[10159]_ ;
  assign \new_[9461]_  = (~\new_[7704]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[19] );
  assign \new_[9462]_  = (~\new_[11177]_  | ~\new_[10186]_ ) & (~\new_[7960]_  | ~\new_[10245]_ );
  assign \new_[9463]_  = (~\new_[7749]_  | ~\new_[10188]_ ) & (~\new_[8355]_  | ~\new_[10249]_ );
  assign \new_[9464]_  = (~\new_[7743]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[31] );
  assign \new_[9465]_  = (~\new_[7741]_  | ~\new_[10188]_ ) & (~\new_[8232]_  | ~\new_[10249]_ );
  assign \new_[9466]_  = (~\new_[7926]_  | ~\new_[10186]_ ) & (~\new_[7833]_  | ~\new_[10245]_ );
  assign \new_[9467]_  = (~\new_[7745]_  | ~\new_[10188]_ ) & (~\new_[8400]_  | ~\new_[10249]_ );
  assign \new_[9468]_  = (~\new_[11173]_  | ~\new_[10186]_ ) & (~\new_[11008]_  | ~\new_[10245]_ );
  assign \new_[9469]_  = (~\new_[7927]_  | ~\new_[10186]_ ) & (~\new_[7723]_  | ~\new_[10245]_ );
  assign \new_[9470]_  = (~\new_[7934]_  | ~\new_[10186]_ ) & (~\new_[10245]_  | ~\new_[7850]_ );
  assign \new_[9471]_  = (~\new_[7972]_  | ~\new_[10186]_ ) & (~\new_[10245]_  | ~\new_[7828]_ );
  assign \new_[9472]_  = (~\new_[7620]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[17] );
  assign \new_[9473]_  = (~\new_[7622]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[12] );
  assign \new_[9474]_  = (~\new_[8078]_  | ~\new_[10242]_ ) & (~\new_[10188]_  | ~\new_[7616]_ );
  assign \new_[9475]_  = (~\new_[7735]_  | ~\new_[10188]_ ) & (~\new_[8352]_  | ~\new_[10249]_ );
  assign n5101 = \wb_data_i[6]  ? \new_[10221]_  : n5486;
  assign n4966 = \wb_data_i[9]  ? \new_[10221]_  : n5586;
  assign n4951 = \wb_data_i[7]  ? \new_[10221]_  : n5566;
  assign \new_[9479]_  = ~\new_[9954]_ ;
  assign n5076 = \wb_data_i[22]  ? \new_[10221]_  : n5546;
  assign n4956 = \wb_data_i[24]  ? \new_[10221]_  : n5661;
  assign n4986 = \wb_data_i[26]  ? \new_[10221]_  : n5506;
  assign n5131 = \wb_data_i[2]  ? \new_[10221]_  : n5581;
  assign n5006 = \wb_data_i[19]  ? \new_[10221]_  : n5491;
  assign n5116 = \wb_data_i[23]  ? \new_[10221]_  : n5601;
  assign n5031 = \wb_data_i[15]  ? \new_[10221]_  : n5626;
  assign n5121 = \wb_data_i[12]  ? \new_[10221]_  : n5641;
  assign n5036 = \wb_data_i[10]  ? \new_[10221]_  : n5611;
  assign \new_[9489]_  = ~\new_[10417]_  & ~\new_[10673]_ ;
  assign n5051 = \wb_data_i[21]  ? \new_[10221]_  : n5561;
  assign n4976 = \wb_data_i[20]  ? \new_[10221]_  : n5571;
  assign n5061 = \wb_data_i[31]  ? \new_[10221]_  : n5496;
  assign \new_[9493]_  = ~u4_rfr_en_reg;
  assign \new_[9494]_  = ~\new_[9959]_ ;
  assign \new_[9495]_  = ~\new_[10096]_  | ~\new_[10034]_ ;
  assign \new_[9496]_  = ~\new_[9973]_  | ~\new_[10145]_ ;
  assign \new_[9497]_  = ~\new_[10131]_  | ~\new_[10014]_ ;
  assign \new_[9498]_  = ~\new_[10073]_  | ~\new_[10067]_ ;
  assign \new_[9499]_  = ~\new_[10100]_  | ~\new_[10142]_ ;
  assign \new_[9500]_  = (~\new_[12607]_  | ~\new_[4339]_ ) & (~\new_[12670]_  | ~\new_[4528]_ );
  assign \new_[9501]_  = (~\new_[11800]_  | ~\new_[4401]_ ) & (~\new_[11802]_  | ~\new_[4426]_ );
  assign \new_[9502]_  = (~\new_[11800]_  | ~\new_[4415]_ ) & (~\new_[11802]_  | ~\new_[4440]_ );
  assign \new_[9503]_  = (~\new_[11800]_  | ~\new_[4416]_ ) & (~\new_[11792]_  | ~\new_[4391]_ );
  assign \new_[9504]_  = (~\new_[11792]_  | ~\new_[4182]_ ) & (~\new_[12670]_  | ~\new_[4353]_ );
  assign \new_[9505]_  = (~\new_[11802]_  | ~\new_[4430]_ ) & (~\new_[11792]_  | ~\new_[4379]_ );
  assign \new_[9506]_  = (~\new_[11800]_  | ~\new_[4410]_ ) & (~\new_[11802]_  | ~\new_[4434]_ );
  assign \new_[9507]_  = (~\new_[11800]_  | ~\new_[4417]_ ) & (~\new_[11802]_  | ~\new_[4443]_ );
  assign \new_[9508]_  = (~\new_[11792]_  | ~\new_[4371]_ ) & (~\new_[12670]_  | ~\new_[4346]_ );
  assign \new_[9509]_  = (~\new_[11800]_  | ~\new_[4396]_ ) & (~\new_[11802]_  | ~\new_[4421]_ );
  assign \new_[9510]_  = (~\new_[11800]_  | ~\new_[4395]_ ) & (~\new_[11802]_  | ~\new_[4419]_ );
  assign \new_[9511]_  = (~\new_[11792]_  | ~\new_[4385]_ ) & (~\new_[11790]_  | ~\new_[4358]_ );
  assign \new_[9512]_  = (~\new_[11800]_  | ~\new_[4289]_ ) & (~\new_[11802]_  | ~\new_[4420]_ );
  assign \new_[9513]_  = (~\new_[11800]_  | ~\new_[4399]_ ) & (~\new_[11802]_  | ~\new_[4424]_ );
  assign \new_[9514]_  = (~\new_[11802]_  | ~\new_[4438]_ ) & (~\new_[12607]_  | ~\new_[4388]_ );
  assign \new_[9515]_  = (~\new_[11792]_  | ~\new_[4380]_ ) & (~\new_[12670]_  | ~\new_[4532]_ );
  assign \new_[9516]_  = (~\new_[11802]_  | ~\new_[4427]_ ) & (~\new_[11790]_  | ~\new_[4349]_ );
  assign \new_[9517]_  = (~\new_[11800]_  | ~\new_[4404]_ ) & (~\new_[11802]_  | ~\new_[4429]_ );
  assign \new_[9518]_  = (~\new_[11800]_  | ~\new_[4408]_ ) & (~\new_[11802]_  | ~\new_[4433]_ );
  assign \new_[9519]_  = (~\new_[11800]_  | ~\new_[4278]_ ) & (~\new_[11802]_  | ~\new_[4535]_ );
  assign \new_[9520]_  = (~\new_[11792]_  | ~\new_[4494]_ ) & (~\new_[11790]_  | ~\new_[4188]_ );
  assign \new_[9521]_  = (~\new_[11800]_  | ~\new_[4411]_ ) & (~\new_[11802]_  | ~\new_[4436]_ );
  assign \new_[9522]_  = (~\new_[11800]_  | ~\new_[4405]_ ) & (~\new_[11790]_  | ~\new_[4352]_ );
  assign \new_[9523]_  = (~\new_[11802]_  | ~\new_[4425]_ ) & (~\new_[11792]_  | ~\new_[4374]_ );
  assign \new_[9524]_  = (~\new_[11800]_  | ~\new_[4191]_ ) & (~\new_[11802]_  | ~\new_[4509]_ );
  assign \new_[9525]_  = (~\new_[11800]_  | ~\new_[4409]_ ) & (~\new_[11802]_  | ~\new_[4506]_ );
  assign \new_[9526]_  = (~\new_[11792]_  | ~\new_[4377]_ ) & (~\new_[12670]_  | ~\new_[4351]_ );
  assign \new_[9527]_  = (~\new_[11800]_  | ~\new_[4533]_ ) & (~\new_[11802]_  | ~\new_[4442]_ );
  assign \new_[9528]_  = (~\new_[11800]_  | ~\new_[4249]_ ) & (~\new_[11802]_  | ~\new_[4517]_ );
  assign \new_[9529]_  = (~\new_[11792]_  | ~\new_[4295]_ ) & (~\new_[12670]_  | ~\new_[4364]_ );
  assign \new_[9530]_  = (~\new_[12607]_  | ~\new_[4383]_ ) & (~\new_[11790]_  | ~\new_[4356]_ );
  assign \new_[9531]_  = (~\new_[11792]_  | ~\new_[4373]_ ) & (~\new_[12670]_  | ~\new_[4347]_ );
  assign \new_[9532]_  = (~\new_[11792]_  | ~\new_[4369]_ ) & (~\new_[11790]_  | ~\new_[4344]_ );
  assign \new_[9533]_  = (~\new_[11800]_  | ~\new_[4407]_ ) & (~\new_[11802]_  | ~\new_[4432]_ );
  assign \new_[9534]_  = (~\new_[11792]_  | ~\new_[4510]_ ) & (~\new_[12670]_  | ~\new_[4199]_ );
  assign \new_[9535]_  = (~\new_[11802]_  | ~\new_[4515]_ ) & (~\new_[11790]_  | ~\new_[4354]_ );
  assign \new_[9536]_  = (~\new_[11800]_  | ~\new_[4195]_ ) & (~\new_[11792]_  | ~\new_[4381]_ );
  assign \new_[9537]_  = (~\new_[11800]_  | ~\new_[4406]_ ) & (~\new_[11802]_  | ~\new_[4431]_ );
  assign \new_[9538]_  = (~\new_[11800]_  | ~\new_[4414]_ ) & (~\new_[11802]_  | ~\new_[4439]_ );
  assign \new_[9539]_  = (~\new_[11800]_  | ~\new_[4521]_ ) & (~\new_[11802]_  | ~\new_[4495]_ );
  assign \new_[9540]_  = (~\new_[11792]_  | ~\new_[4303]_ ) & (~\new_[11790]_  | ~\new_[4480]_ );
  assign \new_[9541]_  = (~\new_[11802]_  | ~\new_[4418]_ ) & (~\new_[11792]_  | ~\new_[4365]_ );
  assign \new_[9542]_  = (~\new_[12607]_  | ~\new_[4389]_ ) & (~\new_[11790]_  | ~\new_[4362]_ );
  assign \new_[9543]_  = (~\new_[11800]_  | ~\new_[4400]_ ) & (~\new_[11790]_  | ~\new_[4189]_ );
  assign \new_[9544]_  = (~\new_[11800]_  | ~\new_[4403]_ ) & (~\new_[11802]_  | ~\new_[4428]_ );
  assign \new_[9545]_  = (~\new_[11800]_  | ~\new_[4205]_ ) & (~\new_[11802]_  | ~\new_[4527]_ );
  assign \new_[9546]_  = (~\new_[11800]_  | ~\new_[4412]_ ) & (~\new_[11802]_  | ~\new_[4437]_ );
  assign \new_[9547]_  = (~\new_[11800]_  | ~\new_[4398]_ ) & (~\new_[11802]_  | ~\new_[4423]_ );
  assign \new_[9548]_  = (~\new_[11800]_  | ~\new_[4185]_ ) & (~\new_[11790]_  | ~\new_[4523]_ );
  assign \new_[9549]_  = (~\new_[11792]_  | ~\new_[4366]_ ) & (~\new_[12670]_  | ~\new_[4343]_ );
  assign \new_[9550]_  = (~\new_[11792]_  | ~\new_[4378]_ ) & (~\new_[11790]_  | ~\new_[4181]_ );
  assign \new_[9551]_  = (~\new_[11800]_  | ~\new_[4198]_ ) & (~\new_[11802]_  | ~\new_[4512]_ );
  assign \new_[9552]_  = (~\new_[12607]_  | ~\new_[4375]_ ) & (~\new_[11790]_  | ~\new_[4186]_ );
  assign \new_[9553]_  = (~\new_[12607]_  | ~\new_[4386]_ ) & (~\new_[12670]_  | ~\new_[4359]_ );
  assign \new_[9554]_  = (~\new_[11792]_  | ~\new_[4368]_ ) & (~\new_[11790]_  | ~\new_[4190]_ );
  assign \new_[9555]_  = (~\new_[11800]_  | ~\new_[4413]_ ) & (~\new_[12670]_  | ~\new_[4361]_ );
  assign \new_[9556]_  = u5_lookup_ready1_reg;
  assign \new_[9557]_  = ~\new_[10412]_  | ~\new_[10851]_ ;
  assign n4946 = ~\new_[11354]_  | ~\new_[11387]_ ;
  assign \new_[9559]_  = ~\new_[9712]_ ;
  assign \new_[9560]_  = \new_[10253]_  & \new_[10872]_ ;
  assign \new_[9561]_  = \new_[10473]_  & \new_[12444]_ ;
  assign \new_[9562]_  = \new_[10253]_  & \new_[11317]_ ;
  assign \new_[9563]_  = ~\new_[8809]_  & ~\new_[9988]_ ;
  assign \new_[9564]_  = ~\new_[12669]_  | ~\new_[9972]_ ;
  assign \new_[9565]_  = ~\new_[12038]_  | ~\new_[10000]_ ;
  assign \new_[9566]_  = ~\new_[12469]_  & ~\new_[10108]_ ;
  assign \new_[9567]_  = ~\new_[9859]_ ;
  assign \new_[9568]_  = ~\new_[10040]_  | ~\new_[10846]_ ;
  assign \new_[9569]_  = \\u0_spec_req_cs_reg[0] ;
  assign \new_[9570]_  = \new_[10391]_  & \new_[11351]_ ;
  assign \new_[9571]_  = ~\new_[10393]_  | ~\new_[10551]_ ;
  assign n5001 = ~\new_[11573]_ ;
  assign \new_[9573]_  = \new_[10572]_  & \new_[11323]_ ;
  assign \new_[9574]_  = ~\new_[10529]_  & ~\new_[10328]_ ;
  assign \new_[9575]_  = \new_[10062]_  & \new_[10846]_ ;
  assign \new_[9576]_  = ~\new_[10125]_  | ~\new_[11227]_ ;
  assign \new_[9577]_  = \new_[9975]_  & \new_[10846]_ ;
  assign \new_[9578]_  = ~\new_[9823]_ ;
  assign \new_[9579]_  = \new_[9969]_  & \new_[10846]_ ;
  assign \new_[9580]_  = ~\new_[11833]_  & ~\new_[11735]_ ;
  assign \new_[9581]_  = ~\new_[4147]_  & ~\new_[11393]_ ;
  assign \new_[9582]_  = ~\new_[9927]_ ;
  assign \new_[9583]_  = ~\new_[7850]_  | (~\new_[10194]_  & ~\new_[10515]_ );
  assign \new_[9584]_  = ~\new_[10088]_  & ~\new_[10698]_ ;
  assign \new_[9585]_  = ~\new_[10088]_  & ~\new_[11317]_ ;
  assign \new_[9586]_  = ~\new_[10417]_  & ~\new_[10704]_ ;
  assign \new_[9587]_  = ~\new_[10088]_  & ~\new_[12184]_ ;
  assign \new_[9588]_  = ~\new_[10088]_  & ~\new_[11349]_ ;
  assign \new_[9589]_  = ~\new_[10088]_  & ~\new_[12555]_ ;
  assign \new_[9590]_  = ~\new_[9936]_ ;
  assign \new_[9591]_  = ~\new_[10417]_  & ~\new_[10747]_ ;
  assign \new_[9592]_  = ~\new_[10088]_  & ~\new_[11737]_ ;
  assign \new_[9593]_  = ~\new_[10088]_  & ~\new_[11321]_ ;
  assign \new_[9594]_  = ~\new_[11062]_  & ~\new_[12045]_ ;
  assign \new_[9595]_  = ~\new_[9743]_ ;
  assign \new_[9596]_  = ~\new_[10417]_  & ~\new_[11889]_ ;
  assign \new_[9597]_  = (~\new_[11048]_  | ~\new_[10186]_ ) & (~\new_[11089]_  | ~\new_[10245]_ );
  assign \new_[9598]_  = ~\new_[4147]_  & ~\new_[12094]_ ;
  assign \new_[9599]_  = ~\new_[9921]_ ;
  assign \new_[9600]_  = (~\new_[12607]_  | ~\new_[4387]_ ) & (~\new_[12670]_  | ~\new_[4360]_ );
  assign \new_[9601]_  = ~\new_[10088]_  & ~\new_[10872]_ ;
  assign \new_[9602]_  = ~\new_[10088]_  & ~\new_[10591]_ ;
  assign \new_[9603]_  = ~\new_[10417]_  & ~\new_[11344]_ ;
  assign \new_[9604]_  = ~\new_[9925]_ ;
  assign \new_[9605]_  = (~\new_[11011]_  | ~\new_[10186]_ ) & (~\new_[7702]_  | ~\new_[10245]_ );
  assign \new_[9606]_  = ~\new_[10511]_  & ~\new_[10552]_ ;
  assign \new_[9607]_  = ~\new_[9894]_ ;
  assign \new_[9608]_  = ~\new_[10511]_  & ~\new_[10754]_ ;
  assign \new_[9609]_  = ~\new_[10148]_  & ~\new_[11324]_ ;
  assign \new_[9610]_  = ~\new_[11062]_  & ~\new_[10658]_ ;
  assign \new_[9611]_  = ~\new_[9956]_ ;
  assign \new_[9612]_  = ~\new_[10088]_  & ~\new_[10752]_ ;
  assign \new_[9613]_  = ~\new_[10148]_  & ~\new_[11338]_ ;
  assign \new_[9614]_  = ~\new_[10088]_  & ~\new_[10724]_ ;
  assign \new_[9615]_  = ~\new_[10088]_  & ~\new_[11881]_ ;
  assign \new_[9616]_  = ~\new_[10417]_  & ~\new_[10575]_ ;
  assign \new_[9617]_  = ~\new_[10111]_ ;
  assign \new_[9618]_  = ~\new_[9742]_ ;
  assign \new_[9619]_  = ~\new_[9714]_ ;
  assign \new_[9620]_  = ~\new_[10511]_  & ~\new_[10485]_ ;
  assign \new_[9621]_  = ~\new_[4147]_  & ~\new_[11012]_ ;
  assign \new_[9622]_  = ~\new_[11973]_ ;
  assign \new_[9623]_  = ~\new_[10097]_ ;
  assign \new_[9624]_  = ~\new_[10874]_  | ~\new_[8809]_  | ~\new_[10075]_  | ~\new_[10823]_ ;
  assign \new_[9625]_  = ~\new_[8197]_  & ~\new_[12045]_ ;
  assign \new_[9626]_  = ~\new_[8197]_  & ~\new_[11299]_ ;
  assign \new_[9627]_  = ~\new_[9774]_ ;
  assign \new_[9628]_  = ~\new_[8197]_  & ~\new_[10485]_ ;
  assign \new_[9629]_  = ~\new_[8197]_  & ~\new_[12274]_ ;
  assign \new_[9630]_  = ~\new_[8197]_  & ~\new_[10673]_ ;
  assign \new_[9631]_  = ~\new_[10367]_  & ~\new_[11526]_ ;
  assign \new_[9632]_  = ~\new_[8197]_  & ~\new_[10348]_ ;
  assign \new_[9633]_  = ~\new_[8197]_  & ~\new_[11368]_ ;
  assign \new_[9634]_  = ~\new_[10326]_  & ~\new_[9968]_ ;
  assign \new_[9635]_  = ~\new_[8197]_  & ~\new_[11317]_ ;
  assign \new_[9636]_  = (~\new_[11800]_  | ~\new_[4393]_ ) & (~\new_[11790]_  | ~\new_[4342]_ );
  assign \new_[9637]_  = (~\new_[11200]_  | ~\new_[10186]_ ) & (~\new_[10978]_  | ~\new_[10245]_ );
  assign \new_[9638]_  = ~\new_[10300]_  | ~\new_[10785]_ ;
  assign \new_[9639]_  = ~\new_[8809]_  | ~\new_[10133]_  | ~\new_[10969]_ ;
  assign \new_[9640]_  = \new_[10064]_  & \new_[10846]_ ;
  assign \new_[9641]_  = ~\new_[9866]_ ;
  assign \new_[9642]_  = ~\new_[10102]_  | ~\new_[10846]_ ;
  assign \new_[9643]_  = ~\new_[10092]_  & ~\new_[10369]_ ;
  assign \new_[9644]_  = ~\new_[9836]_ ;
  assign \new_[9645]_  = (~\new_[7706]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[20] );
  assign \new_[9646]_  = \new_[10084]_  & \new_[10846]_ ;
  assign \new_[9647]_  = ~\new_[10809]_ ;
  assign \new_[9648]_  = ~\new_[12555]_ ;
  assign \new_[9649]_  = ~\new_[10511]_  & ~\new_[10160]_ ;
  assign \new_[9650]_  = (~\new_[11061]_  | ~\new_[10186]_ ) & (~\new_[11198]_  | ~\new_[10245]_ );
  assign \new_[9651]_  = ~\new_[10529]_  & ~\new_[11575]_ ;
  assign \new_[9652]_  = (~\new_[11802]_  | ~\new_[4441]_ ) & (~\new_[11790]_  | ~\new_[4519]_ );
  assign \new_[9653]_  = ~\new_[9950]_ ;
  assign \new_[9654]_  = (~\new_[7613]_  | ~\new_[10188]_ ) & (~\new_[10236]_  | ~\poc_o[15] );
  assign \new_[9655]_  = ~\new_[10150]_ ;
  assign \new_[9656]_  = (~\new_[11117]_  | ~\new_[10186]_ ) & (~\new_[11190]_  | ~\new_[10245]_ );
  assign \new_[9657]_  = \new_[9950]_ ;
  assign \new_[9658]_  = ~\new_[9902]_ ;
  assign \new_[9659]_  = ~\new_[10148]_  & ~\new_[11314]_ ;
  assign \new_[9660]_  = ~\new_[9908]_ ;
  assign \new_[9661]_  = ~\new_[9867]_ ;
  assign n5126 = \wb_data_i[4]  ? \new_[10221]_  : n5631;
  assign \new_[9663]_  = ~\new_[4147]_  & ~\new_[12611]_ ;
  assign \new_[9664]_  = ~\new_[10047]_  | ~\new_[10846]_ ;
  assign \new_[9665]_  = ~\new_[9899]_ ;
  assign \new_[9666]_  = (~\new_[11792]_  | ~\new_[4384]_ ) & (~\new_[11790]_  | ~\new_[4357]_ );
  assign \new_[9667]_  = (~\new_[11800]_  | ~\new_[4183]_ ) & (~\new_[11802]_  | ~\new_[4511]_ );
  assign \new_[9668]_  = ~\new_[10511]_  & ~\new_[11881]_ ;
  assign \new_[9669]_  = ~\new_[10881]_  | ~\new_[10945]_  | ~\new_[10225]_ ;
  assign \new_[9670]_  = ~\new_[10106]_  & (~\new_[3388]_  | ~\new_[10425]_ );
  assign n4996 = \wb_data_i[1]  ? \new_[10221]_  : n5676;
  assign n4981 = \wb_data_i[3]  ? \new_[10221]_  : n5606;
  assign \new_[9673]_  = (~\new_[11800]_  | ~\new_[4397]_ ) & (~\new_[11802]_  | ~\new_[4422]_ );
  assign \new_[9674]_  = ~\new_[12052]_ ;
  assign \new_[9675]_  = ~\new_[9918]_ ;
  assign n5086 = \wb_data_i[17]  ? \new_[10221]_  : n5666;
  assign \new_[9677]_  = (~\new_[11792]_  | ~\new_[4372]_ ) & (~\new_[11790]_  | ~\new_[4180]_ );
  assign \new_[9678]_  = ~\new_[10088]_  & ~\new_[11341]_ ;
  assign n5091 = \wb_data_i[30]  ? \new_[10221]_  : n5536;
  assign \new_[9680]_  = ~\new_[9838]_ ;
  assign \new_[9681]_  = \new_[10304]_  & \new_[12444]_ ;
  assign \new_[9682]_  = ~\new_[9860]_ ;
  assign n5026 = \wb_data_i[29]  ? \new_[10221]_  : n5636;
  assign \new_[9684]_  = ~\new_[9911]_ ;
  assign \new_[9685]_  = \new_[10488]_  | \new_[11015]_ ;
  assign n5066 = \wb_data_i[28]  ? \new_[10221]_  : n5516;
  assign \new_[9687]_  = (~\new_[11792]_  | ~\new_[4392]_ ) & (~\new_[12670]_  | ~\new_[4514]_ );
  assign \new_[9688]_  = (~\new_[11792]_  | ~\new_[4390]_ ) & (~\new_[11790]_  | ~\new_[4516]_ );
  assign n5016 = \wb_data_i[18]  ? \new_[10221]_  : n5521;
  assign \new_[9690]_  = ~\new_[10886]_  | ~\new_[8809]_  | ~\new_[10035]_  | ~\new_[10974]_ ;
  assign \new_[9691]_  = ~\new_[10154]_  | ~\new_[12093]_ ;
  assign \new_[9692]_  = \\u1_u0_out_r_reg[2] ;
  assign \new_[9693]_  = \new_[12668]_  & \new_[11344]_ ;
  assign \new_[9694]_  = ~\new_[10511]_  & ~\new_[10397]_ ;
  assign \new_[9695]_  = ~\new_[10861]_  | ~\new_[10431]_  | ~\new_[10881]_ ;
  assign n4991 = \wb_data_i[16]  ? \new_[10221]_  : n5551;
  assign n5096 = \wb_data_i[14]  ? \new_[10221]_  : n5591;
  assign \new_[9698]_  = (~\new_[11800]_  | ~\new_[4402]_ ) & (~\new_[11792]_  | ~\new_[4376]_ );
  assign n5011 = \wb_data_i[13]  ? \new_[10221]_  : n5596;
  assign n4971 = \wb_data_i[0]  ? \new_[10221]_  : n5656;
  assign \new_[9701]_  = ~\new_[12442]_  | ~\new_[10304]_ ;
  assign n4961 = \wb_data_i[25]  ? \new_[10221]_  : n5616;
  assign n5056 = \wb_data_i[27]  ? \new_[10221]_  : n5621;
  assign n5081 = \wb_data_i[5]  ? \new_[10221]_  : n5531;
  assign n5111 = \wb_data_i[8]  ? \new_[10221]_  : n5471;
  assign \new_[9706]_  = ~\new_[9752]_ ;
  assign \new_[9707]_  = ~\new_[9955]_ ;
  assign \new_[9708]_  = (~\new_[11802]_  | ~\new_[4504]_ ) & (~\new_[11792]_  | ~\new_[4313]_ );
  assign \new_[9709]_  = ~\new_[9905]_ ;
  assign \new_[9710]_  = ~\new_[9868]_ ;
  assign \new_[9711]_  = \new_[10907]_  | \new_[1611]_  | \new_[10173]_  | \new_[2070]_ ;
  assign \new_[9712]_  = ~\new_[11921]_  | ~\new_[10486]_  | ~\new_[11920]_ ;
  assign \new_[9713]_  = ~\new_[10137]_ ;
  assign \new_[9714]_  = ~\new_[10154]_  | ~\new_[1488]_ ;
  assign \new_[9715]_  = ~\new_[10154]_  | ~\new_[12756]_ ;
  assign \new_[9716]_  = ~\new_[10162]_  & ~\new_[2056]_ ;
  assign \new_[9717]_  = ~\new_[10154]_  | ~\new_[12609]_ ;
  assign \new_[9718]_  = ~\new_[10154]_  | ~\new_[10827]_ ;
  assign n5241 = \new_[9366]_  ? \new_[10851]_  : \wb_addr_i[21] ;
  assign \new_[9720]_  = ~\new_[10159]_  & (~\new_[10414]_  | ~\new_[1539]_ );
  assign \new_[9721]_  = ~\new_[10853]_  | ~\new_[10261]_  | ~\new_[10505]_ ;
  assign \new_[9722]_  = ~\new_[8049]_  | ~\new_[8075]_  | ~\new_[10230]_  | ~\new_[10834]_ ;
  assign \new_[9723]_  = (~\new_[3048]_  | ~\new_[10371]_ ) & (~\new_[10896]_  | ~\new_[10956]_ );
  assign \new_[9724]_  = \new_[1611]_  ^ \new_[10350]_ ;
  assign \new_[9725]_  = \new_[1657]_  ^ \new_[10341]_ ;
  assign \new_[9726]_  = ~\new_[10176]_  & ~\new_[11098]_ ;
  assign \new_[9727]_  = ~\new_[10230]_  | ~\new_[8049]_ ;
  assign \new_[9728]_  = ~\new_[10307]_  | ~\new_[10480]_  | ~\new_[10426]_ ;
  assign n5231 = \new_[9362]_  ? \new_[10851]_  : \wb_addr_i[14] ;
  assign \new_[9730]_  = \new_[10214]_  & \new_[10554]_ ;
  assign n5196 = \new_[9337]_  ? \new_[10851]_  : \wb_addr_i[10] ;
  assign \new_[9732]_  = ~\new_[1433]_  | ~\new_[10526]_ ;
  assign \new_[9733]_  = ~\new_[10331]_  | ~\new_[10448]_  | ~\new_[10403]_ ;
  assign \new_[9734]_  = \new_[10253]_  & \new_[10676]_ ;
  assign \new_[9735]_  = (~\new_[3049]_  | ~\new_[10371]_ ) & (~\new_[10828]_  | ~\new_[10956]_ );
  assign \new_[9736]_  = u5_mc_adv_r_reg;
  assign \new_[9737]_  = ~\new_[11062]_  & ~\new_[10809]_ ;
  assign \new_[9738]_  = ~\new_[9987]_ ;
  assign \new_[9739]_  = ~\new_[10154]_  | ~\new_[10933]_ ;
  assign n5211 = \new_[9347]_  ? \new_[10851]_  : \wb_addr_i[9] ;
  assign \new_[9741]_  = (~\new_[3709]_  | ~\new_[10371]_ ) & (~\new_[10852]_  | ~\new_[10956]_ );
  assign \new_[9742]_  = ~\new_[10517]_  | ~\new_[10950]_ ;
  assign \new_[9743]_  = ~\new_[9980]_ ;
  assign \new_[9744]_  = ~\new_[11335]_  | ~\new_[10252]_ ;
  assign \new_[9745]_  = \new_[2070]_  ^ \new_[10317]_ ;
  assign \new_[9746]_  = ~\new_[10417]_  & ~\new_[10348]_ ;
  assign \new_[9747]_  = \new_[7284]_  ^ \new_[10298]_ ;
  assign \new_[9748]_  = ~\new_[8197]_  & ~\new_[11314]_ ;
  assign \new_[9749]_  = (~\new_[10296]_  | ~\new_[10434]_ ) & (~\new_[10338]_  | ~\new_[10422]_ );
  assign \new_[9750]_  = \new_[10231]_  & \new_[10934]_ ;
  assign \new_[9751]_  = ~\new_[10206]_  & (~\new_[10939]_  | ~\new_[10956]_ );
  assign \new_[9752]_  = ~\new_[10004]_ ;
  assign n5156 = ~\new_[10174]_  & ~\new_[11033]_ ;
  assign \new_[9754]_  = ~\new_[10236]_  | ~\poc_o[10] ;
  assign \new_[9755]_  = ~\new_[10222]_  & ~\new_[10646]_ ;
  assign \new_[9756]_  = ~\new_[10187]_  & ~\new_[10619]_ ;
  assign \new_[9757]_  = ~\new_[10236]_  | ~\poc_o[27] ;
  assign \new_[9758]_  = ~\new_[10236]_  | ~\poc_o[8] ;
  assign \new_[9759]_  = ~\new_[10236]_  | ~\poc_o[24] ;
  assign \new_[9760]_  = ~\new_[10236]_  | ~\poc_o[25] ;
  assign \new_[9761]_  = ~\new_[10236]_  | ~\poc_o[29] ;
  assign \new_[9762]_  = ~\new_[10191]_  & ~\new_[10570]_ ;
  assign \new_[9763]_  = ~\new_[10192]_  & ~\new_[10643]_ ;
  assign \new_[9764]_  = ~\new_[10189]_  & ~\new_[10779]_ ;
  assign \new_[9765]_  = ~\new_[10158]_  & ~\new_[10757]_ ;
  assign \new_[9766]_  = ~\new_[10249]_  | ~\new_[8365]_ ;
  assign \new_[9767]_  = ~\new_[8390]_  | ~\new_[10249]_ ;
  assign \new_[9768]_  = ~\new_[11082]_  | ~\new_[10242]_ ;
  assign \new_[9769]_  = ~\new_[11234]_  | ~\new_[10242]_ ;
  assign \new_[9770]_  = ~\new_[11028]_  | ~\new_[10242]_ ;
  assign \new_[9771]_  = ~\new_[10249]_  | ~mc_vpen_pad_o;
  assign \new_[9772]_  = ~\new_[10092]_ ;
  assign \new_[9773]_  = ~\new_[11220]_  | ~\new_[10242]_ ;
  assign \new_[9774]_  = ~\new_[10367]_  & ~\new_[10818]_ ;
  assign \new_[9775]_  = ~\new_[11223]_  | ~\new_[10242]_ ;
  assign \new_[9776]_  = ~\new_[10264]_  & ~\new_[10613]_ ;
  assign \new_[9777]_  = ~\new_[11253]_  | ~\new_[10249]_ ;
  assign \new_[9778]_  = ~\new_[10249]_  | ~\new_[8387]_ ;
  assign \new_[9779]_  = ~\new_[11243]_  | ~\new_[10242]_ ;
  assign \new_[9780]_  = ~\new_[11042]_  | ~\new_[10249]_ ;
  assign \new_[9781]_  = ~\new_[10341]_  & (~\new_[10601]_  | ~\new_[1644]_ );
  assign \new_[9782]_  = ~\new_[11188]_  | ~\new_[10242]_ ;
  assign \new_[9783]_  = ~\new_[11250]_  | ~\new_[10242]_ ;
  assign \new_[9784]_  = ~\new_[11093]_  | ~\new_[10242]_ ;
  assign \new_[9785]_  = ~\new_[10397]_ ;
  assign \new_[9786]_  = ~\new_[11066]_  | ~\new_[10242]_ ;
  assign \new_[9787]_  = ~\new_[11245]_  | ~\new_[10242]_ ;
  assign \new_[9788]_  = ~\new_[10306]_  | ~\new_[10422]_  | ~\new_[10421]_ ;
  assign \new_[9789]_  = ~\new_[10226]_  & ~\new_[10515]_ ;
  assign \new_[9790]_  = ~\new_[10308]_  | ~\new_[10429]_  | ~\new_[10443]_ ;
  assign \new_[9791]_  = ~\new_[10389]_  | ~\new_[10415]_  | ~\new_[10424]_ ;
  assign \new_[9792]_  = (~\new_[3043]_  | ~\new_[10371]_ ) & (~\new_[10817]_  | ~\new_[10956]_ );
  assign \new_[9793]_  = (~\new_[3697]_  | ~\new_[10371]_ ) & (~\new_[10844]_  | ~\new_[10956]_ );
  assign \new_[9794]_  = (~\new_[3707]_  | ~\new_[10371]_ ) & (~\new_[10869]_  | ~\new_[10956]_ );
  assign \new_[9795]_  = (~\new_[3045]_  | ~\new_[10371]_ ) & (~\new_[10885]_  | ~\new_[10956]_ );
  assign \new_[9796]_  = (~\new_[2971]_  | ~\new_[10371]_ ) & (~\new_[10825]_  | ~\new_[10956]_ );
  assign \new_[9797]_  = (~\new_[3706]_  | ~\new_[10371]_ ) & (~\new_[10968]_  | ~\new_[10956]_ );
  assign \new_[9798]_  = (~\new_[3711]_  | ~\new_[10371]_ ) & (~\new_[10833]_  | ~\new_[10956]_ );
  assign \new_[9799]_  = (~\new_[3710]_  | ~\new_[10371]_ ) & (~\new_[10819]_  | ~\new_[10956]_ );
  assign \new_[9800]_  = (~\new_[3705]_  | ~\new_[10371]_ ) & (~\new_[10845]_  | ~\new_[10956]_ );
  assign \new_[9801]_  = (~\new_[3046]_  | ~\new_[10371]_ ) & (~\new_[10878]_  | ~\new_[10956]_ );
  assign \new_[9802]_  = ~\new_[11240]_  | ~\new_[10242]_ ;
  assign \new_[9803]_  = \new_[10163]_  | \new_[11141]_ ;
  assign \new_[9804]_  = \new_[10168]_  & \new_[11341]_ ;
  assign \new_[9805]_  = \new_[10253]_  & \new_[11335]_ ;
  assign \new_[9806]_  = ~wb_cyc_i | ~\new_[10151]_  | ~\new_[11258]_ ;
  assign \new_[9807]_  = ~\new_[10358]_  & ~\new_[10872]_ ;
  assign \new_[9808]_  = (~\new_[3887]_  | ~\new_[10598]_ ) & (~\new_[10972]_  | ~\new_[10956]_ );
  assign \new_[9809]_  = ~\new_[10224]_  & (~\new_[10947]_  | ~\new_[10956]_ );
  assign \new_[9810]_  = ~\new_[10070]_ ;
  assign \new_[9811]_  = ~\new_[10169]_  & (~\new_[10835]_  | ~\new_[10956]_ );
  assign \new_[9812]_  = (~\new_[3876]_  | ~\new_[10598]_ ) & (~\new_[10814]_  | ~\new_[10956]_ );
  assign \new_[9813]_  = ~\new_[10771]_  | ~\new_[9913]_  | ~\new_[11299]_ ;
  assign \new_[9814]_  = \new_[10920]_  & \new_[10216]_ ;
  assign \new_[9815]_  = \new_[10552]_  & \new_[10211]_ ;
  assign \new_[9816]_  = ~\new_[9978]_ ;
  assign \new_[9817]_  = \new_[10572]_  & \new_[10938]_ ;
  assign \new_[9818]_  = ~\new_[10417]_  & ~\new_[11311]_ ;
  assign \new_[9819]_  = ~\new_[10959]_  | ~\new_[10157]_  | ~\new_[10771]_ ;
  assign \new_[9820]_  = ~\new_[8197]_  & ~\new_[11393]_ ;
  assign \new_[9821]_  = \new_[10572]_  & \new_[10922]_ ;
  assign \new_[9822]_  = ~\new_[11062]_  & ~\new_[11575]_ ;
  assign \new_[9823]_  = \new_[10210]_  & \new_[10846]_ ;
  assign \new_[9824]_  = ~\new_[10417]_  & ~\new_[12599]_ ;
  assign n5251 = \new_[9373]_  ? \new_[10851]_  : \wb_addr_i[19] ;
  assign n5151 = \new_[9207]_  ? \new_[10851]_  : \wb_addr_i[22] ;
  assign n5216 = \new_[9350]_  ? \new_[10851]_  : \wb_addr_i[17] ;
  assign n5166 = \new_[9306]_  ? \new_[10851]_  : \wb_addr_i[25] ;
  assign n5221 = \new_[9351]_  ? \new_[10851]_  : \wb_addr_i[16] ;
  assign n5136 = \new_[9176]_  ? \new_[10851]_  : \wb_addr_i[7] ;
  assign n5186 = \new_[9334]_  ? \new_[10851]_  : \wb_addr_i[2] ;
  assign n5206 = \new_[9342]_  ? \new_[10851]_  : \wb_addr_i[15] ;
  assign n5246 = \new_[9369]_  ? \new_[10851]_  : \wb_addr_i[24] ;
  assign n5256 = \new_[9380]_  ? \new_[10851]_  : \wb_addr_i[11] ;
  assign \new_[9835]_  = \new_[8079]_  ^ \new_[10359]_ ;
  assign \new_[9836]_  = ~\new_[10154]_  | ~\new_[10164]_ ;
  assign \new_[9837]_  = ~\new_[10417]_  & ~\new_[10676]_ ;
  assign \new_[9838]_  = ~\new_[10154]_  | ~\new_[10177]_ ;
  assign \new_[9839]_  = ~\new_[11062]_  & ~\new_[12555]_ ;
  assign \new_[9840]_  = ~\new_[10417]_  & ~\new_[11329]_ ;
  assign \new_[9841]_  = ~\new_[11062]_  & ~\new_[12564]_ ;
  assign \new_[9842]_  = ~\new_[10417]_  & ~\new_[10920]_ ;
  assign \new_[9843]_  = ~\new_[11062]_  & ~\new_[11364]_ ;
  assign \new_[9844]_  = ~\new_[10417]_  & ~\new_[12757]_ ;
  assign \new_[9845]_  = ~\new_[10254]_ ;
  assign \new_[9846]_  = ~\new_[10378]_  & ~\new_[12052]_ ;
  assign \new_[9847]_  = ~\new_[11062]_  & ~\new_[12599]_ ;
  assign \new_[9848]_  = ~\new_[11062]_  & ~\new_[10551]_ ;
  assign \new_[9849]_  = ~\new_[11062]_  & ~\new_[10920]_ ;
  assign \new_[9850]_  = ~\new_[10417]_  & ~\new_[10767]_ ;
  assign \new_[9851]_  = ~\new_[9979]_ ;
  assign \new_[9852]_  = ~\new_[10618]_  & ~\new_[10202]_ ;
  assign \new_[9853]_  = ~\new_[10101]_ ;
  assign \new_[9854]_  = ~\new_[11062]_  & ~\new_[11334]_ ;
  assign \new_[9855]_  = ~\new_[10417]_  & ~\new_[10897]_ ;
  assign \new_[9856]_  = ~\new_[10378]_  & ~\new_[12094]_ ;
  assign \new_[9857]_  = ~\new_[10417]_  & ~\new_[12052]_ ;
  assign \new_[9858]_  = ~\new_[11043]_  | ~\new_[10242]_ ;
  assign \new_[9859]_  = ~\new_[10517]_  | ~\new_[11310]_ ;
  assign \new_[9860]_  = ~\new_[10517]_  | ~\new_[9674]_ ;
  assign \new_[9861]_  = ~\new_[10517]_  | ~\new_[10743]_ ;
  assign \new_[9862]_  = ~\new_[10417]_  & ~\new_[10579]_ ;
  assign \new_[9863]_  = ~\new_[10417]_  & ~\new_[10783]_ ;
  assign \new_[9864]_  = \new_[12577]_  & \new_[12089]_ ;
  assign \new_[9865]_  = ~\new_[10417]_  & ~\new_[12564]_ ;
  assign \new_[9866]_  = ~\new_[10154]_  | ~\new_[9913]_ ;
  assign \new_[9867]_  = ~\new_[1433]_  | ~\new_[11348]_ ;
  assign \new_[9868]_  = ~\new_[10083]_ ;
  assign \new_[9869]_  = ~\new_[11241]_  | ~\new_[10242]_ ;
  assign \new_[9870]_  = ~\new_[10378]_  & ~\new_[11368]_ ;
  assign \new_[9871]_  = ~\new_[11062]_  & ~\new_[11324]_ ;
  assign \new_[9872]_  = ~\new_[10378]_  & ~\new_[12611]_ ;
  assign \new_[9873]_  = (~\new_[10371]_  | ~\new_[3044]_ ) & (~\new_[10956]_  | ~\new_[10908]_ );
  assign \new_[9874]_  = ~\new_[10417]_  & ~\new_[10754]_ ;
  assign \new_[9875]_  = ~\new_[11013]_  | ~\new_[10242]_ ;
  assign \new_[9876]_  = ~\new_[11249]_  | ~\new_[10242]_ ;
  assign \new_[9877]_  = \new_[11045]_  & \new_[12089]_ ;
  assign \new_[9878]_  = ~\new_[8197]_  & ~\new_[11324]_ ;
  assign \new_[9879]_  = ~\new_[10922]_  & ~\new_[10827]_ ;
  assign \new_[9880]_  = ~\new_[11062]_  & ~\new_[11344]_ ;
  assign \new_[9881]_  = ~\new_[10991]_  | ~\new_[10242]_ ;
  assign \new_[9882]_  = \new_[10253]_  & \new_[10638]_ ;
  assign \new_[9883]_  = ~\new_[10023]_ ;
  assign \new_[9884]_  = ~\new_[10238]_  & (~\new_[10879]_  | ~\new_[10956]_ );
  assign \new_[9885]_  = \new_[10228]_  & \new_[11917]_ ;
  assign \new_[9886]_  = ~\new_[10219]_  & (~\new_[10867]_  | ~\new_[10956]_ );
  assign \new_[9887]_  = ~\new_[11022]_  | ~\new_[10242]_ ;
  assign n5191 = \new_[9335]_  ? \new_[10851]_  : \wb_addr_i[18] ;
  assign \new_[9889]_  = ~\new_[9997]_ ;
  assign \new_[9890]_  = \new_[10302]_  & \new_[10175]_ ;
  assign \new_[9891]_  = ~\new_[11203]_  | ~\new_[10249]_ ;
  assign \new_[9892]_  = \new_[10572]_  & \new_[11353]_ ;
  assign \new_[9893]_  = ~\new_[10986]_  | ~\new_[10242]_ ;
  assign \new_[9894]_  = ~\new_[10154]_  | ~\new_[10962]_ ;
  assign \new_[9895]_  = ~\new_[10218]_  | ~\wb_addr_i[11] ;
  assign \new_[9896]_  = ~\new_[10010]_ ;
  assign n5146 = \new_[9184]_  ? \new_[10851]_  : \wb_addr_i[20] ;
  assign \new_[9898]_  = ~\new_[11226]_  | ~\new_[10242]_ ;
  assign \new_[9899]_  = ~\new_[10154]_  | ~\new_[10960]_ ;
  assign \new_[9900]_  = ~\new_[11074]_  | ~\new_[10242]_ ;
  assign \new_[9901]_  = ~\new_[11213]_  | ~\new_[10249]_ ;
  assign \new_[9902]_  = ~\new_[10743]_ ;
  assign \new_[9903]_  = ~\new_[10704]_ ;
  assign \new_[9904]_  = ~\new_[10378]_  & ~\new_[10704]_ ;
  assign \new_[9905]_  = ~\new_[10517]_  | ~\new_[11328]_ ;
  assign \new_[9906]_  = ~\new_[10417]_  & ~\new_[11364]_ ;
  assign \new_[9907]_  = ~\new_[10236]_  | ~\poc_o[7] ;
  assign \new_[9908]_  = ~\new_[10154]_  | ~\new_[11320]_ ;
  assign \new_[9909]_  = ~\new_[10236]_  | ~\poc_o[0] ;
  assign \new_[9910]_  = ~\new_[10236]_  | ~\poc_o[26] ;
  assign \new_[9911]_  = ~\new_[10517]_  | ~\new_[11361]_ ;
  assign \new_[9912]_  = ~\new_[11062]_  & ~\new_[12184]_ ;
  assign \new_[9913]_  = ~\new_[10872]_ ;
  assign \new_[9914]_  = \new_[10396]_  & \new_[10246]_ ;
  assign \new_[9915]_  = \new_[10163]_  | \new_[11153]_ ;
  assign \new_[9916]_  = \new_[10253]_  & \new_[10584]_ ;
  assign n5176 = \new_[9332]_  ? \new_[10851]_  : \wb_addr_i[4] ;
  assign \new_[9918]_  = ~\new_[10154]_  | ~\new_[10955]_ ;
  assign \new_[9919]_  = ~\new_[10236]_  | ~\poc_o[28] ;
  assign \new_[9920]_  = ~\new_[10236]_  | ~\poc_o[30] ;
  assign \new_[9921]_  = ~\new_[10154]_  | ~\new_[10419]_ ;
  assign \new_[9922]_  = ~\new_[10011]_ ;
  assign n5171 = \new_[9331]_  ? \new_[10851]_  : \wb_addr_i[13] ;
  assign \new_[9924]_  = ~\new_[10517]_  | ~\new_[10938]_ ;
  assign \new_[9925]_  = ~\new_[10154]_  | ~\new_[11526]_ ;
  assign \new_[9926]_  = ~\new_[10724]_ ;
  assign \new_[9927]_  = ~\new_[10154]_  | ~\new_[11363]_ ;
  assign n5141 = \new_[9179]_  ? \new_[10851]_  : \wb_addr_i[8] ;
  assign \new_[9929]_  = ~\new_[10417]_  & ~\new_[10809]_ ;
  assign \new_[9930]_  = ~\new_[10057]_ ;
  assign n5226 = \new_[9354]_  ? \new_[10851]_  : \wb_addr_i[3] ;
  assign \new_[9932]_  = ~\new_[10412]_ ;
  assign \new_[9933]_  = ~\new_[10417]_  & ~\new_[10722]_ ;
  assign \new_[9934]_  = ~\new_[10171]_  & ~\new_[1712]_ ;
  assign \new_[9935]_  = (~\new_[3047]_  | ~\new_[10371]_ ) & (~\new_[10901]_  | ~\new_[10956]_ );
  assign \new_[9936]_  = ~\new_[10367]_  & ~\new_[10397]_ ;
  assign \new_[9937]_  = ~\new_[10417]_  & ~\new_[10397]_ ;
  assign \new_[9938]_  = \new_[12577]_  & \new_[10922]_ ;
  assign \new_[9939]_  = ~u6_rmw_r_reg;
  assign \new_[9940]_  = ~\new_[10114]_ ;
  assign \new_[9941]_  = ~\new_[10126]_ ;
  assign \new_[9942]_  = ~\new_[10018]_ ;
  assign \new_[9943]_  = ~\new_[10388]_  | ~\new_[10524]_  | ~\new_[10271]_ ;
  assign \new_[9944]_  = \new_[10412]_  | wb_err_o;
  assign n5236 = \new_[9364]_  ? \new_[10851]_  : \wb_addr_i[6] ;
  assign \new_[9946]_  = ~\new_[10767]_ ;
  assign \new_[9947]_  = ~\new_[10202]_  & ~n5416;
  assign n5181 = \new_[9333]_  ? \new_[10851]_  : \wb_addr_i[12] ;
  assign \new_[9949]_  = \new_[1580]_  | \new_[10880]_  | \new_[10193]_  | \new_[1463]_ ;
  assign \new_[9950]_  = ~\new_[10367]_  & ~\new_[12555]_ ;
  assign \new_[9951]_  = ~\new_[10215]_  & ~\new_[12089]_ ;
  assign n5201 = \new_[9339]_  ? \new_[10851]_  : \wb_addr_i[5] ;
  assign \new_[9953]_  = ~\new_[11062]_  & ~\new_[11889]_ ;
  assign \new_[9954]_  = ~\new_[10517]_  | ~\new_[10411]_ ;
  assign \new_[9955]_  = ~\new_[10517]_  | ~\new_[11313]_ ;
  assign \new_[9956]_  = ~\new_[10154]_  | ~n5021;
  assign \new_[9957]_  = \new_[10516]_  & \new_[10239]_ ;
  assign \new_[9958]_  = ~\new_[11776]_  & ~\new_[10897]_ ;
  assign \new_[9959]_  = \new_[10175]_  & \new_[11119]_ ;
  assign \new_[9960]_  = ~\new_[10417]_  & ~\new_[11334]_ ;
  assign \new_[9961]_  = ~\new_[9992]_ ;
  assign \new_[9962]_  = ~\new_[10156]_  & (~\new_[10935]_  | ~\new_[10956]_ );
  assign \new_[9963]_  = ~\new_[10146]_ ;
  assign n5161 = \new_[9257]_  ? \new_[10851]_  : \wb_addr_i[23] ;
  assign \new_[9965]_  = ~\new_[10378]_  & ~\new_[10897]_ ;
  assign \new_[9966]_  = (~\new_[3708]_  | ~\new_[10371]_ ) & (~\new_[10916]_  | ~\new_[10956]_ );
  assign \new_[9967]_  = ~\new_[11062]_  & ~\new_[11338]_ ;
  assign \new_[9968]_  = ~\new_[12555]_ ;
  assign \new_[9969]_  = ~\new_[10417]_  & ~\new_[10658]_ ;
  assign \new_[9970]_  = ~\new_[10511]_  & ~\new_[12757]_ ;
  assign \new_[9971]_  = ~\new_[10833]_  | ~\new_[10598]_ ;
  assign \new_[9972]_  = ~\new_[12445]_ ;
  assign \new_[9973]_  = ~\new_[10968]_  | ~\new_[10491]_ ;
  assign n5271 = ~\new_[10390]_  | (~\new_[8185]_  & ~\new_[11153]_ );
  assign \new_[9975]_  = ~\new_[10417]_  & ~\new_[10551]_ ;
  assign n5266 = ~\new_[10151]_ ;
  assign n5261 = ~\new_[10394]_  | ~\new_[10451]_ ;
  assign \new_[9978]_  = ~\new_[11776]_  & ~\new_[11338]_ ;
  assign \new_[9979]_  = ~\new_[10367]_  & ~\new_[10747]_ ;
  assign \new_[9980]_  = ~\new_[10714]_  & ~\new_[12599]_ ;
  assign \new_[9981]_  = ~\new_[10261]_ ;
  assign \new_[9982]_  = ~\new_[10968]_  | ~\new_[10598]_ ;
  assign \new_[9983]_  = \new_[10650]_  | \new_[10727]_  | \new_[10795]_  | \new_[10642]_ ;
  assign \new_[9984]_  = ~\new_[10919]_  | ~\new_[11920]_  | ~\new_[12045]_ ;
  assign \new_[9985]_  = \new_[10594]_  & \new_[10922]_ ;
  assign \new_[9986]_  = ~\new_[12507]_ ;
  assign \new_[9987]_  = ~\new_[11776]_  & ~\new_[10591]_ ;
  assign \new_[9988]_  = ~\new_[10488]_  | ~wb_we_i;
  assign \new_[9989]_  = ~\new_[10166]_ ;
  assign \new_[9990]_  = ~\new_[10166]_ ;
  assign \new_[9991]_  = \new_[12052]_  & \new_[10552]_ ;
  assign \new_[9992]_  = ~\new_[10267]_ ;
  assign \new_[9993]_  = ~\new_[10819]_  | ~\new_[10491]_ ;
  assign \new_[9994]_  = \new_[3388]_  ^ \new_[10446]_ ;
  assign \new_[9995]_  = ~\new_[10155]_ ;
  assign \new_[9996]_  = ~\new_[10237]_ ;
  assign \new_[9997]_  = \new_[10963]_ ;
  assign \new_[9998]_  = ~\new_[10747]_ ;
  assign \new_[9999]_  = ~\new_[10230]_ ;
  assign \new_[10000]_  = ~\new_[12036]_ ;
  assign \new_[10001]_  = ~\new_[10356]_  & ~\new_[10325]_ ;
  assign \new_[10002]_  = ~\new_[10350]_  & (~\new_[10669]_  | ~\new_[1519]_ );
  assign \new_[10003]_  = ~\new_[10342]_  & (~\new_[11033]_  | ~\new_[10910]_ );
  assign \new_[10004]_  = ~\new_[10235]_ ;
  assign \new_[10005]_  = ~\new_[10343]_  & (~\new_[10944]_  | ~\new_[1462]_ );
  assign \new_[10006]_  = \new_[10615]_  | \new_[10800]_  | \new_[10647]_  | \new_[10753]_ ;
  assign \new_[10007]_  = \new_[10602]_  | \new_[10729]_  | \new_[10796]_  | \new_[10680]_ ;
  assign \new_[10008]_  = \new_[10600]_  | \new_[10763]_  | \new_[10725]_  | \new_[10775]_ ;
  assign \new_[10009]_  = ~u6_write_go_r_reg;
  assign \new_[10010]_  = ~\new_[10325]_  | ~\new_[10821]_ ;
  assign \new_[10011]_  = ~\new_[10714]_  & ~\new_[11334]_ ;
  assign \new_[10012]_  = ~\new_[10299]_  | ~\poc_o[3] ;
  assign \new_[10013]_  = ~\new_[10309]_  & (~\new_[3440]_  | ~\new_[10936]_ );
  assign \new_[10014]_  = (~\new_[10845]_  | ~\new_[10598]_ ) & (~\new_[10942]_  | ~\new_[10956]_ );
  assign \new_[10015]_  = ~\new_[11062]_  & ~\new_[10579]_ ;
  assign \new_[10016]_  = \new_[11387]_  & \new_[10809]_ ;
  assign \new_[10017]_  = \new_[11881]_  & \new_[10322]_ ;
  assign \new_[10018]_  = \new_[11881]_  & \new_[10320]_ ;
  assign \new_[10019]_  = ~\new_[10255]_ ;
  assign \new_[10020]_  = \new_[11324]_  & \new_[10322]_ ;
  assign \new_[10021]_  = ~\new_[12089]_  & ~\new_[10334]_ ;
  assign \new_[10022]_  = \new_[11323]_  & \new_[10322]_ ;
  assign \new_[10023]_  = \new_[10318]_  & \new_[10274]_ ;
  assign \new_[10024]_  = ~\new_[11327]_  & ~\new_[11575]_ ;
  assign \new_[10025]_  = ~\new_[10819]_  | ~\new_[10598]_ ;
  assign \new_[10026]_  = (~\new_[11055]_  | ~\new_[10576]_ ) & (~\new_[11199]_  | ~\new_[10463]_ );
  assign \new_[10027]_  = ~\new_[10916]_  | ~\new_[10598]_ ;
  assign \new_[10028]_  = ~\new_[10176]_ ;
  assign \new_[10029]_  = \new_[10319]_  & \new_[10486]_ ;
  assign \new_[10030]_  = ~\new_[11218]_  | ~\new_[11920]_  | ~\new_[12044]_ ;
  assign \new_[10031]_  = ~\new_[10208]_ ;
  assign \new_[10032]_  = ~\new_[10844]_  | ~\new_[10491]_ ;
  assign \new_[10033]_  = ~\new_[10491]_  | ~\new_[10908]_ ;
  assign \new_[10034]_  = (~\new_[3884]_  | ~\new_[10598]_ ) & (~\new_[10943]_  | ~\new_[10956]_ );
  assign \new_[10035]_  = ~\new_[10339]_  & ~\new_[10858]_ ;
  assign \new_[10036]_  = ~\new_[10239]_ ;
  assign \new_[10037]_  = ~\new_[10199]_ ;
  assign \new_[10038]_  = (~\new_[3885]_  | ~\new_[10598]_ ) & (~\new_[10860]_  | ~\new_[10956]_ );
  assign \new_[10039]_  = ~\new_[10258]_ ;
  assign \new_[10040]_  = ~\new_[10417]_  & ~\new_[11493]_ ;
  assign \new_[10041]_  = ~\\u0_u0_addr_r_reg[2] ;
  assign \new_[10042]_  = \\u0_u1_addr_r_reg[2] ;
  assign \new_[10043]_  = ~\new_[11062]_  & ~\new_[10767]_ ;
  assign \new_[10044]_  = ~\new_[11062]_  & ~\new_[11329]_ ;
  assign \new_[10045]_  = \new_[10594]_  & \new_[12089]_ ;
  assign \new_[10046]_  = ~\new_[11062]_  & ~\new_[11737]_ ;
  assign \new_[10047]_  = ~\new_[10417]_  & ~\new_[12045]_ ;
  assign \new_[10048]_  = ~\new_[11062]_  & ~\new_[10799]_ ;
  assign \new_[10049]_  = ~\new_[11062]_  & ~\new_[11311]_ ;
  assign \new_[10050]_  = ~\new_[11062]_  & ~\new_[10771]_ ;
  assign \new_[10051]_  = ~\new_[10378]_  & ~\new_[11393]_ ;
  assign \new_[10052]_  = ~\new_[10262]_ ;
  assign \new_[10053]_  = ~\new_[10358]_  & ~\new_[10722]_ ;
  assign \new_[10054]_  = ~\new_[10358]_  & ~\new_[10698]_ ;
  assign \new_[10055]_  = ~\new_[11062]_  & ~\new_[10749]_ ;
  assign \new_[10056]_  = ~\new_[10378]_  & ~\new_[11314]_ ;
  assign \new_[10057]_  = ~\new_[10517]_  | ~\new_[11492]_ ;
  assign \new_[10058]_  = ~\new_[8185]_  | ~\new_[10458]_  | ~\new_[10494]_ ;
  assign \new_[10059]_  = ~\new_[10378]_  & ~\new_[12401]_ ;
  assign \new_[10060]_  = ~\new_[12054]_  & ~\new_[10704]_ ;
  assign \new_[10061]_  = ~\new_[10378]_  & ~\new_[11012]_ ;
  assign \new_[10062]_  = ~\new_[4147]_  & ~\new_[12400]_ ;
  assign \new_[10063]_  = ~\new_[10511]_  & ~\new_[10783]_ ;
  assign \new_[10064]_  = ~\new_[10417]_  & ~\new_[11299]_ ;
  assign \new_[10065]_  = ~\new_[10358]_  & ~\new_[11349]_ ;
  assign \new_[10066]_  = ~\new_[10834]_  | ~\new_[10849]_  | ~\new_[10534]_ ;
  assign \new_[10067]_  = (~\new_[3917]_  | ~\new_[10598]_ ) & (~\new_[10847]_  | ~\new_[10956]_ );
  assign \new_[10068]_  = ~\new_[10839]_  & ~\new_[12567]_ ;
  assign \new_[10069]_  = ~\new_[10869]_  | ~\new_[10598]_ ;
  assign \new_[10070]_  = (~\new_[11207]_  | ~\new_[10576]_ ) & (~\new_[11111]_  | ~\new_[10463]_ );
  assign \new_[10071]_  = ~\new_[10358]_  & ~\new_[11317]_ ;
  assign \new_[10072]_  = u5_mc_le_reg;
  assign \new_[10073]_  = ~\new_[10916]_  | ~\new_[10491]_ ;
  assign \new_[10074]_  = \new_[10604]_  | \new_[10740]_  | \new_[10644]_  | \new_[10764]_ ;
  assign \new_[10075]_  = ~\new_[10392]_  & ~\new_[10876]_ ;
  assign \new_[10076]_  = (~\new_[10844]_  | ~\new_[10598]_ ) & (~\new_[10923]_  | ~\new_[10956]_ );
  assign \new_[10077]_  = (~\new_[3889]_  | ~\new_[10598]_ ) & (~\new_[10843]_  | ~\new_[10956]_ );
  assign \new_[10078]_  = ~\new_[11062]_  & ~\new_[10752]_ ;
  assign \new_[10079]_  = ~\new_[12035]_ ;
  assign \new_[10080]_  = ~\new_[10576]_  | ~\new_[10444]_  | ~\new_[10442]_ ;
  assign \new_[10081]_  = ~\new_[10358]_  & ~\new_[11341]_ ;
  assign \new_[10082]_  = ~\new_[10358]_  & ~\new_[11321]_ ;
  assign \new_[10083]_  = ~\new_[10367]_  & ~\new_[11324]_ ;
  assign \new_[10084]_  = ~\new_[10417]_  & ~\new_[12454]_ ;
  assign \new_[10085]_  = \new_[10560]_  | \new_[10693]_  | \new_[10636]_  | \new_[10694]_ ;
  assign \new_[10086]_  = \new_[11357]_  & \new_[10827]_ ;
  assign \new_[10087]_  = ~\new_[10378]_  & ~\new_[10352]_ ;
  assign \new_[10088]_  = ~\new_[12577]_ ;
  assign \new_[10089]_  = ~\new_[11062]_  & ~\new_[10348]_ ;
  assign \new_[10090]_  = ~\new_[10159]_ ;
  assign \new_[10091]_  = ~\new_[10805]_ ;
  assign \new_[10092]_  = \new_[10325]_  | \new_[10549]_ ;
  assign \new_[10093]_  = \new_[10407]_  ? \new_[10883]_  : \new_[7730]_ ;
  assign \new_[10094]_  = \new_[10474]_  ? \new_[10898]_  : \new_[7706]_ ;
  assign \new_[10095]_  = ~\new_[10536]_  | ~\new_[10946]_  | ~\new_[10816]_ ;
  assign \new_[10096]_  = ~\new_[10845]_  | ~\new_[10491]_ ;
  assign \new_[10097]_  = ~\new_[10714]_  & ~\new_[11393]_ ;
  assign \new_[10098]_  = ~\new_[10332]_  & ~\new_[1541]_ ;
  assign \new_[10099]_  = ~\new_[10229]_ ;
  assign \new_[10100]_  = ~\new_[10852]_  | ~\new_[10491]_ ;
  assign \new_[10101]_  = ~\new_[10154]_  | ~\new_[12567]_ ;
  assign \new_[10102]_  = ~\new_[10417]_  & ~\new_[12274]_ ;
  assign \new_[10103]_  = \new_[10405]_  ? \new_[10887]_  : \new_[7960]_ ;
  assign \new_[10104]_  = ~\new_[10234]_ ;
  assign \new_[10105]_  = \new_[8081]_  ^ \new_[10483]_ ;
  assign \new_[10106]_  = ~\new_[10203]_ ;
  assign \new_[10107]_  = ~\new_[10358]_  & ~\new_[10715]_ ;
  assign \new_[10108]_  = ~\new_[10160]_ ;
  assign \new_[10109]_  = \new_[10750]_  | \new_[10695]_  | \new_[10723]_  | \new_[10620]_ ;
  assign \new_[10110]_  = \new_[11357]_  & \new_[11348]_ ;
  assign \new_[10111]_  = ~\new_[11776]_  & ~\new_[11299]_ ;
  assign \new_[10112]_  = ~\new_[10519]_  | ~\new_[10313]_ ;
  assign \new_[10113]_  = \new_[10456]_  & \new_[11335]_ ;
  assign \new_[10114]_  = \new_[10280]_  | \new_[1712]_ ;
  assign \new_[10115]_  = ~\new_[10172]_ ;
  assign \new_[10116]_  = \new_[10284]_  & \new_[10733]_ ;
  assign n5276 = \new_[3114]_  ^ \new_[10538]_ ;
  assign \new_[10118]_  = ~\new_[11062]_  & ~\new_[10724]_ ;
  assign \new_[10119]_  = ~\new_[10200]_ ;
  assign \new_[10120]_  = ~\new_[10299]_  | ~\poc_o[2] ;
  assign \new_[10121]_  = \new_[11053]_  ^ \new_[10490]_ ;
  assign \new_[10122]_  = ~\new_[10468]_  | ~\new_[10905]_  | ~\new_[10749]_ ;
  assign \new_[10123]_  = ~\new_[10920]_  & ~\new_[10288]_ ;
  assign \new_[10124]_  = ~\new_[10805]_ ;
  assign \new_[10125]_  = ~\new_[10218]_ ;
  assign \new_[10126]_  = ~\new_[11776]_  & ~\new_[11881]_ ;
  assign \new_[10127]_  = ~\new_[10378]_  & ~\new_[12400]_ ;
  assign \new_[10128]_  = ~\new_[10256]_ ;
  assign \new_[10129]_  = ~\new_[10394]_  & ~\new_[10811]_ ;
  assign \new_[10130]_  = ~\new_[11062]_  & ~\new_[10673]_ ;
  assign \new_[10131]_  = ~\new_[10817]_  | ~\new_[10491]_ ;
  assign \new_[10132]_  = ~u0_rst_r3_reg;
  assign \new_[10133]_  = ~\\u0_wb_addr_r_reg[2] ;
  assign \new_[10134]_  = ~\new_[10852]_  | ~\new_[10598]_ ;
  assign \new_[10135]_  = u6_rmw_en_reg;
  assign \new_[10136]_  = ~\new_[10167]_ ;
  assign \new_[10137]_  = ~\new_[10714]_  & ~\new_[10767]_ ;
  assign \new_[10138]_  = (~\new_[11109]_  | ~\new_[10508]_ ) & (~\new_[11176]_  | ~\new_[10502]_ );
  assign \new_[10139]_  = ~\new_[3438]_  & ~\new_[10325]_ ;
  assign \new_[10140]_  = ~\new_[11062]_  & ~\new_[11529]_ ;
  assign \new_[10141]_  = ~\new_[10587]_  & ~\new_[10364]_ ;
  assign \new_[10142]_  = (~\new_[3888]_  | ~\new_[10598]_ ) & (~\new_[10832]_  | ~\new_[10956]_ );
  assign \new_[10143]_  = \new_[12559]_  & \new_[10531]_ ;
  assign \new_[10144]_  = ~\new_[10869]_  | ~\new_[10491]_ ;
  assign \new_[10145]_  = (~\new_[3886]_  | ~\new_[10598]_ ) & (~\new_[10868]_  | ~\new_[10956]_ );
  assign \new_[10146]_  = ~\new_[10154]_  | ~\new_[10928]_ ;
  assign \new_[10147]_  = ~\new_[10285]_  & ~\new_[10592]_ ;
  assign \new_[10148]_  = ~\new_[12577]_ ;
  assign \new_[10149]_  = ~\new_[10833]_  | ~\new_[10491]_ ;
  assign \new_[10150]_  = ~\new_[10154]_  | ~\new_[12453]_ ;
  assign \new_[10151]_  = ~n5766 | ~\new_[10488]_ ;
  assign \new_[10152]_  = \new_[11359]_  & \new_[11361]_ ;
  assign \new_[10153]_  = ~\new_[10378]_  & ~\new_[12454]_ ;
  assign \new_[10154]_  = ~\new_[11776]_ ;
  assign \new_[10155]_  = ~\new_[10154]_  | ~\new_[10808]_ ;
  assign \new_[10156]_  = \new_[10896]_  & \new_[10491]_ ;
  assign \new_[10157]_  = ~\new_[10955]_  & ~\new_[10933]_ ;
  assign \new_[10158]_  = ~\new_[10528]_  | ~\new_[10508]_ ;
  assign \new_[10159]_  = ~\new_[10414]_  & ~\new_[1539]_ ;
  assign \new_[10160]_  = ~\new_[10326]_ ;
  assign \new_[10161]_  = ~\new_[11772]_ ;
  assign \new_[10162]_  = \new_[10856]_  | \new_[1454]_  | \new_[1453]_  | \new_[2070]_ ;
  assign \new_[10163]_  = ~\new_[10476]_  | ~\new_[11816]_ ;
  assign \new_[10164]_  = ~\new_[10658]_ ;
  assign \new_[10165]_  = \new_[11012]_  & \new_[11990]_ ;
  assign \new_[10166]_  = ~\new_[10154]_  | ~\new_[10964]_ ;
  assign \new_[10167]_  = ~\new_[10517]_  | ~\new_[10634]_ ;
  assign \new_[10168]_  = \new_[10473]_  & \new_[11346]_ ;
  assign \new_[10169]_  = \new_[10901]_  & \new_[10491]_ ;
  assign \new_[10170]_  = \new_[10856]_  | \new_[2056]_  | \new_[10669]_  | \new_[2070]_ ;
  assign \new_[10171]_  = ~\new_[10341]_ ;
  assign \new_[10172]_  = ~\new_[10154]_  | ~\new_[11366]_ ;
  assign \new_[10173]_  = ~\new_[10350]_ ;
  assign \new_[10174]_  = \new_[10910]_  | \new_[11053]_ ;
  assign \new_[10175]_  = \new_[10538]_  & \new_[3114]_ ;
  assign \new_[10176]_  = ~\new_[10536]_  | ~\new_[7284]_ ;
  assign \new_[10177]_  = ~\new_[10752]_ ;
  assign \new_[10178]_  = \new_[10585]_  ^ \new_[10614]_ ;
  assign \new_[10179]_  = \new_[10559]_  ^ \new_[10624]_ ;
  assign \new_[10180]_  = \new_[10612]_  ^ \new_[10631]_ ;
  assign \new_[10181]_  = \new_[10652]_  ^ \new_[10654]_ ;
  assign \new_[10182]_  = \new_[10776]_  ^ \new_[10662]_ ;
  assign \new_[10183]_  = \new_[10651]_  ^ \new_[10564]_ ;
  assign \new_[10184]_  = \new_[10699]_  ^ \new_[10711]_ ;
  assign \new_[10185]_  = \new_[10768]_  ^ \new_[10558]_ ;
  assign \new_[10186]_  = ~\new_[10428]_  & ~\new_[10979]_ ;
  assign \new_[10187]_  = ~\new_[10436]_  | ~\new_[10502]_ ;
  assign \new_[10188]_  = ~\new_[10477]_  & ~\wb_addr_i[2] ;
  assign \new_[10189]_  = ~\new_[10430]_  | ~\new_[10508]_ ;
  assign \new_[10190]_  = ~\new_[10533]_  | ~\new_[3036]_ ;
  assign \new_[10191]_  = ~\new_[10406]_  | ~\new_[10463]_ ;
  assign \new_[10192]_  = ~\new_[10513]_  | ~\new_[10463]_ ;
  assign \new_[10193]_  = \new_[1465]_  | \new_[10954]_  | \new_[1541]_  | \new_[1462]_ ;
  assign \new_[10194]_  = ~\new_[10460]_  | (~\new_[10904]_  & ~\new_[7694]_ );
  assign \new_[10195]_  = ~\new_[10283]_ ;
  assign \new_[10196]_  = \new_[10450]_  & \new_[12757]_ ;
  assign \new_[10197]_  = ~\new_[10473]_  | ~\new_[10418]_ ;
  assign \new_[10198]_  = ~\new_[11067]_  | ~\new_[10508]_ ;
  assign \new_[10199]_  = ~\new_[10154]_  | ~\new_[10919]_ ;
  assign \new_[10200]_  = \new_[10278]_ ;
  assign \new_[10201]_  = ~\new_[10433]_  | ~\new_[10398]_ ;
  assign \new_[10202]_  = ~\new_[11119]_  | ~\new_[10836]_  | ~\new_[3183]_  | ~\new_[3114]_ ;
  assign \new_[10203]_  = \new_[3388]_  | \new_[10425]_ ;
  assign \new_[10204]_  = ~\new_[11334]_  & ~\new_[10912]_ ;
  assign \new_[10205]_  = ~\new_[10313]_ ;
  assign \new_[10206]_  = \new_[10885]_  & \new_[10491]_ ;
  assign \new_[10207]_  = ~\new_[10276]_ ;
  assign \new_[10208]_  = ~\new_[10517]_  | ~\new_[10922]_ ;
  assign \new_[10209]_  = ~\new_[10316]_ ;
  assign \new_[10210]_  = ~\new_[10417]_  & ~\new_[10749]_ ;
  assign \new_[10211]_  = ~\new_[10738]_ ;
  assign \new_[10212]_  = ~\new_[11299]_  | ~\new_[12564]_ ;
  assign \new_[10213]_  = ~\new_[10747]_  | ~\new_[10402]_ ;
  assign \new_[10214]_  = ~\new_[11310]_  & ~\new_[1488]_ ;
  assign \new_[10215]_  = ~\new_[10591]_  | ~\new_[10897]_ ;
  assign \new_[10216]_  = ~\new_[10288]_ ;
  assign \new_[10217]_  = \new_[10326]_ ;
  assign \new_[10218]_  = \new_[11167]_  ? \new_[10804]_  : \new_[10851]_ ;
  assign \new_[10219]_  = \new_[10825]_  & \new_[10491]_ ;
  assign n5286 = ~\new_[12429]_ ;
  assign \new_[10221]_  = ~\new_[10398]_  & ~\new_[11167]_ ;
  assign \new_[10222]_  = ~\new_[10520]_  | ~\new_[10502]_ ;
  assign \new_[10223]_  = \new_[10553]_  & \new_[10549]_ ;
  assign \new_[10224]_  = \new_[10828]_  & \new_[10491]_ ;
  assign \new_[10225]_  = \new_[10431]_  & \new_[10861]_ ;
  assign \new_[10226]_  = ~\new_[10506]_  | (~\new_[10904]_  & ~\new_[7598]_ );
  assign \new_[10227]_  = ~\new_[10455]_  | (~\new_[10864]_  & ~\new_[7621]_ );
  assign \new_[10228]_  = ~\new_[10526]_  & ~\new_[10919]_ ;
  assign \new_[10229]_  = ~\new_[10517]_  | ~\new_[11355]_ ;
  assign \new_[10230]_  = \new_[10534]_  & \new_[8079]_ ;
  assign \new_[10231]_  = ~\new_[10356]_ ;
  assign \new_[10232]_  = \\u1_u0_out_r_reg[1] ;
  assign \new_[10233]_  = ~\new_[11991]_  | ~\new_[10584]_ ;
  assign \new_[10234]_  = ~\new_[10154]_  | ~\new_[10963]_ ;
  assign \new_[10235]_  = ~\new_[10638]_  | ~\new_[10514]_ ;
  assign \new_[10236]_  = ~\new_[10478]_  & ~\new_[10979]_ ;
  assign \new_[10237]_  = ~\new_[11776]_  & ~\new_[10673]_ ;
  assign \new_[10238]_  = \new_[10878]_  & \new_[10491]_ ;
  assign \new_[10239]_  = ~\new_[11348]_  & ~\new_[10928]_ ;
  assign \new_[10240]_  = \new_[11346]_  & \new_[10752]_ ;
  assign n5281 = \new_[9736]_  ? n5306 : \new_[11121]_ ;
  assign \new_[10242]_  = ~\new_[10477]_  & ~\new_[10979]_ ;
  assign \new_[10243]_  = ~\new_[10673]_ ;
  assign \new_[10244]_  = ~\new_[11062]_  & ~\new_[11493]_ ;
  assign \new_[10245]_  = ~\new_[10428]_  & ~\wb_addr_i[2] ;
  assign \new_[10246]_  = ~\new_[11526]_  & ~\new_[12044]_ ;
  assign \new_[10247]_  = ~\new_[11360]_  | ~\new_[12399]_ ;
  assign \new_[10248]_  = ~\new_[10409]_  | ~\new_[10532]_ ;
  assign \new_[10249]_  = ~\new_[10478]_  & ~\wb_addr_i[2] ;
  assign \new_[10250]_  = ~\new_[10552]_ ;
  assign \new_[10251]_  = ~\new_[12052]_  & ~\new_[10950]_ ;
  assign \new_[10252]_  = ~\new_[10334]_ ;
  assign \new_[10253]_  = \new_[10344]_ ;
  assign \new_[10254]_  = ~\new_[10154]_  | ~\new_[11340]_ ;
  assign \new_[10255]_  = ~\new_[1433]_  | ~\new_[10902]_ ;
  assign \new_[10256]_  = ~\new_[10517]_  | ~\new_[11576]_ ;
  assign \new_[10257]_  = ~u5_cke_o_del_reg;
  assign \new_[10258]_  = ~\new_[10154]_  | ~\new_[12273]_ ;
  assign \new_[10259]_  = \new_[12577]_  | \new_[10468]_ ;
  assign \new_[10260]_  = \new_[10414]_  | \new_[10525]_ ;
  assign \new_[10261]_  = ~\new_[10440]_  & ~\new_[10414]_ ;
  assign \new_[10262]_  = ~\new_[10287]_ ;
  assign \new_[10263]_  = ~\new_[10340]_ ;
  assign \new_[10264]_  = ~\new_[10487]_  | ~\new_[10576]_ ;
  assign \new_[10265]_  = ~\new_[10378]_  & ~\new_[12274]_ ;
  assign \new_[10266]_  = ~\new_[10708]_  | ~\new_[10930]_  | ~\new_[7416]_ ;
  assign \new_[10267]_  = ~\new_[11336]_  | ~\new_[10500]_ ;
  assign \new_[10268]_  = ~\new_[10511]_ ;
  assign \new_[10269]_  = ~\new_[10497]_  | (~\new_[10864]_  & ~\new_[7738]_ );
  assign \new_[10270]_  = ~\new_[1465]_  & ~\new_[10525]_ ;
  assign \new_[10271]_  = ~\new_[10550]_  & ~\new_[10656]_ ;
  assign \new_[10272]_  = ~\new_[10590]_  & ~\new_[10761]_ ;
  assign \new_[10273]_  = \new_[10917]_  ? \new_[10913]_  : \new_[7601]_ ;
  assign \new_[10274]_  = \new_[12454]_  & \new_[10575]_ ;
  assign \new_[10275]_  = ~\new_[10452]_ ;
  assign \new_[10276]_  = ~\new_[12184]_  & ~\new_[10922]_ ;
  assign \new_[10277]_  = \\u0_spec_req_cs_reg[5] ;
  assign \new_[10278]_  = ~\new_[10522]_ ;
  assign \new_[10279]_  = \\u0_cs_reg[6] ;
  assign \new_[10280]_  = ~\new_[10895]_  | ~\new_[10861]_  | ~\new_[11071]_ ;
  assign \new_[10281]_  = ~\new_[10649]_  & ~\new_[10639]_ ;
  assign \new_[10282]_  = u0_u1_rst_r2_reg;
  assign \new_[10283]_  = ~\new_[10420]_ ;
  assign \new_[10284]_  = \new_[10842]_  & \new_[10979]_ ;
  assign \new_[10285]_  = \new_[6409]_  ^ \new_[2721]_ ;
  assign \new_[10286]_  = ~\new_[10704]_  | ~\new_[12555]_ ;
  assign \new_[10287]_  = ~\new_[11776]_  & ~\new_[11317]_ ;
  assign \new_[10288]_  = ~\new_[10475]_ ;
  assign \new_[10289]_  = \\u0_spec_req_cs_reg[4] ;
  assign \new_[10291]_  = ~\new_[10402]_ ;
  assign n5311 = u0_rst_r2_reg;
  assign \new_[10293]_  = ~\new_[10545]_  & ~\new_[10700]_ ;
  assign \new_[10294]_  = ~\new_[10621]_  & ~\new_[10625]_ ;
  assign \new_[10295]_  = ~\new_[10745]_  & ~\new_[10803]_ ;
  assign \new_[10296]_  = \new_[10875]_  ? \new_[10973]_  : \new_[7703]_ ;
  assign \new_[10297]_  = \new_[3440]_  ^ \new_[10857]_ ;
  assign \new_[10298]_  = ~\new_[10536]_ ;
  assign \new_[10299]_  = u0_u0_rst_r2_reg;
  assign \new_[10300]_  = ~\new_[10412]_ ;
  assign \new_[10301]_  = \new_[10786]_  & \new_[11321]_ ;
  assign \new_[10302]_  = ~\new_[10617]_  & ~\new_[3184]_ ;
  assign \new_[10303]_  = ~\new_[10671]_  & ~\new_[10736]_ ;
  assign \new_[10304]_  = ~\new_[11955]_  & ~\new_[10772]_ ;
  assign \new_[10305]_  = ~\new_[10553]_  | ~\new_[10583]_ ;
  assign \new_[10306]_  = ~\new_[8179]_  | ~\new_[10713]_  | ~\new_[7620]_ ;
  assign \new_[10307]_  = \new_[10801]_  | \new_[10883]_ ;
  assign \new_[10308]_  = ~\new_[8198]_  | ~\new_[10543]_  | ~\new_[7737]_ ;
  assign \new_[10309]_  = ~\new_[10425]_ ;
  assign \new_[10310]_  = ~\new_[3036]_ ;
  assign \new_[10311]_  = \\u0_cs_reg[7] ;
  assign n5321 = ~\new_[10510]_ ;
  assign \new_[10313]_  = ~\\u0_wb_addr_r_reg[3] ;
  assign \new_[10314]_  = ~\new_[10441]_ ;
  assign \new_[10315]_  = ~\new_[10563]_  & ~\new_[10611]_ ;
  assign \new_[10316]_  = ~\new_[11338]_  | ~\new_[10677]_  | ~\new_[12611]_ ;
  assign \new_[10317]_  = ~\new_[10669]_  & ~\new_[10856]_ ;
  assign \new_[10318]_  = \new_[10676]_  & \new_[11364]_ ;
  assign \new_[10319]_  = ~\new_[10743]_  & ~\new_[10892]_ ;
  assign \new_[10320]_  = \new_[10418]_ ;
  assign \new_[10321]_  = ~\new_[10599]_  & ~\new_[10697]_ ;
  assign \new_[10322]_  = \new_[10409]_ ;
  assign \new_[10323]_  = ~\new_[10658]_  | ~\new_[11364]_ ;
  assign \new_[10324]_  = \\u0_cs_reg[4] ;
  assign \new_[10325]_  = ~\new_[3036]_  & ~\new_[10583]_ ;
  assign \new_[10326]_  = \new_[10906]_ ;
  assign \new_[10327]_  = \\u0_spec_req_cs_reg[7] ;
  assign \new_[10328]_  = ~\new_[10634]_ ;
  assign \new_[10329]_  = ~\new_[10568]_  & ~\new_[10692]_ ;
  assign \new_[10330]_  = \\u0_cs_reg[3] ;
  assign \new_[10331]_  = ~\new_[8196]_  | ~\new_[10748]_  | ~\new_[7812]_ ;
  assign \new_[10332]_  = ~\new_[11219]_  | ~\new_[11209]_  | ~\new_[11129]_  | ~\new_[10853]_ ;
  assign \new_[10333]_  = \\u0_spec_req_cs_reg[6] ;
  assign \new_[10334]_  = ~\new_[10500]_ ;
  assign \new_[10335]_  = ~\new_[10773]_  & (~\new_[1541]_  | ~\new_[1465]_ );
  assign \new_[10336]_  = ~\new_[10666]_  & ~\new_[12564]_ ;
  assign \new_[10337]_  = \new_[10966]_  ? \new_[10973]_  : \new_[7704]_ ;
  assign \new_[10338]_  = \new_[10889]_  ? \new_[10854]_  : \new_[7702]_ ;
  assign \new_[10339]_  = ~\\u0_u1_addr_r_reg[3] ;
  assign \new_[10340]_  = ~\new_[10154]_  | ~\new_[11343]_ ;
  assign \new_[10341]_  = ~\new_[10601]_  & ~\new_[1644]_ ;
  assign \new_[10342]_  = ~\new_[10490]_ ;
  assign \new_[10343]_  = ~\new_[10414]_ ;
  assign \new_[10344]_  = ~\new_[10666]_  & ~\new_[10689]_ ;
  assign \new_[10345]_  = ~\new_[11492]_  & ~\new_[11341]_ ;
  assign \new_[10346]_  = \new_[10677]_  & \new_[10554]_ ;
  assign \new_[10347]_  = \\u0_cs_reg[2] ;
  assign \new_[10348]_  = ~\new_[10933]_ ;
  assign \new_[10349]_  = ~\new_[10682]_  & (~\new_[4145]_  | ~\new_[3881]_ );
  assign \new_[10350]_  = ~\new_[10669]_  & ~\new_[1519]_ ;
  assign \new_[10351]_  = \\u0_spec_req_cs_reg[3] ;
  assign \new_[10352]_  = ~\new_[10411]_ ;
  assign \new_[10353]_  = ~\new_[7278]_  | ~\new_[7416]_  | ~\new_[7265]_ ;
  assign \new_[10354]_  = \\u1_u0_out_r_reg[0] ;
  assign \new_[10355]_  = ~\new_[10640]_  & ~\new_[10257]_ ;
  assign \new_[10356]_  = \new_[10549]_  | \new_[10369]_ ;
  assign \new_[10357]_  = ~\new_[10574]_  & ~\new_[10742]_ ;
  assign \new_[10358]_  = ~\new_[8862]_ ;
  assign \new_[10359]_  = ~\new_[10534]_ ;
  assign \new_[10360]_  = \\u0_cs_reg[5] ;
  assign \new_[10361]_  = ~\new_[10617]_  & ~\new_[10736]_ ;
  assign \new_[10362]_  = ~\new_[10701]_  & ~\new_[10760]_ ;
  assign \new_[10363]_  = ~\new_[10709]_  & ~\new_[10678]_ ;
  assign \new_[10364]_  = \new_[6644]_  ^ \new_[2721]_ ;
  assign \new_[10365]_  = ~\new_[10696]_  & ~\new_[10686]_ ;
  assign \new_[10366]_  = ~\new_[10555]_  & ~\new_[10739]_ ;
  assign \new_[10367]_  = ~\new_[10517]_ ;
  assign \new_[10368]_  = \\u0_spec_req_cs_reg[2] ;
  assign \new_[10369]_  = u0_init_req_reg;
  assign \new_[10370]_  = ~\new_[10670]_  & ~\new_[7618]_ ;
  assign \new_[10371]_  = ~\new_[10841]_  | ~\new_[10665]_ ;
  assign \new_[10372]_  = ~\new_[10582]_  & ~\new_[10635]_ ;
  assign \new_[10373]_  = ~\new_[10595]_  & ~\new_[10781]_ ;
  assign \new_[10374]_  = ~\new_[11329]_  & ~\new_[11366]_ ;
  assign \new_[10375]_  = ~\new_[10626]_  & ~\new_[10810]_ ;
  assign \new_[10376]_  = ~\new_[10629]_  & ~\new_[10655]_ ;
  assign \new_[10377]_  = ~\new_[10788]_  & ~\new_[10645]_ ;
  assign \new_[10378]_  = ~\new_[10594]_ ;
  assign \new_[10379]_  = ~\new_[10794]_  & ~\new_[10597]_ ;
  assign \new_[10380]_  = ~\new_[10687]_  & ~\new_[10593]_ ;
  assign \new_[10381]_  = ~\new_[10734]_  & ~\new_[1955]_ ;
  assign \new_[10382]_  = ~\new_[10784]_  & ~\new_[10792]_ ;
  assign \new_[10383]_  = ~\new_[12097]_ ;
  assign \new_[10384]_  = ~\new_[10573]_  & ~\new_[10610]_ ;
  assign \new_[10385]_  = ~\new_[10720]_  & ~\new_[10769]_ ;
  assign \new_[10386]_  = ~\new_[10703]_  & ~\new_[10681]_ ;
  assign \new_[10387]_  = ~\new_[10588]_  & ~\new_[10806]_ ;
  assign \new_[10388]_  = ~\new_[10780]_  & ~\new_[10628]_ ;
  assign \new_[10389]_  = \new_[10542]_  | \new_[10887]_ ;
  assign \new_[10390]_  = ~\new_[10571]_  | ~\new_[8185]_ ;
  assign \new_[10391]_  = ~\new_[10728]_  & ~\new_[10758]_ ;
  assign \new_[10392]_  = \\u0_u0_addr_r_reg[3] ;
  assign \new_[10393]_  = ~\new_[10529]_ ;
  assign \new_[10394]_  = \new_[10608]_  | \new_[10893]_ ;
  assign \new_[10395]_  = ~\new_[11241]_  | ~\new_[10949]_ ;
  assign \new_[10396]_  = ~\new_[10964]_  & ~\new_[10960]_ ;
  assign \new_[10397]_  = ~\new_[10892]_ ;
  assign \new_[10398]_  = \new_[10813]_  | \new_[2494]_ ;
  assign \new_[10399]_  = ~\new_[8061]_  | ~\new_[10949]_ ;
  assign \new_[10400]_  = ~\new_[10891]_  & ~\wb_addr_i[31] ;
  assign \new_[10401]_  = ~\new_[10578]_ ;
  assign \new_[10402]_  = ~\new_[1480]_ ;
  assign \new_[10403]_  = ~\new_[10913]_  | ~\new_[11065]_ ;
  assign \new_[10404]_  = ~\new_[11493]_  & ~\new_[11340]_ ;
  assign \new_[10405]_  = ~\new_[7960]_  | ~\new_[8201]_ ;
  assign \new_[10406]_  = ~\new_[10848]_  | (~\new_[6417]_  & ~\new_[2841]_ );
  assign \new_[10407]_  = ~\new_[7730]_  | ~\new_[8199]_ ;
  assign \new_[10408]_  = \new_[11063]_  ^ \new_[2769]_ ;
  assign \new_[10409]_  = ~\new_[10562]_ ;
  assign \new_[10410]_  = ~\new_[8068]_  | ~\new_[10949]_ ;
  assign \new_[10411]_  = ~\new_[10676]_ ;
  assign \new_[10412]_  = \new_[10829]_  | \wb_addr_i[31] ;
  assign \new_[10413]_  = \new_[11139]_  ^ \new_[2769]_ ;
  assign \new_[10414]_  = \new_[10944]_  | \new_[1462]_ ;
  assign \new_[10415]_  = ~\new_[10887]_  | ~\new_[11031]_ ;
  assign \new_[10416]_  = ~\new_[10857]_  | ~\new_[10936]_ ;
  assign \new_[10417]_  = ~\new_[12577]_ ;
  assign \new_[10418]_  = ~\new_[10641]_ ;
  assign \new_[10419]_  = ~\new_[10771]_ ;
  assign \new_[10420]_  = ~\new_[10804]_ ;
  assign \new_[10421]_  = ~\new_[10854]_  | ~\new_[11030]_ ;
  assign \new_[10422]_  = ~\new_[10854]_  | ~\new_[11214]_ ;
  assign \new_[10423]_  = ~\new_[11093]_  | ~\new_[10949]_ ;
  assign \new_[10424]_  = ~\new_[10887]_  | ~\new_[11130]_ ;
  assign \new_[10425]_  = \new_[3440]_  | \new_[10936]_ ;
  assign \new_[10426]_  = ~\new_[10883]_  | ~\new_[11174]_ ;
  assign \new_[10427]_  = \new_[11180]_  ^ \new_[11133]_ ;
  assign \new_[10428]_  = ~\wb_addr_i[4]  | ~\new_[10842]_  | ~\wb_addr_i[3] ;
  assign \new_[10429]_  = ~\new_[10898]_  | ~\new_[11108]_ ;
  assign \new_[10430]_  = ~\new_[10862]_  | (~\new_[6446]_  & ~\new_[2843]_ );
  assign \new_[10431]_  = ~\new_[1644]_  & ~\new_[1657]_ ;
  assign \new_[10432]_  = ~\new_[10728]_ ;
  assign \new_[10433]_  = ~\new_[2478]_  | ~\new_[11159]_  | ~\new_[11073]_ ;
  assign \new_[10434]_  = ~\new_[10973]_  | ~\new_[11029]_ ;
  assign \new_[10435]_  = \new_[11025]_  ^ \new_[11133]_ ;
  assign \new_[10436]_  = ~\new_[10903]_  | (~\new_[6529]_  & ~\new_[2841]_ );
  assign \new_[10437]_  = ~\new_[8072]_  | ~\new_[10949]_ ;
  assign \new_[10438]_  = ~\new_[11737]_  & ~\new_[10962]_ ;
  assign \new_[10439]_  = \\u0_csr_r_reg[0] ;
  assign \new_[10440]_  = \new_[1582]_  | \new_[10954]_ ;
  assign \new_[10441]_  = ~\new_[10657]_ ;
  assign \new_[10442]_  = ~\new_[10953]_  | (~\new_[6331]_  & ~\new_[2841]_ );
  assign \new_[10443]_  = ~\new_[10898]_  | ~\new_[11181]_ ;
  assign \new_[10444]_  = ~\new_[10870]_  | (~\new_[6471]_  & ~\new_[2830]_ );
  assign \new_[10445]_  = ~u6_read_go_r_reg;
  assign \new_[10446]_  = \new_[10857]_  | \new_[11148]_ ;
  assign \new_[10447]_  = ~\new_[10864]_  & ~\new_[8200]_ ;
  assign \new_[10448]_  = ~\new_[10913]_  | ~\new_[11072]_ ;
  assign \new_[10449]_  = \new_[10927]_  & \new_[10914]_ ;
  assign \new_[10450]_  = ~\new_[10568]_ ;
  assign \new_[10451]_  = ~\new_[7382]_  | ~\new_[10890]_  | ~\new_[11192]_ ;
  assign \new_[10452]_  = \new_[12184]_  & \new_[10922]_ ;
  assign \new_[10453]_  = ~\new_[8023]_  | ~\new_[10949]_ ;
  assign \new_[10454]_  = \new_[10822]_  & \new_[10816]_ ;
  assign \new_[10455]_  = ~\new_[8200]_  | ~\new_[10864]_  | ~\new_[7621]_ ;
  assign \new_[10456]_  = ~\new_[10906]_  & ~\new_[10897]_ ;
  assign \new_[10457]_  = \new_[11147]_  ^ \new_[2769]_ ;
  assign \new_[10458]_  = ~\new_[10837]_  & (~\new_[7617]_  | ~\new_[10369]_ );
  assign \new_[10459]_  = \new_[11004]_  ^ \new_[2769]_ ;
  assign \new_[10460]_  = ~\new_[7694]_  | ~\new_[10904]_  | ~\new_[8149]_ ;
  assign \new_[10461]_  = ~\new_[10805]_ ;
  assign \new_[10462]_  = ~\new_[11043]_  | ~\new_[10949]_ ;
  assign \new_[10463]_  = ~\new_[2719]_  & ~\new_[11179]_ ;
  assign \new_[10464]_  = ~\new_[11082]_  | ~\new_[10949]_ ;
  assign \new_[10465]_  = ~\new_[11028]_  | ~\new_[10949]_ ;
  assign \new_[10466]_  = ~\new_[10758]_ ;
  assign \new_[10467]_  = \new_[7624]_  & \new_[10949]_ ;
  assign \new_[10468]_  = ~\new_[10689]_ ;
  assign \new_[10469]_  = \new_[10872]_  & \new_[11300]_ ;
  assign \new_[10470]_  = ~\new_[10666]_ ;
  assign \new_[10471]_  = ~\new_[10731]_ ;
  assign \new_[10472]_  = \new_[7595]_  & \new_[10949]_ ;
  assign \new_[10473]_  = ~\new_[10556]_ ;
  assign \new_[10474]_  = ~\new_[7706]_  | ~\new_[8198]_ ;
  assign \new_[10475]_  = ~\new_[10807]_ ;
  assign \new_[10476]_  = u0_lmr_ack_r_reg;
  assign \new_[10477]_  = ~\wb_addr_i[4]  | ~\new_[10842]_  | ~\new_[11189]_ ;
  assign \new_[10478]_  = ~\new_[10824]_  | ~\new_[10842]_ ;
  assign \new_[10479]_  = \new_[7625]_  & \new_[10949]_ ;
  assign \new_[10480]_  = ~\new_[10883]_  | ~\new_[11246]_ ;
  assign \new_[10481]_  = ~wb_we_i | ~\new_[10851]_ ;
  assign \new_[10482]_  = \new_[11183]_  ^ \new_[2769]_ ;
  assign \new_[10483]_  = ~\new_[8071]_  | ~\new_[7977]_  | ~\new_[10849]_  | ~\new_[8077]_ ;
  assign \new_[10484]_  = \new_[11123]_  ^ \new_[2769]_ ;
  assign \new_[10485]_  = ~\new_[10743]_ ;
  assign \new_[10486]_  = ~\new_[10561]_ ;
  assign \new_[10487]_  = ~\new_[10909]_  | (~\new_[6434]_  & ~\new_[2841]_ );
  assign \new_[10488]_  = ~\new_[10735]_ ;
  assign \new_[10489]_  = ~\new_[11234]_  | ~\new_[10949]_ ;
  assign \new_[10490]_  = \new_[11033]_  | \new_[10910]_ ;
  assign \new_[10491]_  = ~\new_[10665]_ ;
  assign \new_[10492]_  = ~\new_[11223]_  | ~\new_[10949]_ ;
  assign \new_[10493]_  = ~\new_[11334]_  | ~\new_[10912]_ ;
  assign \new_[10494]_  = ~\new_[10571]_ ;
  assign \new_[10495]_  = ~\new_[8809]_  | ~\new_[10948]_ ;
  assign \new_[10496]_  = ~\new_[10575]_ ;
  assign \new_[10497]_  = ~\new_[8200]_  | ~\new_[10864]_  | ~\new_[7738]_ ;
  assign \new_[10498]_  = ~\new_[3225]_  | ~\new_[3176]_  | ~\new_[3169]_  | ~\new_[3177]_ ;
  assign \new_[10499]_  = ~\new_[10888]_  | ~\new_[8410]_ ;
  assign \new_[10500]_  = ~\new_[10623]_ ;
  assign \new_[10501]_  = u0_lmr_req_reg;
  assign \new_[10502]_  = ~\new_[2719]_  & ~\new_[2767]_ ;
  assign \new_[10503]_  = ~\new_[11329]_  | ~\new_[11366]_ ;
  assign \new_[10504]_  = ~\new_[11105]_  & ~\new_[10899]_ ;
  assign \new_[10505]_  = ~\new_[1580]_  & ~\new_[1581]_ ;
  assign \new_[10506]_  = ~\new_[7598]_  | ~\new_[10904]_  | ~\new_[8149]_ ;
  assign \new_[10507]_  = ~\new_[10861]_  & (~\new_[1841]_  | ~\new_[1656]_ );
  assign \new_[10508]_  = ~\new_[11080]_  & ~\new_[2767]_ ;
  assign \new_[10509]_  = ~\new_[10754]_ ;
  assign \new_[10510]_  = ~wb_ack_o & (~\new_[10135]_  | ~wb_cyc_i);
  assign \new_[10511]_  = ~\new_[8862]_ ;
  assign \new_[10512]_  = \new_[10934]_  & \new_[10369]_ ;
  assign \new_[10513]_  = ~\new_[10815]_  | (~\new_[6385]_  & ~\new_[2841]_ );
  assign \new_[10514]_  = ~\new_[10746]_ ;
  assign \new_[10515]_  = ~\new_[10904]_  & ~\new_[8149]_ ;
  assign \new_[10516]_  = ~\new_[10963]_  & ~\new_[11576]_ ;
  assign \new_[10517]_  = ~\new_[10714]_ ;
  assign \new_[10518]_  = ~\new_[10859]_  & (~\new_[1453]_  | ~\new_[1454]_ );
  assign \new_[10519]_  = ~\new_[10958]_  & ~\new_[10840]_ ;
  assign \new_[10520]_  = ~\new_[10951]_  | (~\new_[6523]_  & ~\new_[2841]_ );
  assign \new_[10521]_  = \new_[10952]_  & \new_[10971]_ ;
  assign \new_[10522]_  = ~\new_[2055]_ ;
  assign \new_[10523]_  = ~\new_[10893]_  & ~\new_[7813]_ ;
  assign \new_[10524]_  = ~\new_[10894]_  | (~\new_[7966]_  & ~\new_[8390]_ );
  assign \new_[10525]_  = \new_[10880]_  | \new_[10954]_ ;
  assign \new_[10526]_  = ~\new_[10715]_ ;
  assign n5021 = ~\new_[10749]_ ;
  assign \new_[10528]_  = ~\new_[10924]_  | (~\new_[6424]_  & ~\new_[2842]_ );
  assign \new_[10529]_  = ~\new_[10657]_ ;
  assign n5331 = u5_cke_o_r2_reg;
  assign \new_[10531]_  = \new_[10989]_  & \new_[12094]_ ;
  assign \new_[10532]_  = ~\new_[10738]_ ;
  assign \new_[10533]_  = ~u5_cs_le_r_reg;
  assign \new_[10534]_  = \new_[8077]_  & \new_[8071]_ ;
  assign \new_[10535]_  = \new_[8077]_  ^ \new_[8071]_ ;
  assign \new_[10536]_  = \new_[7416]_  & \new_[7285]_ ;
  assign \new_[10537]_  = \new_[7416]_  ^ \new_[7285]_ ;
  assign \new_[10538]_  = \new_[3182]_  & \new_[3183]_ ;
  assign n5326 = \new_[3182]_  ^ \new_[3183]_ ;
  assign \new_[10540]_  = ~\new_[8051]_  | ~\new_[11238]_ ;
  assign n5336 = ~\new_[8185]_  & ~\new_[11185]_ ;
  assign \new_[10542]_  = \new_[11130]_  | \new_[11031]_ ;
  assign \new_[10543]_  = ~\new_[10898]_ ;
  assign \mc_data_pad_o[8]  = \\u7_mc_data_o_reg[8] ;
  assign \new_[10545]_  = \new_[6412]_  ^ \new_[2829]_ ;
  assign \mc_dp_pad_o[3]  = \\u7_mc_dp_o_reg[3] ;
  assign \mc_dp_pad_o[2]  = \\u7_mc_dp_o_reg[2] ;
  assign \mc_data_pad_o[6]  = \\u7_mc_data_o_reg[6] ;
  assign \new_[10549]_  = ~\new_[10821]_ ;
  assign \new_[10550]_  = \new_[8378]_  ^ \new_[8049]_ ;
  assign \new_[10551]_  = ~\new_[10818]_ ;
  assign \new_[10552]_  = ~\new_[10873]_ ;
  assign \new_[10553]_  = ~\new_[3438]_  & ~\new_[10369]_ ;
  assign \new_[10554]_  = \new_[11314]_  & \new_[12401]_ ;
  assign \new_[10555]_  = \new_[6582]_  ^ \new_[2721]_ ;
  assign \new_[10556]_  = ~\new_[11322]_  | ~\new_[11165]_ ;
  assign n5406 = ~n5766 & ~\new_[11161]_ ;
  assign \new_[10558]_  = \wb_data_i[23]  ^ \wb_data_i[16] ;
  assign \new_[10559]_  = \wb_data_i[6]  ^ \wb_data_i[1] ;
  assign \new_[10560]_  = \new_[6542]_  ^ \new_[2839]_ ;
  assign \new_[10561]_  = ~\new_[11150]_  | ~\new_[11252]_ ;
  assign \new_[10562]_  = ~\new_[11330]_  | ~\new_[11369]_ ;
  assign \new_[10563]_  = \new_[6401]_  ^ \new_[2830]_ ;
  assign \new_[10564]_  = \wb_data_i[31]  ^ \wb_data_i[24] ;
  assign \mc_data_pad_o[19]  = \\u7_mc_data_o_reg[19] ;
  assign \mc_data_pad_o[31]  = \\u7_mc_data_o_reg[31] ;
  assign \new_[10567]_  = ~\new_[11245]_  | ~\new_[11238]_ ;
  assign \new_[10568]_  = ~\new_[12600]_  | ~\new_[12612]_ ;
  assign n5421 = ~n5766 & ~\new_[11135]_ ;
  assign \new_[10570]_  = \new_[6513]_  ^ \new_[2842]_ ;
  assign \new_[10571]_  = \new_[7626]_  ? \new_[10369]_  : \new_[7280]_ ;
  assign \new_[10572]_  = ~u5_resume_req_r_reg;
  assign \new_[10573]_  = \new_[6425]_  ^ \new_[2845]_ ;
  assign \new_[10574]_  = \new_[6575]_  ^ \new_[2830]_ ;
  assign \new_[10575]_  = ~\new_[10866]_ ;
  assign \new_[10576]_  = ~\new_[11080]_  & ~\new_[11179]_ ;
  assign \new_[10577]_  = ~\new_[8048]_  | ~\new_[11238]_ ;
  assign \new_[10578]_  = ~\new_[10990]_  | ~\new_[11124]_ ;
  assign \new_[10579]_  = ~\new_[10955]_ ;
  assign n5391 = ~n5766 & ~\new_[11052]_ ;
  assign \mc_data_pad_o[26]  = \\u7_mc_data_o_reg[26] ;
  assign \new_[10582]_  = \new_[6445]_  ^ \new_[2842]_ ;
  assign \new_[10583]_  = ~u5_susp_req_r_reg;
  assign \new_[10584]_  = \new_[11039]_  & \new_[11078]_ ;
  assign \new_[10585]_  = \wb_data_i[12]  ^ \wb_data_i[10] ;
  assign \mc_data_pad_o[28]  = \\u7_mc_data_o_reg[28] ;
  assign \new_[10587]_  = \new_[6614]_  ^ \new_[2845]_ ;
  assign \new_[10588]_  = \new_[6403]_  ^ \new_[2768]_ ;
  assign \mc_data_pad_o[18]  = \\u7_mc_data_o_reg[18] ;
  assign \new_[10590]_  = \new_[6382]_  ^ \new_[2768]_ ;
  assign \new_[10591]_  = ~\new_[10906]_ ;
  assign \new_[10592]_  = \new_[6414]_  ^ \new_[2768]_ ;
  assign \new_[10593]_  = \new_[6386]_  ^ \new_[2830]_ ;
  assign \new_[10594]_  = ~\new_[11062]_ ;
  assign \new_[10595]_  = \new_[6413]_  ^ \new_[2842]_ ;
  assign n5411 = ~\new_[8185]_  & ~\new_[11057]_ ;
  assign \new_[10597]_  = \new_[6454]_  ^ \new_[2845]_ ;
  assign \new_[10598]_  = ~\new_[10841]_ ;
  assign \new_[10599]_  = \new_[6550]_  ^ \new_[2720]_ ;
  assign \new_[10600]_  = \new_[6330]_  ^ \new_[2839]_ ;
  assign \new_[10601]_  = ~\new_[10861]_ ;
  assign \new_[10602]_  = \new_[6467]_  ^ \new_[2839]_ ;
  assign n5361 = u0_rst_r1_reg;
  assign \new_[10604]_  = \new_[6562]_  ^ \new_[2839]_ ;
  assign \new_[10605]_  = ~\new_[11249]_  | ~\new_[11238]_ ;
  assign n5386 = ~\new_[8185]_  & ~\new_[10977]_ ;
  assign \mc_data_pad_o[5]  = \\u7_mc_data_o_reg[5] ;
  assign \new_[10608]_  = ~\new_[11257]_  | ~\new_[7850]_ ;
  assign \mc_data_pad_o[30]  = \\u7_mc_data_o_reg[30] ;
  assign \new_[10610]_  = \new_[6420]_  ^ \new_[2720]_ ;
  assign \new_[10611]_  = \new_[6435]_  ^ \new_[2843]_ ;
  assign \new_[10612]_  = \wb_data_i[22]  ^ \wb_data_i[17] ;
  assign \new_[10613]_  = \new_[6404]_  ^ \new_[2842]_ ;
  assign \new_[10614]_  = \wb_data_i[15]  ^ \wb_data_i[8] ;
  assign \new_[10615]_  = \new_[6653]_  ^ \new_[2833]_ ;
  assign \new_[10616]_  = ~\new_[11188]_  | ~\new_[11238]_ ;
  assign \new_[10617]_  = ~\new_[11146]_  | ~\new_[11100]_ ;
  assign \new_[10618]_  = ~\new_[3182]_  | ~\new_[11100]_ ;
  assign \new_[10619]_  = \new_[6429]_  ^ \new_[2842]_ ;
  assign \new_[10620]_  = \new_[6439]_  ^ \new_[2839]_ ;
  assign \new_[10621]_  = \new_[6408]_  ^ \new_[2720]_ ;
  assign \new_[10622]_  = ~\new_[8067]_  | ~\new_[11238]_ ;
  assign \new_[10623]_  = ~\new_[11184]_  | ~\new_[11034]_ ;
  assign \new_[10624]_  = \wb_data_i[5]  ^ \wb_data_i[3] ;
  assign \new_[10625]_  = \new_[6633]_  ^ \new_[2845]_ ;
  assign \new_[10626]_  = \new_[6335]_  ^ \new_[2768]_ ;
  assign n5351 = ~\new_[8185]_  & ~\new_[11255]_ ;
  assign \new_[10628]_  = \new_[8352]_  ^ \new_[8077]_ ;
  assign \new_[10629]_  = \new_[6458]_  ^ \new_[2720]_ ;
  assign n5366 = u0_u0_rst_r1_reg;
  assign \new_[10631]_  = \wb_data_i[21]  ^ \wb_data_i[19] ;
  assign \mc_data_pad_o[22]  = \\u7_mc_data_o_reg[22] ;
  assign \mc_data_pad_o[16]  = \\u7_mc_data_o_reg[16] ;
  assign \new_[10634]_  = ~\new_[11889]_ ;
  assign \new_[10635]_  = \new_[6444]_  ^ \new_[2841]_ ;
  assign \new_[10636]_  = \new_[6490]_  ^ \new_[2829]_ ;
  assign \mc_data_pad_o[11]  = \\u7_mc_data_o_reg[11] ;
  assign \new_[10638]_  = \new_[11378]_  & \new_[11195]_ ;
  assign \new_[10639]_  = \new_[6518]_  ^ \new_[2830]_ ;
  assign \new_[10640]_  = ~\new_[11058]_  | ~\new_[3036]_ ;
  assign \new_[10641]_  = ~\new_[11494]_  | ~\new_[11342]_ ;
  assign \new_[10642]_  = \new_[6341]_  ^ \new_[2829]_ ;
  assign \new_[10643]_  = \new_[6387]_  ^ \new_[2843]_ ;
  assign \new_[10644]_  = \new_[6427]_  ^ \new_[2829]_ ;
  assign \new_[10645]_  = \new_[6453]_  ^ \new_[2843]_ ;
  assign \new_[10646]_  = \new_[6451]_  ^ \new_[2842]_ ;
  assign \new_[10647]_  = \new_[6647]_  ^ \new_[2840]_ ;
  assign \new_[10648]_  = \new_[8260]_  ^ \new_[7977]_ ;
  assign \new_[10649]_  = \new_[6537]_  ^ \new_[2843]_ ;
  assign \new_[10650]_  = \new_[6443]_  ^ \new_[2840]_ ;
  assign \new_[10651]_  = \wb_data_i[28]  ^ \wb_data_i[26] ;
  assign \new_[10652]_  = \wb_data_i[29]  ^ \wb_data_i[27] ;
  assign \new_[10653]_  = \new_[8400]_  ^ \new_[8081]_ ;
  assign \new_[10654]_  = \wb_data_i[30]  ^ \wb_data_i[25] ;
  assign \new_[10655]_  = \new_[6430]_  ^ \new_[2721]_ ;
  assign \new_[10656]_  = \new_[8071]_  ^ \new_[8296]_ ;
  assign \new_[10657]_  = ~\new_[10957]_ ;
  assign \new_[10658]_  = ~\new_[10905]_ ;
  assign \mc_data_pad_o[21]  = \\u7_mc_data_o_reg[21] ;
  assign \mc_data_pad_o[7]  = \\u7_mc_data_o_reg[7] ;
  assign n5371 = ~n5766 & ~\new_[11158]_ ;
  assign \new_[10662]_  = \wb_data_i[14]  ^ \wb_data_i[9] ;
  assign \new_[10663]_  = ~\new_[11022]_  | ~\new_[11238]_ ;
  assign n5396 = ~\new_[8185]_  & ~\new_[11231]_ ;
  assign \new_[10665]_  = ~\new_[2316]_  | ~\new_[10996]_ ;
  assign \new_[10666]_  = ~\new_[11193]_  | ~\new_[10989]_ ;
  assign \new_[10667]_  = ~\new_[11240]_  | ~\new_[11238]_ ;
  assign n5426 = ~\new_[8185]_  & ~\new_[11040]_ ;
  assign \new_[10669]_  = ~\new_[10859]_ ;
  assign \new_[10670]_  = ~\new_[10890]_ ;
  assign \new_[10671]_  = ~\new_[11205]_  | ~\new_[11051]_ ;
  assign \new_[10672]_  = ~\new_[8078]_  | ~\new_[11238]_ ;
  assign \new_[10673]_  = ~\new_[10871]_ ;
  assign \new_[10674]_  = ~\new_[8043]_  | ~\new_[11238]_ ;
  assign \mc_data_pad_o[20]  = \\u7_mc_data_o_reg[20] ;
  assign \new_[10676]_  = ~\new_[1526]_ ;
  assign \new_[10677]_  = \new_[12599]_  & \new_[12757]_ ;
  assign \new_[10678]_  = \new_[6329]_  ^ \new_[2720]_ ;
  assign \new_[10679]_  = ~\new_[10310]_ ;
  assign \new_[10680]_  = \new_[6405]_  ^ \new_[2840]_ ;
  assign \new_[10681]_  = \new_[6407]_  ^ \new_[2833]_ ;
  assign \new_[10682]_  = ~\new_[10910]_ ;
  assign \new_[10683]_  = ~\new_[3181]_ ;
  assign \new_[10684]_  = \new_[8232]_  ^ \new_[8075]_ ;
  assign \new_[10685]_  = \new_[3398]_  ^ \new_[3439]_ ;
  assign \new_[10686]_  = \new_[6419]_  ^ \new_[2768]_ ;
  assign \new_[10687]_  = \new_[6388]_  ^ \new_[2842]_ ;
  assign n5346 = u0_u1_rst_r1_reg;
  assign \new_[10689]_  = ~\new_[12560]_  | ~\new_[12095]_ ;
  assign \new_[10690]_  = ~\new_[11318]_  | ~\new_[12178]_ ;
  assign \new_[10691]_  = ~\new_[10826]_ ;
  assign \new_[10692]_  = ~\new_[12758]_  | ~\new_[11339]_ ;
  assign \new_[10693]_  = \new_[6455]_  ^ \new_[2833]_ ;
  assign \new_[10694]_  = \new_[6544]_  ^ \new_[2840]_ ;
  assign \new_[10695]_  = \new_[6437]_  ^ \new_[2833]_ ;
  assign \new_[10696]_  = \new_[6415]_  ^ \new_[2720]_ ;
  assign \new_[10697]_  = \new_[6428]_  ^ \new_[2721]_ ;
  assign \new_[10698]_  = ~\new_[10827]_ ;
  assign \new_[10699]_  = \wb_data_i[7]  ^ \wb_data_i[0] ;
  assign \new_[10700]_  = \new_[6410]_  ^ \new_[2839]_ ;
  assign \new_[10701]_  = \new_[6423]_  ^ \new_[2841]_ ;
  assign \mc_data_pad_o[2]  = \\u7_mc_data_o_reg[2] ;
  assign \new_[10703]_  = \new_[6411]_  ^ \new_[2840]_ ;
  assign \new_[10704]_  = ~\new_[10950]_ ;
  assign \new_[10705]_  = ~\new_[8063]_  | ~\new_[11238]_ ;
  assign \mc_data_pad_o[9]  = \\u7_mc_data_o_reg[9] ;
  assign \mc_data_pad_o[14]  = \\u7_mc_data_o_reg[14] ;
  assign \new_[10708]_  = ~\new_[11098]_  & ~\new_[10975]_ ;
  assign \new_[10709]_  = \new_[6447]_  ^ \new_[2721]_ ;
  assign \new_[10710]_  = ~\new_[3184]_ ;
  assign \new_[10711]_  = \wb_data_i[4]  ^ \wb_data_i[2] ;
  assign \new_[10712]_  = ~\new_[11312]_  | ~\new_[11315]_ ;
  assign \new_[10713]_  = ~\new_[10854]_ ;
  assign \new_[10714]_  = ~\new_[1433]_ ;
  assign \new_[10715]_  = ~\new_[10965]_ ;
  assign \mc_data_pad_o[13]  = \\u7_mc_data_o_reg[13] ;
  assign \mc_data_pad_o[23]  = \\u7_mc_data_o_reg[23] ;
  assign n5381 = ~n5766 & ~\new_[11020]_ ;
  assign \new_[10719]_  = ~\new_[8052]_  | ~\new_[11238]_ ;
  assign \new_[10720]_  = \new_[6438]_  ^ \new_[2721]_ ;
  assign \new_[10721]_  = ~\new_[11243]_  | ~\new_[11238]_ ;
  assign \new_[10722]_  = ~\new_[10928]_ ;
  assign \new_[10723]_  = \new_[6440]_  ^ \new_[2829]_ ;
  assign \new_[10724]_  = ~\new_[10902]_ ;
  assign \new_[10725]_  = \new_[6450]_  ^ \new_[2829]_ ;
  assign \mc_data_pad_o[3]  = \\u7_mc_data_o_reg[3] ;
  assign \new_[10727]_  = \new_[6362]_  ^ \new_[2839]_ ;
  assign \new_[10728]_  = ~\new_[12556]_  | ~\new_[11079]_ ;
  assign \new_[10729]_  = \new_[6390]_  ^ \new_[2833]_ ;
  assign \mc_data_pad_o[10]  = \\u7_mc_data_o_reg[10] ;
  assign \new_[10731]_  = ~\new_[11168]_  | ~\new_[11140]_ ;
  assign n5341 = ~n5766 & ~\new_[11254]_ ;
  assign \new_[10733]_  = ~\new_[11189]_  & ~\wb_addr_i[4] ;
  assign \new_[10734]_  = ~\new_[10895]_ ;
  assign \new_[10735]_  = ~\new_[10948]_ ;
  assign \new_[10736]_  = ~\new_[11202]_  | ~\new_[11131]_ ;
  assign \new_[10737]_  = ~\new_[11066]_  | ~\new_[11238]_ ;
  assign \new_[10738]_  = ~\new_[11394]_  | ~\new_[11326]_ ;
  assign \new_[10739]_  = \new_[6426]_  ^ \new_[2768]_ ;
  assign \new_[10740]_  = \new_[6570]_  ^ \new_[2833]_ ;
  assign \new_[10741]_  = ~\new_[11345]_  | ~\new_[11212]_ ;
  assign \new_[10742]_  = \new_[6418]_  ^ \new_[2843]_ ;
  assign \new_[10743]_  = ~\new_[11105]_ ;
  assign \mc_data_pad_o[25]  = \\u7_mc_data_o_reg[25] ;
  assign \new_[10745]_  = \new_[6326]_  ^ \new_[2845]_ ;
  assign \new_[10746]_  = ~\new_[11365]_  | ~\new_[11107]_ ;
  assign \new_[10747]_  = ~\new_[10838]_ ;
  assign \new_[10748]_  = ~\new_[10913]_ ;
  assign \new_[10749]_  = ~\new_[10839]_ ;
  assign \new_[10750]_  = \new_[6389]_  ^ \new_[2840]_ ;
  assign \new_[10751]_  = ~\new_[11250]_  | ~\new_[11238]_ ;
  assign \new_[10752]_  = ~\new_[10912]_ ;
  assign \new_[10753]_  = \new_[6645]_  ^ \new_[2829]_ ;
  assign \new_[10754]_  = ~\new_[10964]_ ;
  assign \mc_data_pad_o[27]  = \\u7_mc_data_o_reg[27] ;
  assign \mc_data_pad_o[15]  = \\u7_mc_data_o_reg[15] ;
  assign \new_[10757]_  = \new_[6588]_  ^ \new_[2843]_ ;
  assign \new_[10758]_  = ~\new_[12053]_  | ~\new_[11041]_ ;
  assign \new_[10759]_  = ~\new_[10826]_ ;
  assign \new_[10760]_  = \new_[6552]_  ^ \new_[2830]_ ;
  assign \new_[10761]_  = \new_[6323]_  ^ \new_[2845]_ ;
  assign \new_[10762]_  = \new_[8382]_  & \new_[11145]_ ;
  assign \new_[10763]_  = \new_[6333]_  ^ \new_[2833]_ ;
  assign \new_[10764]_  = \new_[6422]_  ^ \new_[2840]_ ;
  assign \mc_data_pad_o[4]  = \\u7_mc_data_o_reg[4] ;
  assign \mc_data_pad_o[29]  = \\u7_mc_data_o_reg[29] ;
  assign \new_[10767]_  = ~\new_[10959]_ ;
  assign \new_[10768]_  = \wb_data_i[20]  ^ \wb_data_i[18] ;
  assign \new_[10769]_  = \new_[6441]_  ^ \new_[2768]_ ;
  assign \mc_data_pad_o[12]  = \\u7_mc_data_o_reg[12] ;
  assign \new_[10771]_  = ~\new_[10899]_ ;
  assign \new_[10772]_  = ~\new_[11951]_  | ~\new_[11817]_ ;
  assign \new_[10773]_  = ~\new_[10944]_ ;
  assign \mc_dp_pad_o[0]  = \\u7_mc_dp_o_reg[0] ;
  assign \new_[10775]_  = \new_[6643]_  ^ \new_[2840]_ ;
  assign \new_[10776]_  = \wb_data_i[13]  ^ \wb_data_i[11] ;
  assign n5356 = u5_rsts1_reg;
  assign \mc_data_pad_o[0]  = \\u7_mc_data_o_reg[0] ;
  assign \new_[10779]_  = \new_[6334]_  ^ \new_[2830]_ ;
  assign \new_[10780]_  = \new_[8355]_  ^ \new_[8079]_ ;
  assign \new_[10781]_  = \new_[6318]_  ^ \new_[2843]_ ;
  assign \new_[10782]_  = ~\new_[11220]_  | ~\new_[11238]_ ;
  assign \new_[10783]_  = ~\new_[10919]_ ;
  assign \new_[10784]_  = \new_[6370]_  ^ \new_[2845]_ ;
  assign \new_[10785]_  = ~wb_we_i & ~\new_[11000]_ ;
  assign \new_[10786]_  = \new_[11012]_  & \new_[11881]_ ;
  assign \new_[10787]_  = ~\new_[12185]_  | ~\new_[10988]_ ;
  assign \new_[10788]_  = \new_[6452]_  ^ \new_[2830]_ ;
  assign \mc_data_pad_o[24]  = \\u7_mc_data_o_reg[24] ;
  assign \mc_data_pad_o[17]  = \\u7_mc_data_o_reg[17] ;
  assign n5431 = \new_[7280]_  | \new_[11182]_ ;
  assign \new_[10792]_  = \new_[6392]_  ^ \new_[2720]_ ;
  assign \new_[10793]_  = ~\new_[8382]_  & ~\new_[11145]_ ;
  assign \new_[10794]_  = \new_[6606]_  ^ \new_[2768]_ ;
  assign \new_[10795]_  = \new_[6324]_  ^ \new_[2833]_ ;
  assign \new_[10796]_  = \new_[6433]_  ^ \new_[2829]_ ;
  assign \new_[10797]_  = ~\new_[11350]_  | ~\new_[11091]_ ;
  assign \mc_dp_pad_o[1]  = \\u7_mc_dp_o_reg[1] ;
  assign \new_[10799]_  = ~\new_[10960]_ ;
  assign \new_[10800]_  = \new_[6651]_  ^ \new_[2839]_ ;
  assign \new_[10801]_  = \new_[11174]_  | \new_[11246]_ ;
  assign \new_[10802]_  = ~\new_[10897]_ ;
  assign \new_[10803]_  = \new_[6368]_  ^ \new_[2721]_ ;
  assign \new_[10804]_  = ~\new_[2606]_ ;
  assign \new_[10805]_  = ~\new_[4242]_ ;
  assign \new_[10806]_  = \new_[6436]_  ^ \new_[2845]_ ;
  assign \new_[10807]_  = ~\new_[11760]_  | ~\new_[11070]_ ;
  assign \new_[10808]_  = ~\new_[10920]_ ;
  assign \new_[10809]_  = ~\new_[10962]_ ;
  assign \new_[10810]_  = \new_[6442]_  ^ \new_[2720]_ ;
  assign \new_[10811]_  = \new_[11113]_  & \new_[11097]_ ;
  assign \mc_data_pad_o[1]  = \\u7_mc_data_o_reg[1] ;
  assign \new_[10813]_  = \new_[2479]_  | \new_[2478]_ ;
  assign \new_[10814]_  = \\u7_mc_data_ir_reg[23] ;
  assign \new_[10815]_  = ~\new_[6385]_  | ~\new_[2841]_ ;
  assign \new_[10816]_  = \new_[7284]_  & \new_[7265]_ ;
  assign \new_[10817]_  = \\u7_mc_data_ir_reg[8] ;
  assign \new_[10818]_  = ~\new_[11150]_ ;
  assign \new_[10819]_  = \\u7_mc_data_ir_reg[6] ;
  assign \new_[10820]_  = \new_[11202]_ ;
  assign \new_[10821]_  = ~\new_[10501]_  | ~\new_[8813]_ ;
  assign \new_[10822]_  = \new_[7285]_  & \new_[8399]_ ;
  assign \new_[10823]_  = ~\\u0_u0_addr_r_reg[6] ;
  assign \new_[10824]_  = ~\wb_addr_i[3]  & ~\wb_addr_i[4] ;
  assign \new_[10825]_  = \\u7_mc_data_ir_reg[13] ;
  assign \new_[10826]_  = n5766 | wb_we_i;
  assign \new_[10827]_  = ~\new_[11091]_ ;
  assign \new_[10828]_  = \\u7_mc_data_ir_reg[14] ;
  assign \new_[10829]_  = \wb_addr_i[30]  | \wb_addr_i[29] ;
  assign \new_[10830]_  = ~\\u7_mc_dqm_r2_reg[3] ;
  assign \new_[10831]_  = \\u7_mc_data_ir_reg[35] ;
  assign \new_[10832]_  = \\u7_mc_data_ir_reg[21] ;
  assign \new_[10833]_  = \\u7_mc_data_ir_reg[7] ;
  assign \new_[10834]_  = \new_[8081]_  & \new_[7977]_ ;
  assign \new_[10835]_  = \\u7_mc_data_ir_reg[28] ;
  assign \new_[10836]_  = \new_[11146]_ ;
  assign \new_[10837]_  = ~\new_[7390]_  & ~\new_[10369]_ ;
  assign \new_[10838]_  = ~\new_[11259]_ ;
  assign \new_[10839]_  = ~\new_[10989]_ ;
  assign \new_[10840]_  = \\u0_wb_addr_r_reg[5] ;
  assign \new_[10841]_  = \new_[2316]_  | \new_[2315]_ ;
  assign \new_[10842]_  = ~\wb_addr_i[5]  & ~\wb_addr_i[6] ;
  assign \new_[10843]_  = \\u7_mc_data_ir_reg[22] ;
  assign \new_[10844]_  = \\u7_mc_data_ir_reg[1] ;
  assign \new_[10845]_  = \\u7_mc_data_ir_reg[0] ;
  assign \new_[10846]_  = ~u7_mc_ack_r_reg;
  assign \new_[10847]_  = \\u7_mc_data_ir_reg[19] ;
  assign \new_[10848]_  = ~\new_[6417]_  | ~\new_[2841]_ ;
  assign \new_[10849]_  = \new_[8079]_  & \new_[8049]_ ;
  assign n5466 = u5_cs_le_r1_reg;
  assign \new_[10851]_  = ~\new_[11000]_ ;
  assign \new_[10852]_  = \\u7_mc_data_ir_reg[5] ;
  assign \new_[10853]_  = ~\new_[1463]_  & ~\new_[1464]_ ;
  assign \new_[10854]_  = ~\new_[8179]_  | ~\wb_addr_i[22] ;
  assign \new_[10855]_  = ~\new_[3388]_ ;
  assign \new_[10856]_  = \new_[1611]_  | \new_[1519]_ ;
  assign \new_[10857]_  = ~\new_[3439]_  | ~\new_[3398]_ ;
  assign \new_[10858]_  = ~\\u0_u1_addr_r_reg[4] ;
  assign \new_[10859]_  = ~\new_[1453]_  & ~\new_[1454]_ ;
  assign \new_[10860]_  = \\u7_mc_data_ir_reg[17] ;
  assign \new_[10861]_  = ~\new_[1841]_  & ~\new_[1656]_ ;
  assign \new_[10862]_  = ~\new_[6446]_  | ~\new_[2843]_ ;
  assign \new_[10863]_  = \new_[10501]_  | \new_[10369]_ ;
  assign \new_[10864]_  = \new_[8200]_  & \wb_addr_i[27] ;
  assign \new_[10865]_  = ~\\u7_mc_dqm_r2_reg[2] ;
  assign \new_[10866]_  = ~\new_[11107]_ ;
  assign \new_[10867]_  = \\u7_mc_data_ir_reg[29] ;
  assign \new_[10868]_  = \\u7_mc_data_ir_reg[18] ;
  assign \new_[10869]_  = \\u7_mc_data_ir_reg[4] ;
  assign \new_[10870]_  = ~\new_[6471]_  | ~\new_[2830]_ ;
  assign \new_[10871]_  = ~\new_[11165]_ ;
  assign \new_[10872]_  = \new_[11078]_ ;
  assign \new_[10873]_  = ~\new_[11079]_ ;
  assign \new_[10874]_  = ~\\u0_u0_addr_r_reg[5] ;
  assign \new_[10875]_  = ~\new_[7703]_  | ~\new_[8229]_ ;
  assign \new_[10876]_  = ~\\u0_u0_addr_r_reg[4] ;
  assign \new_[10877]_  = \new_[3041]_  & \new_[3042]_ ;
  assign \new_[10878]_  = \\u7_mc_data_ir_reg[11] ;
  assign \new_[10879]_  = \\u7_mc_data_ir_reg[27] ;
  assign \new_[10880]_  = \new_[1582]_  | \new_[1581]_ ;
  assign \new_[10881]_  = ~\new_[1712]_  & ~\new_[1796]_ ;
  assign n5441 = u7_mc_sts_ir_reg;
  assign \new_[10883]_  = ~\wb_addr_i[26]  | ~\new_[8199]_ ;
  assign \new_[10884]_  = ~\new_[8734]_  | ~wb_cyc_i;
  assign \new_[10885]_  = \\u7_mc_data_ir_reg[10] ;
  assign \new_[10886]_  = ~\\u0_u1_addr_r_reg[5] ;
  assign \new_[10887]_  = ~\wb_addr_i[28]  | ~\new_[8201]_ ;
  assign \new_[10888]_  = ~wb_err_o & ~wb_ack_o;
  assign \new_[10889]_  = ~\new_[7702]_  | ~\new_[8179]_ ;
  assign \new_[10890]_  = ~\new_[7732]_  & ~\new_[7616]_ ;
  assign \new_[10891]_  = ~\wb_addr_i[30]  | ~\wb_addr_i[29] ;
  assign \new_[10892]_  = ~\new_[11019]_ ;
  assign \new_[10893]_  = \new_[7851]_  | \new_[7828]_ ;
  assign \new_[10894]_  = ~\new_[7966]_  | ~\new_[8390]_ ;
  assign \new_[10895]_  = ~\new_[1796]_  & ~\new_[1657]_ ;
  assign \new_[10896]_  = \\u7_mc_data_ir_reg[15] ;
  assign \new_[10897]_  = \new_[11034]_ ;
  assign \new_[10898]_  = ~\new_[8198]_  | ~\wb_addr_i[25] ;
  assign \new_[10899]_  = ~\new_[11086]_ ;
  assign \new_[10900]_  = \\u7_mc_data_ir_reg[34] ;
  assign \new_[10901]_  = \\u7_mc_data_ir_reg[12] ;
  assign \new_[10902]_  = ~\new_[11252]_ ;
  assign \new_[10903]_  = ~\new_[6529]_  | ~\new_[2841]_ ;
  assign \new_[10904]_  = \new_[8149]_  & \wb_addr_i[21] ;
  assign \new_[10905]_  = ~\new_[11193]_ ;
  assign \new_[10906]_  = ~\new_[11184]_ ;
  assign \new_[10907]_  = \new_[2056]_  | \new_[2138]_ ;
  assign \new_[10908]_  = \\u7_mc_data_ir_reg[9] ;
  assign \new_[10909]_  = ~\new_[6434]_  | ~\new_[2841]_ ;
  assign \new_[10910]_  = \new_[4145]_  | \new_[3881]_ ;
  assign \new_[10911]_  = \\u7_mc_data_ir_reg[33] ;
  assign \new_[10912]_  = ~\new_[11070]_ ;
  assign \new_[10913]_  = ~\new_[8196]_  | ~\wb_addr_i[23] ;
  assign \new_[10914]_  = ~\new_[8355]_  & ~\new_[8378]_ ;
  assign \new_[10915]_  = \new_[8382]_  & \new_[8365]_ ;
  assign \new_[10916]_  = \\u7_mc_data_ir_reg[3] ;
  assign \new_[10917]_  = ~\new_[7601]_  | ~\new_[8196]_ ;
  assign \new_[10918]_  = \new_[7275]_  & \new_[7278]_ ;
  assign \new_[10919]_  = ~\new_[11218]_ ;
  assign \new_[10920]_  = \new_[11212]_ ;
  assign \new_[10921]_  = ~\\u7_mc_dqm_r2_reg[0] ;
  assign \new_[10922]_  = ~\new_[10988]_ ;
  assign \new_[10923]_  = \\u7_mc_data_ir_reg[25] ;
  assign \new_[10924]_  = ~\new_[6424]_  | ~\new_[2842]_ ;
  assign n5461 = u5_cke_o_r1_reg;
  assign \new_[10926]_  = ~\new_[2138]_  & ~\new_[2137]_ ;
  assign \new_[10927]_  = ~\new_[8296]_  & ~\new_[8352]_ ;
  assign \new_[10928]_  = ~\new_[11817]_ ;
  assign \new_[10929]_  = ~\new_[8382]_  & ~\new_[8365]_ ;
  assign \new_[10930]_  = \new_[7285]_  & \new_[7284]_ ;
  assign \new_[10931]_  = \new_[3145]_  & \new_[3041]_ ;
  assign \new_[10932]_  = ~\new_[1582]_  & ~\new_[1579]_ ;
  assign \new_[10933]_  = ~\new_[11124]_ ;
  assign \new_[10934]_  = ~\new_[3438]_ ;
  assign \new_[10935]_  = \\u7_mc_data_ir_reg[31] ;
  assign \new_[10936]_  = \new_[3439]_  | \new_[3398]_ ;
  assign \new_[10937]_  = ~\\u7_mc_dqm_r2_reg[1] ;
  assign \new_[10938]_  = ~\new_[11012]_ ;
  assign \new_[10939]_  = \\u7_mc_data_ir_reg[26] ;
  assign \new_[10940]_  = ~\new_[1843]_  & ~\new_[1842]_ ;
  assign \new_[10941]_  = \new_[3179]_  & \new_[3145]_ ;
  assign \new_[10942]_  = \\u7_mc_data_ir_reg[24] ;
  assign \new_[10943]_  = \\u7_mc_data_ir_reg[16] ;
  assign \new_[10944]_  = \new_[1541]_  | \new_[1465]_ ;
  assign \new_[10945]_  = ~\new_[1955]_  & ~\new_[1843]_ ;
  assign \new_[10946]_  = \new_[7279]_  & \new_[7275]_ ;
  assign \new_[10947]_  = \\u7_mc_data_ir_reg[30] ;
  assign \new_[10948]_  = wb_cyc_i & wb_stb_i;
  assign \new_[10949]_  = ~\new_[11153]_ ;
  assign \new_[10950]_  = ~\new_[11041]_ ;
  assign \new_[10951]_  = ~\new_[6523]_  | ~\new_[2841]_ ;
  assign \new_[10952]_  = ~\new_[8260]_  & ~\new_[8400]_ ;
  assign \new_[10953]_  = ~\new_[6331]_  | ~\new_[2841]_ ;
  assign \new_[10954]_  = \new_[1579]_  | \new_[1539]_ ;
  assign \new_[10955]_  = ~\new_[11151]_ ;
  assign \new_[10956]_  = ~\new_[10996]_ ;
  assign \new_[10957]_  = ~u7_mc_br_r_reg;
  assign \new_[10958]_  = \\u0_wb_addr_r_reg[6] ;
  assign \new_[10959]_  = ~\new_[11140]_ ;
  assign \new_[10960]_  = ~\new_[10990]_ ;
  assign \new_[10961]_  = \new_[3176]_  & \new_[3179]_ ;
  assign \new_[10962]_  = ~\new_[11954]_ ;
  assign \new_[10963]_  = ~\new_[11737]_ ;
  assign \new_[10964]_  = ~\new_[11168]_ ;
  assign \new_[10965]_  = ~\new_[11197]_ ;
  assign \new_[10966]_  = ~\new_[7704]_  | ~\new_[8229]_ ;
  assign n5456 = \new_[7626]_  | \new_[7390]_ ;
  assign \new_[10968]_  = \\u7_mc_data_ir_reg[2] ;
  assign \new_[10969]_  = ~\\u0_wb_addr_r_reg[4] ;
  assign \new_[10970]_  = \\u7_mc_data_ir_reg[32] ;
  assign \new_[10971]_  = ~\new_[8232]_  & ~\new_[8390]_ ;
  assign \new_[10972]_  = \\u7_mc_data_ir_reg[20] ;
  assign \new_[10973]_  = ~\new_[8229]_  | ~\wb_addr_i[24] ;
  assign \new_[10974]_  = ~\\u0_u1_addr_r_reg[6] ;
  assign \new_[10975]_  = ~\new_[7279]_ ;
  assign n5546 = ~\new_[9138]_ ;
  assign \new_[10977]_  = ~\new_[10327]_ ;
  assign \new_[10978]_  = ~\new_[7746]_ ;
  assign \new_[10979]_  = ~\wb_addr_i[2] ;
  assign \new_[10980]_  = ~\new_[7984]_ ;
  assign \new_[10981]_  = ~\new_[7972]_ ;
  assign \new_[10982]_  = ~\new_[7938]_ ;
  assign \new_[10983]_  = ~\new_[7981]_ ;
  assign n5536 = ~\new_[9148]_ ;
  assign \new_[10985]_  = ~\new_[2082]_ ;
  assign \new_[10986]_  = ~\new_[8082]_ ;
  assign n5646 = ~\new_[8718]_ ;
  assign \new_[10988]_  = ~\new_[1557]_ ;
  assign \new_[10989]_  = ~\new_[1497]_ ;
  assign \new_[10990]_  = ~\new_[1537]_ ;
  assign \new_[10991]_  = ~\new_[8066]_ ;
  assign n5521 = ~\new_[9100]_ ;
  assign \new_[10993]_  = ~\new_[2128]_ ;
  assign \new_[10994]_  = ~\new_[2366]_ ;
  assign \new_[10995]_  = ~\new_[7950]_ ;
  assign \new_[10996]_  = ~\new_[2315]_ ;
  assign n5666 = ~\new_[9147]_ ;
  assign n5556 = ~\new_[9127]_ ;
  assign \new_[10999]_  = ~\new_[7974]_ ;
  assign \new_[11000]_  = ~wb_stb_i;
  assign \new_[11001]_  = ~\new_[2120]_ ;
  assign \new_[11002]_  = ~\new_[2100]_ ;
  assign n5581 = ~\new_[9171]_ ;
  assign \new_[11004]_  = ~\new_[6378]_ ;
  assign \new_[11005]_  = ~\new_[2096]_ ;
  assign \new_[11006]_  = ~\new_[2111]_ ;
  assign \new_[11007]_  = ~\new_[7936]_ ;
  assign \new_[11008]_  = ~\new_[7929]_ ;
  assign n5531 = ~\new_[9143]_ ;
  assign \new_[11010]_  = ~\new_[7970]_ ;
  assign \new_[11011]_  = ~\new_[7941]_ ;
  assign \new_[11012]_  = ~\new_[1542]_ ;
  assign \new_[11013]_  = ~\new_[8076]_ ;
  assign \new_[11014]_  = ~\new_[2095]_ ;
  assign \new_[11015]_  = ~\new_[8810]_ ;
  assign \new_[11016]_  = ~wb_ack_o;
  assign n5506 = ~\new_[9036]_ ;
  assign \new_[11018]_  = ~\new_[7968]_ ;
  assign \new_[11019]_  = ~\new_[1559]_ ;
  assign \new_[11020]_  = ~\new_[10324]_ ;
  assign n5516 = ~\new_[9135]_ ;
  assign \new_[11022]_  = ~\new_[8065]_ ;
  assign \new_[11023]_  = ~\new_[7942]_ ;
  assign \new_[11024]_  = ~\new_[2122]_ ;
  assign \new_[11025]_  = ~\new_[6416]_ ;
  assign \new_[11026]_  = ~\new_[3113]_ ;
  assign \new_[11027]_  = ~\new_[2139]_ ;
  assign \new_[11028]_  = ~\new_[8055]_ ;
  assign \new_[11029]_  = ~\new_[8229]_ ;
  assign \new_[11030]_  = ~\new_[7620]_ ;
  assign \new_[11031]_  = ~\new_[8201]_ ;
  assign \new_[11032]_  = ~\new_[7937]_ ;
  assign \new_[11033]_  = ~\new_[3882]_ ;
  assign \new_[11034]_  = ~\new_[1524]_ ;
  assign \new_[11035]_  = ~\new_[2102]_ ;
  assign \new_[11036]_  = ~\new_[7748]_ ;
  assign \new_[11037]_  = ~\new_[2117]_ ;
  assign \new_[11038]_  = ~\new_[2132]_ ;
  assign \new_[11039]_  = ~\new_[1542]_ ;
  assign \new_[11040]_  = ~\new_[10368]_ ;
  assign \new_[11041]_  = ~\new_[1543]_ ;
  assign \new_[11042]_  = ~\new_[8364]_ ;
  assign \new_[11043]_  = ~\new_[8058]_ ;
  assign \new_[11044]_  = ~\new_[2089]_ ;
  assign \new_[11045]_  = ~\new_[8197]_ ;
  assign \new_[11046]_  = ~\new_[7985]_ ;
  assign \new_[11047]_  = ~\new_[2125]_ ;
  assign \new_[11048]_  = ~\new_[7917]_ ;
  assign \new_[11050]_  = ~\new_[3180]_ ;
  assign \new_[11051]_  = ~\new_[3112]_ ;
  assign \new_[11052]_  = ~\new_[10330]_ ;
  assign \new_[11053]_  = ~\new_[4126]_ ;
  assign \new_[11054]_  = ~\new_[7971]_ ;
  assign \new_[11055]_  = ~\new_[2354]_ ;
  assign \new_[11056]_  = ~\new_[7943]_ ;
  assign \new_[11057]_  = ~\new_[10351]_ ;
  assign \new_[11058]_  = ~\new_[2927]_ ;
  assign \new_[11059]_  = ~\new_[3308]_ ;
  assign \new_[11060]_  = ~\new_[2367]_ ;
  assign \new_[11061]_  = ~\new_[7932]_ ;
  assign \new_[11062]_  = ~\new_[8862]_ ;
  assign \new_[11063]_  = ~\new_[6548]_ ;
  assign \new_[11064]_  = ~\new_[2115]_ ;
  assign \new_[11065]_  = ~\new_[7812]_ ;
  assign \new_[11066]_  = ~\new_[8034]_ ;
  assign \new_[11067]_  = ~\new_[2359]_ ;
  assign \new_[11068]_  = ~\new_[2721]_ ;
  assign n5416 = ~\new_[3182]_ ;
  assign \new_[11070]_  = ~\new_[1490]_ ;
  assign \new_[11071]_  = ~\new_[1644]_ ;
  assign \new_[11072]_  = ~\new_[8196]_ ;
  assign \new_[11073]_  = ~\new_[2479]_ ;
  assign \new_[11074]_  = ~\new_[8045]_ ;
  assign n5491 = ~\new_[9061]_ ;
  assign \new_[11076]_  = ~\new_[2091]_ ;
  assign \new_[11077]_  = ~\new_[7982]_ ;
  assign \new_[11078]_  = ~\new_[1498]_ ;
  assign \new_[11079]_  = ~\new_[1562]_ ;
  assign \new_[11080]_  = ~\new_[2719]_ ;
  assign \new_[11081]_  = ~\new_[4341]_ ;
  assign \new_[11082]_  = ~\new_[8073]_ ;
  assign \new_[11083]_  = ~\new_[2074]_ ;
  assign \new_[11084]_  = ~\new_[2105]_ ;
  assign n5591 = ~\new_[9150]_ ;
  assign \new_[11086]_  = ~\new_[1469]_ ;
  assign n5631 = ~\new_[9167]_ ;
  assign \new_[11088]_  = ~\new_[7740]_ ;
  assign \new_[11089]_  = ~\new_[7709]_ ;
  assign \new_[11090]_  = ~\new_[2092]_ ;
  assign \new_[11091]_  = ~\new_[1483]_ ;
  assign \new_[11092]_  = ~\new_[7739]_ ;
  assign \new_[11093]_  = ~\new_[8060]_ ;
  assign n5306 = ~\new_[10072]_ ;
  assign n5571 = ~\new_[9027]_ ;
  assign \new_[11096]_  = ~\new_[7919]_ ;
  assign \new_[11097]_  = ~\new_[4242]_ ;
  assign \new_[11098]_  = ~\new_[7265]_ ;
  assign \new_[11099]_  = ~\new_[2365]_ ;
  assign \new_[11100]_  = ~\new_[3185]_ ;
  assign \new_[11101]_  = ~\new_[2078]_ ;
  assign \new_[11102]_  = ~\new_[3077]_ ;
  assign \new_[11103]_  = ~\new_[2124]_ ;
  assign \new_[11104]_  = ~\new_[2130]_ ;
  assign \new_[11105]_  = ~\new_[1460]_ ;
  assign \new_[11106]_  = ~\new_[2119]_ ;
  assign \new_[11107]_  = ~\new_[1560]_ ;
  assign \new_[11108]_  = ~\new_[8198]_ ;
  assign \new_[11109]_  = ~\new_[2388]_ ;
  assign n5596 = ~\new_[9076]_ ;
  assign \new_[11111]_  = ~\new_[2358]_ ;
  assign n5566 = ~\new_[8979]_ ;
  assign \new_[11113]_  = ~\new_[4691]_ ;
  assign \new_[11114]_  = ~\new_[2837]_ ;
  assign n5496 = ~\new_[9130]_ ;
  assign n5561 = ~\new_[9128]_ ;
  assign \new_[11117]_  = ~\new_[7973]_ ;
  assign \new_[11118]_  = ~\new_[7944]_ ;
  assign \new_[11119]_  = ~\new_[3184]_ ;
  assign \new_[11120]_  = ~\new_[2118]_ ;
  assign \new_[11121]_  = ~\new_[4146]_ ;
  assign \new_[11122]_  = ~\new_[2093]_ ;
  assign \new_[11123]_  = ~\new_[6366]_ ;
  assign \new_[11124]_  = ~\new_[1535]_ ;
  assign n5486 = ~\new_[9152]_ ;
  assign \new_[11126]_  = ~\new_[8350]_ ;
  assign \new_[11127]_  = ~\new_[7969]_ ;
  assign \new_[11128]_  = ~\new_[2106]_ ;
  assign \new_[11129]_  = ~\new_[1462]_ ;
  assign \new_[11130]_  = ~\new_[7734]_ ;
  assign \new_[11131]_  = ~\new_[3167]_ ;
  assign \new_[11132]_  = ~\new_[2104]_ ;
  assign \new_[11133]_  = ~\new_[2769]_ ;
  assign \new_[11134]_  = ~\new_[7922]_ ;
  assign \new_[11135]_  = ~\new_[10360]_ ;
  assign \new_[11136]_  = ~\new_[2097]_ ;
  assign \new_[11137]_  = ~\new_[2099]_ ;
  assign n5481 = ~\new_[8717]_ ;
  assign \new_[11139]_  = ~\new_[6421]_ ;
  assign \new_[11140]_  = ~\new_[1536]_ ;
  assign \new_[11141]_  = ~\new_[9136]_ ;
  assign \new_[11142]_  = ~\new_[2133]_ ;
  assign \new_[11143]_  = ~\new_[2112]_ ;
  assign n5601 = ~\new_[9155]_ ;
  assign \new_[11145]_  = ~\new_[8365]_ ;
  assign \new_[11146]_  = ~\new_[3153]_ ;
  assign \new_[11147]_  = ~\new_[6448]_ ;
  assign \new_[11148]_  = ~\new_[3440]_ ;
  assign \new_[11149]_  = ~\new_[7945]_ ;
  assign \new_[11150]_  = ~\new_[1455]_ ;
  assign \new_[11151]_  = ~\new_[1529]_ ;
  assign \new_[11152]_  = ~\new_[7983]_ ;
  assign \new_[11153]_  = ~\new_[9569]_ ;
  assign \new_[11154]_  = ~\new_[2134]_ ;
  assign \new_[11155]_  = ~\new_[2135]_ ;
  assign \new_[11156]_  = ~\new_[7736]_ ;
  assign \new_[11157]_  = ~\new_[7927]_ ;
  assign \new_[11158]_  = ~\new_[10311]_ ;
  assign \new_[11159]_  = ~\new_[2494]_ ;
  assign \new_[11160]_  = ~\new_[2113]_ ;
  assign \new_[11161]_  = ~\new_[10347]_ ;
  assign \new_[11162]_  = ~\new_[4236]_ ;
  assign \new_[11163]_  = ~\new_[7926]_ ;
  assign \new_[11164]_  = ~\new_[6120]_ ;
  assign \new_[11165]_  = ~\new_[1494]_ ;
  assign \new_[11166]_  = ~\new_[7933]_ ;
  assign \new_[11167]_  = ~\new_[1646]_ ;
  assign \new_[11168]_  = ~\new_[1504]_ ;
  assign \new_[11169]_  = ~\new_[2123]_ ;
  assign \new_[11170]_  = ~\new_[2136]_ ;
  assign \new_[11171]_  = ~\new_[2073]_ ;
  assign \new_[11172]_  = ~\new_[7975]_ ;
  assign \new_[11173]_  = ~\new_[7935]_ ;
  assign \new_[11174]_  = ~\new_[7697]_ ;
  assign \new_[11175]_  = ~\new_[7710]_ ;
  assign \new_[11176]_  = ~\new_[2356]_ ;
  assign \new_[11177]_  = ~\new_[7939]_ ;
  assign \new_[11178]_  = ~\new_[2372]_ ;
  assign \new_[11179]_  = ~\new_[2767]_ ;
  assign \new_[11180]_  = ~\new_[6332]_ ;
  assign \new_[11181]_  = ~\new_[7737]_ ;
  assign \new_[11182]_  = ~\new_[7617]_ ;
  assign \new_[11183]_  = ~\new_[6431]_ ;
  assign \new_[11184]_  = ~\new_[1481]_ ;
  assign \new_[11185]_  = ~\new_[10277]_ ;
  assign \new_[11186]_  = ~\new_[7839]_ ;
  assign n5661 = ~\new_[8984]_ ;
  assign \new_[11188]_  = ~\new_[8032]_ ;
  assign \new_[11189]_  = ~\wb_addr_i[3] ;
  assign \new_[11190]_  = ~\new_[7751]_ ;
  assign n5671 = ~\new_[8721]_ ;
  assign \new_[11192]_  = ~\new_[7618]_ ;
  assign \new_[11193]_  = ~\new_[1501]_ ;
  assign \new_[11194]_  = ~\new_[2098]_ ;
  assign \new_[11195]_  = ~\new_[1507]_ ;
  assign n5551 = ~\new_[9050]_ ;
  assign \new_[11197]_  = ~\new_[1506]_ ;
  assign \new_[11198]_  = ~\new_[7979]_ ;
  assign \new_[11199]_  = ~\new_[2355]_ ;
  assign \new_[11200]_  = ~\new_[7914]_ ;
  assign \new_[11201]_  = ~\new_[2361]_ ;
  assign \new_[11202]_  = ~\new_[3186]_ ;
  assign \new_[11203]_  = ~\new_[8389]_ ;
  assign n5586 = ~\new_[8986]_ ;
  assign \new_[11205]_  = ~\new_[3181]_ ;
  assign \new_[11206]_  = ~\new_[2114]_ ;
  assign \new_[11207]_  = ~\new_[2357]_ ;
  assign n5621 = ~\new_[9129]_ ;
  assign \new_[11209]_  = ~\new_[1482]_ ;
  assign n5606 = ~\new_[9029]_ ;
  assign n5641 = ~\new_[9166]_ ;
  assign \new_[11212]_  = ~\new_[1467]_ ;
  assign \new_[11213]_  = ~\new_[8380]_ ;
  assign \new_[11214]_  = ~\new_[8179]_ ;
  assign \new_[11215]_  = ~\new_[2126]_ ;
  assign \new_[11216]_  = ~\new_[2101]_ ;
  assign \new_[11217]_  = ~\new_[7934]_ ;
  assign \new_[11218]_  = ~\new_[1505]_ ;
  assign \new_[11219]_  = ~\new_[1580]_ ;
  assign \new_[11220]_  = ~\new_[8056]_ ;
  assign \new_[11221]_  = ~\new_[8168]_ ;
  assign n5476 = ~\new_[8704]_ ;
  assign \new_[11223]_  = ~\new_[8059]_ ;
  assign \new_[11224]_  = ~\new_[2360]_ ;
  assign \new_[11225]_  = ~\new_[2129]_ ;
  assign \new_[11226]_  = ~\new_[8053]_ ;
  assign \new_[11227]_  = ~\new_[3050]_ ;
  assign n5656 = ~\new_[9004]_ ;
  assign n5611 = ~\new_[9119]_ ;
  assign n5616 = ~\new_[8985]_ ;
  assign \new_[11231]_  = ~\new_[10333]_ ;
  assign \new_[11232]_  = ~\new_[2090]_ ;
  assign \new_[11233]_  = ~\new_[8197]_ ;
  assign \new_[11234]_  = ~\new_[8080]_ ;
  assign \new_[11235]_  = ~\new_[3178]_ ;
  assign n5626 = ~\new_[9116]_ ;
  assign n5636 = ~\new_[9106]_ ;
  assign \new_[11238]_  = \new_[9569]_ ;
  assign n5676 = ~\new_[9052]_ ;
  assign \new_[11240]_  = ~\new_[8064]_ ;
  assign \new_[11241]_  = ~\new_[8074]_ ;
  assign n5471 = ~\new_[9154]_ ;
  assign \new_[11243]_  = ~\new_[8047]_ ;
  assign \new_[11244]_  = ~\new_[2107]_ ;
  assign \new_[11245]_  = ~\new_[8057]_ ;
  assign \new_[11246]_  = ~\new_[8199]_ ;
  assign \new_[11247]_  = ~\new_[7718]_ ;
  assign \new_[11248]_  = ~\new_[2362]_ ;
  assign \new_[11249]_  = ~\new_[8054]_ ;
  assign \new_[11250]_  = ~\new_[8083]_ ;
  assign \new_[11251]_  = ~\new_[2109]_ ;
  assign \new_[11252]_  = ~\new_[1500]_ ;
  assign \new_[11253]_  = ~\new_[8396]_ ;
  assign \new_[11254]_  = ~\new_[10279]_ ;
  assign \new_[11255]_  = ~\new_[10289]_ ;
  assign \new_[11256]_  = ~\new_[8399]_ ;
  assign \new_[11257]_  = ~\new_[7813]_ ;
  assign \new_[11258]_  = ~\new_[6543]_ ;
  assign \new_[11259]_  = ~\new_[1452]_ ;
  assign \new_[11260]_  = ~\new_[2121]_ ;
  assign \new_[11261]_  = ~\new_[2110]_ ;
  assign \new_[11262]_  = ~\new_[2127]_ ;
  assign \new_[11263]_  = \new_[7688]_ ;
  assign \new_[11264]_  = \new_[7701]_ ;
  assign n661 = ~\new_[11266]_ ;
  assign \new_[11266]_  = \new_[12224]_ ;
  assign \new_[11267]_  = \new_[12420]_ ;
  assign \new_[11268]_  = \new_[12420]_ ;
  assign \new_[11269]_  = ~\new_[11270]_ ;
  assign \new_[11270]_  = ~\new_[4995]_ ;
  assign \new_[11271]_  = ~\new_[11270]_ ;
  assign \new_[11272]_  = ~\new_[11273]_ ;
  assign \new_[11273]_  = ~\new_[11277]_ ;
  assign \new_[11274]_  = \new_[11277]_ ;
  assign \new_[11275]_  = ~\new_[12531]_ ;
  assign \new_[11276]_  = ~\new_[12531]_ ;
  assign \new_[11277]_  = ~\new_[12531]_ ;
  assign \new_[11278]_  = ~\new_[12532]_ ;
  assign \new_[11279]_  = ~\new_[11386]_ ;
  assign \new_[11280]_  = ~\new_[11283]_ ;
  assign \new_[11281]_  = ~\new_[11283]_ ;
  assign \new_[11282]_  = ~\new_[11283]_ ;
  assign \new_[11283]_  = \new_[11287]_ ;
  assign \new_[11284]_  = ~\new_[11285]_ ;
  assign \new_[11285]_  = \new_[11287]_ ;
  assign \new_[11286]_  = ~\new_[11287]_ ;
  assign \new_[11287]_  = ~\new_[11291]_ ;
  assign \new_[11288]_  = ~\new_[11290]_ ;
  assign \new_[11289]_  = ~\new_[11290]_ ;
  assign \new_[11290]_  = ~\new_[11291]_ ;
  assign \new_[11291]_  = ~\new_[11384]_ ;
  assign \new_[11292]_  = ~\new_[12280]_ ;
  assign \new_[11293]_  = ~\new_[11296]_ ;
  assign \new_[11294]_  = ~\new_[11296]_ ;
  assign \new_[11295]_  = ~\new_[11296]_ ;
  assign \new_[11296]_  = ~\new_[11578]_ ;
  assign \new_[11297]_  = ~\new_[11503]_ ;
  assign \new_[11298]_  = ~\new_[11299]_ ;
  assign \new_[11299]_  = \new_[11300]_ ;
  assign \new_[11300]_  = ~\new_[1521]_ ;
  assign \new_[11301]_  = \new_[11302]_ ;
  assign \new_[11302]_  = \new_[11306]_ ;
  assign \new_[11303]_  = \new_[11306]_ ;
  assign \new_[11304]_  = \new_[11306]_ ;
  assign \new_[11305]_  = \new_[11306]_ ;
  assign \new_[11306]_  = \new_[11307]_ ;
  assign \new_[11307]_  = ~\new_[7179]_ ;
  assign \new_[11308]_  = ~\new_[11309]_ ;
  assign \new_[11309]_  = ~\new_[11876]_ ;
  assign \new_[11310]_  = ~\new_[11311]_ ;
  assign \new_[11311]_  = \new_[11312]_ ;
  assign \new_[11312]_  = ~\new_[1532]_ ;
  assign \new_[11313]_  = ~\new_[11314]_ ;
  assign \new_[11314]_  = \new_[11315]_ ;
  assign \new_[11315]_  = ~\new_[1533]_ ;
  assign \new_[11316]_  = ~\new_[11317]_ ;
  assign \new_[11317]_  = \new_[11318]_ ;
  assign \new_[11318]_  = ~\new_[1496]_ ;
  assign \new_[11319]_  = ~\new_[12216]_ ;
  assign \new_[11320]_  = ~\new_[11321]_ ;
  assign \new_[11321]_  = \new_[11322]_ ;
  assign \new_[11322]_  = ~\new_[1495]_ ;
  assign \new_[11323]_  = ~\new_[11324]_ ;
  assign \new_[11324]_  = \new_[11325]_ ;
  assign \new_[11325]_  = \new_[11326]_ ;
  assign \new_[11326]_  = ~\new_[1456]_ ;
  assign \new_[11327]_  = ~\new_[11762]_ ;
  assign \new_[11328]_  = ~\new_[11329]_ ;
  assign \new_[11329]_  = \new_[11330]_ ;
  assign \new_[11330]_  = ~\new_[1503]_ ;
  assign \new_[11331]_  = ~\new_[11334]_ ;
  assign \new_[11332]_  = ~\new_[11334]_ ;
  assign \new_[11333]_  = ~\new_[11334]_ ;
  assign \new_[11334]_  = \new_[11761]_ ;
  assign \new_[11335]_  = \new_[11336]_ ;
  assign \new_[11336]_  = ~\new_[10690]_ ;
  assign \new_[11337]_  = ~\new_[11338]_ ;
  assign \new_[11338]_  = \new_[11339]_ ;
  assign \new_[11339]_  = ~\new_[1468]_ ;
  assign \new_[11340]_  = ~\new_[11341]_ ;
  assign \new_[11341]_  = \new_[11342]_ ;
  assign \new_[11342]_  = ~\new_[1493]_ ;
  assign \new_[11343]_  = ~\new_[11344]_ ;
  assign \new_[11344]_  = \new_[11345]_ ;
  assign \new_[11345]_  = ~\new_[1491]_ ;
  assign \new_[11346]_  = \new_[11347]_ ;
  assign \new_[11347]_  = ~\new_[10741]_ ;
  assign \new_[11348]_  = ~\new_[11349]_ ;
  assign \new_[11349]_  = \new_[11350]_ ;
  assign \new_[11350]_  = ~\new_[1466]_ ;
  assign \new_[11351]_  = \new_[11352]_ ;
  assign \new_[11352]_  = ~\new_[10248]_ ;
  assign \new_[11353]_  = ~\new_[11393]_ ;
  assign \new_[11354]_  = \new_[11950]_ ;
  assign \new_[11355]_  = ~\new_[12184]_ ;
  assign \new_[11356]_  = ~\new_[12400]_ ;
  assign \new_[11357]_  = \new_[11358]_ ;
  assign \new_[11358]_  = ~\new_[10787]_ ;
  assign \new_[11359]_  = \new_[11360]_ ;
  assign \new_[11360]_  = ~\new_[10712]_ ;
  assign \new_[11361]_  = ~\new_[12401]_ ;
  assign \new_[11362]_  = ~\new_[10797]_ ;
  assign \new_[11363]_  = ~\new_[11364]_ ;
  assign \new_[11364]_  = \new_[11365]_ ;
  assign \new_[11365]_  = ~\new_[1499]_ ;
  assign \new_[11366]_  = ~\new_[11368]_ ;
  assign \new_[11367]_  = ~\new_[11368]_ ;
  assign \new_[11368]_  = \new_[11369]_ ;
  assign \new_[11369]_  = ~\new_[1530]_ ;
  assign \new_[11370]_  = \new_[12467]_  | \new_[11406]_ ;
  assign \new_[11371]_  = ~\new_[11418]_ ;
  assign \new_[11372]_  = ~\new_[11406]_  & ~\new_[12468]_ ;
  assign \new_[11373]_  = ~\new_[11409]_  & ~\new_[12468]_ ;
  assign \new_[11374]_  = ~\new_[11375]_  & ~\new_[12050]_ ;
  assign \new_[11375]_  = ~\new_[11378]_  | ~\new_[12053]_  | ~\new_[11376]_  | ~\new_[11041]_ ;
  assign \new_[11376]_  = \new_[11377]_  & \new_[12454]_ ;
  assign \new_[11377]_  = ~\new_[12554]_  & ~\new_[10866]_ ;
  assign \new_[11378]_  = ~\new_[1526]_ ;
  assign \new_[11379]_  = ~\new_[11382]_  & (~\new_[11380]_  | ~\new_[11381]_ );
  assign \new_[11380]_  = ~\new_[11054]_  & ~\new_[11286]_ ;
  assign \new_[11381]_  = ~\new_[9569]_  & ~\new_[11141]_ ;
  assign \new_[11382]_  = ~\new_[11383]_  & ~\new_[11291]_ ;
  assign \new_[11383]_  = ~\new_[10949]_  | ~\new_[11013]_ ;
  assign \new_[11384]_  = ~\new_[2632]_  | ~\new_[10495]_ ;
  assign \new_[11385]_  = ~\new_[11386]_ ;
  assign \new_[11386]_  = ~\new_[11291]_ ;
  assign \new_[11387]_  = \new_[11761]_  & \new_[11817]_ ;
  assign \new_[11388]_  = ~\new_[11389]_ ;
  assign \new_[11389]_  = ~\new_[12564]_  | ~\new_[12585]_  | ~\new_[10470]_ ;
  assign \new_[11390]_  = \new_[11391]_  | \new_[11395]_ ;
  assign \new_[11391]_  = ~\new_[11393]_  | ~\new_[11329]_  | ~\new_[11392]_  | ~\new_[10450]_ ;
  assign \new_[11392]_  = \new_[11325]_  & \new_[12757]_ ;
  assign \new_[11393]_  = \new_[11394]_ ;
  assign \new_[11394]_  = ~\new_[1531]_ ;
  assign \new_[11395]_  = ~\new_[11396]_  | ~\new_[11338]_ ;
  assign \new_[11396]_  = \new_[11368]_  & \new_[12733]_ ;
  assign \new_[11397]_  = ~\new_[11398]_  | ~\new_[11399]_ ;
  assign \new_[11398]_  = ~\new_[8171]_ ;
  assign \new_[11399]_  = ~\new_[8170]_ ;
  assign \new_[11400]_  = ~\new_[11401]_  | ~\new_[11402]_ ;
  assign \new_[11401]_  = \new_[10451]_  ? \new_[10811]_  : \new_[8351]_ ;
  assign \new_[11402]_  = ~\new_[10129]_  & (~\new_[8354]_  | ~\new_[10811]_ );
  assign \new_[11403]_  = \new_[11402]_ ;
  assign \new_[11404]_  = \new_[11401]_ ;
  assign \new_[11405]_  = ~\new_[12467]_  & ~\new_[11406]_ ;
  assign \new_[11406]_  = ~\new_[8474]_  | ~\new_[8471]_ ;
  assign \new_[11407]_  = \new_[8473]_  & \new_[8470]_ ;
  assign \new_[11408]_  = ~\new_[11406]_  & ~\new_[12467]_ ;
  assign \new_[11409]_  = ~\new_[11407]_ ;
  assign \new_[11410]_  = ~\new_[11411]_ ;
  assign \new_[11411]_  = \new_[11412]_  & \new_[12506]_ ;
  assign \new_[11412]_  = ~\new_[4237]_ ;
  assign \new_[11413]_  = ~\new_[12182]_  | ~\new_[9736]_  | ~\new_[11164]_ ;
  assign \new_[11414]_  = ~\new_[9121]_  | ~\new_[7672]_  | ~\new_[10355]_ ;
  assign \new_[11415]_  = ~\new_[11481]_ ;
  assign \new_[11416]_  = ~\new_[12591]_  & ~\new_[11417]_ ;
  assign \new_[11417]_  = \new_[11215]_  ? \new_[12622]_  : \new_[11084]_ ;
  assign \new_[11418]_  = ~\new_[12499]_  & (~\new_[11407]_  | ~\new_[11408]_ );
  assign \new_[11419]_  = ~\new_[7875]_  | ~\new_[10899]_  | ~\new_[11105]_ ;
  assign \new_[11420]_  = ~\new_[10438]_  | ~\new_[12446]_  | ~\new_[12437]_  | ~\new_[8714]_ ;
  assign n1156 = ~\new_[11429]_  | ~\new_[11422]_  | ~\new_[11425]_ ;
  assign \new_[11422]_  = ~\new_[11423]_  | ~\new_[11424]_ ;
  assign \new_[11423]_  = ~\new_[2253]_  | ~\new_[8361]_ ;
  assign \new_[11424]_  = ~\new_[12397]_ ;
  assign \new_[11425]_  = \new_[11426]_  & \new_[11427]_ ;
  assign \new_[11426]_  = ~\new_[12396]_  | (~\new_[12755]_  & ~\new_[9902]_ );
  assign \new_[11427]_  = ~\new_[12397]_  | ~\new_[11428]_  | ~\new_[8713]_ ;
  assign \new_[11428]_  = ~\new_[10553]_  | ~\new_[3800]_  | ~\new_[9772]_ ;
  assign \new_[11429]_  = \new_[11430]_  | \new_[11431]_ ;
  assign \new_[11430]_  = ~\new_[11428]_ ;
  assign \new_[11431]_  = ~\new_[12396]_ ;
  assign \new_[11432]_  = ~\new_[11895]_ ;
  assign \new_[11433]_  = \new_[12274]_  & \new_[10838]_ ;
  assign \new_[11434]_  = ~\new_[7543]_  & ~\new_[11813]_ ;
  assign \new_[11435]_  = ~\new_[12286]_ ;
  assign \new_[11436]_  = \new_[10811]_ ;
  assign \new_[11437]_  = ~\new_[4150]_  | ~\new_[11438]_ ;
  assign \new_[11438]_  = ~\new_[11987]_  & ~\new_[11439]_ ;
  assign \new_[11439]_  = ~\new_[7180]_  | ~\new_[7174]_ ;
  assign \new_[11440]_  = \new_[11441]_  | \new_[6464]_ ;
  assign \new_[11441]_  = ~\new_[12486]_  | ~\new_[11442]_ ;
  assign \new_[11442]_  = ~\new_[2606]_  & ~\new_[7019]_ ;
  assign \new_[11443]_  = ~\new_[6073]_  | ~\new_[4815]_  | ~\new_[6367]_  | ~\new_[5246]_ ;
  assign n1121 = \new_[12615]_  | \new_[11446]_  | \new_[11445]_  | \new_[11437]_ ;
  assign \new_[11445]_  = ~\new_[12486]_  | ~\new_[5246]_  | ~\new_[4815]_ ;
  assign \new_[11446]_  = ~\new_[6073]_  | ~\new_[11447]_  | ~\new_[6367]_ ;
  assign \new_[11447]_  = ~\new_[7019]_  & ~\new_[6464]_ ;
  assign \new_[11448]_  = ~\new_[11786]_  | ~\new_[11452]_ ;
  assign \new_[11449]_  = \new_[11419]_  & \new_[11420]_ ;
  assign \new_[11450]_  = ~\new_[11451]_  | ~\new_[7531]_  | ~\new_[10320]_ ;
  assign \new_[11451]_  = \new_[11321]_  & \new_[10871]_ ;
  assign \new_[11452]_  = ~\new_[10575]_  & ~\new_[10511]_ ;
  assign \new_[11453]_  = \new_[11454]_  & \new_[11456]_ ;
  assign \new_[11454]_  = ~\new_[11472]_ ;
  assign \new_[11455]_  = ~\new_[12213]_  & ~\new_[11714]_ ;
  assign \new_[11456]_  = ~\new_[11510]_  | ~\new_[11062]_ ;
  assign \new_[11457]_  = ~\new_[11458]_  | ~\new_[7428]_ ;
  assign \new_[11458]_  = ~\new_[4754]_  | ~\new_[9643]_ ;
  assign \new_[11459]_  = \new_[11460]_  & \new_[11461]_ ;
  assign \new_[11460]_  = ~\new_[12523]_  | ~\new_[11720]_  | ~\new_[8030]_ ;
  assign \new_[11461]_  = \new_[11462]_  & \new_[11463]_ ;
  assign \new_[11462]_  = ~\new_[11435]_  | ~\new_[7911]_  | ~\new_[7298]_  | ~\new_[11415]_ ;
  assign \new_[11463]_  = ~\new_[11878]_  & ~\new_[11464]_ ;
  assign \new_[11464]_  = ~\new_[11465]_  | ~\new_[7871]_ ;
  assign \new_[11465]_  = \new_[11466]_  | \new_[11554]_ ;
  assign \new_[11466]_  = ~\new_[3438]_  | ~\new_[1643]_ ;
  assign \new_[11467]_  = \new_[11468]_ ;
  assign \new_[11468]_  = ~\new_[11469]_ ;
  assign \new_[11469]_  = ~\new_[11470]_  | ~\new_[11473]_ ;
  assign \new_[11470]_  = ~\new_[11471]_  | ~\new_[11807]_ ;
  assign \new_[11471]_  = \new_[11472]_ ;
  assign \new_[11472]_  = ~\new_[11433]_  | ~\new_[11455]_  | ~\new_[11914]_ ;
  assign \new_[11473]_  = \new_[7782]_  | \new_[11471]_ ;
  assign \new_[11474]_  = \new_[11468]_ ;
  assign \new_[11475]_  = ~\new_[12090]_  | ~\new_[12392]_ ;
  assign \new_[11476]_  = ~\new_[7151]_ ;
  assign \new_[11477]_  = ~\new_[11478]_ ;
  assign \new_[11478]_  = ~\new_[11479]_ ;
  assign \new_[11479]_  = \new_[5977]_  & \new_[11480]_ ;
  assign \new_[11480]_  = ~\new_[11481]_  & ~\new_[11482]_ ;
  assign \new_[11481]_  = ~\new_[12283]_  | ~\new_[11510]_ ;
  assign \new_[11482]_  = ~\new_[11483]_  | ~\new_[7525]_  | ~\new_[10471]_ ;
  assign \new_[11483]_  = \new_[10960]_  & \new_[11124]_ ;
  assign \new_[11484]_  = ~\new_[11492]_  | ~\new_[11485]_  | ~\new_[11491]_ ;
  assign \new_[11485]_  = \new_[11486]_ ;
  assign \new_[11486]_  = \new_[11487]_  & \new_[11489]_ ;
  assign \new_[11487]_  = ~\new_[11488]_  & ~\new_[11475]_ ;
  assign \new_[11488]_  = ~\new_[11763]_  | ~\new_[10383]_ ;
  assign \new_[11489]_  = ~\new_[12172]_  & ~\new_[11490]_ ;
  assign \new_[11490]_  = ~\new_[9361]_  & ~\new_[10203]_ ;
  assign \new_[11491]_  = \new_[12523]_ ;
  assign \new_[11492]_  = ~\new_[11493]_ ;
  assign \new_[11493]_  = \new_[11494]_ ;
  assign \new_[11494]_  = ~\new_[1558]_ ;
  assign \new_[11495]_  = \new_[11496]_  & \new_[11779]_ ;
  assign \new_[11496]_  = ~\new_[12634]_  & ~\new_[11497]_  & ~\new_[8708]_ ;
  assign \new_[11497]_  = ~\new_[5977]_ ;
  assign \new_[11498]_  = ~\new_[8708]_  & ~\new_[12634]_ ;
  assign \new_[11499]_  = ~\new_[11500]_  | ~\new_[11504]_ ;
  assign \new_[11500]_  = \new_[11501]_ ;
  assign \new_[11501]_  = ~\new_[11502]_  | ~\new_[11503]_ ;
  assign \new_[11502]_  = ~\new_[9814]_  | ~\new_[9311]_  | ~\new_[7788]_  | ~\new_[8714]_ ;
  assign \new_[11503]_  = \new_[11983]_ ;
  assign \new_[11504]_  = ~\new_[11062]_  & ~\new_[11299]_ ;
  assign \new_[11505]_  = ~\new_[2055]_  & ~\new_[11506]_ ;
  assign \new_[11506]_  = ~\new_[11507]_  & ~\new_[11510]_ ;
  assign \new_[11507]_  = ~\new_[11508]_ ;
  assign \new_[11508]_  = ~\new_[11509]_  | ~\new_[12500]_ ;
  assign \new_[11509]_  = ~\new_[11405]_  | ~\new_[11407]_ ;
  assign \new_[11510]_  = \new_[2258]_  ? \new_[12765]_  : \new_[2363]_ ;
  assign \new_[11511]_  = ~\new_[5914]_  | ~\new_[3426]_  | ~\new_[11512]_ ;
  assign \new_[11512]_  = ~\new_[11513]_  & ~\new_[11516]_ ;
  assign \new_[11513]_  = ~\new_[11514]_  | ~\new_[5864]_  | ~\new_[7450]_ ;
  assign \new_[11514]_  = (~\new_[9107]_  | ~\new_[7060]_ ) & (~\new_[12385]_  | ~\new_[11515]_ );
  assign \new_[11515]_  = ~\new_[10417]_  & ~\new_[10552]_ ;
  assign \new_[11516]_  = ~\new_[11517]_  | ~\new_[11518]_ ;
  assign \new_[11517]_  = ~\new_[11777]_  | ~\new_[12628]_  | ~\new_[10250]_ ;
  assign \new_[11518]_  = (~\new_[8889]_  | ~\new_[7109]_ ) & (~\new_[6826]_  | ~\new_[11519]_ );
  assign \new_[11519]_  = \new_[11776]_  | \new_[10250]_ ;
  assign \new_[11520]_  = ~\new_[11522]_  & (~\new_[11976]_  | ~\new_[11521]_ );
  assign \new_[11521]_  = ~\new_[11529]_  & ~\new_[10088]_ ;
  assign \new_[11522]_  = ~\new_[11523]_  | ~\new_[11527]_ ;
  assign \new_[11523]_  = ~\new_[11526]_  | ~\new_[12702]_  | ~\new_[12673]_ ;
  assign \new_[11524]_  = ~\new_[11525]_  | ~\new_[7177]_ ;
  assign \new_[11525]_  = ~\new_[10203]_  | ~\new_[11779]_ ;
  assign \new_[11526]_  = \new_[1470]_ ;
  assign \new_[11527]_  = ~\new_[11526]_  | ~\new_[12655]_  | ~\new_[11528]_ ;
  assign \new_[11528]_  = ~\new_[11525]_ ;
  assign \new_[11529]_  = ~\new_[11526]_ ;
  assign \new_[11530]_  = ~\new_[1470]_ ;
  assign n761 = ~\new_[11536]_  | ~\new_[11532]_  | ~\new_[11534]_ ;
  assign \new_[11532]_  = ~\new_[2696]_  & ~\new_[11533]_ ;
  assign \new_[11533]_  = ~\new_[1701]_ ;
  assign \new_[11534]_  = ~\new_[11535]_ ;
  assign \new_[11535]_  = ~\new_[4251]_  | ~\new_[3287]_  | ~\new_[6168]_  | ~\new_[2907]_ ;
  assign \new_[11536]_  = ~\new_[11537]_  & ~\new_[2776]_ ;
  assign \new_[11537]_  = ~\new_[6127]_  | ~\new_[11538]_  | ~\new_[1968]_ ;
  assign \new_[11538]_  = \new_[2033]_  & \new_[5517]_ ;
  assign n776 = ~\new_[11544]_  | ~\new_[11540]_  | ~\new_[11543]_ ;
  assign \new_[11540]_  = ~\new_[11541]_  & ~\new_[2797]_ ;
  assign \new_[11541]_  = ~\new_[6148]_  | ~\new_[11542]_  | ~\new_[1943]_ ;
  assign \new_[11542]_  = \new_[2014]_  & \new_[5597]_ ;
  assign \new_[11543]_  = \new_[1705]_  & \new_[6191]_ ;
  assign \new_[11544]_  = ~\new_[11545]_  & ~\new_[2763]_ ;
  assign \new_[11545]_  = ~\new_[2918]_  | ~\new_[11546]_ ;
  assign \new_[11546]_  = \new_[3151]_  & \new_[4601]_ ;
  assign n781 = ~\new_[11550]_  | ~\new_[1706]_  | ~\new_[11548]_  | ~\new_[11549]_ ;
  assign \new_[11548]_  = ~\new_[2798]_  & ~\new_[2832]_ ;
  assign \new_[11549]_  = \new_[6196]_  & \new_[6149]_ ;
  assign \new_[11550]_  = ~\new_[11551]_  & ~\new_[11552]_ ;
  assign \new_[11551]_  = ~\new_[4259]_  | ~\new_[3134]_  | ~\new_[3302]_ ;
  assign \new_[11552]_  = ~\new_[5602]_  | ~\new_[1945]_  | ~\new_[2015]_ ;
  assign \new_[11553]_  = ~\new_[12573]_ ;
  assign \new_[11554]_  = ~\new_[7875]_  | ~\new_[10504]_ ;
  assign \new_[11555]_  = ~\new_[11556]_ ;
  assign \new_[11556]_  = \new_[11557]_  | \new_[11558]_ ;
  assign \new_[11557]_  = \new_[7302]_  | \new_[7295]_ ;
  assign \new_[11558]_  = ~\new_[12532]_  | ~\new_[11559]_ ;
  assign \new_[11559]_  = ~\new_[10325]_  & ~\new_[7861]_ ;
  assign \new_[11560]_  = ~\new_[12533]_ ;
  assign n766 = ~\new_[11567]_  | ~\new_[11562]_  | ~\new_[11564]_ ;
  assign \new_[11562]_  = ~\new_[2699]_  & ~\new_[11563]_ ;
  assign \new_[11563]_  = ~\new_[1702]_ ;
  assign \new_[11564]_  = ~\new_[11565]_  & ~\new_[2681]_ ;
  assign \new_[11565]_  = ~\new_[6136]_  | ~\new_[11566]_  | ~\new_[1976]_ ;
  assign \new_[11566]_  = \new_[2036]_  & \new_[5539]_ ;
  assign \new_[11567]_  = ~\new_[11568]_ ;
  assign \new_[11568]_  = ~\new_[4588]_  | ~\new_[3293]_  | ~\new_[6175]_  | ~\new_[2909]_ ;
  assign \new_[11569]_  = ~\new_[10029]_  | ~\new_[2605]_  | ~\new_[11570]_ ;
  assign \new_[11570]_  = ~\new_[11571]_  & ~\new_[11574]_ ;
  assign \new_[11571]_  = ~\new_[11572]_  | ~\new_[11573]_ ;
  assign \new_[11572]_  = ~\new_[10962]_  & ~\new_[11333]_ ;
  assign \new_[11573]_  = \new_[10320]_  & \new_[10673]_ ;
  assign \new_[11574]_  = ~\new_[11575]_  | ~\new_[10157]_  | ~\new_[10301]_  | ~\new_[10240]_ ;
  assign \new_[11575]_  = \new_[11951]_ ;
  assign \new_[11576]_  = ~\new_[11575]_ ;
  assign \new_[11577]_  = ~\new_[12210]_  & ~\new_[12211]_ ;
  assign \new_[11578]_  = ~\new_[11586]_  | (~\new_[11579]_  & ~\new_[11584]_ );
  assign \new_[11579]_  = ~\new_[2145]_  | ~\new_[11580]_  | ~\new_[2144]_  | ~\new_[6497]_ ;
  assign \new_[11580]_  = \new_[6108]_  & \new_[11581]_ ;
  assign \new_[11581]_  = ~\new_[11582]_  & ~\new_[11583]_ ;
  assign \new_[11582]_  = ~\new_[7998]_  | ~\new_[7679]_  | ~\new_[7309]_  | ~\new_[12382]_ ;
  assign \new_[11583]_  = ~\new_[7323]_ ;
  assign \new_[11584]_  = ~\new_[2606]_  | ~\new_[11585]_  | ~\new_[5880]_ ;
  assign \new_[11585]_  = ~\new_[10001]_  | ~\new_[6015]_  | ~\new_[7432]_ ;
  assign \new_[11586]_  = \new_[2606]_  | n2936;
  assign n2936 = \new_[12506]_ ;
  assign \new_[11588]_  = ~\new_[2144]_  | ~\new_[11585]_  | ~\new_[11589]_  | ~\new_[11590]_ ;
  assign \new_[11589]_  = \new_[6497]_  & \new_[11580]_ ;
  assign \new_[11590]_  = \new_[2145]_  & \new_[5880]_ ;
  assign n846 = ~\new_[11597]_  | ~\new_[11595]_  | ~\new_[11592]_  | ~\new_[11594]_ ;
  assign \new_[11592]_  = ~\new_[11593]_ ;
  assign \new_[11593]_  = ~\new_[5924]_  | ~\new_[1734]_ ;
  assign \new_[11594]_  = ~\new_[2791]_ ;
  assign \new_[11595]_  = ~\new_[11596]_  & ~\new_[2746]_ ;
  assign \new_[11596]_  = ~\new_[4031]_  | ~\new_[2998]_  | ~\new_[3371]_ ;
  assign \new_[11597]_  = ~\new_[11598]_ ;
  assign \new_[11598]_  = ~\new_[6621]_  | ~\new_[6131]_  | ~\new_[1972]_  | ~\new_[2034]_ ;
  assign n811 = ~\new_[11604]_  | ~\new_[11602]_  | ~\new_[11600]_  | ~\new_[11601]_ ;
  assign \new_[11600]_  = \new_[6169]_  & \new_[1732]_ ;
  assign \new_[11601]_  = ~\new_[2788]_ ;
  assign \new_[11602]_  = ~\new_[11603]_  & ~\new_[2687]_ ;
  assign \new_[11603]_  = ~\new_[5921]_  | ~\new_[1969]_  | ~\new_[2007]_ ;
  assign \new_[11604]_  = ~\new_[11605]_ ;
  assign \new_[11605]_  = ~\new_[4252]_  | ~\new_[6128]_  | ~\new_[2908]_  | ~\new_[3288]_ ;
  assign n831 = ~\new_[11611]_  | ~\new_[11607]_  | ~\new_[11610]_ ;
  assign \new_[11607]_  = ~\new_[11608]_  & ~\new_[2792]_ ;
  assign \new_[11608]_  = ~\new_[6132]_  | ~\new_[11609]_  | ~\new_[1973]_ ;
  assign \new_[11609]_  = \new_[2009]_  & \new_[5530]_ ;
  assign \new_[11610]_  = \new_[6172]_  & \new_[1735]_ ;
  assign \new_[11611]_  = ~\new_[11612]_  & ~\new_[2747]_ ;
  assign \new_[11612]_  = ~\new_[3027]_  | ~\new_[11613]_ ;
  assign \new_[11613]_  = \new_[3291]_  & \new_[4254]_ ;
  assign n866 = ~\new_[11620]_  | ~\new_[11617]_  | ~\new_[11615]_  | ~\new_[11616]_ ;
  assign \new_[11615]_  = \new_[6183]_  & \new_[1743]_ ;
  assign \new_[11616]_  = ~\new_[2703]_ ;
  assign \new_[11617]_  = ~\new_[11618]_  & ~\new_[2671]_ ;
  assign \new_[11618]_  = ~\new_[2914]_  | ~\new_[11619]_ ;
  assign \new_[11619]_  = \new_[3297]_  & \new_[4257]_ ;
  assign \new_[11620]_  = ~\new_[11621]_ ;
  assign \new_[11621]_  = ~\new_[5557]_  | ~\new_[6141]_  | ~\new_[1926]_  | ~\new_[1983]_ ;
  assign n876 = ~\new_[11623]_  | ~\new_[11629]_ ;
  assign \new_[11623]_  = \new_[11624]_  & \new_[11627]_ ;
  assign \new_[11624]_  = ~\new_[11625]_  & ~\new_[2750]_ ;
  assign \new_[11625]_  = ~\new_[2912]_  | ~\new_[11626]_ ;
  assign \new_[11626]_  = \new_[3296]_  & \new_[4594]_ ;
  assign \new_[11627]_  = ~\new_[11628]_ ;
  assign \new_[11628]_  = ~\new_[5553]_  | ~\new_[6140]_  | ~\new_[1925]_  | ~\new_[1982]_ ;
  assign \new_[11629]_  = ~\new_[2734]_  & ~\new_[11630]_ ;
  assign \new_[11630]_  = ~\new_[6180]_  | ~\new_[1742]_ ;
  assign n911 = ~\new_[11636]_  | ~\new_[11632]_  | ~\new_[11634]_ ;
  assign \new_[11632]_  = ~\new_[2800]_  & ~\new_[11633]_ ;
  assign \new_[11633]_  = ~\new_[1756]_ ;
  assign \new_[11634]_  = ~\new_[11635]_ ;
  assign \new_[11635]_  = ~\new_[4261]_  | ~\new_[3037]_  | ~\new_[6184]_  | ~\new_[2921]_ ;
  assign \new_[11636]_  = ~\new_[11637]_  & ~\new_[2738]_ ;
  assign \new_[11637]_  = ~\new_[6151]_  | ~\new_[11638]_  | ~\new_[1949]_ ;
  assign \new_[11638]_  = \new_[2017]_  & \new_[5975]_ ;
  assign n801 = ~\new_[11644]_  | ~\new_[11640]_  | ~\new_[11642]_ ;
  assign \new_[11640]_  = ~\new_[2775]_  & ~\new_[11641]_ ;
  assign \new_[11641]_  = ~\new_[1730]_ ;
  assign \new_[11642]_  = ~\new_[11643]_  & ~\new_[2694]_ ;
  assign \new_[11643]_  = ~\new_[5510]_  | ~\new_[6125]_  | ~\new_[1964]_  | ~\new_[2005]_ ;
  assign \new_[11644]_  = ~\new_[11645]_ ;
  assign \new_[11645]_  = ~\new_[4248]_  | ~\new_[3286]_  | ~\new_[6167]_  | ~\new_[2906]_ ;
  assign n841 = ~\new_[11651]_  | ~\new_[11649]_  | ~\new_[11647]_  | ~\new_[11648]_ ;
  assign \new_[11647]_  = \new_[6174]_  & \new_[1737]_ ;
  assign \new_[11648]_  = ~\new_[2793]_ ;
  assign \new_[11649]_  = ~\new_[11650]_  & ~\new_[2698]_ ;
  assign \new_[11650]_  = ~\new_[5926]_  | ~\new_[1975]_  | ~\new_[2010]_ ;
  assign \new_[11651]_  = ~\new_[11652]_ ;
  assign \new_[11652]_  = ~\new_[6135]_  | ~\new_[4604]_  | ~\new_[3251]_  | ~\new_[3292]_ ;
  assign n851 = ~\new_[11659]_  | ~\new_[11656]_  | ~\new_[11654]_  | ~\new_[11655]_ ;
  assign \new_[11654]_  = \new_[6177]_  & \new_[1738]_ ;
  assign \new_[11655]_  = ~\new_[2794]_ ;
  assign \new_[11656]_  = ~\new_[11657]_  & ~\new_[2700]_ ;
  assign \new_[11657]_  = ~\new_[11658]_  | ~\new_[3128]_ ;
  assign \new_[11658]_  = \new_[3295]_  & \new_[4256]_ ;
  assign \new_[11659]_  = ~\new_[11660]_ ;
  assign \new_[11660]_  = ~\new_[5542]_  | ~\new_[6137]_  | ~\new_[1978]_  | ~\new_[2038]_ ;
  assign n861 = ~\new_[11662]_  | ~\new_[11668]_ ;
  assign \new_[11662]_  = \new_[11663]_  & \new_[11666]_ ;
  assign \new_[11663]_  = ~\new_[11664]_  & ~\new_[2749]_ ;
  assign \new_[11664]_  = ~\new_[2911]_  | ~\new_[11665]_ ;
  assign \new_[11665]_  = \new_[3141]_  & \new_[4591]_ ;
  assign \new_[11666]_  = ~\new_[11667]_ ;
  assign \new_[11667]_  = ~\new_[5548]_  | ~\new_[6139]_  | ~\new_[1981]_  | ~\new_[2041]_ ;
  assign \new_[11668]_  = ~\new_[2733]_  & ~\new_[11669]_ ;
  assign \new_[11669]_  = ~\new_[6179]_  | ~\new_[1740]_ ;
  assign \new_[11670]_  = \new_[3303]_  & \new_[4260]_ ;
  assign n836 = ~\new_[11676]_  | ~\new_[11672]_  | ~\new_[11675]_ ;
  assign \new_[11672]_  = ~\new_[11673]_  & ~\new_[2643]_ ;
  assign \new_[11673]_  = ~\new_[6134]_  | ~\new_[11674]_  | ~\new_[1974]_ ;
  assign \new_[11674]_  = \new_[2035]_  & \new_[5534]_ ;
  assign \new_[11675]_  = \new_[6173]_  & \new_[1736]_ ;
  assign \new_[11676]_  = ~\new_[11677]_  & ~\new_[2748]_ ;
  assign \new_[11677]_  = ~\new_[3127]_  | ~\new_[11678]_ ;
  assign \new_[11678]_  = \new_[3139]_  & \new_[4587]_ ;
  assign n856 = ~\new_[11686]_  | ~\new_[11683]_  | ~\new_[11680]_  | ~\new_[11682]_ ;
  assign \new_[11680]_  = ~\new_[11681]_ ;
  assign \new_[11681]_  = ~\new_[6178]_  | ~\new_[1739]_ ;
  assign \new_[11682]_  = ~\new_[2701]_ ;
  assign \new_[11683]_  = ~\new_[2672]_  & ~\new_[11684]_ ;
  assign \new_[11684]_  = ~\new_[2910]_  | ~\new_[11685]_ ;
  assign \new_[11685]_  = \new_[3140]_  & \new_[4590]_ ;
  assign \new_[11686]_  = ~\new_[11687]_ ;
  assign \new_[11687]_  = ~\new_[5545]_  | ~\new_[6138]_  | ~\new_[1980]_  | ~\new_[2040]_ ;
  assign n886 = ~\new_[11692]_  | ~\new_[11689]_  | ~\new_[11691]_ ;
  assign \new_[11689]_  = ~\new_[11690]_ ;
  assign \new_[11690]_  = ~\new_[6142]_  | ~\new_[1748]_  | ~\new_[6189]_ ;
  assign \new_[11691]_  = ~\new_[2712]_  & ~\new_[2629]_ ;
  assign \new_[11692]_  = ~\new_[11693]_  & ~\new_[11694]_ ;
  assign \new_[11693]_  = ~\new_[5577]_  | ~\new_[1932]_  | ~\new_[1985]_ ;
  assign \new_[11694]_  = ~\new_[4597]_  | ~\new_[2916]_  | ~\new_[3298]_ ;
  assign n816 = ~\new_[11701]_  | ~\new_[11696]_  | ~\new_[11698]_  | ~\new_[11697]_ ;
  assign \new_[11696]_  = ~\new_[2789]_ ;
  assign \new_[11697]_  = \new_[1733]_  & \new_[6170]_ ;
  assign \new_[11698]_  = ~\new_[11699]_  & ~\new_[2697]_ ;
  assign \new_[11699]_  = ~\new_[3126]_  | ~\new_[11700]_ ;
  assign \new_[11700]_  = \new_[3124]_  & \new_[4585]_ ;
  assign \new_[11701]_  = ~\new_[11702]_ ;
  assign \new_[11702]_  = ~\new_[5922]_  | ~\new_[6129]_  | ~\new_[1970]_  | ~\new_[2008]_ ;
  assign \new_[11703]_  = ~\new_[11704]_  & ~\new_[11705]_ ;
  assign \new_[11704]_  = ~\new_[11833]_  & (~\new_[8402]_  | ~\new_[10018]_ );
  assign \new_[11705]_  = \new_[11706]_  & \new_[11833]_ ;
  assign \new_[11706]_  = ~\new_[11831]_  | ~\new_[11707]_ ;
  assign \new_[11707]_  = (~\new_[11251]_  | ~\new_[12622]_ ) & (~\new_[12621]_  | ~\new_[11104]_ );
  assign \new_[11708]_  = ~\new_[11761]_  | ~\new_[11950]_  | ~\new_[11838]_ ;
  assign \new_[11709]_  = ~\new_[11259]_  | ~\new_[12275]_ ;
  assign \new_[11710]_  = ~\new_[11711]_  | ~\new_[11712]_ ;
  assign \new_[11711]_  = ~\new_[12213]_ ;
  assign \new_[11712]_  = \new_[12037]_ ;
  assign \new_[11713]_  = ~\new_[11709]_ ;
  assign \new_[11714]_  = ~\new_[11712]_ ;
  assign \new_[11715]_  = \new_[11716]_  | \new_[11719]_ ;
  assign \new_[11716]_  = \new_[11717]_  & \new_[7373]_ ;
  assign \new_[11717]_  = ~\new_[11718]_  & ~\new_[7717]_ ;
  assign \new_[11718]_  = \new_[11224]_  ? \new_[12623]_  : \new_[11060]_ ;
  assign \new_[11719]_  = ~\new_[7714]_  & ~\new_[7118]_ ;
  assign \new_[11720]_  = ~\new_[11721]_  & ~\new_[11722]_ ;
  assign \new_[11721]_  = ~\new_[12599]_  | ~\new_[9570]_  | ~\new_[9266]_ ;
  assign \new_[11722]_  = ~\new_[12463]_  | ~\new_[12609]_ ;
  assign \new_[11723]_  = ~\new_[12463]_ ;
  assign \new_[11724]_  = ~\new_[12096]_ ;
  assign \new_[11725]_  = \new_[11726]_  & \new_[7373]_ ;
  assign \new_[11726]_  = \new_[7717]_  & \new_[7714]_ ;
  assign \new_[11727]_  = ~\new_[11728]_  | ~\new_[11731]_ ;
  assign \new_[11728]_  = ~\new_[11729]_  | (~\new_[12623]_  & ~\new_[2315]_ );
  assign \new_[11729]_  = ~\new_[12623]_  | ~\new_[11730]_ ;
  assign \new_[11730]_  = ~\new_[2381]_ ;
  assign \new_[11731]_  = ~\new_[11732]_ ;
  assign \new_[11732]_  = (~\new_[2316]_  | ~\new_[12624]_ ) & (~\new_[12623]_  | ~\new_[2364]_ );
  assign \new_[11733]_  = ~\new_[11726]_ ;
  assign \new_[11734]_  = ~\new_[11735]_  | ~\new_[12695]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[11735]_  = ~\new_[11881]_ ;
  assign \new_[11736]_  = ~\new_[12552]_  | ~\new_[10522]_ ;
  assign \new_[11737]_  = \new_[11953]_ ;
  assign \new_[11738]_  = ~\new_[11824]_  & ~\new_[11825]_ ;
  assign \new_[11739]_  = ~\new_[12676]_  | ~\new_[2486]_ ;
  assign \new_[11740]_  = ~\new_[11824]_ ;
  assign \new_[11741]_  = ~\new_[11748]_  | (~\new_[11742]_  & ~\new_[11743]_ );
  assign \new_[11742]_  = \new_[6282]_  & \new_[1759]_ ;
  assign \new_[11743]_  = ~\new_[11744]_  | ~\new_[11940]_ ;
  assign \new_[11744]_  = \new_[11745]_  & \new_[4293]_ ;
  assign \new_[11745]_  = ~\new_[11746]_  & ~\new_[5839]_ ;
  assign \new_[11746]_  = ~\new_[11747]_ ;
  assign \new_[11747]_  = \new_[7747]_  | \new_[12664]_ ;
  assign \new_[11748]_  = ~\new_[11749]_ ;
  assign \new_[11749]_  = ~\new_[11750]_  & ~\new_[11941]_ ;
  assign \new_[11750]_  = \new_[11106]_  ? \new_[12622]_  : \new_[11136]_ ;
  assign \new_[11751]_  = ~\new_[11752]_ ;
  assign \new_[11752]_  = \new_[8847]_ ;
  assign \new_[11753]_  = \new_[12392]_  & \new_[11752]_ ;
  assign \new_[11754]_  = ~\new_[12071]_  | ~\new_[12237]_ ;
  assign \new_[11755]_  = ~\new_[11984]_  | ~\new_[11985]_ ;
  assign \new_[11756]_  = ~\new_[11843]_ ;
  assign \new_[11757]_  = ~\new_[7875]_  | ~\new_[10504]_ ;
  assign \new_[11758]_  = ~\new_[11951]_ ;
  assign \new_[11759]_  = ~\new_[11760]_ ;
  assign \new_[11760]_  = ~\new_[1489]_ ;
  assign \new_[11761]_  = ~\new_[11759]_ ;
  assign \new_[11762]_  = ~\new_[11955]_ ;
  assign \new_[11763]_  = ~\new_[12098]_ ;
  assign \new_[11764]_  = ~\new_[11769]_  | ~\new_[11765]_  | ~\new_[11768]_ ;
  assign \new_[11765]_  = ~\new_[11766]_  | ~\new_[11767]_ ;
  assign \new_[11766]_  = ~\new_[2002]_  | ~\new_[2147]_ ;
  assign \new_[11767]_  = ~\new_[1433]_  & ~\new_[7078]_ ;
  assign \new_[11768]_  = ~\new_[11993]_  & ~\new_[4589]_ ;
  assign \new_[11769]_  = ~\new_[11770]_  & (~\new_[12789]_  | ~\new_[9571]_ );
  assign \new_[11770]_  = ~\new_[11771]_  | ~\new_[11775]_ ;
  assign \new_[11771]_  = (~\new_[11772]_  | ~\new_[11773]_ ) & (~\new_[11864]_  | ~\new_[11772]_ );
  assign \new_[11772]_  = ~\new_[10551]_  & ~\new_[11776]_ ;
  assign \new_[11773]_  = ~\new_[11774]_ ;
  assign \new_[11774]_  = \new_[12211]_  | \new_[9984]_ ;
  assign \new_[11775]_  = (~\new_[9300]_  | ~\new_[7109]_ ) & (~\new_[7327]_  | ~\new_[11772]_ );
  assign \new_[11776]_  = ~\new_[1433]_ ;
  assign \new_[11777]_  = ~\new_[11778]_  | ~\new_[3036]_ ;
  assign \new_[11778]_  = ~\new_[11779]_ ;
  assign \new_[11779]_  = ~\new_[12429]_  | ~\new_[9939]_  | ~n5291;
  assign n5291 = ~\new_[10785]_  & ~\new_[10884]_ ;
  assign \new_[11781]_  = ~\new_[11782]_  | (~\new_[1869]_  & ~\new_[5639]_ );
  assign \new_[11782]_  = ~\new_[11783]_  & ~\new_[11788]_ ;
  assign \new_[11783]_  = ~\new_[11785]_  | ~\new_[11784]_  | ~\new_[11994]_  | ~\new_[5251]_ ;
  assign \new_[11784]_  = (~\new_[9383]_  | ~\new_[7060]_ ) & (~\new_[7109]_  | ~\new_[9048]_ );
  assign \new_[11785]_  = ~\new_[11786]_  | ~\new_[11787]_ ;
  assign \new_[11786]_  = ~\new_[12061]_ ;
  assign \new_[11787]_  = ~\new_[10402]_  & ~\new_[11062]_ ;
  assign \new_[11788]_  = ~\new_[7564]_  & (~\new_[2049]_  | ~\new_[11777]_ );
  assign \new_[11789]_  = (~\new_[4531]_  | ~\new_[12670]_ ) & (~\new_[11792]_  | ~\new_[4448]_ );
  assign \new_[11790]_  = ~\new_[11791]_  & ~\new_[7152]_  & ~\new_[7119]_  & ~\new_[7151]_ ;
  assign \new_[11791]_  = ~\new_[7150]_ ;
  assign \new_[11792]_  = ~\new_[11793]_  & ~\new_[7151]_  & ~\new_[7119]_  & ~\new_[7150]_ ;
  assign \new_[11793]_  = ~\new_[7152]_ ;
  assign \new_[11794]_  = \new_[7119]_ ;
  assign \new_[11795]_  = ~\new_[7119]_ ;
  assign \new_[11796]_  = \new_[12581]_  | \new_[11409]_ ;
  assign \new_[11797]_  = ~\new_[11801]_  | ~\new_[11798]_  | ~\new_[11799]_ ;
  assign \new_[11798]_  = (~\new_[4350]_  | ~\new_[11790]_ ) & (~\new_[11792]_  | ~\new_[4474]_ );
  assign \new_[11799]_  = ~\new_[11800]_  | ~\new_[4231]_ ;
  assign \new_[11800]_  = ~\new_[11476]_  & ~\new_[7119]_  & ~\new_[7152]_  & ~\new_[7150]_ ;
  assign \new_[11801]_  = ~\new_[11802]_  | ~\new_[4518]_ ;
  assign \new_[11802]_  = \new_[11803]_ ;
  assign \new_[11803]_  = \new_[11804]_  & \new_[11805]_ ;
  assign \new_[11804]_  = ~\new_[11795]_  & ~\new_[7150]_ ;
  assign \new_[11805]_  = ~\new_[7151]_  & ~\new_[7152]_ ;
  assign \new_[11806]_  = n5041 & \new_[7908]_ ;
  assign \new_[11807]_  = ~\new_[11810]_  | ~\new_[12728]_  | ~\new_[11808]_  | ~\new_[11809]_ ;
  assign \new_[11808]_  = ~\new_[9058]_  | ~\new_[8877]_  | ~\new_[7590]_  | ~\new_[8714]_ ;
  assign \new_[11809]_  = ~\new_[11432]_  & ~\new_[7543]_ ;
  assign \new_[11810]_  = ~\new_[11811]_  | ~\new_[11812]_ ;
  assign \new_[11811]_  = \new_[12091]_  & \new_[9681]_ ;
  assign \new_[11812]_  = ~\new_[8869]_  & ~\new_[12447]_ ;
  assign \new_[11813]_  = ~\new_[11810]_ ;
  assign \new_[11814]_  = ~\new_[12513]_ ;
  assign \new_[11815]_  = ~\new_[11816]_  | ~\new_[11817]_ ;
  assign \new_[11816]_  = ~n5451;
  assign \new_[11817]_  = ~\new_[1485]_ ;
  assign \new_[11818]_  = ~\new_[11953]_  | ~\new_[11954]_ ;
  assign \new_[11819]_  = \new_[12585]_  & \new_[10336]_ ;
  assign \new_[11820]_  = ~\new_[11821]_  & ~\new_[11823]_ ;
  assign \new_[11821]_  = (~\new_[11826]_  | ~\new_[2486]_ ) & (~\new_[12724]_  | ~\new_[11822]_ );
  assign \new_[11822]_  = ~\new_[7602]_  | ~\new_[7605]_ ;
  assign \new_[11823]_  = ~\new_[11826]_  & ~\new_[2486]_ ;
  assign \new_[11824]_  = ~\new_[7602]_  & ~\new_[11828]_ ;
  assign \new_[11825]_  = ~\new_[7605]_  & ~\new_[11828]_ ;
  assign \new_[11826]_  = ~\new_[11827]_  & ~\new_[11828]_ ;
  assign \new_[11827]_  = \new_[11171]_  ? \new_[12622]_  : \new_[11132]_ ;
  assign \new_[11828]_  = ~\new_[12725]_  | ~\new_[12579]_  | ~\new_[11845]_ ;
  assign \new_[11829]_  = ~\new_[11834]_  & (~\new_[11830]_  | ~\new_[11833]_ );
  assign \new_[11830]_  = ~\new_[11831]_  | ~\new_[11832]_ ;
  assign \new_[11831]_  = ~\new_[12590]_ ;
  assign \new_[11832]_  = (~\new_[11128]_  | ~\new_[12622]_ ) & (~\new_[12621]_  | ~\new_[10993]_ );
  assign \new_[11833]_  = ~\new_[12184]_  | ~\new_[11575]_  | ~\new_[11334]_  | ~\new_[12274]_ ;
  assign \new_[11834]_  = ~\new_[11833]_  & (~\new_[8491]_  | ~\new_[10018]_ );
  assign \new_[11835]_  = \new_[2478]_  ? \new_[12617]_  : \new_[2390]_ ;
  assign \new_[11836]_  = ~\new_[11818]_ ;
  assign \new_[11837]_  = ~\new_[11759]_  & ~\new_[11758]_ ;
  assign \new_[11838]_  = ~\new_[11815]_ ;
  assign \new_[11839]_  = ~\new_[12054]_  | ~\new_[12695]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[11840]_  = ~\new_[12547]_ ;
  assign \new_[11841]_  = ~\new_[12513]_ ;
  assign \new_[11842]_  = \new_[11843]_ ;
  assign \new_[11843]_  = ~\new_[11983]_  | ~\new_[11757]_ ;
  assign \new_[11844]_  = \new_[3438]_  ? \new_[12588]_  : \new_[4242]_ ;
  assign \new_[11845]_  = ~\new_[11842]_  | ~\new_[11844]_ ;
  assign \new_[11846]_  = ~\new_[11842]_ ;
  assign \new_[11847]_  = ~\new_[11848]_  | ~\new_[11850]_ ;
  assign \new_[11848]_  = ~\new_[11849]_  & (~\new_[12751]_  | ~\new_[9841]_ );
  assign \new_[11849]_  = ~\new_[7424]_  & ~\new_[12704]_ ;
  assign \new_[11850]_  = ~\new_[11851]_  & (~\new_[7540]_  | ~\new_[9865]_ );
  assign \new_[11851]_  = \new_[5473]_  | \new_[6538]_  | \new_[7678]_  | \new_[11852]_ ;
  assign \new_[11852]_  = ~\new_[11853]_ ;
  assign \new_[11853]_  = (~\new_[9865]_  | ~\new_[7873]_ ) & (~\new_[12657]_  | ~\new_[11854]_ );
  assign \new_[11854]_  = ~\new_[12564]_  & ~\new_[8408]_ ;
  assign \new_[11855]_  = ~\new_[11856]_  & ~\new_[11862]_ ;
  assign \new_[11856]_  = ~\new_[7237]_  | ~\new_[11861]_  | ~\new_[5989]_  | ~\new_[11857]_ ;
  assign \new_[11857]_  = ~\new_[11858]_  & (~\new_[6656]_  | ~\new_[10045]_ );
  assign \new_[11858]_  = ~\new_[11859]_ ;
  assign \new_[11859]_  = (~\new_[11485]_  | ~\new_[8274]_ ) & (~\new_[7067]_  | ~\new_[11860]_ );
  assign \new_[11860]_  = \new_[10154]_  & \new_[12089]_ ;
  assign \new_[11861]_  = ~\new_[7056]_ ;
  assign \new_[11862]_  = \new_[5461]_  | \new_[3397]_ ;
  assign \new_[11863]_  = ~\new_[11864]_  | ~\new_[11860]_ ;
  assign \new_[11864]_  = ~\new_[12109]_ ;
  assign \new_[11865]_  = ~\new_[11860]_ ;
  assign \new_[11866]_  = ~\new_[11867]_  | ~\new_[11870]_ ;
  assign \new_[11867]_  = ~\new_[11868]_  & ~\new_[11869]_ ;
  assign \new_[11868]_  = n4501 | \new_[10735]_  | wb_we_i | \new_[2370]_ ;
  assign \new_[11869]_  = \new_[1837]_  & \new_[7632]_ ;
  assign \new_[11870]_  = ~\new_[11874]_  | ~\new_[11873]_  | ~\new_[11871]_  | ~\new_[11872]_ ;
  assign \new_[11871]_  = ~\new_[7378]_  | ~\wb_sel_i[0] ;
  assign \new_[11872]_  = ~\new_[7377]_  | ~\wb_sel_i[2] ;
  assign \new_[11873]_  = ~\new_[7379]_  | ~\wb_sel_i[3] ;
  assign \new_[11874]_  = ~\wb_sel_i[1]  | ~\new_[7380]_ ;
  assign n1151 = ~n4501 & ~\new_[11869]_ ;
  assign \new_[11876]_  = ~\new_[11877]_ ;
  assign \new_[11877]_  = ~\new_[11836]_  | ~\new_[11837]_  | ~\new_[11838]_ ;
  assign \new_[11878]_  = ~\new_[11879]_  & ~\new_[11880]_ ;
  assign \new_[11879]_  = ~\new_[11299]_  | ~\new_[8945]_  | ~\new_[9916]_ ;
  assign \new_[11880]_  = ~\new_[12389]_  | ~\new_[11735]_ ;
  assign \new_[11881]_  = \new_[11882]_ ;
  assign \new_[11882]_  = ~\new_[1461]_ ;
  assign \new_[11883]_  = ~\new_[12054]_  | ~\new_[11884]_  | ~\new_[12239]_ ;
  assign \new_[11884]_  = \new_[11885]_ ;
  assign \new_[11885]_  = ~\new_[12549]_ ;
  assign \new_[11886]_  = ~\new_[11709]_  & ~\new_[11710]_ ;
  assign \new_[11887]_  = ~\new_[11888]_ ;
  assign \new_[11888]_  = ~\new_[11890]_  | ~\new_[12040]_  | ~\new_[10634]_ ;
  assign \new_[11889]_  = ~\new_[1540]_ ;
  assign \new_[11890]_  = ~\new_[1480]_ ;
  assign \new_[11891]_  = ~\new_[11886]_ ;
  assign \new_[11892]_  = ~\new_[11919]_ ;
  assign \new_[11893]_  = \new_[11720]_  | \new_[7220]_ ;
  assign \new_[11894]_  = ~\new_[11895]_ ;
  assign \new_[11895]_  = ~\new_[12153]_  | ~\new_[12156]_  | ~\new_[12157]_ ;
  assign \new_[11896]_  = ~\new_[4242]_ ;
  assign \new_[11897]_  = ~\new_[11898]_  | ~\new_[2055]_ ;
  assign \new_[11898]_  = ~\new_[11900]_  | ~\new_[12573]_  | ~\new_[11899]_ ;
  assign \new_[11899]_  = ~\new_[11893]_ ;
  assign \new_[11900]_  = ~\new_[6688]_  & ~\new_[7010]_ ;
  assign \new_[11901]_  = ~\new_[11902]_ ;
  assign \new_[11902]_  = ~\new_[11903]_  | (~\new_[4755]_  & ~\new_[12694]_ );
  assign \new_[11903]_  = ~\new_[11904]_  & (~\new_[7599]_  | ~\new_[2055]_ );
  assign \new_[11904]_  = \new_[11894]_  & \new_[4242]_ ;
  assign \new_[11905]_  = ~\new_[11906]_  | ~\new_[11912]_ ;
  assign \new_[11906]_  = ~\new_[1747]_  & ~\new_[11907]_ ;
  assign \new_[11907]_  = ~\new_[3594]_  | ~\new_[11908]_  | ~\new_[11909]_ ;
  assign \new_[11908]_  = ~\new_[11363]_  | ~\new_[12638]_  | ~\new_[12603]_ ;
  assign \new_[11909]_  = ~\new_[11910]_  & ~\new_[11911]_ ;
  assign \new_[11910]_  = ~\new_[6558]_  | ~\new_[5888]_ ;
  assign \new_[11911]_  = ~\new_[6728]_  | ~\new_[5057]_  | ~\new_[5945]_ ;
  assign \new_[11912]_  = ~\new_[11913]_  & (~\new_[12628]_  | ~\new_[8501]_ );
  assign \new_[11913]_  = ~\new_[7451]_  | ~\new_[3364]_  | ~\new_[4966]_ ;
  assign \new_[11914]_  = \new_[12040]_  & \new_[11917]_ ;
  assign \new_[11915]_  = ~\new_[11218]_  | ~\new_[12046]_ ;
  assign \new_[11916]_  = ~\new_[11530]_  | ~\new_[11197]_ ;
  assign \new_[11917]_  = ~\new_[11918]_ ;
  assign \new_[11918]_  = ~\new_[11890]_  | ~\new_[11889]_ ;
  assign \new_[11919]_  = ~\new_[12040]_ ;
  assign \new_[11920]_  = ~\new_[11916]_ ;
  assign \new_[11921]_  = ~\new_[11915]_ ;
  assign \new_[11922]_  = ~\new_[11929]_  | ~\new_[11923]_  | ~\new_[11924]_ ;
  assign \new_[11923]_  = ~\new_[4921]_ ;
  assign \new_[11924]_  = \new_[11925]_  & \new_[11927]_ ;
  assign \new_[11925]_  = (~\new_[9665]_  | ~\new_[6807]_ ) & (~\new_[12792]_  | ~\new_[11926]_ );
  assign \new_[11926]_  = \new_[10960]_  & \new_[10314]_ ;
  assign \new_[11927]_  = (~\new_[11928]_  | ~\new_[12308]_ ) & (~\new_[11976]_  | ~\new_[11928]_ );
  assign \new_[11928]_  = ~\new_[10799]_  & ~\new_[10417]_ ;
  assign \new_[11929]_  = ~\new_[11930]_ ;
  assign \new_[11930]_  = ~\new_[11932]_  | (~\new_[12700]_  & ~\new_[11931]_ );
  assign \new_[11931]_  = \new_[10799]_  | \new_[12672]_ ;
  assign \new_[11932]_  = \new_[11933]_  | \new_[12651]_ ;
  assign \new_[11933]_  = \new_[10799]_  | \new_[8499]_ ;
  assign \new_[11934]_  = \new_[12459]_  & \new_[10251]_ ;
  assign \new_[11935]_  = ~\new_[11942]_  | (~\new_[11936]_  & ~\new_[11938]_ );
  assign \new_[11936]_  = \new_[1824]_  & \new_[11937]_ ;
  assign \new_[11937]_  = \new_[6336]_  | \new_[6282]_ ;
  assign \new_[11938]_  = ~\new_[11939]_ ;
  assign \new_[11939]_  = \new_[11940]_  & \new_[11941]_ ;
  assign \new_[11940]_  = ~\new_[2389]_  | ~\new_[6639]_ ;
  assign \new_[11941]_  = \new_[4293]_  & \new_[11747]_ ;
  assign \new_[11942]_  = \new_[11943]_  | \new_[11941]_ ;
  assign \new_[11943]_  = \new_[11260]_  ? \new_[12619]_  : \new_[11194]_ ;
  assign \new_[11944]_  = ~\new_[11941]_ ;
  assign n5446 = \new_[8688]_  & wb_cyc_i;
  assign \new_[11946]_  = \new_[12426]_  & \new_[9939]_ ;
  assign \new_[11947]_  = ~\new_[11948]_  | ~\new_[11949]_ ;
  assign \new_[11948]_  = ~\new_[11309]_  | ~\new_[2368]_ ;
  assign \new_[11949]_  = ~\new_[12627]_  | ~\new_[2479]_ ;
  assign \new_[11950]_  = ~\new_[11758]_  & ~\new_[11952]_ ;
  assign \new_[11951]_  = ~\new_[1487]_ ;
  assign \new_[11952]_  = ~\new_[11953]_  | ~\new_[11954]_ ;
  assign \new_[11953]_  = ~\new_[1486]_ ;
  assign \new_[11954]_  = ~\new_[1492]_ ;
  assign \new_[11955]_  = ~\new_[11954]_  | ~\new_[11953]_ ;
  assign \new_[11956]_  = ~\new_[11963]_  | ~\new_[11957]_  | ~\new_[11958]_ ;
  assign \new_[11957]_  = ~\new_[4917]_ ;
  assign \new_[11958]_  = \new_[11959]_  & \new_[11961]_ ;
  assign \new_[11959]_  = (~\new_[9684]_  | ~\new_[7238]_ ) & (~\new_[12792]_  | ~\new_[11960]_ );
  assign \new_[11960]_  = \new_[11361]_  & \new_[10657]_ ;
  assign \new_[11961]_  = (~\new_[11962]_  | ~\new_[7684]_ ) & (~\new_[11976]_  | ~\new_[11962]_ );
  assign \new_[11962]_  = ~\new_[12401]_  & ~\new_[4147]_ ;
  assign \new_[11963]_  = ~\new_[11964]_ ;
  assign \new_[11964]_  = ~\new_[11966]_  | (~\new_[12700]_  & ~\new_[11965]_ );
  assign \new_[11965]_  = \new_[12401]_  | \new_[12672]_ ;
  assign \new_[11966]_  = \new_[11967]_  | \new_[12654]_ ;
  assign \new_[11967]_  = \new_[12401]_  | \new_[8499]_ ;
  assign \new_[11968]_  = ~\new_[11969]_  | ~\new_[11978]_ ;
  assign \new_[11969]_  = ~\new_[11970]_  & ~\new_[4637]_ ;
  assign \new_[11970]_  = ~\new_[11975]_  | ~\new_[11974]_  | ~\new_[11971]_  | ~\new_[11972]_ ;
  assign \new_[11971]_  = ~\new_[7076]_  | ~\new_[10115]_ ;
  assign \new_[11972]_  = ~\new_[7683]_  | ~\new_[11973]_ ;
  assign \new_[11973]_  = ~\new_[10417]_  & ~\new_[11368]_ ;
  assign \new_[11974]_  = ~\new_[10657]_  | ~\new_[12792]_  | ~\new_[11367]_ ;
  assign \new_[11975]_  = ~\new_[11976]_  | ~\new_[11973]_ ;
  assign \new_[11976]_  = ~\new_[11977]_ ;
  assign \new_[11977]_  = \new_[12170]_  & \new_[12493]_ ;
  assign \new_[11978]_  = ~\new_[11979]_ ;
  assign \new_[11979]_  = ~\new_[11981]_  | (~\new_[12713]_  & ~\new_[11980]_ );
  assign \new_[11980]_  = \new_[11368]_  | \new_[12672]_ ;
  assign \new_[11981]_  = \new_[11982]_  | \new_[12654]_ ;
  assign \new_[11982]_  = \new_[11368]_  | \new_[8499]_ ;
  assign \new_[11983]_  = ~\new_[11984]_  | ~\new_[11985]_ ;
  assign \new_[11984]_  = ~\new_[11151]_  & ~\new_[9712]_ ;
  assign \new_[11985]_  = ~\new_[11986]_  & ~\new_[12214]_ ;
  assign \new_[11986]_  = ~\new_[11019]_  | ~\new_[10079]_  | ~\new_[12038]_ ;
  assign \new_[11987]_  = ~\new_[11988]_  & ~\new_[11989]_ ;
  assign \new_[11988]_  = ~\new_[12392]_  | ~\new_[12395]_ ;
  assign \new_[11989]_  = ~\new_[10938]_  | ~\new_[11990]_  | ~\new_[9560]_  | ~\new_[8945]_ ;
  assign \new_[11990]_  = \new_[11300]_  & \new_[11882]_ ;
  assign \new_[11991]_  = \new_[11300]_  & \new_[11882]_ ;
  assign \new_[11992]_  = ~\new_[11988]_ ;
  assign \new_[11993]_  = ~\new_[12166]_ ;
  assign \new_[11994]_  = ~\new_[11995]_ ;
  assign \new_[11995]_  = ~\new_[11996]_  | ~\new_[12001]_ ;
  assign \new_[11996]_  = ~\new_[11997]_  | ~\new_[12000]_ ;
  assign \new_[11997]_  = \new_[11998]_ ;
  assign \new_[11998]_  = ~\new_[12386]_  | ~\new_[11999]_ ;
  assign \new_[11999]_  = \new_[12464]_  | \new_[8696]_ ;
  assign \new_[12000]_  = ~\new_[10402]_  & ~\new_[4147]_ ;
  assign \new_[12001]_  = ~\new_[12002]_  | ~\new_[9383]_ ;
  assign \new_[12002]_  = ~\new_[12234]_ ;
  assign \new_[12003]_  = \new_[10402]_  | \new_[10714]_ ;
  assign n946 = ~\new_[12005]_  | ~\new_[12008]_ ;
  assign \new_[12005]_  = ~\new_[12174]_  & ~\new_[12006]_ ;
  assign \new_[12006]_  = ~\new_[2862]_  | ~\new_[2691]_  | ~\new_[12007]_ ;
  assign \new_[12007]_  = ~\new_[1813]_ ;
  assign \new_[12008]_  = \new_[11855]_  & \new_[12009]_ ;
  assign \new_[12009]_  = ~\new_[12010]_  & ~\new_[12011]_ ;
  assign \new_[12010]_  = ~\new_[8005]_  | ~\new_[6726]_  | ~\new_[6185]_  | ~\new_[5935]_ ;
  assign \new_[12011]_  = ~\new_[11863]_  | ~\new_[3938]_  | ~\new_[6272]_ ;
  assign n941 = ~\new_[12017]_  | ~\new_[12015]_  | ~\new_[12013]_  | ~\new_[2913]_ ;
  assign \new_[12013]_  = ~\new_[12014]_ ;
  assign \new_[12014]_  = ~\new_[4595]_  | ~\new_[6271]_  | ~\new_[2690]_  | ~\new_[3144]_ ;
  assign \new_[12015]_  = ~\new_[1811]_  & ~\new_[12016]_ ;
  assign \new_[12016]_  = ~\new_[2861]_ ;
  assign \new_[12017]_  = ~\new_[12019]_  & (~\new_[12018]_  | ~\new_[12636]_ );
  assign \new_[12018]_  = \new_[12603]_  & \new_[11298]_ ;
  assign \new_[12019]_  = ~\new_[12023]_  | ~\new_[5556]_  | ~\new_[12020]_  | ~\new_[12022]_ ;
  assign \new_[12020]_  = ~\new_[12021]_ ;
  assign \new_[12021]_  = ~\new_[12388]_  | ~\new_[5933]_  | ~\new_[6181]_  | ~\new_[6725]_ ;
  assign \new_[12022]_  = ~\new_[11777]_  | ~\new_[12628]_  | ~\new_[11298]_ ;
  assign \new_[12023]_  = ~\new_[12064]_  | ~\new_[11504]_ ;
  assign \new_[12024]_  = ~\new_[12027]_  | (~\new_[12025]_  & ~\new_[12026]_ );
  assign \new_[12025]_  = ~\new_[4151]_  & ~\new_[2066]_ ;
  assign \new_[12026]_  = ~\new_[2240]_  | ~\new_[12337]_ ;
  assign \new_[12027]_  = ~\new_[12030]_  & (~\new_[12028]_  | ~\new_[12338]_ );
  assign \new_[12028]_  = ~\new_[12029]_  | (~\new_[2554]_  & ~\new_[11740]_ );
  assign \new_[12029]_  = ~\new_[2554]_  | ~\new_[11740]_ ;
  assign \new_[12030]_  = ~\new_[12340]_ ;
  assign \new_[12031]_  = ~\new_[12032]_ ;
  assign \new_[12032]_  = ~\new_[11713]_  | ~\new_[12033]_  | ~\new_[11917]_ ;
  assign \new_[12033]_  = ~\new_[11916]_  & ~\new_[11915]_ ;
  assign \new_[12034]_  = ~\new_[12035]_  & ~\new_[12036]_ ;
  assign \new_[12035]_  = ~\new_[10401]_  | ~\new_[10471]_ ;
  assign \new_[12036]_  = ~\new_[10486]_  | ~\new_[12153]_ ;
  assign \new_[12037]_  = ~\new_[12035]_  & ~\new_[12036]_ ;
  assign \new_[12038]_  = ~\new_[12039]_ ;
  assign \new_[12039]_  = ~\new_[11713]_  | ~\new_[11917]_ ;
  assign \new_[12040]_  = ~\new_[11916]_  & ~\new_[11915]_ ;
  assign \new_[12041]_  = \new_[12042]_  | \new_[1817]_ ;
  assign \new_[12042]_  = ~\new_[12048]_  | ~\new_[12047]_  | ~\new_[12043]_ ;
  assign \new_[12043]_  = ~\new_[12044]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[12044]_  = ~\new_[12045]_ ;
  assign \new_[12045]_  = \new_[12046]_ ;
  assign \new_[12046]_  = ~\new_[1534]_ ;
  assign \new_[12047]_  = ~\new_[12044]_  | ~\new_[12635]_  | ~\new_[12606]_ ;
  assign \new_[12048]_  = ~\new_[12064]_  | ~\new_[9594]_ ;
  assign \new_[12049]_  = \new_[12050]_  ? \new_[12052]_  : \new_[12051]_ ;
  assign \new_[12050]_  = \new_[11390]_  | \new_[10873]_ ;
  assign \new_[12051]_  = (~\new_[10873]_  | ~\new_[8457]_ ) & (~\new_[8671]_  | ~\new_[9815]_ );
  assign \new_[12052]_  = \new_[12053]_ ;
  assign \new_[12053]_  = ~\new_[1502]_ ;
  assign \new_[12054]_  = ~\new_[12052]_ ;
  assign \new_[12055]_  = ~\new_[12063]_  | ~\new_[12056]_  | ~\new_[12057]_ ;
  assign \new_[12056]_  = \new_[5639]_  | \new_[1764]_ ;
  assign \new_[12057]_  = ~\new_[12058]_  & ~\new_[3389]_ ;
  assign \new_[12058]_  = ~\new_[12062]_  | ~\new_[4760]_  | ~\new_[12059]_ ;
  assign \new_[12059]_  = (~\new_[12060]_  | ~\new_[6656]_ ) & (~\new_[11786]_  | ~\new_[12060]_ );
  assign \new_[12060]_  = ~\new_[10747]_  & ~\new_[11062]_ ;
  assign \new_[12061]_  = \new_[11449]_  & \new_[11450]_ ;
  assign \new_[12062]_  = ~\new_[7052]_  & (~\new_[7067]_  | ~\new_[9979]_ );
  assign \new_[12063]_  = ~\new_[12645]_  | ~\new_[10838]_  | ~\new_[12602]_ ;
  assign \new_[12064]_  = ~\new_[12061]_ ;
  assign n1686 = ~\new_[12067]_  | ~\new_[12066]_  | ~\new_[11457]_  | ~\new_[11459]_ ;
  assign \new_[12066]_  = ~\new_[6841]_  | ~\new_[3036]_ ;
  assign \new_[12067]_  = ~\new_[12068]_  & ~\new_[7132]_ ;
  assign \new_[12068]_  = ~\new_[12069]_  | ~\new_[12070]_ ;
  assign \new_[12069]_  = ~\new_[10110]_  | ~\new_[8874]_  | ~\new_[11811]_  | ~\new_[8175]_ ;
  assign \new_[12070]_  = \new_[12071]_ ;
  assign \new_[12071]_  = ~\new_[11711]_  | ~\new_[12072]_ ;
  assign \new_[12072]_  = ~\new_[8866]_  & ~\new_[12073]_ ;
  assign \new_[12073]_  = \new_[12275]_  | \new_[11714]_ ;
  assign \new_[12074]_  = ~\new_[12070]_ ;
  assign \new_[12075]_  = ~\new_[12069]_ ;
  assign n1076 = ~\new_[12088]_  | ~\new_[12085]_  | ~\new_[12077]_  | ~\new_[12080]_ ;
  assign \new_[12077]_  = \new_[12078]_  & \new_[12079]_ ;
  assign \new_[12078]_  = ~\new_[2751]_ ;
  assign \new_[12079]_  = ~\new_[3441]_  & ~\new_[5502]_ ;
  assign \new_[12080]_  = \new_[12081]_  & \new_[12082]_ ;
  assign \new_[12081]_  = \new_[3228]_  & \new_[2972]_ ;
  assign \new_[12082]_  = ~\new_[12083]_  & ~\new_[12084]_ ;
  assign \new_[12083]_  = ~\new_[7679]_  | ~\new_[7998]_  | ~\new_[4621]_  | ~\new_[6163]_ ;
  assign \new_[12084]_  = ~\new_[1927]_ ;
  assign \new_[12085]_  = \new_[12086]_  & \new_[12087]_ ;
  assign \new_[12086]_  = ~\new_[4170]_ ;
  assign \new_[12087]_  = ~\new_[11268]_  | ~\new_[8504]_ ;
  assign \new_[12088]_  = ~\new_[1744]_ ;
  assign \new_[12089]_  = ~\new_[12177]_ ;
  assign \new_[12090]_  = ~\new_[12448]_ ;
  assign \new_[12091]_  = ~\new_[12440]_ ;
  assign \new_[12092]_  = ~\new_[6554]_  | ~\new_[5884]_ ;
  assign \new_[12093]_  = \new_[1523]_ ;
  assign \new_[12094]_  = ~\new_[12093]_ ;
  assign \new_[12095]_  = ~\new_[1523]_ ;
  assign \new_[12096]_  = ~\new_[12097]_  & ~\new_[12098]_ ;
  assign \new_[12097]_  = ~\new_[11105]_  | ~\new_[11086]_ ;
  assign \new_[12098]_  = \new_[12099]_ ;
  assign \new_[12099]_  = ~\new_[12100]_ ;
  assign \new_[12100]_  = ~\new_[12101]_ ;
  assign \new_[12101]_  = ~\new_[10344]_  | ~\new_[12586]_  | ~\new_[10004]_ ;
  assign \new_[12102]_  = ~\new_[4176]_  | ~\new_[12103]_  | ~\new_[3681]_ ;
  assign \new_[12103]_  = ~\new_[12104]_  & ~\new_[3405]_ ;
  assign \new_[12104]_  = ~\new_[12112]_  | ~\new_[12111]_  | ~\new_[12105]_  | ~\new_[6005]_ ;
  assign \new_[12105]_  = ~\new_[5498]_  & ~\new_[12106]_ ;
  assign \new_[12106]_  = ~\new_[12108]_  | ~\new_[12107]_  | ~\new_[7244]_ ;
  assign \new_[12107]_  = ~\new_[7058]_ ;
  assign \new_[12108]_  = ~\new_[11864]_  | ~\new_[12110]_ ;
  assign \new_[12109]_  = \new_[12381]_ ;
  assign \new_[12110]_  = ~\new_[12045]_  & ~\new_[10714]_ ;
  assign \new_[12111]_  = ~\new_[6656]_  | ~\new_[9594]_ ;
  assign \new_[12112]_  = (~\new_[11485]_  | ~\new_[8147]_ ) & (~\new_[7067]_  | ~\new_[12110]_ );
  assign \new_[12113]_  = ~\new_[12110]_ ;
  assign \new_[12114]_  = ~\new_[12120]_  | ~\new_[12119]_  | ~\new_[12115]_  | ~\new_[12118]_ ;
  assign \new_[12115]_  = ~\new_[12116]_  & (~\new_[12628]_  | ~\new_[8506]_ );
  assign \new_[12116]_  = ~\new_[12605]_  & ~\new_[12117]_ ;
  assign \new_[12117]_  = ~\new_[12093]_  | ~\new_[12635]_ ;
  assign \new_[12118]_  = ~\new_[1768]_ ;
  assign \new_[12119]_  = ~\new_[12092]_  & ~\new_[3005]_ ;
  assign \new_[12120]_  = ~\new_[2984]_ ;
  assign \new_[12121]_  = ~\new_[12127]_  | ~\new_[3271]_  | ~\new_[12122]_  | ~\new_[12126]_ ;
  assign \new_[12122]_  = ~\new_[12123]_  & ~\new_[1770]_ ;
  assign \new_[12123]_  = \new_[12124]_  | \new_[12125]_ ;
  assign \new_[12124]_  = ~\new_[6613]_  | ~\new_[7454]_  | ~\new_[5572]_  | ~\new_[5047]_ ;
  assign \new_[12125]_  = ~\new_[5889]_  | ~\new_[3595]_  | ~\new_[6559]_  | ~\new_[5058]_ ;
  assign \new_[12126]_  = ~\new_[12644]_  | ~\new_[10411]_  | ~\new_[12603]_ ;
  assign \new_[12127]_  = ~\new_[12628]_  | ~\new_[8510]_ ;
  assign \new_[12128]_  = ~\new_[12133]_  | ~\new_[12132]_  | ~\new_[12129]_  | ~\new_[3275]_ ;
  assign \new_[12129]_  = ~\new_[12130]_  & ~\new_[1775]_ ;
  assign \new_[12130]_  = ~\new_[6622]_  | ~\new_[5593]_  | ~\new_[12131]_  | ~\new_[3600]_ ;
  assign \new_[12131]_  = ~\new_[11267]_  | ~\new_[8513]_ ;
  assign \new_[12132]_  = ~\new_[12641]_  | ~\new_[10955]_  | ~\new_[12602]_ ;
  assign \new_[12133]_  = ~\new_[12134]_  & ~\new_[12135]_ ;
  assign \new_[12134]_  = ~\new_[6564]_  | ~\new_[5899]_ ;
  assign \new_[12135]_  = ~\new_[7468]_  | ~\new_[5076]_  | ~\new_[5450]_ ;
  assign \new_[12136]_  = ~\new_[12141]_  | ~\new_[12140]_  | ~\new_[12137]_  | ~\new_[3278]_ ;
  assign \new_[12137]_  = ~\new_[12138]_  & ~\new_[1777]_ ;
  assign \new_[12138]_  = ~\new_[6627]_  | ~\new_[5598]_  | ~\new_[12139]_  | ~\new_[3603]_ ;
  assign \new_[12139]_  = ~\new_[12420]_  | ~\new_[8518]_ ;
  assign \new_[12140]_  = ~\new_[12644]_  | ~\new_[11310]_  | ~\new_[12604]_ ;
  assign \new_[12141]_  = ~\new_[12142]_  & ~\new_[12143]_ ;
  assign \new_[12142]_  = ~\new_[6567]_  | ~\new_[5902]_ ;
  assign \new_[12143]_  = ~\new_[7472]_  | ~\new_[5080]_  | ~\new_[5491]_ ;
  assign \new_[12144]_  = ~\new_[12149]_  | ~\new_[12145]_  | ~\new_[12148]_ ;
  assign \new_[12145]_  = ~\new_[12146]_  & (~\new_[12628]_  | ~\new_[8505]_ );
  assign \new_[12146]_  = ~\new_[6601]_  | ~\new_[5564]_  | ~\new_[3269]_  | ~\new_[12147]_ ;
  assign \new_[12147]_  = \new_[4964]_  & \new_[7460]_ ;
  assign \new_[12148]_  = ~\new_[12639]_  | ~\new_[10802]_  | ~\new_[12603]_ ;
  assign \new_[12149]_  = ~\new_[12150]_  & ~\new_[1767]_ ;
  assign \new_[12150]_  = ~\new_[5883]_  | ~\new_[6553]_  | ~\new_[5052]_  | ~\new_[3590]_ ;
  assign \new_[12151]_  = \new_[12152]_  | \new_[12154]_ ;
  assign \new_[12152]_  = ~\new_[11150]_  | ~\new_[9261]_  | ~\new_[12153]_ ;
  assign \new_[12153]_  = \new_[11151]_  & \new_[11019]_ ;
  assign \new_[12154]_  = ~\new_[10079]_  | ~\new_[12155]_  | ~\new_[12038]_ ;
  assign \new_[12155]_  = ~\new_[12215]_ ;
  assign \new_[12156]_  = ~\new_[12154]_ ;
  assign \new_[12157]_  = \new_[9261]_  & \new_[11150]_ ;
  assign \new_[12158]_  = ~\new_[12164]_  | ~\new_[3281]_  | ~\new_[12159]_  | ~\new_[12163]_ ;
  assign \new_[12159]_  = ~\new_[12160]_  & ~\new_[1779]_ ;
  assign \new_[12160]_  = ~\new_[12161]_ ;
  assign \new_[12161]_  = ~\new_[12162]_  & (~\new_[11267]_  | ~\new_[8498]_ );
  assign \new_[12162]_  = ~\new_[6629]_  | ~\new_[5905]_  | ~\new_[6569]_  | ~\new_[5560]_ ;
  assign \new_[12163]_  = ~\new_[12639]_  | ~\new_[10933]_  | ~\new_[12603]_ ;
  assign \new_[12164]_  = ~\new_[12165]_ ;
  assign \new_[12165]_  = ~\new_[7449]_  | ~\new_[5495]_  | ~\new_[3605]_  | ~\new_[5082]_ ;
  assign \new_[12166]_  = \new_[12167]_  | \new_[8695]_ ;
  assign \new_[12167]_  = ~\new_[12168]_  | ~\new_[12096]_ ;
  assign \new_[12168]_  = \new_[12090]_  & \new_[12392]_ ;
  assign \new_[12169]_  = ~\new_[10839]_  | ~\new_[10468]_  | ~\new_[8019]_  | ~\new_[10658]_ ;
  assign \new_[12170]_  = ~\new_[11388]_  | ~\new_[12389]_  | ~\new_[9201]_ ;
  assign \new_[12171]_  = \new_[12167]_  | \new_[12172]_ ;
  assign \new_[12172]_  = ~\new_[12598]_  | ~\new_[12611]_  | ~\new_[9570]_  | ~\new_[9266]_ ;
  assign \new_[12173]_  = ~\new_[12168]_  | ~\new_[12096]_ ;
  assign \new_[12174]_  = ~\new_[12175]_  | ~\new_[12179]_  | ~\new_[12176]_ ;
  assign \new_[12175]_  = ~\new_[4327]_  & (~\new_[12747]_  | ~\new_[10045]_ );
  assign \new_[12176]_  = ~\new_[12089]_  | ~\new_[12628]_  | ~\new_[11777]_ ;
  assign \new_[12177]_  = \new_[12178]_ ;
  assign \new_[12178]_  = ~\new_[1522]_ ;
  assign \new_[12179]_  = ~\new_[12180]_  & (~\new_[12064]_  | ~\new_[10045]_ );
  assign \new_[12180]_  = ~\new_[12181]_ ;
  assign \new_[12181]_  = ~\new_[12089]_  | ~\new_[12647]_  | ~\new_[12606]_ ;
  assign \new_[12182]_  = ~\new_[8699]_  & ~\new_[12464]_ ;
  assign \new_[12183]_  = ~\new_[11355]_  | ~\new_[12695]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[12184]_  = \new_[12185]_ ;
  assign \new_[12185]_  = ~\new_[1484]_ ;
  assign \new_[12186]_  = ~\new_[12194]_  | ~\new_[12190]_  | ~\new_[12187]_  | ~\new_[12189]_ ;
  assign \new_[12187]_  = ~\new_[1753]_  & ~\new_[12188]_ ;
  assign \new_[12188]_  = ~\new_[3277]_ ;
  assign \new_[12189]_  = ~\new_[11356]_  | ~\new_[12635]_  | ~\new_[12603]_ ;
  assign \new_[12190]_  = ~\new_[12191]_  & ~\new_[12193]_ ;
  assign \new_[12191]_  = ~\new_[7309]_  | ~\new_[12192]_  | ~\new_[5596]_  | ~\new_[5489]_ ;
  assign \new_[12192]_  = \new_[7471]_  & \new_[6625]_ ;
  assign \new_[12193]_  = ~\new_[2693]_  | ~\new_[6342]_ ;
  assign \new_[12194]_  = ~\new_[12195]_  & (~\new_[11267]_  | ~\new_[8500]_ );
  assign \new_[12195]_  = ~\new_[3602]_  | ~\new_[5079]_ ;
  assign n1541 = ~\new_[12201]_  | (~\new_[12197]_  & ~\new_[12200]_ );
  assign \new_[12197]_  = ~\new_[12198]_  | ~\new_[12199]_ ;
  assign \new_[12198]_  = ~\new_[6948]_  | ~\new_[10576]_ ;
  assign \new_[12199]_  = ~\new_[2354]_  & ~\new_[10461]_ ;
  assign \new_[12200]_  = \new_[2627]_ ;
  assign \new_[12201]_  = ~\new_[7771]_  | ~\new_[10576]_ ;
  assign \new_[12202]_  = ~\new_[10461]_  & ~\new_[2627]_ ;
  assign n1556 = ~\new_[12208]_  | (~\new_[12204]_  & ~\new_[12207]_ );
  assign \new_[12204]_  = ~\new_[12205]_  | ~\new_[12206]_ ;
  assign \new_[12205]_  = ~\new_[6949]_  | ~\new_[10576]_ ;
  assign \new_[12206]_  = ~\new_[2357]_  & ~\new_[10461]_ ;
  assign \new_[12207]_  = \new_[2628]_ ;
  assign \new_[12208]_  = ~\new_[7773]_  | ~\new_[10576]_ ;
  assign \new_[12209]_  = ~\new_[10461]_  & ~\new_[2628]_ ;
  assign \new_[12210]_  = ~\new_[11530]_  | ~\new_[11921]_  | ~\new_[10965]_ ;
  assign \new_[12211]_  = ~\new_[12038]_  | ~\new_[12212]_  | ~\new_[11712]_ ;
  assign \new_[12212]_  = ~\new_[12213]_ ;
  assign \new_[12213]_  = \new_[12214]_ ;
  assign \new_[12214]_  = \new_[12215]_ ;
  assign \new_[12215]_  = ~\new_[12393]_  | ~\new_[8847]_  | ~\new_[12100]_ ;
  assign \new_[12216]_  = ~\new_[12212]_ ;
  assign \new_[12217]_  = ~\new_[12218]_  & ~\new_[12219]_ ;
  assign \new_[12218]_  = \new_[12590]_ ;
  assign \new_[12219]_  = \new_[11262]_  ? \new_[12622]_  : \new_[11090]_ ;
  assign \new_[12220]_  = ~\new_[12221]_  | ~\new_[12222]_ ;
  assign \new_[12221]_  = ~\new_[11436]_  | ~\new_[7696]_ ;
  assign \new_[12222]_  = ~\new_[11400]_  & (~\new_[11397]_  | ~\new_[11436]_ );
  assign \new_[12223]_  = \new_[11435]_  & \new_[8813]_ ;
  assign \new_[12224]_  = ~\new_[12225]_  | ~\new_[12228]_ ;
  assign \new_[12225]_  = ~\new_[12227]_  | ~\new_[12616]_  | ~\new_[12226]_ ;
  assign \new_[12226]_  = ~\new_[11443]_ ;
  assign \new_[12227]_  = ~\new_[11440]_  & ~\new_[11437]_ ;
  assign \new_[12228]_  = ~\new_[10420]_  | ~\new_[12229]_ ;
  assign \new_[12229]_  = ~\new_[1552]_ ;
  assign \new_[12230]_  = ~\new_[12236]_  | ~\new_[12235]_  | ~\new_[12231]_  | ~\new_[12234]_ ;
  assign \new_[12231]_  = ~\new_[12232]_  | ~\new_[12233]_ ;
  assign \new_[12232]_  = ~\new_[2072]_  | ~\new_[12512]_ ;
  assign \new_[12233]_  = \new_[11887]_  & \new_[11886]_ ;
  assign \new_[12234]_  = ~\new_[11934]_  | ~\new_[7859]_  | ~\new_[8797]_ ;
  assign \new_[12235]_  = ~\new_[10020]_  | ~\new_[12543]_  | ~\new_[7859]_  | ~\new_[8796]_ ;
  assign \new_[12236]_  = \new_[12237]_ ;
  assign \new_[12237]_  = \new_[8335]_  | \new_[8790]_  | \new_[12097]_  | \new_[9376]_ ;
  assign \new_[12238]_  = ~\new_[12235]_ ;
  assign \new_[12239]_  = ~\new_[12240]_ ;
  assign \new_[12240]_  = ~\new_[12233]_ ;
  assign n806 = ~\new_[1731]_  | ~\new_[12242]_  | ~\new_[12245]_  | ~\new_[12244]_ ;
  assign \new_[12242]_  = ~\new_[12243]_  & ~\new_[2695]_ ;
  assign \new_[12243]_  = ~\new_[6161]_  | ~\new_[1967]_  | ~\new_[2032]_ ;
  assign \new_[12244]_  = ~\new_[2787]_ ;
  assign \new_[12245]_  = \new_[12246]_  & \new_[12248]_ ;
  assign \new_[12246]_  = ~\new_[12247]_ ;
  assign \new_[12247]_  = ~\new_[4250]_  | ~\new_[3125]_  | ~\new_[3123]_ ;
  assign \new_[12248]_  = \new_[5919]_  & \new_[6126]_ ;
  assign n1046 = ~\new_[1916]_  | ~\new_[12257]_  | ~\new_[12250]_  | ~\new_[12252]_ ;
  assign \new_[12250]_  = ~\new_[1690]_  & ~\new_[12251]_ ;
  assign \new_[12251]_  = ~\new_[4592]_  | ~\new_[5931]_  | ~\new_[2849]_  | ~\new_[3268]_ ;
  assign \new_[12252]_  = \new_[12253]_  & \new_[1924]_ ;
  assign \new_[12253]_  = ~\new_[12254]_  & ~\new_[5370]_ ;
  assign \new_[12254]_  = ~\new_[12256]_  | ~\new_[4566]_  | ~\new_[12255]_  | ~\new_[5551]_ ;
  assign \new_[12255]_  = ~\new_[4677]_ ;
  assign \new_[12256]_  = ~\new_[11500]_  | ~\new_[10061]_ ;
  assign \new_[12257]_  = \new_[12258]_  & \new_[12259]_ ;
  assign \new_[12258]_  = ~\new_[2879]_ ;
  assign \new_[12259]_  = ~\new_[3116]_  | ~\new_[6985]_ ;
  assign n1051 = ~\new_[1917]_  | ~\new_[12268]_  | ~\new_[12261]_  | ~\new_[12263]_ ;
  assign \new_[12261]_  = ~\new_[1691]_  & ~\new_[12262]_ ;
  assign \new_[12262]_  = ~\new_[4598]_  | ~\new_[5579]_  | ~\new_[2855]_  | ~\new_[3272]_ ;
  assign \new_[12263]_  = \new_[12264]_  & \new_[1933]_ ;
  assign \new_[12264]_  = ~\new_[12265]_  & ~\new_[5372]_ ;
  assign \new_[12265]_  = ~\new_[12267]_  | ~\new_[4571]_  | ~\new_[12266]_  | ~\new_[5580]_ ;
  assign \new_[12266]_  = ~\new_[4701]_ ;
  assign \new_[12267]_  = ~\new_[11500]_  | ~\new_[9904]_ ;
  assign \new_[12268]_  = \new_[12269]_  & \new_[12270]_ ;
  assign \new_[12269]_  = ~\new_[2881]_ ;
  assign \new_[12270]_  = ~\new_[3119]_  | ~\new_[6985]_ ;
  assign \new_[12271]_  = ~\new_[5654]_ ;
  assign \new_[12272]_  = ~\new_[12273]_  | ~\new_[4926]_  | ~\new_[5242]_ ;
  assign \new_[12273]_  = ~\new_[12274]_ ;
  assign \new_[12274]_  = \new_[12275]_ ;
  assign \new_[12275]_  = ~\new_[1459]_ ;
  assign \new_[12276]_  = ~\new_[6112]_  & (~\new_[7577]_  | ~\new_[10265]_ );
  assign \new_[12277]_  = ~\new_[12273]_  | ~\new_[12695]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[12278]_  = ~\new_[12452]_ ;
  assign \new_[12279]_  = ~\new_[12567]_  | ~\new_[12695]_  | ~\new_[12661]_  | ~\new_[11292]_ ;
  assign \new_[12280]_  = \new_[12452]_ ;
  assign \new_[12281]_  = ~\new_[1645]_  & ~\new_[12282]_ ;
  assign \new_[12282]_  = ~\new_[12283]_ ;
  assign \new_[12283]_  = ~\new_[12284]_  | ~\new_[12285]_ ;
  assign \new_[12284]_  = \new_[12523]_  | \new_[9191]_ ;
  assign \new_[12285]_  = \new_[11000]_  & wb_cyc_i;
  assign \new_[12286]_  = ~\new_[12284]_ ;
  assign \new_[12287]_  = ~\new_[12288]_  | ~\new_[12290]_ ;
  assign \new_[12288]_  = ~\new_[5308]_  & ~\new_[12289]_ ;
  assign \new_[12289]_  = ~\new_[12738]_  & ~\new_[10256]_ ;
  assign \new_[12290]_  = ~\new_[12291]_  & ~\new_[12294]_ ;
  assign \new_[12291]_  = ~\new_[7524]_  | ~\new_[12292]_ ;
  assign \new_[12292]_  = ~\new_[12492]_  | ~\new_[12293]_ ;
  assign \new_[12293]_  = ~\new_[11575]_  & ~\new_[10417]_ ;
  assign \new_[12294]_  = ~\new_[12297]_  | ~\new_[12295]_  | ~\new_[12296]_ ;
  assign \new_[12295]_  = ~\new_[12750]_  | (~\new_[8830]_  & ~\new_[9822]_ );
  assign \new_[12296]_  = (~\new_[10128]_  | ~\new_[7077]_ ) & (~\new_[12792]_  | ~\new_[9651]_ );
  assign \new_[12297]_  = ~\new_[7873]_  | ~\new_[12293]_ ;
  assign \new_[12298]_  = ~\new_[12299]_  | ~\new_[12301]_ ;
  assign \new_[12299]_  = ~\new_[12300]_  & ~\new_[4810]_ ;
  assign \new_[12300]_  = ~\new_[9861]_  & ~\new_[12738]_ ;
  assign \new_[12301]_  = \new_[5622]_  & \new_[12302]_ ;
  assign \new_[12302]_  = ~\new_[12303]_  & (~\new_[7077]_  | ~\new_[9388]_ );
  assign \new_[12303]_  = ~\new_[12304]_  | ~\new_[12305]_ ;
  assign \new_[12304]_  = ~\new_[10657]_  | ~\new_[12792]_  | ~\new_[10743]_ ;
  assign \new_[12305]_  = (~\new_[12306]_  | ~\new_[12307]_ ) & (~\new_[11976]_  | ~\new_[12306]_ );
  assign \new_[12306]_  = ~\new_[10485]_  & ~\new_[4147]_ ;
  assign \new_[12307]_  = \new_[12308]_ ;
  assign \new_[12308]_  = ~\new_[12383]_ ;
  assign \new_[12309]_  = ~\new_[12310]_  | ~\new_[10531]_  | ~\new_[8637]_ ;
  assign \new_[12310]_  = ~\new_[12311]_  & ~\new_[12313]_ ;
  assign \new_[12311]_  = ~\new_[12555]_  | ~\new_[9991]_  | ~\new_[12312]_ ;
  assign \new_[12312]_  = \new_[10274]_  & \new_[10704]_ ;
  assign \new_[12313]_  = ~\new_[9804]_  | ~\new_[12317]_  | ~\new_[12314]_  | ~\new_[10786]_ ;
  assign \new_[12314]_  = ~\new_[12315]_ ;
  assign \new_[12315]_  = ~\new_[12316]_  | ~\new_[11493]_ ;
  assign \new_[12316]_  = \new_[10318]_  & \new_[12559]_ ;
  assign \new_[12317]_  = \new_[9992]_  & \new_[10469]_ ;
  assign \new_[12318]_  = \new_[9991]_  & \new_[12555]_ ;
  assign \new_[12319]_  = ~\new_[12317]_  | ~\new_[10531]_ ;
  assign \new_[12320]_  = ~\new_[11844]_  | ~\new_[11842]_ ;
  assign \new_[12321]_  = ~\new_[12596]_  | ~\new_[11756]_  | ~\new_[11754]_ ;
  assign \new_[12322]_  = ~\new_[12323]_  | ~\new_[12587]_ ;
  assign \new_[12323]_  = ~\new_[11843]_  & ~\new_[11896]_ ;
  assign \new_[12324]_  = ~\new_[11370]_  & ~\new_[11796]_ ;
  assign n916 = ~\new_[12326]_  | ~\new_[12329]_ ;
  assign \new_[12326]_  = ~\new_[12327]_  & ~\new_[12328]_ ;
  assign \new_[12327]_  = ~\new_[5608]_  | ~\new_[6150]_  | ~\new_[1947]_  | ~\new_[1990]_ ;
  assign \new_[12328]_  = ~\new_[5377]_  | ~\new_[3024]_  | ~\new_[11670]_  | ~\new_[2919]_ ;
  assign \new_[12329]_  = ~\new_[12330]_ ;
  assign \new_[12330]_  = ~\new_[12331]_  | ~\new_[2947]_  | ~\new_[1754]_ ;
  assign \new_[12331]_  = ~\new_[12332]_  & ~\new_[12333]_ ;
  assign \new_[12332]_  = ~\new_[4287]_  | ~\new_[5976]_ ;
  assign \new_[12333]_  = ~\new_[5612]_  | ~\new_[5613]_  | ~\new_[4887]_ ;
  assign \new_[12334]_  = ~\new_[12339]_  | (~\new_[12335]_  & ~\new_[12336]_ );
  assign \new_[12335]_  = ~\new_[4151]_  & ~\new_[2067]_ ;
  assign \new_[12336]_  = ~\new_[2241]_  | ~\new_[12337]_ ;
  assign \new_[12337]_  = ~\new_[12338]_ ;
  assign \new_[12338]_  = ~\new_[11889]_  | ~\new_[10783]_ ;
  assign \new_[12339]_  = ~\new_[12030]_  & ~\new_[12342]_ ;
  assign \new_[12340]_  = ~\new_[12341]_  & ~\new_[11555]_ ;
  assign \new_[12341]_  = \new_[11553]_  & \new_[12665]_ ;
  assign \new_[12342]_  = \new_[12343]_  ? \new_[2222]_  : \new_[12344]_ ;
  assign \new_[12343]_  = ~\new_[12337]_  & ~\new_[11738]_ ;
  assign \new_[12344]_  = \new_[11738]_  & \new_[12338]_ ;
  assign \new_[12345]_  = ~\new_[12346]_  & ~\new_[12350]_ ;
  assign \new_[12346]_  = ~\new_[2905]_  | ~\new_[12347]_ ;
  assign \new_[12347]_  = ~\new_[12348]_  & ~\new_[12349]_ ;
  assign \new_[12348]_  = ~\new_[12276]_  | ~\new_[12272]_  | ~\new_[12271]_ ;
  assign \new_[12349]_  = ~\new_[6571]_  | ~\new_[6166]_  | ~\new_[6269]_ ;
  assign \new_[12350]_  = ~\new_[12277]_  | ~\new_[12351]_  | ~\new_[3135]_ ;
  assign \new_[12351]_  = ~\new_[12352]_  & (~\new_[2021]_  | ~\new_[12603]_ );
  assign \new_[12352]_  = ~\new_[12354]_  | ~\new_[6160]_  | ~\new_[4582]_  | ~\new_[12353]_ ;
  assign \new_[12353]_  = ~\new_[12628]_  | ~\new_[8503]_ ;
  assign \new_[12354]_  = (~\new_[10265]_  | ~\new_[7065]_ ) & (~\new_[7226]_  | ~\new_[10039]_ );
  assign \new_[12355]_  = ~\new_[12356]_  & ~\new_[12359]_ ;
  assign \new_[12356]_  = ~\new_[3146]_  | ~\new_[12357]_  | ~\new_[3130]_ ;
  assign \new_[12357]_  = ~\new_[12358]_  & (~\new_[2023]_  | ~\new_[12606]_ );
  assign \new_[12358]_  = ~\new_[2044]_  | ~\new_[4596]_  | ~\new_[5563]_ ;
  assign \new_[12359]_  = ~\new_[1892]_  | ~\new_[12360]_ ;
  assign \new_[12360]_  = ~\new_[12361]_  & ~\new_[12365]_ ;
  assign \new_[12361]_  = ~\new_[8001]_  | ~\new_[12362]_  | ~\new_[3991]_  | ~\new_[5678]_ ;
  assign \new_[12362]_  = ~\new_[12363]_  & ~\new_[12364]_ ;
  assign \new_[12363]_  = (~\new_[11419]_  & ~\new_[9327]_ ) | (~\new_[12236]_  & ~\new_[9738]_ );
  assign \new_[12364]_  = ~\new_[9327]_  & ~\new_[6394]_ ;
  assign \new_[12365]_  = ~\new_[6273]_  | ~\new_[6188]_  | ~\new_[6599]_ ;
  assign \new_[12366]_  = ~\new_[12367]_  & ~\new_[12374]_ ;
  assign \new_[12367]_  = ~\new_[5552]_  | ~\new_[2043]_  | ~\new_[12368]_  | ~\new_[4593]_ ;
  assign \new_[12368]_  = ~\new_[12369]_  & ~\new_[12373]_ ;
  assign \new_[12369]_  = ~\new_[7871]_  | ~\new_[12370]_  | ~\new_[3986]_  | ~\new_[5672]_ ;
  assign \new_[12370]_  = ~\new_[12371]_  & ~\new_[12372]_ ;
  assign \new_[12371]_  = (~\new_[11419]_  & ~\new_[9303]_ ) | (~\new_[12236]_  & ~\new_[9941]_ );
  assign \new_[12372]_  = ~\new_[9303]_  & ~\new_[6394]_ ;
  assign \new_[12373]_  = ~\new_[6270]_  | ~\new_[6551]_  | ~\new_[6591]_ ;
  assign \new_[12374]_  = ~\new_[12375]_  | ~\new_[11734]_  | ~\new_[3129]_  | ~\new_[3143]_ ;
  assign \new_[12375]_  = ~\new_[2022]_  | ~\new_[12603]_ ;
  assign \new_[12376]_  = ~\new_[12377]_  | ~\new_[12381]_ ;
  assign \new_[12377]_  = ~\new_[12457]_  & ~\new_[12378]_ ;
  assign \new_[12378]_  = \new_[12379]_  | \new_[12380]_ ;
  assign \new_[12379]_  = ~\new_[12633]_  & ~\new_[8953]_ ;
  assign \new_[12380]_  = ~\new_[12210]_  & ~\new_[12211]_ ;
  assign \new_[12381]_  = ~\new_[10024]_  | ~\new_[8876]_  | ~\new_[12437]_  | ~\new_[8175]_ ;
  assign \new_[12382]_  = ~\new_[12457]_ ;
  assign \new_[12383]_  = ~\new_[12379]_ ;
  assign \new_[12384]_  = ~\new_[12385]_  | ~\new_[4147]_ ;
  assign \new_[12385]_  = ~\new_[12386]_ ;
  assign \new_[12386]_  = ~\new_[1507]_  | ~\new_[9734]_  | ~\new_[12389]_  | ~\new_[12387]_ ;
  assign \new_[12387]_  = \new_[12585]_  & \new_[10514]_ ;
  assign \new_[12388]_  = ~\new_[10165]_  | ~\new_[8945]_  | ~\new_[12632]_  | ~\new_[12394]_ ;
  assign \new_[12389]_  = ~\new_[11751]_  & ~\new_[12390]_  & ~\new_[12391]_ ;
  assign \new_[12390]_  = \new_[12448]_ ;
  assign \new_[12391]_  = ~\new_[12392]_ ;
  assign \new_[12392]_  = \new_[12393]_ ;
  assign \new_[12393]_  = ~\new_[9701]_  & ~\new_[9564]_ ;
  assign \new_[12394]_  = \new_[10253]_  & \new_[9913]_ ;
  assign \new_[12395]_  = ~\new_[12390]_  & ~\new_[11751]_ ;
  assign \new_[12396]_  = \new_[12642]_  & \new_[12397]_ ;
  assign \new_[12397]_  = (~\new_[10743]_  | ~\new_[12755]_ ) & (~\new_[12754]_  | ~\new_[10485]_ );
  assign \new_[12398]_  = \new_[12523]_ ;
  assign \new_[12399]_  = ~\new_[1538]_  & ~\new_[1488]_ ;
  assign \new_[12400]_  = ~\new_[1488]_ ;
  assign \new_[12401]_  = ~\new_[1538]_ ;
  assign \new_[12402]_  = ~\new_[12403]_ ;
  assign \new_[12403]_  = ~\new_[10818]_  | ~\new_[9059]_  | ~\new_[12153]_ ;
  assign n976 = ~\new_[12408]_  | ~\new_[2713]_  | ~\new_[12405]_ ;
  assign \new_[12405]_  = ~\new_[12406]_  & ~\new_[12407]_ ;
  assign \new_[12406]_  = ~\new_[5959]_  | ~\new_[3242]_  | ~\new_[3149]_ ;
  assign \new_[12407]_  = ~\new_[4127]_  | ~\new_[3011]_  | ~\new_[5734]_ ;
  assign \new_[12408]_  = ~\new_[12409]_  & ~\new_[1773]_ ;
  assign \new_[12409]_  = ~\new_[5896]_  | ~\new_[6561]_  | ~\new_[12410]_  | ~\new_[12411]_ ;
  assign \new_[12410]_  = ~\new_[12610]_  | ~\new_[12647]_  | ~\new_[12604]_ ;
  assign \new_[12411]_  = ~\new_[12420]_  | ~\new_[8512]_ ;
  assign \new_[12412]_  = ~\new_[12422]_  | ~\new_[12417]_  | ~\new_[12413]_  | ~\new_[12416]_ ;
  assign \new_[12413]_  = ~\new_[12415]_  & (~\new_[12414]_  | ~\new_[12636]_ );
  assign \new_[12414]_  = \new_[12606]_  & \new_[11361]_ ;
  assign \new_[12415]_  = ~\new_[5776]_  | ~\new_[5293]_ ;
  assign \new_[12416]_  = ~\new_[2988]_  & ~\new_[2991]_ ;
  assign \new_[12417]_  = ~\new_[12418]_ ;
  assign \new_[12418]_  = ~\new_[12419]_  | ~\new_[1907]_  | ~\new_[4014]_ ;
  assign \new_[12419]_  = ~\new_[11777]_  | ~\new_[12420]_  | ~\new_[11361]_ ;
  assign \new_[12420]_  = ~\new_[12421]_ ;
  assign \new_[12421]_  = ~\new_[2218]_  | ~\new_[2229]_ ;
  assign \new_[12422]_  = \new_[6195]_  & \new_[5904]_ ;
  assign \new_[12423]_  = ~\new_[2218]_  | ~\new_[2229]_ ;
  assign \new_[12424]_  = ~\new_[12465]_  | (~\new_[9170]_  & ~\new_[12425]_ );
  assign \new_[12425]_  = \new_[10507]_  | \new_[12469]_ ;
  assign \new_[12426]_  = ~\new_[10948]_  | ~\new_[12427]_  | ~\new_[11015]_ ;
  assign \new_[12427]_  = ~\new_[12428]_ ;
  assign \new_[12428]_  = ~wb_we_i | ~\new_[10135]_ ;
  assign \new_[12429]_  = ~\new_[10948]_  | ~\new_[12427]_  | ~\new_[11015]_ ;
  assign \new_[12430]_  = ~\new_[12432]_  | ~\new_[12431]_  | ~\new_[11897]_  | ~\new_[11901]_ ;
  assign \new_[12431]_  = ~\new_[7013]_  | ~\new_[10278]_ ;
  assign \new_[12432]_  = ~\new_[12433]_  & ~\new_[12435]_ ;
  assign \new_[12433]_  = ~\new_[12434]_  | (~\new_[7174]_  & ~\new_[7677]_ );
  assign \new_[12434]_  = ~\new_[12455]_  | ~\new_[2577]_ ;
  assign \new_[12435]_  = ~\new_[12436]_  | (~\new_[10522]_  & ~\new_[7865]_ );
  assign \new_[12436]_  = ~\new_[2577]_  | ~\new_[7298]_  | ~\new_[7686]_ ;
  assign \new_[12437]_  = ~\new_[12438]_ ;
  assign \new_[12438]_  = ~\new_[12444]_  | ~\new_[12439]_  | ~\new_[12441]_ ;
  assign \new_[12439]_  = ~\new_[12440]_ ;
  assign \new_[12440]_  = \new_[12097]_  | \new_[8335]_ ;
  assign \new_[12441]_  = \new_[12442]_ ;
  assign \new_[12442]_  = ~\new_[12443]_ ;
  assign \new_[12443]_  = ~\new_[11362]_  | ~\new_[11358]_ ;
  assign \new_[12444]_  = ~\new_[12445]_ ;
  assign \new_[12445]_  = ~\new_[11347]_  | ~\new_[10475]_ ;
  assign \new_[12446]_  = ~\new_[10772]_  & ~\new_[12666]_ ;
  assign \new_[12447]_  = \new_[12448]_ ;
  assign \new_[12448]_  = ~\new_[12034]_  | ~\new_[12031]_ ;
  assign \new_[12449]_  = ~\new_[10809]_  & ~\new_[10963]_ ;
  assign \new_[12450]_  = ~\new_[12453]_  | ~\new_[12695]_  | ~\new_[11840]_  | ~\new_[12451]_ ;
  assign \new_[12451]_  = ~\new_[12452]_ ;
  assign \new_[12452]_  = \new_[12552]_ ;
  assign \new_[12453]_  = ~\new_[12454]_ ;
  assign \new_[12454]_  = ~\new_[1507]_ ;
  assign \new_[12455]_  = \new_[12156]_  & \new_[12402]_ ;
  assign \new_[12456]_  = ~\new_[12464]_  & ~\new_[8700]_ ;
  assign \new_[12457]_  = ~\new_[12458]_  & ~\new_[12462]_ ;
  assign \new_[12458]_  = ~\new_[12461]_  | ~\new_[12459]_  | ~\new_[12460]_ ;
  assign \new_[12459]_  = \new_[11351]_  & \new_[10329]_ ;
  assign \new_[12460]_  = ~\new_[10250]_  & ~\new_[12730]_ ;
  assign \new_[12461]_  = ~\new_[10758]_  & ~\new_[12555]_ ;
  assign \new_[12462]_  = ~\new_[12168]_  | ~\new_[12096]_ ;
  assign \new_[12463]_  = ~\new_[12462]_ ;
  assign \new_[12464]_  = ~\new_[12168]_  | ~\new_[12096]_ ;
  assign \new_[12465]_  = ~\new_[12466]_  | ~\new_[12469]_ ;
  assign \new_[12466]_  = \new_[12467]_  | \new_[12468]_ ;
  assign \new_[12467]_  = ~\new_[8469]_  | ~\new_[8472]_ ;
  assign \new_[12468]_  = \new_[12590]_ ;
  assign \new_[12469]_  = ~\new_[10872]_  | ~\new_[10470]_  | ~\new_[10897]_ ;
  assign \new_[12470]_  = ~\new_[12476]_  | ~\new_[12737]_  | ~\new_[12471]_  | ~\new_[12474]_ ;
  assign \new_[12471]_  = ~\new_[12473]_  & ~\new_[12472]_ ;
  assign \new_[12472]_  = ~\new_[8174]_  & ~\new_[7368]_ ;
  assign \new_[12473]_  = ~\new_[7998]_  | ~\new_[8002]_ ;
  assign \new_[12474]_  = ~\new_[12475]_  & ~\new_[7573]_ ;
  assign \new_[12475]_  = ~\new_[11482]_  | ~\new_[12386]_ ;
  assign \new_[12476]_  = ~\new_[12182]_  & ~\new_[7420]_ ;
  assign \new_[12477]_  = ~\new_[12606]_  & ~\new_[12734]_ ;
  assign \new_[12478]_  = ~\new_[7998]_  | ~\new_[12386]_ ;
  assign \new_[12479]_  = ~\new_[8002]_  | ~\new_[12680]_ ;
  assign \new_[12480]_  = ~\new_[12481]_  | ~\new_[12484]_  | ~\new_[12483]_  | ~\new_[12482]_ ;
  assign \new_[12481]_  = ~\new_[12755]_  | ~\new_[11884]_  | ~\new_[5638]_ ;
  assign \new_[12482]_  = ~\new_[5691]_  & (~\new_[7226]_  | ~\new_[9391]_ );
  assign \new_[12483]_  = ~\new_[12064]_  | ~\new_[9970]_ ;
  assign \new_[12484]_  = ~\new_[12755]_  | ~\new_[12695]_  | ~\new_[12661]_  | ~\new_[12278]_ ;
  assign \new_[12485]_  = ~\new_[12233]_  | ~\new_[11814]_  | ~\new_[12722]_  | ~\new_[12549]_ ;
  assign \new_[12486]_  = ~\new_[12487]_  & ~\new_[12488]_ ;
  assign \new_[12487]_  = ~\new_[12166]_  | ~\new_[12171]_ ;
  assign \new_[12488]_  = ~\new_[12489]_  | ~\new_[12490]_ ;
  assign \new_[12489]_  = \new_[12169]_  & \new_[12170]_ ;
  assign \new_[12490]_  = ~\new_[12491]_  & ~\new_[12492]_ ;
  assign \new_[12491]_  = ~\new_[10122]_  & ~\new_[8150]_ ;
  assign \new_[12492]_  = ~\new_[12493]_ ;
  assign \new_[12493]_  = ~\new_[12494]_  | ~\new_[11992]_  | ~\new_[11819]_ ;
  assign \new_[12494]_  = \new_[9706]_  & \new_[12094]_ ;
  assign \new_[12495]_  = ~\new_[12490]_ ;
  assign \new_[12496]_  = \new_[12497]_  | \new_[12487]_ ;
  assign \new_[12497]_  = ~\new_[12498]_ ;
  assign \new_[12498]_  = \new_[12169]_  & \new_[12170]_ ;
  assign \new_[12499]_  = ~\new_[12500]_ ;
  assign \new_[12500]_  = (~\new_[2075]_  | ~\new_[11876]_ ) & (~\new_[12617]_  | ~\new_[2085]_ );
  assign \new_[12501]_  = ~\new_[11836]_  | ~\new_[11837]_  | ~\new_[11838]_ ;
  assign n2186 = ~\new_[12507]_  & (~\new_[12503]_  | ~\new_[12504]_ );
  assign \new_[12503]_  = \new_[4236]_  | n2936;
  assign \new_[12504]_  = ~\new_[12505]_  | ~\new_[12506]_ ;
  assign \new_[12505]_  = ~\new_[4340]_ ;
  assign \new_[12506]_  = ~\new_[11413]_  | ~\new_[11414]_ ;
  assign \new_[12507]_  = ~\new_[10481]_  | ~wb_cyc_i;
  assign \new_[12508]_  = ~\new_[12513]_  | ~\new_[12550]_  | ~\new_[12512]_ ;
  assign \new_[12509]_  = ~\new_[12510]_  | ~\new_[8143]_ ;
  assign \new_[12510]_  = ~\new_[7290]_ ;
  assign \new_[12511]_  = ~\new_[7290]_  | ~\new_[1711]_ ;
  assign \new_[12512]_  = ~\new_[11371]_  | ~\new_[10679]_ ;
  assign \new_[12513]_  = ~\new_[11507]_  & ~\new_[3036]_ ;
  assign \new_[12514]_  = ~\new_[12550]_ ;
  assign \new_[12515]_  = ~\new_[12509]_ ;
  assign \new_[12516]_  = ~\new_[12511]_ ;
  assign \new_[12517]_  = ~\new_[12518]_  & ~\new_[12519]_ ;
  assign \new_[12518]_  = ~n5446 | ~\new_[12426]_  | ~\new_[9939]_ ;
  assign \new_[12519]_  = ~\new_[12520]_ ;
  assign \new_[12520]_  = ~\new_[12552]_ ;
  assign n5041 = ~\new_[10270]_  | ~\new_[10098]_ ;
  assign \new_[12522]_  = ~\new_[12324]_  | ~\new_[12322]_  | ~\new_[12320]_  | ~\new_[12321]_ ;
  assign \new_[12523]_  = ~\new_[12518]_ ;
  assign \new_[12524]_  = ~\new_[12530]_  | ~\new_[12525]_  | ~\new_[12526]_ ;
  assign \new_[12525]_  = ~\new_[12453]_  | ~\new_[11277]_  | ~\new_[10441]_ ;
  assign \new_[12526]_  = \new_[12527]_  | \new_[12529]_ ;
  assign \new_[12527]_  = \new_[12528]_ ;
  assign \new_[12528]_  = ~\new_[12220]_  | ~\new_[12223]_ ;
  assign \new_[12529]_  = (~\new_[7509]_  | ~\new_[11306]_ ) & (~\new_[6767]_  | ~\new_[7825]_ );
  assign \new_[12530]_  = ~\new_[12453]_  | ~\new_[4758]_  | ~\new_[11233]_ ;
  assign \new_[12531]_  = ~\new_[12528]_ ;
  assign \new_[12532]_  = ~\new_[12528]_ ;
  assign \new_[12533]_  = ~\new_[12220]_  | ~\new_[12223]_ ;
  assign \new_[12534]_  = \new_[12535]_ ;
  assign \new_[12535]_  = ~\new_[12536]_  | ~\new_[12537]_ ;
  assign \new_[12536]_  = ~\new_[12455]_  & ~\new_[12456]_ ;
  assign \new_[12537]_  = ~\new_[12540]_  | ~\new_[12538]_  | ~\new_[12539]_ ;
  assign \new_[12538]_  = ~\new_[10503]_  & ~\new_[8477]_ ;
  assign \new_[12539]_  = ~\new_[11724]_ ;
  assign \new_[12540]_  = ~\new_[12541]_  & ~\new_[12391]_ ;
  assign \new_[12541]_  = ~\new_[12542]_  | ~\new_[12543]_ ;
  assign \new_[12542]_  = \new_[12731]_  & \new_[10211]_ ;
  assign \new_[12543]_  = \new_[12544]_ ;
  assign \new_[12544]_  = ~\new_[12545]_ ;
  assign \new_[12545]_  = ~\new_[10391]_  | ~\new_[10329]_ ;
  assign \new_[12546]_  = ~\new_[12554]_  | ~\new_[12553]_  | ~\new_[11840]_  | ~\new_[12278]_ ;
  assign \new_[12547]_  = ~\new_[12551]_  | ~\new_[12548]_  | ~\new_[12549]_ ;
  assign \new_[12548]_  = \new_[11841]_  & \new_[12233]_ ;
  assign \new_[12549]_  = \new_[12550]_ ;
  assign \new_[12550]_  = ~\new_[12509]_  | ~\new_[12511]_ ;
  assign \new_[12551]_  = ~\new_[11806]_  | ~\new_[12522]_  | ~\new_[11418]_ ;
  assign \new_[12552]_  = ~n5041 | ~\new_[12522]_ ;
  assign \new_[12553]_  = ~\new_[12523]_  | ~\new_[7908]_ ;
  assign \new_[12554]_  = \new_[1527]_ ;
  assign \new_[12555]_  = ~\new_[12554]_ ;
  assign \new_[12556]_  = ~\new_[1527]_ ;
  assign \new_[12557]_  = ~\new_[12561]_  & (~\new_[7277]_  | ~\new_[12558]_ );
  assign \new_[12558]_  = \new_[10023]_  & \new_[12559]_ ;
  assign \new_[12559]_  = \new_[12560]_  & \new_[11193]_ ;
  assign \new_[12560]_  = ~\new_[1525]_ ;
  assign \new_[12561]_  = (~\new_[7282]_  & ~\new_[12562]_ ) | (~\new_[7282]_  & ~\new_[12565]_ );
  assign \new_[12562]_  = (~\new_[12563]_  | ~\new_[11364]_ ) & (~\new_[11363]_  | ~\new_[12559]_ );
  assign \new_[12563]_  = \new_[10905]_  & \new_[12564]_ ;
  assign \new_[12564]_  = \new_[12560]_ ;
  assign \new_[12565]_  = \new_[12564]_  | \new_[10323]_ ;
  assign \new_[12566]_  = ~\new_[10323]_  & ~\new_[7282]_ ;
  assign \new_[12567]_  = ~\new_[12564]_ ;
  assign \new_[12568]_  = ~\new_[12574]_  | ~\new_[12571]_  | ~\new_[12569]_  | ~\new_[12570]_ ;
  assign \new_[12569]_  = ~\new_[7588]_  | ~\new_[10594]_ ;
  assign \new_[12570]_  = ~\new_[7572]_ ;
  assign \new_[12571]_  = ~\new_[12074]_  & ~\new_[12572]_ ;
  assign \new_[12572]_  = ~\new_[12573]_ ;
  assign \new_[12573]_  = ~\new_[10374]_  | ~\new_[12542]_  | ~\new_[7859]_  | ~\new_[12543]_ ;
  assign \new_[12574]_  = ~\new_[12788]_  | ~\new_[12577]_ ;
  assign \new_[12575]_  = ~\new_[8797]_  | ~\new_[7698]_  | ~\new_[12576]_ ;
  assign \new_[12576]_  = \new_[10060]_  & \new_[12459]_ ;
  assign \new_[12577]_  = ~\new_[4147]_ ;
  assign \new_[12578]_  = ~\new_[12074]_  & ~\new_[7572]_ ;
  assign \new_[12579]_  = ~\new_[12581]_  & (~\new_[12580]_  | ~\new_[12587]_ );
  assign \new_[12580]_  = ~\new_[11896]_  & ~\new_[11843]_ ;
  assign \new_[12581]_  = ~\new_[10811]_  | ~n1681;
  assign \new_[12582]_  = ~\new_[11844]_  | ~\new_[11842]_ ;
  assign \new_[12583]_  = ~\new_[12449]_  | ~\new_[8714]_  | ~\new_[12437]_  | ~\new_[12446]_ ;
  assign \new_[12584]_  = ~\new_[12449]_  | ~\new_[8714]_  | ~\new_[12437]_  | ~\new_[12446]_ ;
  assign \new_[12585]_  = ~\new_[10267]_  & ~\new_[12719]_ ;
  assign \new_[12586]_  = ~\new_[10267]_  & ~\new_[10233]_ ;
  assign \new_[12587]_  = ~\new_[11755]_  | ~\new_[12151]_ ;
  assign \new_[12588]_  = ~\new_[11755]_  | ~\new_[12151]_ ;
  assign \new_[12589]_  = \new_[11891]_  | \new_[8794]_ ;
  assign \new_[12590]_  = ~\new_[12726]_  | ~\new_[12579]_  | ~\new_[12582]_ ;
  assign \new_[12591]_  = ~\new_[12726]_  | ~\new_[12582]_  | ~\new_[12579]_ ;
  assign \new_[12592]_  = (~\new_[7689]_  & ~\new_[7990]_ ) | (~\new_[7283]_  & ~\new_[10190]_ );
  assign \new_[12593]_  = (~\new_[7689]_  & ~\new_[7990]_ ) | (~\new_[7283]_  & ~\new_[10190]_ );
  assign \new_[12594]_  = ~\new_[12733]_  | ~\new_[11352]_ ;
  assign \new_[12595]_  = ~\new_[11352]_  | ~\new_[12729]_ ;
  assign \new_[12596]_  = ~\new_[12587]_ ;
  assign \new_[12597]_  = ~\new_[12598]_ ;
  assign \new_[12598]_  = ~\new_[12599]_ ;
  assign \new_[12599]_  = \new_[12600]_ ;
  assign \new_[12600]_  = ~\new_[1544]_ ;
  assign \new_[12601]_  = \new_[7727]_ ;
  assign \new_[12602]_  = \new_[12606]_ ;
  assign \new_[12603]_  = ~\new_[12605]_ ;
  assign \new_[12604]_  = ~\new_[12605]_ ;
  assign \new_[12605]_  = ~\new_[12606]_ ;
  assign \new_[12606]_  = \new_[12182]_ ;
  assign \new_[12607]_  = ~\new_[12608]_ ;
  assign \new_[12608]_  = ~\new_[11792]_ ;
  assign \new_[12609]_  = ~\new_[12611]_ ;
  assign \new_[12610]_  = ~\new_[12611]_ ;
  assign \new_[12611]_  = \new_[12612]_ ;
  assign \new_[12612]_  = ~\new_[1528]_ ;
  assign \new_[12613]_  = \new_[12794]_  | \new_[12753]_ ;
  assign \new_[12614]_  = \new_[12794]_  | \new_[12751]_ ;
  assign \new_[12615]_  = ~\new_[12616]_ ;
  assign \new_[12616]_  = ~\new_[1865]_ ;
  assign \new_[12617]_  = ~\new_[12627]_ ;
  assign \new_[12618]_  = ~\new_[12619]_ ;
  assign \new_[12619]_  = \new_[12620]_ ;
  assign \new_[12620]_  = ~\new_[12621]_ ;
  assign \new_[12621]_  = ~\new_[12622]_ ;
  assign \new_[12622]_  = \new_[12623]_ ;
  assign \new_[12623]_  = ~\new_[12624]_ ;
  assign \new_[12624]_  = \new_[12627]_ ;
  assign \new_[12625]_  = ~\new_[12626]_ ;
  assign \new_[12626]_  = ~\new_[12627]_ ;
  assign \new_[12627]_  = ~\new_[12501]_ ;
  assign \new_[12628]_  = ~\new_[12631]_ ;
  assign \new_[12629]_  = \new_[12630]_ ;
  assign \new_[12630]_  = ~\new_[12631]_ ;
  assign \new_[12631]_  = \new_[12423]_ ;
  assign \new_[12632]_  = ~\new_[12633]_ ;
  assign \new_[12633]_  = ~\new_[12389]_ ;
  assign \new_[12634]_  = ~\new_[7532]_ ;
  assign \new_[12635]_  = ~\new_[12637]_ ;
  assign \new_[12636]_  = ~\new_[12637]_ ;
  assign \new_[12637]_  = ~\new_[12648]_ ;
  assign \new_[12638]_  = \new_[12640]_ ;
  assign \new_[12639]_  = \new_[12640]_ ;
  assign \new_[12640]_  = \new_[12648]_ ;
  assign \new_[12641]_  = \new_[12643]_ ;
  assign \new_[12642]_  = ~\new_[12643]_ ;
  assign \new_[12643]_  = \new_[12648]_ ;
  assign \new_[12644]_  = \new_[12647]_ ;
  assign \new_[12645]_  = \new_[12647]_ ;
  assign \new_[12646]_  = \new_[12647]_ ;
  assign \new_[12647]_  = \new_[12648]_ ;
  assign \new_[12648]_  = \new_[12517]_ ;
  assign \new_[12649]_  = \new_[7788]_ ;
  assign \new_[12650]_  = ~\new_[12658]_ ;
  assign \new_[12651]_  = ~\new_[12655]_ ;
  assign \new_[12652]_  = ~\new_[12655]_ ;
  assign \new_[12653]_  = ~\new_[12654]_ ;
  assign \new_[12654]_  = ~\new_[12655]_ ;
  assign \new_[12655]_  = \new_[12658]_ ;
  assign \new_[12656]_  = ~\new_[12657]_ ;
  assign \new_[12657]_  = \new_[12658]_ ;
  assign \new_[12658]_  = \new_[12380]_ ;
  assign \new_[12659]_  = \new_[12663]_ ;
  assign \new_[12660]_  = \new_[12663]_ ;
  assign \new_[12661]_  = ~\new_[12662]_ ;
  assign \new_[12662]_  = ~\new_[12663]_ ;
  assign \new_[12663]_  = ~\new_[12485]_ ;
  assign \new_[12664]_  = ~\new_[12665]_ ;
  assign \new_[12665]_  = \new_[11554]_ ;
  assign \new_[12666]_  = ~\new_[12667]_ ;
  assign \new_[12667]_  = \new_[12668]_ ;
  assign \new_[12668]_  = \new_[12669]_ ;
  assign \new_[12669]_  = ~\new_[10197]_ ;
  assign \new_[12670]_  = ~\new_[12671]_ ;
  assign \new_[12671]_  = ~\new_[11790]_ ;
  assign \new_[12672]_  = ~\new_[12673]_ ;
  assign \new_[12673]_  = ~\new_[12281]_ ;
  assign \new_[12674]_  = ~\new_[12675]_ ;
  assign \new_[12675]_  = \new_[12676]_ ;
  assign \new_[12676]_  = \new_[11826]_ ;
  assign \new_[12677]_  = ~\new_[12678]_ ;
  assign \new_[12678]_  = ~\new_[12686]_ ;
  assign \new_[12679]_  = ~\new_[12680]_ ;
  assign \new_[12680]_  = \new_[12686]_ ;
  assign \new_[12681]_  = ~\new_[12683]_ ;
  assign \new_[12682]_  = ~\new_[12683]_ ;
  assign \new_[12683]_  = ~\new_[12685]_ ;
  assign \new_[12684]_  = ~\new_[12685]_ ;
  assign \new_[12685]_  = ~\new_[12686]_ ;
  assign \new_[12686]_  = \new_[12687]_ ;
  assign \new_[12687]_  = \new_[11482]_ ;
  assign \new_[12688]_  = ~\new_[12689]_ ;
  assign \new_[12689]_  = ~\new_[12690]_ ;
  assign \new_[12690]_  = \new_[11498]_ ;
  assign \new_[12691]_  = ~\new_[12693]_ ;
  assign \new_[12692]_  = ~\new_[12693]_ ;
  assign \new_[12693]_  = \new_[12694]_ ;
  assign \new_[12694]_  = ~\new_[11498]_ ;
  assign \new_[12695]_  = \new_[12553]_ ;
  assign \new_[12696]_  = ~\new_[12697]_ ;
  assign \new_[12697]_  = \new_[7822]_ ;
  assign \new_[12698]_  = \new_[12699]_ ;
  assign \new_[12699]_  = ~\new_[12703]_ ;
  assign \new_[12700]_  = ~\new_[12703]_ ;
  assign \new_[12701]_  = ~\new_[12703]_ ;
  assign \new_[12702]_  = ~\new_[12700]_ ;
  assign \new_[12703]_  = ~\new_[11524]_ ;
  assign \new_[12704]_  = \new_[12705]_ ;
  assign \new_[12705]_  = ~\new_[12708]_ ;
  assign \new_[12706]_  = ~\new_[12708]_ ;
  assign \new_[12707]_  = ~\new_[12708]_ ;
  assign \new_[12708]_  = \new_[12718]_ ;
  assign \new_[12709]_  = ~\new_[12717]_ ;
  assign \new_[12710]_  = ~\new_[12717]_ ;
  assign \new_[12711]_  = ~\new_[12712]_ ;
  assign \new_[12712]_  = \new_[12717]_ ;
  assign \new_[12713]_  = ~\new_[12717]_ ;
  assign \new_[12714]_  = ~\new_[12715]_ ;
  assign \new_[12715]_  = \new_[12717]_ ;
  assign \new_[12716]_  = ~\new_[12717]_ ;
  assign \new_[12717]_  = \new_[12718]_ ;
  assign \new_[12718]_  = ~\new_[11524]_ ;
  assign \new_[12719]_  = \new_[10233]_ ;
  assign \new_[12720]_  = ~\new_[12721]_ ;
  assign \new_[12721]_  = \new_[12722]_ ;
  assign \new_[12722]_  = \new_[12551]_ ;
  assign \new_[12723]_  = ~\new_[12551]_ ;
  assign \new_[12724]_  = ~\new_[11828]_ ;
  assign \new_[12725]_  = ~\new_[12596]_  | ~\new_[11756]_  | ~\new_[11754]_ ;
  assign \new_[12726]_  = ~\new_[12596]_  | ~\new_[11756]_  | ~\new_[11754]_ ;
  assign \new_[12727]_  = \new_[11891]_  | \new_[8794]_ ;
  assign \new_[12728]_  = \new_[11891]_  | \new_[8794]_ ;
  assign \new_[12729]_  = ~\new_[10247]_ ;
  assign \new_[12730]_  = ~\new_[12731]_ ;
  assign \new_[12731]_  = \new_[12733]_ ;
  assign \new_[12732]_  = ~\new_[12733]_ ;
  assign \new_[12733]_  = ~\new_[10247]_ ;
  assign \new_[12734]_  = ~\new_[12737]_ ;
  assign \new_[12735]_  = ~\new_[12736]_ ;
  assign \new_[12736]_  = \new_[12737]_ ;
  assign \new_[12737]_  = ~\new_[7589]_ ;
  assign \new_[12738]_  = ~\new_[12739]_ ;
  assign \new_[12739]_  = ~\new_[12740]_ ;
  assign \new_[12740]_  = \new_[12589]_ ;
  assign \new_[12741]_  = \new_[12746]_ ;
  assign \new_[12742]_  = ~\new_[12744]_ ;
  assign \new_[12743]_  = ~\new_[12744]_ ;
  assign \new_[12744]_  = ~\new_[12746]_ ;
  assign \new_[12745]_  = \new_[12746]_ ;
  assign \new_[12746]_  = \new_[12589]_ ;
  assign \new_[12747]_  = ~\new_[12752]_ ;
  assign \new_[12748]_  = ~\new_[12752]_ ;
  assign \new_[12749]_  = \new_[12751]_ ;
  assign \new_[12750]_  = \new_[12751]_ ;
  assign \new_[12751]_  = ~\new_[12752]_ ;
  assign \new_[12752]_  = \new_[12583]_ ;
  assign \new_[12753]_  = ~\new_[12583]_ ;
  assign \new_[12754]_  = ~\new_[12755]_ ;
  assign \new_[12755]_  = \new_[12756]_ ;
  assign \new_[12756]_  = ~\new_[12757]_ ;
  assign \new_[12757]_  = \new_[12758]_ ;
  assign \new_[12758]_  = ~\new_[1561]_ ;
  assign \new_[12759]_  = ~\new_[12760]_ ;
  assign \new_[12760]_  = \new_[2431]_ ;
  assign \new_[12761]_  = ~\new_[12762]_ ;
  assign \new_[12762]_  = \new_[2430]_ ;
  assign \new_[12763]_  = ~\new_[12764]_ ;
  assign \new_[12764]_  = ~\new_[12767]_ ;
  assign \new_[12765]_  = ~\new_[12766]_ ;
  assign \new_[12766]_  = \new_[12767]_ ;
  assign \new_[12767]_  = ~\new_[11708]_ ;
  assign \new_[12768]_  = \new_[12779]_ ;
  assign \new_[12769]_  = ~\new_[12772]_ ;
  assign \new_[12770]_  = ~\new_[12772]_ ;
  assign \new_[12771]_  = ~\new_[12772]_ ;
  assign \new_[12772]_  = ~\new_[12779]_ ;
  assign \new_[12773]_  = \new_[12779]_ ;
  assign \new_[12774]_  = \new_[12779]_ ;
  assign \new_[12775]_  = ~\new_[12778]_ ;
  assign \new_[12776]_  = ~\new_[12778]_ ;
  assign \new_[12777]_  = ~\new_[12778]_ ;
  assign \new_[12778]_  = ~\new_[12779]_ ;
  assign \new_[12779]_  = \new_[7173]_ ;
  assign \new_[12780]_  = ~\new_[12781]_ ;
  assign \new_[12781]_  = \new_[11999]_ ;
  assign \new_[12782]_  = ~\new_[12788]_ ;
  assign \new_[12783]_  = \new_[12786]_ ;
  assign \new_[12784]_  = ~\new_[12785]_ ;
  assign \new_[12785]_  = ~\new_[12786]_ ;
  assign \new_[12786]_  = \new_[12787]_ ;
  assign \new_[12787]_  = \new_[12788]_ ;
  assign \new_[12788]_  = ~\new_[12575]_ ;
  assign \new_[12789]_  = \new_[12792]_ ;
  assign \new_[12790]_  = ~\new_[12791]_ ;
  assign \new_[12791]_  = ~\new_[12792]_ ;
  assign \new_[12792]_  = \new_[12794]_ ;
  assign \new_[12793]_  = \new_[12794]_ ;
  assign \new_[12794]_  = \new_[11878]_ ;
  assign suspended_o = n4706;
  assign mc_cke_pad_o_ = n5881;
  assign n1146 = n1151;
  assign n5296 = \wb_addr_i[2] ;
  assign n5301 = \wb_addr_i[2] ;
  assign n5316 = \wb_addr_i[2] ;
  assign n5376 = \wb_addr_i[3] ;
  assign n5401 = \wb_addr_i[3] ;
  assign n5436 = \wb_addr_i[3] ;
  assign n5501 = resume_req_i;
  assign n5511 = susp_req_i;
  assign n5526 = new_u5_rsts1_reg_in_;
  assign n5541 = new_u5_rsts1_reg_in_;
  assign n5576 = new_u5_rsts1_reg_in_;
  assign n5681 = \mc_data_pad_i[23] ;
  assign n5686 = \mc_data_pad_i[8] ;
  assign n5691 = \mc_data_pad_i[6] ;
  assign n5696 = \wb_addr_i[6] ;
  assign n5701 = \mc_data_pad_i[13] ;
  assign n5706 = \mc_data_pad_i[14] ;
  assign n5716 = \mc_dp_pad_i[3] ;
  assign n5721 = \mc_data_pad_i[21] ;
  assign n5726 = \mc_data_pad_i[7] ;
  assign n5731 = \mc_data_pad_i[28] ;
  assign n5736 = \wb_addr_i[5] ;
  assign n5741 = \mc_data_pad_i[22] ;
  assign n5746 = \mc_data_pad_i[1] ;
  assign n5751 = \mc_data_pad_i[0] ;
  assign n5756 = mc_ack_pad_i;
  assign n5761 = \mc_data_pad_i[19] ;
  assign n5771 = \mc_data_pad_i[5] ;
  assign n5776 = \wb_addr_i[4] ;
  assign n5781 = \mc_data_pad_i[17] ;
  assign n5791 = \mc_data_pad_i[29] ;
  assign n5796 = \mc_data_pad_i[18] ;
  assign n5801 = \mc_data_pad_i[4] ;
  assign n5806 = \wb_addr_i[5] ;
  assign n5811 = \wb_addr_i[4] ;
  assign n5816 = \mc_data_pad_i[11] ;
  assign n5821 = \mc_data_pad_i[27] ;
  assign n5826 = mc_sts_pad_i;
  assign n5831 = \mc_data_pad_i[10] ;
  assign n5836 = \wb_addr_i[5] ;
  assign n5841 = \mc_data_pad_i[15] ;
  assign n5846 = \mc_dp_pad_i[2] ;
  assign n5851 = \mc_data_pad_i[12] ;
  assign n5856 = \mc_data_pad_i[9] ;
  assign n5861 = \mc_dp_pad_i[1] ;
  assign n5866 = \mc_data_pad_i[3] ;
  assign n5876 = \mc_data_pad_i[25] ;
  assign n5886 = \mc_data_pad_i[31] ;
  assign n5896 = \mc_data_pad_i[26] ;
  assign n5901 = \mc_data_pad_i[24] ;
  assign n5906 = \mc_data_pad_i[16] ;
  assign n5911 = \mc_data_pad_i[30] ;
  assign n5916 = mc_br_pad_i;
  assign n5921 = \wb_addr_i[6] ;
  assign n5926 = \mc_data_pad_i[2] ;
  assign n5931 = \wb_addr_i[4] ;
  assign n5936 = \mc_dp_pad_i[0] ;
  assign n5941 = \mc_data_pad_i[20] ;
  assign n5946 = \wb_addr_i[6] ;
  assign n5651 = 1'b0;
  always @ (posedge clock) begin
    \\u7_mc_addr_reg[10]  <= n536;
    \\u7_mc_addr_reg[12]  <= n541;
    \\u7_mc_addr_reg[11]  <= n546;
    \\u7_mc_addr_reg[9]  <= n551;
    \\u7_mc_addr_reg[8]  <= n556;
    \\u7_mc_addr_reg[7]  <= n561;
    \\u7_mc_addr_reg[6]  <= n566;
    \\u7_mc_addr_reg[5]  <= n571;
    \\u7_mc_addr_reg[4]  <= n576;
    \\u7_mc_addr_reg[3]  <= n581;
    \\u7_mc_addr_reg[2]  <= n586;
    \\u7_mc_addr_reg[1]  <= n591;
    \\u7_mc_addr_reg[0]  <= n596;
    u7_mc_we__reg <= n601;
    \\u7_mc_cs__reg[1]  <= n606;
    \\u7_mc_cs__reg[0]  <= n611;
    \\u7_mc_cs__reg[7]  <= n616;
    \\u7_mc_cs__reg[6]  <= n621;
    \\u7_mc_cs__reg[5]  <= n626;
    \\u7_mc_cs__reg[4]  <= n631;
    \\u7_mc_cs__reg[3]  <= n636;
    \\u7_mc_cs__reg[2]  <= n641;
    \\u5_cmd_del_reg[0]  <= n646;
    \\u5_cmd_r_reg[0]  <= n651;
    u5_cmd_asserted_reg <= n656;
    u7_mc_cas__reg <= n661;
    \\u7_mc_dqm_reg[2]  <= n666;
    \\u7_mc_dqm_reg[1]  <= n671;
    \\u7_mc_dqm_reg[0]  <= n676;
    \\u7_mc_dqm_reg[3]  <= n681;
    \\u5_cmd_del_reg[3]  <= n686;
    u6_wb_ack_o_reg <= n691;
    \\u5_state_reg[16]  <= n696;
    \\u5_timer_reg[0]  <= n701;
    \\u5_timer_reg[1]  <= n706;
    \\u5_state_reg[2]  <= n711;
    \\u5_state_reg[59]  <= n716;
    \\u5_cmd_r_reg[3]  <= n721;
    \\u5_state_reg[17]  <= n726;
    \\u5_state_reg[1]  <= n731;
    \\u5_state_reg[35]  <= n736;
    \\u5_burst_cnt_reg[2]  <= n741;
    \\u5_burst_cnt_reg[8]  <= n746;
    \\u5_burst_cnt_reg[9]  <= n751;
    \\u5_burst_cnt_reg[0]  <= n756;
    \\u5_state_reg[21]  <= n761;
    \\u5_state_reg[29]  <= n766;
    \\u5_state_reg[57]  <= n771;
    \\u5_state_reg[0]  <= n776;
    \\u5_state_reg[10]  <= n781;
    \\u5_state_reg[15]  <= n786;
    \\u5_state_reg[40]  <= n791;
    \\u5_burst_cnt_reg[10]  <= n796;
    \\u5_state_reg[18]  <= n801;
    \\u5_state_reg[20]  <= n806;
    \\u5_state_reg[22]  <= n811;
    \\u5_state_reg[23]  <= n816;
    \\u5_state_reg[24]  <= n821;
    \\u5_state_reg[62]  <= n826;
    \\u5_state_reg[26]  <= n831;
    \\u5_state_reg[27]  <= n836;
    \\u5_state_reg[28]  <= n841;
    \\u5_state_reg[25]  <= n846;
    \\u5_state_reg[30]  <= n851;
    \\u5_state_reg[32]  <= n856;
    \\u5_state_reg[33]  <= n861;
    \\u5_state_reg[38]  <= n866;
    \\u5_state_reg[43]  <= n871;
    \\u5_state_reg[36]  <= n876;
    \\u5_state_reg[46]  <= n881;
    \\u5_state_reg[4]  <= n886;
    \\u5_state_reg[45]  <= n891;
    \\u5_state_reg[52]  <= n896;
    \\u5_state_reg[60]  <= n901;
    \\u5_state_reg[9]  <= n906;
    \\u5_state_reg[13]  <= n911;
    \\u5_state_reg[12]  <= n916;
    \\u5_state_reg[48]  <= n921;
    u7_mc_data_oe_reg <= n926;
    \\u5_timer_reg[2]  <= n931;
    u6_wb_err_reg <= n936;
    \\u5_state_reg[37]  <= n941;
    \\u5_state_reg[39]  <= n946;
    \\u5_state_reg[42]  <= n951;
    \\u5_state_reg[41]  <= n956;
    \\u5_state_reg[44]  <= n961;
    \\u5_state_reg[47]  <= n966;
    \\u5_state_reg[51]  <= n971;
    \\u5_state_reg[56]  <= n976;
    \\u5_state_reg[5]  <= n981;
    \\u5_state_reg[61]  <= n986;
    \\u5_state_reg[58]  <= n991;
    \\u5_state_reg[63]  <= n996;
    \\u5_state_reg[64]  <= n1001;
    \\u5_state_reg[11]  <= n1006;
    \\u5_state_reg[6]  <= n1011;
    \\u5_state_reg[7]  <= n1016;
    \\u5_state_reg[8]  <= n1021;
    \\u5_state_reg[65]  <= n1026;
    \\u5_burst_cnt_reg[3]  <= n1031;
    \\u5_state_reg[14]  <= n1036;
    \\u5_burst_cnt_reg[1]  <= n1041;
    \\u5_state_reg[34]  <= n1046;
    \\u5_state_reg[50]  <= n1051;
    \\u5_state_reg[55]  <= n1056;
    \\u5_cmd_del_reg[1]  <= n1061;
    \\u5_state_reg[19]  <= n1066;
    \\u5_state_reg[31]  <= n1071;
    \\u5_state_reg[3]  <= n1076;
    \\u5_state_reg[49]  <= n1081;
    \\u5_state_reg[54]  <= n1086;
    \\u5_state_reg[53]  <= n1091;
    u7_mc_oe__reg <= n1096;
    \\u5_burst_cnt_reg[4]  <= n1101;
    \\u5_burst_cnt_reg[7]  <= n1106;
    \\u5_burst_cnt_reg[6]  <= n1111;
    \\u5_burst_cnt_reg[5]  <= n1116;
    \\u5_cmd_r_reg[1]  <= n1121;
    \\u5_timer_reg[3]  <= n1126;
    u5_data_oe_reg <= n1131;
    u5_wb_stb_first_reg <= n1136;
    \\u5_timer2_reg[2]  <= n1141;
    u5_mem_ack_r_reg <= n1146;
    mem_ack_r_reg <= n1151;
    u5_oe__reg <= n1156;
    \\u5_timer2_reg[1]  <= n1161;
    \\u5_timer2_reg[3]  <= n1166;
    u5_cke__reg <= n1171;
    u5_data_oe_r2_reg <= n1176;
    u5_cke_r_reg <= n1181;
    \\u5_timer2_reg[5]  <= n1186;
    u5_data_oe_r_reg <= n1191;
    \\u5_timer2_reg[4]  <= n1196;
    \\u5_timer2_reg[0]  <= n1201;
    \\u5_timer2_reg[8]  <= n1206;
    \\u5_timer2_reg[7]  <= n1211;
    \\u5_timer2_reg[6]  <= n1216;
    u5_ap_en_reg <= n1221;
    \\u5_timer_reg[5]  <= n1226;
    \\u5_timer_reg[4]  <= n1231;
    \\u0_tms_reg[21]  <= n1236;
    \\u0_tms_reg[5]  <= n1241;
    \\u0_tms_reg[9]  <= n1246;
    \\u0_tms_reg[27]  <= n1251;
    \\u0_tms_reg[1]  <= n1256;
    \\u0_tms_reg[16]  <= n1261;
    \\u0_sp_tms_reg[9]  <= n1266;
    \\u0_sp_tms_reg[26]  <= n1271;
    \\u0_sp_tms_reg[5]  <= n1276;
    \\u0_sp_tms_reg[20]  <= n1281;
    \\u0_sp_tms_reg[23]  <= n1286;
    \\u0_sp_tms_reg[11]  <= n1291;
    \\u0_sp_tms_reg[0]  <= n1296;
    \\u0_sp_tms_reg[10]  <= n1301;
    \\u0_sp_tms_reg[12]  <= n1306;
    \\u0_sp_tms_reg[13]  <= n1311;
    \\u0_sp_tms_reg[14]  <= n1316;
    \\u0_sp_tms_reg[15]  <= n1321;
    \\u0_sp_tms_reg[17]  <= n1326;
    \\u0_sp_tms_reg[18]  <= n1331;
    \\u0_sp_tms_reg[19]  <= n1336;
    \\u0_sp_tms_reg[1]  <= n1341;
    \\u0_sp_tms_reg[21]  <= n1346;
    \\u0_sp_tms_reg[22]  <= n1351;
    \\u0_sp_tms_reg[24]  <= n1356;
    \\u0_sp_tms_reg[27]  <= n1361;
    \\u0_sp_tms_reg[2]  <= n1366;
    \\u0_sp_tms_reg[25]  <= n1371;
    \\u0_sp_tms_reg[3]  <= n1376;
    \\u0_sp_tms_reg[4]  <= n1381;
    \\u0_sp_tms_reg[6]  <= n1386;
    \\u0_sp_tms_reg[7]  <= n1391;
    \\u0_sp_tms_reg[8]  <= n1396;
    \\u0_tms_reg[11]  <= n1401;
    \\u0_tms_reg[0]  <= n1406;
    \\u0_tms_reg[10]  <= n1411;
    \\u0_tms_reg[12]  <= n1416;
    \\u0_tms_reg[13]  <= n1421;
    \\u0_tms_reg[15]  <= n1426;
    \\u0_tms_reg[14]  <= n1431;
    \\u0_tms_reg[17]  <= n1436;
    \\u0_tms_reg[18]  <= n1441;
    \\u0_tms_reg[19]  <= n1446;
    \\u0_tms_reg[20]  <= n1451;
    \\u0_tms_reg[22]  <= n1456;
    \\u0_tms_reg[23]  <= n1461;
    \\u0_tms_reg[24]  <= n1466;
    \\u0_tms_reg[26]  <= n1471;
    \\u0_tms_reg[25]  <= n1476;
    \\u0_tms_reg[2]  <= n1481;
    \\u0_tms_reg[3]  <= n1486;
    \\u0_tms_reg[4]  <= n1491;
    \\u0_tms_reg[7]  <= n1496;
    \\u0_tms_reg[8]  <= n1501;
    \\u0_tms_reg[6]  <= n1506;
    \\u5_timer_reg[7]  <= n1511;
    \\u5_timer_reg[6]  <= n1516;
    \\u0_sp_tms_reg[16]  <= n1521;
    \\u0_csc_reg[10]  <= n1526;
    \\u0_csc_reg[5]  <= n1531;
    \\u0_csc_reg[4]  <= n1536;
    u2_u0_bank0_open_reg <= n1541;
    u2_u0_bank1_open_reg <= n1546;
    u2_u0_bank3_open_reg <= n1551;
    u2_u1_bank0_open_reg <= n1556;
    u2_u1_bank1_open_reg <= n1561;
    u2_u1_bank2_open_reg <= n1566;
    \\u0_csc_reg[6]  <= n1571;
    \\u0_csc_reg[7]  <= n1576;
    \\u0_csc_reg[9]  <= n1581;
    \\u0_sp_csc_reg[10]  <= n1586;
    \\u0_sp_csc_reg[4]  <= n1591;
    \\u0_sp_csc_reg[7]  <= n1596;
    \\u0_sp_csc_reg[9]  <= n1601;
    \\u0_sp_csc_reg[6]  <= n1606;
    \\u0_sp_csc_reg[3]  <= n1611;
    \\u0_sp_csc_reg[2]  <= n1616;
    \\u0_csc_reg[11]  <= n1621;
    u2_u1_bank3_open_reg <= n1626;
    \\u0_sp_csc_reg[5]  <= n1631;
    u2_u0_bank2_open_reg <= n1636;
    \\u0_sp_csc_reg[1]  <= n1641;
    \\u0_csc_reg[1]  <= n1646;
    \\u0_csc_reg[3]  <= n1651;
    \\u0_csc_reg[2]  <= n1656;
    u5_cmd_a10_r_reg <= n1661;
    u7_mc_ras__reg <= n1666;
    u7_mc_adsc__reg <= n1671;
    u5_wr_cycle_reg <= n1676;
    u7_mc_c_oe_reg <= n1681;
    u5_cs_le_reg <= n1686;
    \\u5_cmd_del_reg[2]  <= n1691;
    u5_mc_c_oe_reg <= n1696;
    \\u1_bank_adr_reg[0]  <= n1701;
    \\u1_row_adr_reg[10]  <= n1706;
    \\u1_row_adr_reg[11]  <= n1711;
    \\u5_cmd_r_reg[2]  <= n1716;
    \\u1_bank_adr_reg[1]  <= n1721;
    \\u1_row_adr_reg[9]  <= n1726;
    \\u1_row_adr_reg[12]  <= n1731;
    \\u1_row_adr_reg[3]  <= n1736;
    \\u1_row_adr_reg[7]  <= n1741;
    \\u1_row_adr_reg[0]  <= n1746;
    \\u1_acs_addr_reg[23]  <= n1751;
    \\u1_row_adr_reg[1]  <= n1756;
    \\u1_row_adr_reg[2]  <= n1761;
    \\u1_row_adr_reg[4]  <= n1766;
    \\u1_row_adr_reg[5]  <= n1771;
    \\u1_row_adr_reg[6]  <= n1776;
    \\u1_row_adr_reg[8]  <= n1781;
    u5_cnt_reg <= n1786;
    \\u3_byte1_reg[5]  <= n1791;
    u5_wb_cycle_reg <= n1796;
    \\u1_acs_addr_reg[19]  <= n1801;
    \\u1_acs_addr_reg[20]  <= n1806;
    \\u3_byte1_reg[0]  <= n1811;
    \\u3_byte1_reg[1]  <= n1816;
    \\u3_byte1_reg[2]  <= n1821;
    \\u3_byte1_reg[3]  <= n1826;
    \\u3_byte1_reg[4]  <= n1831;
    \\u3_byte1_reg[7]  <= n1836;
    \\u3_byte1_reg[6]  <= n1841;
    \\u1_col_adr_reg[8]  <= n1846;
    \\u1_acs_addr_reg[22]  <= n1851;
    \\u1_acs_addr_reg[9]  <= n1856;
    \\u1_acs_addr_reg[10]  <= n1861;
    \\u1_acs_addr_reg[2]  <= n1866;
    \\u1_acs_addr_reg[21]  <= n1871;
    \\u1_acs_addr_reg[18]  <= n1876;
    \\u1_acs_addr_reg[4]  <= n1881;
    \\u1_acs_addr_reg[7]  <= n1886;
    \\u1_acs_addr_reg[13]  <= n1891;
    \\u1_acs_addr_reg[16]  <= n1896;
    \\u1_acs_addr_reg[14]  <= n1901;
    \\u1_acs_addr_reg[11]  <= n1906;
    \\u1_acs_addr_reg[17]  <= n1911;
    \\u1_acs_addr_reg[12]  <= n1916;
    \\u1_acs_addr_reg[8]  <= n1921;
    \\u1_acs_addr_reg[0]  <= n1926;
    \\u1_acs_addr_reg[1]  <= n1931;
    \\u1_acs_addr_reg[3]  <= n1936;
    \\u1_acs_addr_reg[5]  <= n1941;
    \\u1_acs_addr_reg[6]  <= n1946;
    \\u1_acs_addr_reg[15]  <= n1951;
    \\u1_col_adr_reg[9]  <= n1956;
    \\u5_ack_cnt_reg[3]  <= n1961;
    \\u5_ack_cnt_reg[1]  <= n1966;
    u4_rfr_req_reg <= n1971;
    \\u5_ack_cnt_reg[0]  <= n1976;
    \\u5_ack_cnt_reg[2]  <= n1981;
    \\u3_byte0_reg[1]  <= n1986;
    \\u3_byte0_reg[0]  <= n1991;
    \\u3_byte0_reg[2]  <= n1996;
    \\u3_byte0_reg[4]  <= n2001;
    \\u3_byte0_reg[3]  <= n2006;
    \\u3_byte0_reg[5]  <= n2011;
    \\u3_byte0_reg[6]  <= n2016;
    \\u3_byte0_reg[7]  <= n2021;
    \\u3_byte2_reg[7]  <= n2026;
    u5_lmr_ack_reg <= n2031;
    \\u5_ir_cnt_reg[1]  <= n2036;
    \\u5_ir_cnt_reg[2]  <= n2041;
    \\u7_mc_addr_reg[14]  <= n2046;
    \\u3_byte2_reg[0]  <= n2051;
    \\u3_byte2_reg[1]  <= n2056;
    \\u3_byte2_reg[2]  <= n2061;
    \\u3_byte2_reg[4]  <= n2066;
    \\u3_byte2_reg[5]  <= n2071;
    \\u3_byte2_reg[6]  <= n2076;
    \\u3_byte2_reg[3]  <= n2081;
    \\u7_mc_addr_reg[13]  <= n2086;
    \\u5_ir_cnt_reg[3]  <= n2091;
    \\u5_ir_cnt_reg[0]  <= n2096;
    u5_mc_adv_r1_reg <= n2101;
    u5_tmr2_done_reg <= n2106;
    \\u3_u0_r0_reg[16]  <= n2111;
    \\u3_u0_r0_reg[22]  <= n2116;
    \\u3_u0_r1_reg[26]  <= n2121;
    \\u3_u0_r2_reg[25]  <= n2126;
    \\u3_u0_r2_reg[3]  <= n2131;
    \\u3_u0_r0_reg[1]  <= n2136;
    \\u3_u0_r0_reg[18]  <= n2141;
    \\u3_u0_r0_reg[19]  <= n2146;
    \\u3_u0_r0_reg[10]  <= n2151;
    \\u3_u0_r2_reg[32]  <= n2156;
    \\u3_u0_r2_reg[27]  <= n2161;
    \\u3_u0_r2_reg[29]  <= n2166;
    \\u3_u0_r0_reg[14]  <= n2171;
    \\u3_u0_r2_reg[18]  <= n2176;
    \\u3_u0_r2_reg[21]  <= n2181;
    \\u3_u0_wr_adr_reg[1]  <= n2186;
    \\u3_u0_wr_adr_reg[3]  <= n2191;
    u5_rfr_ack_r_reg <= n2196;
    \\u3_u0_r2_reg[14]  <= n2201;
    \\u3_u0_r2_reg[10]  <= n2206;
    \\u3_u0_r2_reg[12]  <= n2211;
    \\u3_u0_r1_reg[9]  <= n2216;
    \\u3_u0_r1_reg[7]  <= n2221;
    \\u3_u0_r1_reg[3]  <= n2226;
    \\u3_u0_r1_reg[32]  <= n2231;
    \\u3_u0_wr_adr_reg[0]  <= n2236;
    \\u3_u0_wr_adr_reg[2]  <= n2241;
    \\u3_u0_r0_reg[0]  <= n2246;
    \\u3_u0_r0_reg[11]  <= n2251;
    \\u3_u0_r0_reg[12]  <= n2256;
    \\u3_u0_r0_reg[13]  <= n2261;
    \\u3_u0_r0_reg[15]  <= n2266;
    \\u3_u0_r0_reg[17]  <= n2271;
    \\u3_u0_r0_reg[20]  <= n2276;
    \\u3_u0_r0_reg[21]  <= n2281;
    \\u3_u0_r0_reg[23]  <= n2286;
    \\u3_u0_r0_reg[24]  <= n2291;
    \\u3_u0_r0_reg[26]  <= n2296;
    \\u3_u0_r0_reg[27]  <= n2301;
    \\u3_u0_r0_reg[28]  <= n2306;
    \\u3_u0_r0_reg[2]  <= n2311;
    \\u3_u0_r0_reg[30]  <= n2316;
    \\u3_u0_r0_reg[31]  <= n2321;
    \\u3_u0_r0_reg[33]  <= n2326;
    \\u3_u0_r0_reg[34]  <= n2331;
    \\u3_u0_r0_reg[35]  <= n2336;
    \\u3_u0_r0_reg[4]  <= n2341;
    \\u3_u0_r0_reg[9]  <= n2346;
    \\u3_u0_r1_reg[0]  <= n2351;
    \\u3_u0_r1_reg[11]  <= n2356;
    \\u3_u0_r1_reg[10]  <= n2361;
    \\u3_u0_r1_reg[12]  <= n2366;
    \\u3_u0_r1_reg[13]  <= n2371;
    \\u3_u0_r1_reg[15]  <= n2376;
    \\u3_u0_r1_reg[16]  <= n2381;
    \\u3_u0_r1_reg[17]  <= n2386;
    \\u3_u0_r1_reg[19]  <= n2391;
    \\u3_u0_r1_reg[1]  <= n2396;
    \\u3_u0_r1_reg[20]  <= n2401;
    \\u3_u0_r1_reg[23]  <= n2406;
    \\u3_u0_r1_reg[22]  <= n2411;
    \\u3_u0_r1_reg[24]  <= n2416;
    \\u3_u0_r1_reg[25]  <= n2421;
    \\u3_u0_r1_reg[27]  <= n2426;
    \\u3_u0_r1_reg[28]  <= n2431;
    \\u3_u0_r1_reg[2]  <= n2436;
    \\u3_u0_r1_reg[30]  <= n2441;
    \\u3_u0_r1_reg[31]  <= n2446;
    \\u3_u0_r1_reg[33]  <= n2451;
    \\u3_u0_r1_reg[34]  <= n2456;
    \\u3_u0_r1_reg[35]  <= n2461;
    \\u3_u0_r1_reg[4]  <= n2466;
    \\u3_u0_r1_reg[5]  <= n2471;
    \\u3_u0_r1_reg[6]  <= n2476;
    \\u3_u0_r1_reg[8]  <= n2481;
    \\u3_u0_r2_reg[0]  <= n2486;
    \\u3_u0_r2_reg[11]  <= n2491;
    \\u3_u0_r2_reg[13]  <= n2496;
    \\u3_u0_r2_reg[15]  <= n2501;
    \\u3_u0_r2_reg[16]  <= n2506;
    \\u3_u0_r2_reg[17]  <= n2511;
    \\u3_u0_r2_reg[19]  <= n2516;
    \\u3_u0_r2_reg[1]  <= n2521;
    \\u3_u0_r2_reg[20]  <= n2526;
    \\u3_u0_r2_reg[22]  <= n2531;
    \\u3_u0_r2_reg[23]  <= n2536;
    \\u3_u0_r2_reg[24]  <= n2541;
    \\u3_u0_r2_reg[26]  <= n2546;
    \\u3_u0_r2_reg[28]  <= n2551;
    \\u3_u0_r2_reg[2]  <= n2556;
    \\u3_u0_r2_reg[30]  <= n2561;
    \\u3_u0_r2_reg[31]  <= n2566;
    \\u3_u0_r2_reg[33]  <= n2571;
    \\u3_u0_r2_reg[34]  <= n2576;
    \\u3_u0_r2_reg[35]  <= n2581;
    \\u3_u0_r2_reg[4]  <= n2586;
    \\u3_u0_r2_reg[5]  <= n2591;
    \\u3_u0_r2_reg[6]  <= n2596;
    \\u3_u0_r2_reg[8]  <= n2601;
    \\u3_u0_r3_reg[0]  <= n2606;
    \\u3_u0_r3_reg[11]  <= n2611;
    \\u3_u0_r3_reg[12]  <= n2616;
    \\u3_u0_r3_reg[13]  <= n2621;
    \\u3_u0_r3_reg[15]  <= n2626;
    \\u3_u0_r3_reg[16]  <= n2631;
    \\u3_u0_r3_reg[17]  <= n2636;
    \\u3_u0_r3_reg[19]  <= n2641;
    \\u3_u0_r3_reg[1]  <= n2646;
    \\u3_u0_r3_reg[20]  <= n2651;
    \\u3_u0_r3_reg[22]  <= n2656;
    \\u3_u0_r3_reg[23]  <= n2661;
    \\u3_u0_r3_reg[24]  <= n2666;
    \\u3_u0_r3_reg[26]  <= n2671;
    \\u3_u0_r3_reg[28]  <= n2676;
    \\u3_u0_r3_reg[2]  <= n2681;
    \\u3_u0_r3_reg[31]  <= n2686;
    \\u3_u0_r3_reg[33]  <= n2691;
    \\u3_u0_r3_reg[34]  <= n2696;
    \\u3_u0_r3_reg[35]  <= n2701;
    \\u3_u0_r3_reg[4]  <= n2706;
    \\u3_u0_r3_reg[5]  <= n2711;
    \\u3_u0_r3_reg[6]  <= n2716;
    \\u3_u0_r3_reg[9]  <= n2721;
    \\u3_u0_r3_reg[8]  <= n2726;
    \\u3_u0_r1_reg[29]  <= n2731;
    \\u3_u0_r1_reg[21]  <= n2736;
    \\u3_u0_r0_reg[7]  <= n2741;
    \\u3_u0_r1_reg[18]  <= n2746;
    \\u3_u0_r3_reg[7]  <= n2751;
    \\u3_u0_r3_reg[3]  <= n2756;
    \\u3_u0_r3_reg[30]  <= n2761;
    \\u3_u0_r3_reg[32]  <= n2766;
    \\u3_u0_r1_reg[14]  <= n2771;
    \\u3_u0_r3_reg[25]  <= n2776;
    \\u3_u0_r3_reg[29]  <= n2781;
    \\u3_u0_r0_reg[8]  <= n2786;
    \\u3_u0_r3_reg[27]  <= n2791;
    \\u3_u0_r0_reg[5]  <= n2796;
    \\u3_u0_r3_reg[14]  <= n2801;
    \\u3_u0_r3_reg[21]  <= n2806;
    \\u3_u0_r0_reg[6]  <= n2811;
    \\u3_u0_r2_reg[7]  <= n2816;
    u4_rfr_clr_reg <= n2821;
    \\u3_u0_r0_reg[3]  <= n2826;
    \\u3_u0_r3_reg[18]  <= n2831;
    \\u3_u0_r0_reg[32]  <= n2836;
    \\u3_u0_r0_reg[29]  <= n2841;
    \\u3_u0_r0_reg[25]  <= n2846;
    \\u3_u0_r2_reg[9]  <= n2851;
    \\u3_u0_r3_reg[10]  <= n2856;
    \\u7_mc_addr_reg[23]  <= n2861;
    \\u7_mc_addr_reg[17]  <= n2866;
    u7_mc_bg_reg <= n2871;
    u5_susp_sel_r_reg <= n2876;
    \\u7_mc_addr_reg[22]  <= n2881;
    \\u7_mc_addr_reg[21]  <= n2886;
    \\u7_mc_addr_reg[19]  <= n2891;
    \\u7_mc_addr_reg[20]  <= n2896;
    \\u7_mc_addr_reg[18]  <= n2901;
    \\u7_mc_addr_reg[16]  <= n2906;
    \\u7_mc_addr_reg[15]  <= n2911;
    u5_pack_le0_reg <= n2916;
    u7_mc_adv__reg <= n2921;
    u5_pack_le2_reg <= n2926;
    u5_wb_wait_r_reg <= n2931;
    u5_dv_r_reg <= n2936;
    \\u2_u0_b0_last_row_reg[6]  <= n2941;
    \\u2_u0_b3_last_row_reg[8]  <= n2946;
    \\u2_u1_b2_last_row_reg[0]  <= n2951;
    \\u2_u1_b2_last_row_reg[8]  <= n2956;
    \\u2_u1_b3_last_row_reg[10]  <= n2961;
    \\u2_u1_b3_last_row_reg[1]  <= n2966;
    \\u2_u0_b0_last_row_reg[4]  <= n2971;
    \\u2_u0_b0_last_row_reg[12]  <= n2976;
    \\u2_u1_b3_last_row_reg[0]  <= n2981;
    \\u2_u1_b2_last_row_reg[7]  <= n2986;
    \\u2_u1_b2_last_row_reg[9]  <= n2991;
    \\u2_u1_b2_last_row_reg[3]  <= n2996;
    \\u2_u1_b2_last_row_reg[1]  <= n3001;
    \\u2_u1_b2_last_row_reg[12]  <= n3006;
    \\u2_u1_b2_last_row_reg[11]  <= n3011;
    \\u2_u1_b1_last_row_reg[8]  <= n3016;
    \\u2_u1_b1_last_row_reg[12]  <= n3021;
    \\u2_u0_b3_last_row_reg[9]  <= n3026;
    \\u2_u1_b1_last_row_reg[4]  <= n3031;
    \\u2_u1_b1_last_row_reg[7]  <= n3036;
    \\u2_u1_b1_last_row_reg[6]  <= n3041;
    \\u2_u1_b1_last_row_reg[5]  <= n3046;
    \\u2_u1_b1_last_row_reg[2]  <= n3051;
    \\u2_u1_b0_last_row_reg[0]  <= n3056;
    \\u2_u1_b1_last_row_reg[10]  <= n3061;
    \\u2_u1_b0_last_row_reg[7]  <= n3066;
    \\u2_u1_b0_last_row_reg[9]  <= n3071;
    \\u2_u1_b0_last_row_reg[5]  <= n3076;
    \\u2_u1_b0_last_row_reg[2]  <= n3081;
    \\u2_u0_b0_last_row_reg[0]  <= n3086;
    \\u2_u0_b0_last_row_reg[10]  <= n3091;
    \\u2_u0_b0_last_row_reg[11]  <= n3096;
    \\u2_u0_b0_last_row_reg[1]  <= n3101;
    \\u2_u0_b0_last_row_reg[2]  <= n3106;
    \\u2_u0_b0_last_row_reg[3]  <= n3111;
    \\u2_u0_b0_last_row_reg[5]  <= n3116;
    \\u2_u0_b0_last_row_reg[9]  <= n3121;
    \\u2_u0_b1_last_row_reg[10]  <= n3126;
    \\u2_u0_b1_last_row_reg[12]  <= n3131;
    \\u2_u0_b1_last_row_reg[4]  <= n3136;
    \\u2_u0_b1_last_row_reg[6]  <= n3141;
    \\u2_u0_b1_last_row_reg[9]  <= n3146;
    \\u2_u0_b2_last_row_reg[10]  <= n3151;
    \\u2_u0_b2_last_row_reg[12]  <= n3156;
    \\u2_u0_b2_last_row_reg[2]  <= n3161;
    \\u2_u0_b2_last_row_reg[4]  <= n3166;
    \\u2_u0_b2_last_row_reg[5]  <= n3171;
    \\u2_u0_b2_last_row_reg[8]  <= n3176;
    \\u2_u0_b2_last_row_reg[9]  <= n3181;
    \\u2_u0_b2_last_row_reg[3]  <= n3186;
    \\u2_u0_b3_last_row_reg[11]  <= n3191;
    \\u2_u0_b3_last_row_reg[5]  <= n3196;
    \\u2_u1_b0_last_row_reg[11]  <= n3201;
    \\u2_u1_b0_last_row_reg[12]  <= n3206;
    \\u2_u1_b0_last_row_reg[3]  <= n3211;
    \\u2_u1_b0_last_row_reg[4]  <= n3216;
    \\u2_u1_b0_last_row_reg[6]  <= n3221;
    \\u2_u1_b0_last_row_reg[8]  <= n3226;
    \\u2_u1_b1_last_row_reg[0]  <= n3231;
    \\u2_u1_b1_last_row_reg[11]  <= n3236;
    \\u2_u1_b1_last_row_reg[1]  <= n3241;
    \\u2_u1_b1_last_row_reg[3]  <= n3246;
    \\u2_u1_b1_last_row_reg[9]  <= n3251;
    \\u2_u1_b2_last_row_reg[10]  <= n3256;
    \\u2_u1_b2_last_row_reg[2]  <= n3261;
    \\u2_u1_b2_last_row_reg[4]  <= n3266;
    \\u2_u1_b2_last_row_reg[5]  <= n3271;
    \\u2_u1_b2_last_row_reg[6]  <= n3276;
    \\u2_u1_b3_last_row_reg[11]  <= n3281;
    \\u2_u1_b3_last_row_reg[12]  <= n3286;
    \\u2_u1_b3_last_row_reg[3]  <= n3291;
    \\u2_u1_b3_last_row_reg[5]  <= n3296;
    \\u2_u1_b3_last_row_reg[7]  <= n3301;
    \\u2_u1_b3_last_row_reg[6]  <= n3306;
    \\u2_u1_b3_last_row_reg[8]  <= n3311;
    \\u2_u0_b3_last_row_reg[0]  <= n3316;
    \\u2_u1_b0_last_row_reg[10]  <= n3321;
    \\u2_u1_b0_last_row_reg[1]  <= n3326;
    \\u2_u0_b0_last_row_reg[7]  <= n3331;
    \\u2_u0_b3_last_row_reg[3]  <= n3336;
    \\u2_u0_b1_last_row_reg[5]  <= n3341;
    \\u2_u0_b3_last_row_reg[7]  <= n3346;
    \\u2_u1_b3_last_row_reg[4]  <= n3351;
    \\u2_u0_b3_last_row_reg[4]  <= n3356;
    \\u2_u0_b3_last_row_reg[6]  <= n3361;
    \\u2_u0_b3_last_row_reg[1]  <= n3366;
    u0_wp_err_reg <= n3371;
    \\u2_u0_b3_last_row_reg[2]  <= n3376;
    \\u2_u0_b3_last_row_reg[12]  <= n3381;
    \\u2_u0_b3_last_row_reg[10]  <= n3386;
    \\u2_u0_b2_last_row_reg[7]  <= n3391;
    \\u2_u0_b2_last_row_reg[1]  <= n3396;
    \\u2_u0_b2_last_row_reg[0]  <= n3401;
    \\u2_u0_b1_last_row_reg[7]  <= n3406;
    \\u2_u0_b2_last_row_reg[11]  <= n3411;
    \\u2_u0_b2_last_row_reg[6]  <= n3416;
    \\u2_u1_b3_last_row_reg[9]  <= n3421;
    \\u2_u0_b1_last_row_reg[8]  <= n3426;
    \\u2_u0_b0_last_row_reg[8]  <= n3431;
    \\u2_u1_b3_last_row_reg[2]  <= n3436;
    \\u2_u0_b1_last_row_reg[11]  <= n3441;
    \\u2_u0_b1_last_row_reg[3]  <= n3446;
    u5_wb_wait_r2_reg <= n3451;
    \\u2_u0_b1_last_row_reg[2]  <= n3456;
    \\u2_u0_b1_last_row_reg[1]  <= n3461;
    \\u2_u0_b1_last_row_reg[0]  <= n3466;
    \\u0_cs_reg[0]  <= n3471;
    \\u3_u0_rd_adr_reg[3]  <= n3476;
    u2_bank_open_reg <= n3481;
    \\u3_u0_rd_adr_reg[0]  <= n3486;
    \\u3_u0_rd_adr_reg[2]  <= n3491;
    \\u3_u0_rd_adr_reg[1]  <= n3496;
    u2_row_same_reg <= n3501;
    \\u4_rfr_cnt_reg[3]  <= n3506;
    \\u4_rfr_cnt_reg[5]  <= n3511;
    \\u4_rfr_cnt_reg[6]  <= n3516;
    \\u4_rfr_cnt_reg[4]  <= n3521;
    u0_u0_init_req_reg <= n3526;
    \\u4_rfr_cnt_reg[7]  <= n3531;
    \\u4_rfr_cnt_reg[2]  <= n3536;
    \\u4_rfr_cnt_reg[1]  <= n3541;
    \\u0_cs_reg[1]  <= n3546;
    \\u0_u0_csc_reg[0]  <= n3551;
    u0_u1_lmr_req_reg <= n3556;
    \\u4_rfr_cnt_reg[0]  <= n3561;
    \\u0_u0_csc_reg[4]  <= n3566;
    \\u0_u0_csc_reg[7]  <= n3571;
    \\u0_u0_csc_reg[16]  <= n3576;
    \\u0_u0_csc_reg[18]  <= n3581;
    \\u0_u0_csc_reg[13]  <= n3586;
    \\u0_u0_csc_reg[14]  <= n3591;
    \\u0_u0_csc_reg[11]  <= n3596;
    \\u0_u0_csc_reg[15]  <= n3601;
    \\u0_u0_csc_reg[2]  <= n3606;
    u0_u1_init_req_reg <= n3611;
    \\u0_u0_csc_reg[1]  <= n3616;
    \\u0_u0_csc_reg[5]  <= n3621;
    \\u0_u0_csc_reg[17]  <= n3626;
    \\u0_u0_csc_reg[22]  <= n3631;
    \\u0_u0_csc_reg[12]  <= n3636;
    \\u0_u0_csc_reg[8]  <= n3641;
    \\u0_u0_csc_reg[9]  <= n3646;
    \\u0_u0_csc_reg[6]  <= n3651;
    u0_u0_lmr_req_reg <= n3656;
    \\u0_u1_csc_reg[16]  <= n3661;
    \\u0_u0_csc_reg[21]  <= n3666;
    \\u0_u1_csc_reg[17]  <= n3671;
    \\u0_u1_csc_reg[19]  <= n3676;
    \\u0_u0_csc_reg[19]  <= n3681;
    \\u0_u0_csc_reg[20]  <= n3686;
    \\u0_u1_csc_reg[13]  <= n3691;
    \\u0_u1_csc_reg[15]  <= n3696;
    \\u0_u0_csc_reg[10]  <= n3701;
    \\u0_u1_csc_reg[10]  <= n3706;
    \\u0_u1_csc_reg[12]  <= n3711;
    \\u0_u0_csc_reg[27]  <= n3716;
    \\u0_u1_csc_reg[5]  <= n3721;
    \\u0_u1_csc_reg[7]  <= n3726;
    \\u0_u1_csc_reg[9]  <= n3731;
    \\u0_u0_csc_reg[28]  <= n3736;
    \\u0_u1_csc_reg[21]  <= n3741;
    \\u0_u0_csc_reg[3]  <= n3746;
    \\u0_u1_csc_reg[4]  <= n3751;
    \\u0_u0_csc_reg[23]  <= n3756;
    \\u0_u0_csc_reg[25]  <= n3761;
    \\u0_u1_csc_reg[14]  <= n3766;
    \\u0_u1_csc_reg[20]  <= n3771;
    \\u0_u1_csc_reg[22]  <= n3776;
    \\u0_u1_csc_reg[26]  <= n3781;
    \\u0_u1_csc_reg[27]  <= n3786;
    \\u0_u0_csc_reg[30]  <= n3791;
    \\u0_u0_csc_reg[31]  <= n3796;
    \\u0_u0_csc_reg[29]  <= n3801;
    \\u0_u1_csc_reg[30]  <= n3806;
    \\u0_u1_csc_reg[24]  <= n3811;
    \\u0_u0_csc_reg[26]  <= n3816;
    \\u0_u1_csc_reg[31]  <= n3821;
    \\u0_u0_csc_reg[24]  <= n3826;
    \\u1_u0_out_r_reg[11]  <= n3831;
    \\u0_u1_csc_reg[18]  <= n3836;
    \\u0_u1_csc_reg[1]  <= n3841;
    \\u0_u1_csc_reg[2]  <= n3846;
    \\u6_wb_data_o_reg[10]  <= n3851;
    \\u6_wb_data_o_reg[2]  <= n3856;
    \\u0_u1_csc_reg[8]  <= n3861;
    \\u6_wb_data_o_reg[7]  <= n3866;
    \\u6_wb_data_o_reg[3]  <= n3871;
    \\u6_wb_data_o_reg[0]  <= n3876;
    \\u0_u1_csc_reg[25]  <= n3881;
    \\u6_wb_data_o_reg[11]  <= n3886;
    \\u6_wb_data_o_reg[14]  <= n3891;
    \\u6_wb_data_o_reg[1]  <= n3896;
    \\u6_wb_data_o_reg[5]  <= n3901;
    \\u6_wb_data_o_reg[9]  <= n3906;
    \\u6_wb_data_o_reg[6]  <= n3911;
    \\u6_wb_data_o_reg[4]  <= n3916;
    \\u6_wb_data_o_reg[12]  <= n3921;
    \\u6_wb_data_o_reg[15]  <= n3926;
    \\u6_wb_data_o_reg[8]  <= n3931;
    \\u0_u1_csc_reg[0]  <= n3936;
    \\u0_u1_csc_reg[3]  <= n3941;
    \\u6_wb_data_o_reg[13]  <= n3946;
    u5_wb_write_go_r_reg <= n3951;
    \\u0_u1_tms_reg[30]  <= n3956;
    \\u6_wb_data_o_reg[31]  <= n3961;
    \\u0_u1_tms_reg[13]  <= n3966;
    \\u0_u1_tms_reg[27]  <= n3971;
    \\u0_u1_tms_reg[15]  <= n3976;
    \\u6_wb_data_o_reg[24]  <= n3981;
    \\u0_u1_tms_reg[8]  <= n3986;
    \\u0_u1_tms_reg[7]  <= n3991;
    \\u6_wb_data_o_reg[26]  <= n3996;
    \\u0_u1_csc_reg[29]  <= n4001;
    \\u0_u1_tms_reg[28]  <= n4006;
    \\u0_u1_csc_reg[11]  <= n4011;
    \\u0_u1_tms_reg[0]  <= n4016;
    \\u0_u1_tms_reg[29]  <= n4021;
    \\u0_u1_tms_reg[16]  <= n4026;
    \\u0_u1_tms_reg[3]  <= n4031;
    \\u0_u1_tms_reg[10]  <= n4036;
    \\u0_u1_tms_reg[23]  <= n4041;
    \\u0_u1_tms_reg[17]  <= n4046;
    \\u0_u1_tms_reg[24]  <= n4051;
    \\u0_u1_tms_reg[12]  <= n4056;
    \\u0_u1_tms_reg[25]  <= n4061;
    \\u0_u1_tms_reg[5]  <= n4066;
    \\u6_wb_data_o_reg[17]  <= n4071;
    \\u6_wb_data_o_reg[18]  <= n4076;
    \\u0_u1_tms_reg[18]  <= n4081;
    \\u0_u1_csc_reg[6]  <= n4086;
    \\u6_wb_data_o_reg[20]  <= n4091;
    \\u6_wb_data_o_reg[23]  <= n4096;
    \\u6_wb_data_o_reg[19]  <= n4101;
    \\u6_wb_data_o_reg[29]  <= n4106;
    \\u0_u1_csc_reg[23]  <= n4111;
    \\u6_wb_data_o_reg[21]  <= n4116;
    \\u6_wb_data_o_reg[25]  <= n4121;
    \\u6_wb_data_o_reg[16]  <= n4126;
    \\u6_wb_data_o_reg[27]  <= n4131;
    \\u6_wb_data_o_reg[30]  <= n4136;
    \\u4_ps_cnt_reg[7]  <= n4141;
    \\u6_wb_data_o_reg[28]  <= n4146;
    \\u0_u1_tms_reg[11]  <= n4151;
    \\u0_u1_tms_reg[14]  <= n4156;
    \\u0_u1_tms_reg[20]  <= n4161;
    \\u0_u1_tms_reg[26]  <= n4166;
    \\u0_u1_tms_reg[2]  <= n4171;
    \\u0_u1_tms_reg[31]  <= n4176;
    \\u0_u1_tms_reg[4]  <= n4181;
    \\u0_u1_tms_reg[6]  <= n4186;
    \\u4_ps_cnt_reg[4]  <= n4191;
    \\u0_u1_csc_reg[28]  <= n4196;
    \\u6_wb_data_o_reg[22]  <= n4201;
    \\u0_u1_tms_reg[19]  <= n4206;
    \\u0_u1_tms_reg[9]  <= n4211;
    \\u0_u1_tms_reg[1]  <= n4216;
    \\u0_u1_tms_reg[22]  <= n4221;
    \\u0_u1_tms_reg[21]  <= n4226;
    \\u0_u0_tms_reg[8]  <= n4231;
    u0_u0_init_req_we_reg <= n4236;
    \\u0_u0_tms_reg[14]  <= n4241;
    \\u0_u0_tms_reg[12]  <= n4246;
    \\u0_u0_tms_reg[9]  <= n4251;
    \\u0_u0_tms_reg[31]  <= n4256;
    \\u0_u0_tms_reg[11]  <= n4261;
    \\u0_u0_tms_reg[4]  <= n4266;
    \\u4_ps_cnt_reg[3]  <= n4271;
    \\u0_u0_tms_reg[6]  <= n4276;
    \\u0_u0_tms_reg[5]  <= n4281;
    \\u0_u0_tms_reg[30]  <= n4286;
    \\u0_u0_tms_reg[23]  <= n4291;
    \\u0_u0_tms_reg[24]  <= n4296;
    \\u0_u0_tms_reg[17]  <= n4301;
    \\u0_u0_tms_reg[18]  <= n4306;
    \\u0_u0_tms_reg[20]  <= n4311;
    \\u0_u0_tms_reg[19]  <= n4316;
    \\u0_u0_tms_reg[13]  <= n4321;
    \\u0_u0_tms_reg[1]  <= n4326;
    \\u0_u0_tms_reg[0]  <= n4331;
    \\u0_u0_tms_reg[15]  <= n4336;
    \\u0_u0_tms_reg[21]  <= n4341;
    \\u0_u0_tms_reg[29]  <= n4346;
    \\u0_u0_tms_reg[3]  <= n4351;
    \\u0_u0_tms_reg[7]  <= n4356;
    \\u4_ps_cnt_reg[0]  <= n4361;
    \\u0_u0_tms_reg[10]  <= n4366;
    \\u0_u0_tms_reg[16]  <= n4371;
    \\u0_u0_tms_reg[25]  <= n4376;
    \\u4_ps_cnt_reg[6]  <= n4381;
    \\u0_u0_tms_reg[26]  <= n4386;
    \\u4_ps_cnt_reg[1]  <= n4391;
    \\u0_u0_tms_reg[2]  <= n4396;
    \\u4_ps_cnt_reg[2]  <= n4401;
    \\u0_u0_tms_reg[27]  <= n4406;
    \\u4_ps_cnt_reg[5]  <= n4411;
    \\u0_u0_tms_reg[28]  <= n4416;
    \\u0_u0_tms_reg[22]  <= n4421;
    \\u0_csc_mask_r_reg[0]  <= n4426;
    u0_u1_inited_reg <= n4431;
    u0_u0_inited_reg <= n4436;
    \\u0_csc_mask_r_reg[1]  <= n4441;
    u0_sreq_cs_le_reg <= n4446;
    \\u0_csc_mask_r_reg[9]  <= n4451;
    \\u0_csc_mask_r_reg[10]  <= n4456;
    \\u0_csc_mask_r_reg[2]  <= n4461;
    u5_cmd_asserted2_reg <= n4466;
    \\u0_csc_mask_r_reg[4]  <= n4471;
    \\u0_csc_mask_r_reg[5]  <= n4476;
    \\u0_csc_mask_r_reg[6]  <= n4481;
    \\u0_csc_mask_r_reg[7]  <= n4486;
    \\u0_csc_mask_r_reg[8]  <= n4491;
    \\u0_csc_mask_r_reg[3]  <= n4496;
    u5_no_wb_cycle_reg <= n4501;
    \\u0_csr_r2_reg[6]  <= n4506;
    \\u0_csr_r2_reg[4]  <= n4511;
    \\u1_u0_out_r_reg[9]  <= n4516;
    u0_u1_init_req_we_reg <= n4521;
    \\u0_csr_r2_reg[0]  <= n4526;
    \\u0_csr_r_reg[7]  <= n4531;
    \\u0_csr_r2_reg[1]  <= n4536;
    \\u0_csr_r2_reg[2]  <= n4541;
    \\u1_u0_out_r_reg[12]  <= n4546;
    \\u0_csr_r_reg[6]  <= n4551;
    \\u0_csr_r_reg[9]  <= n4556;
    \\u1_u0_out_r_reg[7]  <= n4561;
    u4_rfr_ce_reg <= n4566;
    \\u0_csr_r2_reg[3]  <= n4571;
    \\u0_csr_r_reg[1]  <= n4576;
    \\u0_csr_r_reg[3]  <= n4581;
    \\u0_csr_r_reg[8]  <= n4586;
    \\u0_csr_r_reg[2]  <= n4591;
    \\u0_csr_r_reg[4]  <= n4596;
    \\u0_csr_r2_reg[7]  <= n4601;
    \\u0_csr_r_reg[5]  <= n4606;
    \\u0_csr_r_reg[10]  <= n4611;
    \\u0_csr_r2_reg[5]  <= n4616;
    \\u1_u0_out_r_reg[4]  <= n4621;
    u6_wb_first_r_reg <= n4626;
    \\u1_u0_out_r_reg[10]  <= n4631;
    \\u1_u0_out_r_reg[8]  <= n4636;
    u4_rfr_early_reg <= n4641;
    u7_mc_rp_reg <= n4646;
    u0_u1_lmr_req_we_reg <= n4651;
    u6_read_go_r1_reg <= n4656;
    \\u3_mc_dp_o_reg[3]  <= n4661;
    \\u3_mc_dp_o_reg[2]  <= n4666;
    \\u3_mc_dp_o_reg[0]  <= n4671;
    \\u3_mc_dp_o_reg[1]  <= n4676;
    u6_write_go_r1_reg <= n4681;
    \\u1_u0_out_r_reg[5]  <= n4686;
    u0_u0_lmr_req_we_reg <= n4691;
    u0_rf_we_reg <= n4696;
    u6_wr_hold_reg <= n4701;
    u7_mc_zz_o_reg <= n4706;
    u5_lookup_ready2_reg <= n4711;
    \\u1_u0_out_r_reg[6]  <= n4716;
    \\u0_poc_reg[0]  <= n4721;
    \\u0_poc_reg[22]  <= n4726;
    \\u0_poc_reg[25]  <= n4731;
    \\u7_mc_dqm_r_reg[0]  <= n4736;
    u5_tmr_done_reg <= n4741;
    \\u0_poc_reg[23]  <= n4746;
    \\u0_poc_reg[24]  <= n4751;
    \\u0_poc_reg[26]  <= n4756;
    \\u0_poc_reg[21]  <= n4761;
    \\u1_col_adr_reg[0]  <= n4766;
    \\u0_poc_reg[17]  <= n4771;
    \\u0_poc_reg[13]  <= n4776;
    \\u7_mc_dqm_r_reg[2]  <= n4781;
    \\u0_poc_reg[1]  <= n4786;
    \\u0_poc_reg[28]  <= n4791;
    \\u0_poc_reg[11]  <= n4796;
    \\u0_poc_reg[16]  <= n4801;
    \\u0_poc_reg[19]  <= n4806;
    \\u0_poc_reg[10]  <= n4811;
    \\u0_poc_reg[15]  <= n4816;
    \\u0_poc_reg[18]  <= n4821;
    \\u0_poc_reg[20]  <= n4826;
    \\u0_poc_reg[9]  <= n4831;
    \\u0_poc_reg[31]  <= n4836;
    \\u1_col_adr_reg[7]  <= n4841;
    \\u1_col_adr_reg[5]  <= n4846;
    \\u7_mc_dqm_r_reg[3]  <= n4851;
    \\u7_mc_dqm_r_reg[1]  <= n4856;
    \\u0_poc_reg[14]  <= n4861;
    \\u0_poc_reg[5]  <= n4866;
    \\u0_poc_reg[29]  <= n4871;
    \\u0_poc_reg[27]  <= n4876;
    \\u1_col_adr_reg[6]  <= n4881;
    \\u0_poc_reg[12]  <= n4886;
    \\u0_poc_reg[3]  <= n4891;
    \\u0_poc_reg[2]  <= n4896;
    \\u0_poc_reg[7]  <= n4901;
    \\u0_poc_reg[8]  <= n4906;
    \\u1_col_adr_reg[2]  <= n4911;
    \\u0_poc_reg[6]  <= n4916;
    \\u1_col_adr_reg[4]  <= n4921;
    \\u1_col_adr_reg[3]  <= n4926;
    \\u1_col_adr_reg[1]  <= n4931;
    \\u0_poc_reg[30]  <= n4936;
    \\u0_poc_reg[4]  <= n4941;
    u0_init_ack_r_reg <= n4946;
    \\u3_mc_data_o_reg[7]  <= n4951;
    \\u3_mc_data_o_reg[24]  <= n4956;
    \\u3_mc_data_o_reg[25]  <= n4961;
    \\u3_mc_data_o_reg[9]  <= n4966;
    \\u3_mc_data_o_reg[0]  <= n4971;
    \\u3_mc_data_o_reg[20]  <= n4976;
    \\u3_mc_data_o_reg[3]  <= n4981;
    \\u3_mc_data_o_reg[26]  <= n4986;
    \\u3_mc_data_o_reg[16]  <= n4991;
    \\u3_mc_data_o_reg[1]  <= n4996;
    u5_suspended_reg <= n5001;
    \\u3_mc_data_o_reg[19]  <= n5006;
    \\u3_mc_data_o_reg[13]  <= n5011;
    \\u3_mc_data_o_reg[18]  <= n5016;
    u5_pack_le1_reg <= n5021;
    \\u3_mc_data_o_reg[29]  <= n5026;
    \\u3_mc_data_o_reg[15]  <= n5031;
    \\u3_mc_data_o_reg[10]  <= n5036;
    u5_burst_act_rd_reg <= n5041;
    \\u3_mc_data_o_reg[11]  <= n5046;
    \\u3_mc_data_o_reg[21]  <= n5051;
    \\u3_mc_data_o_reg[27]  <= n5056;
    \\u3_mc_data_o_reg[31]  <= n5061;
    \\u3_mc_data_o_reg[28]  <= n5066;
    \\u0_spec_req_cs_reg[1]  <= n5071;
    \\u3_mc_data_o_reg[22]  <= n5076;
    \\u3_mc_data_o_reg[5]  <= n5081;
    \\u3_mc_data_o_reg[17]  <= n5086;
    \\u3_mc_data_o_reg[30]  <= n5091;
    \\u3_mc_data_o_reg[14]  <= n5096;
    \\u3_mc_data_o_reg[6]  <= n5101;
    \\u1_u0_out_r_reg[3]  <= n5106;
    \\u3_mc_data_o_reg[8]  <= n5111;
    \\u3_mc_data_o_reg[23]  <= n5116;
    \\u3_mc_data_o_reg[12]  <= n5121;
    \\u3_mc_data_o_reg[4]  <= n5126;
    \\u3_mc_data_o_reg[2]  <= n5131;
    \\u1_sram_addr_reg[5]  <= n5136;
    \\u1_sram_addr_reg[6]  <= n5141;
    \\u1_sram_addr_reg[18]  <= n5146;
    \\u1_sram_addr_reg[20]  <= n5151;
    u5_ir_cnt_done_reg <= n5156;
    \\u1_sram_addr_reg[21]  <= n5161;
    \\u1_sram_addr_reg[23]  <= n5166;
    \\u1_sram_addr_reg[11]  <= n5171;
    \\u1_sram_addr_reg[2]  <= n5176;
    \\u1_sram_addr_reg[10]  <= n5181;
    \\u1_sram_addr_reg[0]  <= n5186;
    \\u1_sram_addr_reg[16]  <= n5191;
    \\u1_sram_addr_reg[8]  <= n5196;
    \\u1_sram_addr_reg[3]  <= n5201;
    \\u1_sram_addr_reg[13]  <= n5206;
    \\u1_sram_addr_reg[7]  <= n5211;
    \\u1_sram_addr_reg[15]  <= n5216;
    \\u1_sram_addr_reg[14]  <= n5221;
    \\u1_sram_addr_reg[1]  <= n5226;
    \\u1_sram_addr_reg[12]  <= n5231;
    \\u1_sram_addr_reg[4]  <= n5236;
    \\u1_sram_addr_reg[19]  <= n5241;
    \\u1_sram_addr_reg[22]  <= n5246;
    \\u1_sram_addr_reg[17]  <= n5251;
    \\u1_sram_addr_reg[9]  <= n5256;
    u4_rfr_en_reg <= n5261;
    u5_lookup_ready1_reg <= n5266;
    \\u0_spec_req_cs_reg[0]  <= n5271;
    \\u1_u0_out_r_reg[2]  <= n5276;
    u5_mc_adv_r_reg <= n5281;
    u6_rmw_r_reg <= n5286;
    u6_write_go_r_reg <= n5291;
    \\u0_u0_addr_r_reg[2]  <= n5296;
    \\u0_u1_addr_r_reg[2]  <= n5301;
    u5_mc_le_reg <= n5306;
    u0_rst_r3_reg <= n5311;
    \\u0_wb_addr_r_reg[2]  <= n5316;
    u6_rmw_en_reg <= n5321;
    \\u1_u0_out_r_reg[1]  <= n5326;
    u5_cke_o_del_reg <= n5331;
    \\u0_spec_req_cs_reg[5]  <= n5336;
    \\u0_cs_reg[6]  <= n5341;
    u0_u1_rst_r2_reg <= n5346;
    \\u0_spec_req_cs_reg[4]  <= n5351;
    u5_rsts_reg <= n5356;
    u0_rst_r2_reg <= n5361;
    u0_u0_rst_r2_reg <= n5366;
    \\u0_cs_reg[7]  <= n5371;
    \\u0_wb_addr_r_reg[3]  <= n5376;
    \\u0_cs_reg[4]  <= n5381;
    \\u0_spec_req_cs_reg[7]  <= n5386;
    \\u0_cs_reg[3]  <= n5391;
    \\u0_spec_req_cs_reg[6]  <= n5396;
    \\u0_u1_addr_r_reg[3]  <= n5401;
    \\u0_cs_reg[2]  <= n5406;
    \\u0_spec_req_cs_reg[3]  <= n5411;
    \\u1_u0_out_r_reg[0]  <= n5416;
    \\u0_cs_reg[5]  <= n5421;
    \\u0_spec_req_cs_reg[2]  <= n5426;
    u0_init_req_reg <= n5431;
    \\u0_u0_addr_r_reg[3]  <= n5436;
    \\u0_csr_r_reg[0]  <= n5441;
    u6_read_go_r_reg <= n5446;
    u0_lmr_ack_r_reg <= n5451;
    u0_lmr_req_reg <= n5456;
    u5_cke_o_r2_reg <= n5461;
    u5_cs_le_r_reg <= n5466;
    \\u7_mc_data_o_reg[8]  <= n5471;
    \\u7_mc_dp_o_reg[3]  <= n5476;
    \\u7_mc_dp_o_reg[2]  <= n5481;
    \\u7_mc_data_o_reg[6]  <= n5486;
    \\u7_mc_data_o_reg[19]  <= n5491;
    \\u7_mc_data_o_reg[31]  <= n5496;
    u5_resume_req_r_reg <= n5501;
    \\u7_mc_data_o_reg[26]  <= n5506;
    u5_susp_req_r_reg <= n5511;
    \\u7_mc_data_o_reg[28]  <= n5516;
    \\u7_mc_data_o_reg[18]  <= n5521;
    u0_rst_r1_reg <= n5526;
    \\u7_mc_data_o_reg[5]  <= n5531;
    \\u7_mc_data_o_reg[30]  <= n5536;
    u0_u0_rst_r1_reg <= n5541;
    \\u7_mc_data_o_reg[22]  <= n5546;
    \\u7_mc_data_o_reg[16]  <= n5551;
    \\u7_mc_data_o_reg[11]  <= n5556;
    \\u7_mc_data_o_reg[21]  <= n5561;
    \\u7_mc_data_o_reg[7]  <= n5566;
    \\u7_mc_data_o_reg[20]  <= n5571;
    u0_u1_rst_r1_reg <= n5576;
    \\u7_mc_data_o_reg[2]  <= n5581;
    \\u7_mc_data_o_reg[9]  <= n5586;
    \\u7_mc_data_o_reg[14]  <= n5591;
    \\u7_mc_data_o_reg[13]  <= n5596;
    \\u7_mc_data_o_reg[23]  <= n5601;
    \\u7_mc_data_o_reg[3]  <= n5606;
    \\u7_mc_data_o_reg[10]  <= n5611;
    \\u7_mc_data_o_reg[25]  <= n5616;
    \\u7_mc_data_o_reg[27]  <= n5621;
    \\u7_mc_data_o_reg[15]  <= n5626;
    \\u7_mc_data_o_reg[4]  <= n5631;
    \\u7_mc_data_o_reg[29]  <= n5636;
    \\u7_mc_data_o_reg[12]  <= n5641;
    \\u7_mc_dp_o_reg[0]  <= n5646;
    u5_rsts1_reg <= n5651;
    \\u7_mc_data_o_reg[0]  <= n5656;
    \\u7_mc_data_o_reg[24]  <= n5661;
    \\u7_mc_data_o_reg[17]  <= n5666;
    \\u7_mc_dp_o_reg[1]  <= n5671;
    \\u7_mc_data_o_reg[1]  <= n5676;
    \\u7_mc_data_ir_reg[23]  <= n5681;
    \\u7_mc_data_ir_reg[8]  <= n5686;
    \\u7_mc_data_ir_reg[6]  <= n5691;
    \\u0_u0_addr_r_reg[6]  <= n5696;
    \\u7_mc_data_ir_reg[13]  <= n5701;
    \\u7_mc_data_ir_reg[14]  <= n5706;
    \\u7_mc_dqm_r2_reg[3]  <= n5711;
    \\u7_mc_data_ir_reg[35]  <= n5716;
    \\u7_mc_data_ir_reg[21]  <= n5721;
    \\u7_mc_data_ir_reg[7]  <= n5726;
    \\u7_mc_data_ir_reg[28]  <= n5731;
    \\u0_wb_addr_r_reg[5]  <= n5736;
    \\u7_mc_data_ir_reg[22]  <= n5741;
    \\u7_mc_data_ir_reg[1]  <= n5746;
    \\u7_mc_data_ir_reg[0]  <= n5751;
    u7_mc_ack_r_reg <= n5756;
    \\u7_mc_data_ir_reg[19]  <= n5761;
    u5_cs_le_r1_reg <= n5766;
    \\u7_mc_data_ir_reg[5]  <= n5771;
    \\u0_u1_addr_r_reg[4]  <= n5776;
    \\u7_mc_data_ir_reg[17]  <= n5781;
    \\u7_mc_dqm_r2_reg[2]  <= n5786;
    \\u7_mc_data_ir_reg[29]  <= n5791;
    \\u7_mc_data_ir_reg[18]  <= n5796;
    \\u7_mc_data_ir_reg[4]  <= n5801;
    \\u0_u0_addr_r_reg[5]  <= n5806;
    \\u0_u0_addr_r_reg[4]  <= n5811;
    \\u7_mc_data_ir_reg[11]  <= n5816;
    \\u7_mc_data_ir_reg[27]  <= n5821;
    u7_mc_sts_ir_reg <= n5826;
    \\u7_mc_data_ir_reg[10]  <= n5831;
    \\u0_u1_addr_r_reg[5]  <= n5836;
    \\u7_mc_data_ir_reg[15]  <= n5841;
    \\u7_mc_data_ir_reg[34]  <= n5846;
    \\u7_mc_data_ir_reg[12]  <= n5851;
    \\u7_mc_data_ir_reg[9]  <= n5856;
    \\u7_mc_data_ir_reg[33]  <= n5861;
    \\u7_mc_data_ir_reg[3]  <= n5866;
    \\u7_mc_dqm_r2_reg[0]  <= n5871;
    \\u7_mc_data_ir_reg[25]  <= n5876;
    u5_cke_o_r1_reg <= n5881;
    \\u7_mc_data_ir_reg[31]  <= n5886;
    \\u7_mc_dqm_r2_reg[1]  <= n5891;
    \\u7_mc_data_ir_reg[26]  <= n5896;
    \\u7_mc_data_ir_reg[24]  <= n5901;
    \\u7_mc_data_ir_reg[16]  <= n5906;
    \\u7_mc_data_ir_reg[30]  <= n5911;
    u7_mc_br_r_reg <= n5916;
    \\u0_wb_addr_r_reg[6]  <= n5921;
    \\u7_mc_data_ir_reg[2]  <= n5926;
    \\u0_wb_addr_r_reg[4]  <= n5931;
    \\u7_mc_data_ir_reg[32]  <= n5936;
    \\u7_mc_data_ir_reg[20]  <= n5941;
    \\u0_u1_addr_r_reg[6]  <= n5946;
  end
  initial begin
    \\u7_mc_cs__reg[1]  <= 1'b1;
    \\u7_mc_cs__reg[0]  <= 1'b1;
    \\u7_mc_cs__reg[7]  <= 1'b1;
    \\u7_mc_cs__reg[6]  <= 1'b1;
    \\u7_mc_cs__reg[5]  <= 1'b1;
    \\u7_mc_cs__reg[4]  <= 1'b1;
    \\u7_mc_cs__reg[3]  <= 1'b1;
    \\u7_mc_cs__reg[2]  <= 1'b1;
    \\u5_cmd_del_reg[0]  <= 1'b1;
    \\u5_cmd_r_reg[0]  <= 1'b1;
    u5_cmd_asserted_reg <= 1'b0;
    \\u5_cmd_del_reg[3]  <= 1'b0;
    u6_wb_ack_o_reg <= 1'b0;
    \\u5_state_reg[16]  <= 1'b0;
    \\u5_timer_reg[0]  <= 1'b0;
    \\u5_timer_reg[1]  <= 1'b1;
    \\u5_state_reg[2]  <= 1'b0;
    \\u5_state_reg[59]  <= 1'b0;
    \\u5_cmd_r_reg[3]  <= 1'b0;
    \\u5_state_reg[17]  <= 1'b0;
    \\u5_state_reg[1]  <= 1'b0;
    \\u5_state_reg[35]  <= 1'b0;
    \\u5_state_reg[21]  <= 1'b0;
    \\u5_state_reg[29]  <= 1'b0;
    \\u5_state_reg[57]  <= 1'b0;
    \\u5_state_reg[0]  <= 1'b1;
    \\u5_state_reg[10]  <= 1'b0;
    \\u5_state_reg[15]  <= 1'b0;
    \\u5_state_reg[40]  <= 1'b0;
    \\u5_state_reg[18]  <= 1'b0;
    \\u5_state_reg[20]  <= 1'b0;
    \\u5_state_reg[22]  <= 1'b0;
    \\u5_state_reg[23]  <= 1'b0;
    \\u5_state_reg[24]  <= 1'b0;
    \\u5_state_reg[62]  <= 1'b0;
    \\u5_state_reg[26]  <= 1'b0;
    \\u5_state_reg[27]  <= 1'b0;
    \\u5_state_reg[28]  <= 1'b0;
    \\u5_state_reg[25]  <= 1'b0;
    \\u5_state_reg[30]  <= 1'b0;
    \\u5_state_reg[32]  <= 1'b0;
    \\u5_state_reg[33]  <= 1'b0;
    \\u5_state_reg[38]  <= 1'b0;
    \\u5_state_reg[43]  <= 1'b0;
    \\u5_state_reg[36]  <= 1'b0;
    \\u5_state_reg[46]  <= 1'b0;
    \\u5_state_reg[4]  <= 1'b0;
    \\u5_state_reg[45]  <= 1'b0;
    \\u5_state_reg[52]  <= 1'b0;
    \\u5_state_reg[60]  <= 1'b0;
    \\u5_state_reg[9]  <= 1'b0;
    \\u5_state_reg[13]  <= 1'b0;
    \\u5_state_reg[12]  <= 1'b0;
    \\u5_state_reg[48]  <= 1'b0;
    u7_mc_data_oe_reg <= 1'b0;
    \\u5_timer_reg[2]  <= 1'b0;
    u6_wb_err_reg <= 1'b0;
    \\u5_state_reg[37]  <= 1'b0;
    \\u5_state_reg[39]  <= 1'b0;
    \\u5_state_reg[42]  <= 1'b0;
    \\u5_state_reg[41]  <= 1'b0;
    \\u5_state_reg[44]  <= 1'b0;
    \\u5_state_reg[47]  <= 1'b0;
    \\u5_state_reg[51]  <= 1'b0;
    \\u5_state_reg[56]  <= 1'b0;
    \\u5_state_reg[5]  <= 1'b0;
    \\u5_state_reg[61]  <= 1'b0;
    \\u5_state_reg[58]  <= 1'b0;
    \\u5_state_reg[63]  <= 1'b0;
    \\u5_state_reg[64]  <= 1'b0;
    \\u5_state_reg[11]  <= 1'b0;
    \\u5_state_reg[6]  <= 1'b0;
    \\u5_state_reg[7]  <= 1'b0;
    \\u5_state_reg[8]  <= 1'b0;
    \\u5_state_reg[65]  <= 1'b0;
    \\u5_state_reg[14]  <= 1'b0;
    \\u5_state_reg[34]  <= 1'b0;
    \\u5_state_reg[50]  <= 1'b0;
    \\u5_state_reg[55]  <= 1'b0;
    \\u5_cmd_del_reg[1]  <= 1'b1;
    \\u5_state_reg[19]  <= 1'b0;
    \\u5_state_reg[31]  <= 1'b0;
    \\u5_state_reg[3]  <= 1'b0;
    \\u5_state_reg[49]  <= 1'b0;
    \\u5_state_reg[54]  <= 1'b0;
    \\u5_state_reg[53]  <= 1'b0;
    u7_mc_oe__reg <= 1'b1;
    \\u5_cmd_r_reg[1]  <= 1'b1;
    \\u5_timer_reg[3]  <= 1'b1;
    u5_data_oe_reg <= 1'b0;
    u5_wb_stb_first_reg <= 1'b0;
    u5_mem_ack_r_reg <= 1'b0;
    u5_oe__reg <= 1'b1;
    u5_data_oe_r2_reg <= 1'b0;
    u5_data_oe_r_reg <= 1'b0;
    u5_ap_en_reg <= 1'b0;
    \\u5_timer_reg[5]  <= 1'b1;
    \\u5_timer_reg[4]  <= 1'b1;
    \\u0_tms_reg[21]  <= 1'b1;
    \\u0_tms_reg[5]  <= 1'b1;
    \\u0_tms_reg[9]  <= 1'b1;
    \\u0_tms_reg[27]  <= 1'b1;
    \\u0_tms_reg[1]  <= 1'b1;
    \\u0_tms_reg[16]  <= 1'b1;
    \\u0_sp_tms_reg[9]  <= 1'b1;
    \\u0_sp_tms_reg[26]  <= 1'b1;
    \\u0_sp_tms_reg[5]  <= 1'b1;
    \\u0_sp_tms_reg[20]  <= 1'b1;
    \\u0_sp_tms_reg[23]  <= 1'b1;
    \\u0_sp_tms_reg[11]  <= 1'b1;
    \\u0_sp_tms_reg[0]  <= 1'b1;
    \\u0_sp_tms_reg[10]  <= 1'b1;
    \\u0_sp_tms_reg[12]  <= 1'b1;
    \\u0_sp_tms_reg[13]  <= 1'b1;
    \\u0_sp_tms_reg[14]  <= 1'b1;
    \\u0_sp_tms_reg[15]  <= 1'b1;
    \\u0_sp_tms_reg[17]  <= 1'b1;
    \\u0_sp_tms_reg[18]  <= 1'b1;
    \\u0_sp_tms_reg[19]  <= 1'b1;
    \\u0_sp_tms_reg[1]  <= 1'b1;
    \\u0_sp_tms_reg[21]  <= 1'b1;
    \\u0_sp_tms_reg[22]  <= 1'b1;
    \\u0_sp_tms_reg[24]  <= 1'b1;
    \\u0_sp_tms_reg[27]  <= 1'b1;
    \\u0_sp_tms_reg[2]  <= 1'b1;
    \\u0_sp_tms_reg[25]  <= 1'b1;
    \\u0_sp_tms_reg[3]  <= 1'b1;
    \\u0_sp_tms_reg[4]  <= 1'b1;
    \\u0_sp_tms_reg[6]  <= 1'b1;
    \\u0_sp_tms_reg[7]  <= 1'b1;
    \\u0_sp_tms_reg[8]  <= 1'b1;
    \\u0_tms_reg[11]  <= 1'b1;
    \\u0_tms_reg[0]  <= 1'b1;
    \\u0_tms_reg[10]  <= 1'b1;
    \\u0_tms_reg[12]  <= 1'b1;
    \\u0_tms_reg[13]  <= 1'b1;
    \\u0_tms_reg[15]  <= 1'b1;
    \\u0_tms_reg[14]  <= 1'b1;
    \\u0_tms_reg[17]  <= 1'b1;
    \\u0_tms_reg[18]  <= 1'b1;
    \\u0_tms_reg[19]  <= 1'b1;
    \\u0_tms_reg[20]  <= 1'b1;
    \\u0_tms_reg[22]  <= 1'b1;
    \\u0_tms_reg[23]  <= 1'b1;
    \\u0_tms_reg[24]  <= 1'b1;
    \\u0_tms_reg[26]  <= 1'b1;
    \\u0_tms_reg[25]  <= 1'b1;
    \\u0_tms_reg[2]  <= 1'b1;
    \\u0_tms_reg[3]  <= 1'b1;
    \\u0_tms_reg[4]  <= 1'b1;
    \\u0_tms_reg[7]  <= 1'b1;
    \\u0_tms_reg[8]  <= 1'b1;
    \\u0_tms_reg[6]  <= 1'b1;
    \\u5_timer_reg[7]  <= 1'b1;
    \\u5_timer_reg[6]  <= 1'b1;
    \\u0_sp_tms_reg[16]  <= 1'b1;
    \\u0_csc_reg[10]  <= 1'b0;
    \\u0_csc_reg[5]  <= 1'b0;
    \\u0_csc_reg[4]  <= 1'b0;
    u2_u0_bank0_open_reg <= 1'b0;
    u2_u0_bank1_open_reg <= 1'b0;
    u2_u0_bank3_open_reg <= 1'b0;
    u2_u1_bank0_open_reg <= 1'b0;
    u2_u1_bank1_open_reg <= 1'b0;
    u2_u1_bank2_open_reg <= 1'b0;
    \\u0_csc_reg[6]  <= 1'b0;
    \\u0_csc_reg[7]  <= 1'b0;
    \\u0_csc_reg[9]  <= 1'b0;
    \\u0_sp_csc_reg[10]  <= 1'b0;
    \\u0_sp_csc_reg[4]  <= 1'b0;
    \\u0_sp_csc_reg[7]  <= 1'b0;
    \\u0_sp_csc_reg[9]  <= 1'b0;
    \\u0_sp_csc_reg[6]  <= 1'b0;
    \\u0_sp_csc_reg[3]  <= 1'b0;
    \\u0_sp_csc_reg[2]  <= 1'b0;
    \\u0_csc_reg[11]  <= 1'b0;
    u2_u1_bank3_open_reg <= 1'b0;
    \\u0_sp_csc_reg[5]  <= 1'b0;
    u2_u0_bank2_open_reg <= 1'b0;
    \\u0_sp_csc_reg[1]  <= 1'b0;
    \\u0_csc_reg[1]  <= 1'b0;
    \\u0_csc_reg[3]  <= 1'b0;
    \\u0_csc_reg[2]  <= 1'b0;
    u5_wr_cycle_reg <= 1'b0;
    \\u5_cmd_del_reg[2]  <= 1'b1;
    u5_mc_c_oe_reg <= 1'b0;
    \\u5_cmd_r_reg[2]  <= 1'b1;
    u5_wb_cycle_reg <= 1'b0;
    \\u5_ack_cnt_reg[3]  <= 1'b0;
    \\u5_ack_cnt_reg[1]  <= 1'b0;
    u4_rfr_req_reg <= 1'b0;
    \\u5_ack_cnt_reg[0]  <= 1'b0;
    \\u5_ack_cnt_reg[2]  <= 1'b0;
    u5_mc_adv_r1_reg <= 1'b0;
    u5_tmr2_done_reg <= 1'b0;
    \\u3_u0_wr_adr_reg[1]  <= 1'b0;
    \\u3_u0_wr_adr_reg[3]  <= 1'b0;
    u5_rfr_ack_r_reg <= 1'b0;
    \\u3_u0_wr_adr_reg[0]  <= 1'b1;
    \\u3_u0_wr_adr_reg[2]  <= 1'b0;
    u5_susp_sel_r_reg <= 1'b0;
    u5_dv_r_reg <= 1'b0;
    u0_wp_err_reg <= 1'b0;
    \\u0_cs_reg[0]  <= 1'b0;
    \\u3_u0_rd_adr_reg[3]  <= 1'b0;
    \\u3_u0_rd_adr_reg[0]  <= 1'b1;
    \\u3_u0_rd_adr_reg[2]  <= 1'b0;
    \\u3_u0_rd_adr_reg[1]  <= 1'b0;
    \\u4_rfr_cnt_reg[3]  <= 1'b0;
    \\u4_rfr_cnt_reg[5]  <= 1'b0;
    \\u4_rfr_cnt_reg[6]  <= 1'b0;
    \\u4_rfr_cnt_reg[4]  <= 1'b0;
    u0_u0_init_req_reg <= 1'b0;
    \\u4_rfr_cnt_reg[7]  <= 1'b0;
    \\u4_rfr_cnt_reg[2]  <= 1'b0;
    \\u4_rfr_cnt_reg[1]  <= 1'b0;
    \\u0_cs_reg[1]  <= 1'b0;
    u0_u1_lmr_req_reg <= 1'b0;
    \\u4_rfr_cnt_reg[0]  <= 1'b0;
    u0_u1_init_req_reg <= 1'b0;
    u0_u0_lmr_req_reg <= 1'b0;
    \\u4_ps_cnt_reg[7]  <= 1'b0;
    \\u4_ps_cnt_reg[4]  <= 1'b0;
    u0_u0_init_req_we_reg <= 1'b0;
    \\u4_ps_cnt_reg[3]  <= 1'b0;
    \\u4_ps_cnt_reg[0]  <= 1'b0;
    \\u4_ps_cnt_reg[6]  <= 1'b0;
    \\u4_ps_cnt_reg[1]  <= 1'b0;
    \\u4_ps_cnt_reg[2]  <= 1'b0;
    \\u4_ps_cnt_reg[5]  <= 1'b0;
    \\u0_csc_mask_r_reg[0]  <= 1'b1;
    u0_u1_inited_reg <= 1'b0;
    u0_u0_inited_reg <= 1'b0;
    \\u0_csc_mask_r_reg[1]  <= 1'b1;
    u0_sreq_cs_le_reg <= 1'b0;
    \\u0_csc_mask_r_reg[9]  <= 1'b1;
    \\u0_csc_mask_r_reg[10]  <= 1'b1;
    \\u0_csc_mask_r_reg[2]  <= 1'b1;
    u5_cmd_asserted2_reg <= 1'b0;
    \\u0_csc_mask_r_reg[4]  <= 1'b1;
    \\u0_csc_mask_r_reg[5]  <= 1'b1;
    \\u0_csc_mask_r_reg[6]  <= 1'b1;
    \\u0_csc_mask_r_reg[7]  <= 1'b1;
    \\u0_csc_mask_r_reg[8]  <= 1'b1;
    \\u0_csc_mask_r_reg[3]  <= 1'b1;
    u5_no_wb_cycle_reg <= 1'b0;
    \\u0_csr_r2_reg[6]  <= 1'b0;
    \\u0_csr_r2_reg[4]  <= 1'b0;
    u0_u1_init_req_we_reg <= 1'b0;
    \\u0_csr_r2_reg[0]  <= 1'b0;
    \\u0_csr_r_reg[7]  <= 1'b0;
    \\u0_csr_r2_reg[1]  <= 1'b0;
    \\u0_csr_r2_reg[2]  <= 1'b0;
    \\u0_csr_r_reg[6]  <= 1'b0;
    \\u0_csr_r_reg[9]  <= 1'b0;
    u4_rfr_ce_reg <= 1'b0;
    \\u0_csr_r2_reg[3]  <= 1'b0;
    \\u0_csr_r_reg[1]  <= 1'b0;
    \\u0_csr_r_reg[3]  <= 1'b0;
    \\u0_csr_r_reg[8]  <= 1'b0;
    \\u0_csr_r_reg[2]  <= 1'b0;
    \\u0_csr_r_reg[4]  <= 1'b0;
    \\u0_csr_r2_reg[7]  <= 1'b0;
    \\u0_csr_r_reg[5]  <= 1'b0;
    \\u0_csr_r_reg[10]  <= 1'b0;
    \\u0_csr_r2_reg[5]  <= 1'b0;
    u6_wb_first_r_reg <= 1'b0;
    u4_rfr_early_reg <= 1'b0;
    u0_u1_lmr_req_we_reg <= 1'b0;
    u6_read_go_r1_reg <= 1'b0;
    u6_write_go_r1_reg <= 1'b0;
    u0_u0_lmr_req_we_reg <= 1'b0;
    u0_rf_we_reg <= 1'b0;
    u6_wr_hold_reg <= 1'b0;
    u5_lookup_ready2_reg <= 1'b0;
    u5_tmr_done_reg <= 1'b0;
    u5_suspended_reg <= 1'b0;
    \\u0_spec_req_cs_reg[1]  <= 1'b0;
    u4_rfr_en_reg <= 1'b0;
    u5_lookup_ready1_reg <= 1'b0;
    \\u0_spec_req_cs_reg[0]  <= 1'b0;
    u5_mc_adv_r_reg <= 1'b0;
    u6_rmw_r_reg <= 1'b0;
    u6_write_go_r_reg <= 1'b0;
    u5_mc_le_reg <= 1'b0;
    u0_rst_r3_reg <= 1'b1;
    u6_rmw_en_reg <= 1'b0;
    \\u0_spec_req_cs_reg[5]  <= 1'b0;
    \\u0_cs_reg[6]  <= 1'b0;
    u0_u1_rst_r2_reg <= 1'b1;
    \\u0_spec_req_cs_reg[4]  <= 1'b0;
    u5_rsts_reg <= 1'b1;
    u0_rst_r2_reg <= 1'b1;
    u0_u0_rst_r2_reg <= 1'b1;
    \\u0_cs_reg[7]  <= 1'b0;
    \\u0_cs_reg[4]  <= 1'b0;
    \\u0_spec_req_cs_reg[7]  <= 1'b0;
    \\u0_cs_reg[3]  <= 1'b0;
    \\u0_spec_req_cs_reg[6]  <= 1'b0;
    \\u0_cs_reg[2]  <= 1'b0;
    \\u0_spec_req_cs_reg[3]  <= 1'b0;
    \\u0_cs_reg[5]  <= 1'b0;
    \\u0_spec_req_cs_reg[2]  <= 1'b0;
    u0_init_req_reg <= 1'b0;
    u6_read_go_r_reg <= 1'b0;
    u0_lmr_req_reg <= 1'b0;
    u5_resume_req_r_reg <= 1'b0;
    u5_susp_req_r_reg <= 1'b0;
    u0_rst_r1_reg <= 1'b1;
    u0_u0_rst_r1_reg <= 1'b1;
    u0_u1_rst_r1_reg <= 1'b1;
    u5_rsts1_reg <= 1'b1;
  end
endmodule


