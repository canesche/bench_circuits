// Benchmark "testing" written by ABC on Thu Oct  8 22:16:34 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A39  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A39;
  wire new_n_32_, new_n_33_, new_n_37_, new_n_38_, new_n_39_, new_n_40_,
    new_n_46_, new_n_47_, new_n_48_, new_n_49_, new_n_55_, new_n_56_,
    new_n_57_, new_n_58_, new_n_59_, new_n_60_, new_n_66_, new_n_67_,
    new_n_68_, new_n_69_, new_n_72_, new_n_73_, new_n_74_, new_n_81_,
    new_n_82_, new_n_83_, new_n_84_, new_n_87_, new_n_88_, new_n_91_,
    new_n_94_, new_n_97_, new_n_98_, new_n_99_, new_n_104_, new_n_105_,
    new_n_106_, new_n_107_, new_n_108_, new_n_109_, new_n_114_, new_n_120_,
    new_n_121_, new_n_122_, new_n_123_, new_n_126_, new_n_127_, new_n_128_,
    new_n_129_, new_n_130_, new_n_135_, new_n_136_, new_n_140_, new_n_141_,
    new_n_142_, new_n_143_, new_n_149_, new_n_150_, new_n_151_, new_n_152_,
    new_n_158_, new_n_159_, new_n_160_, new_n_161_, new_n_165_, new_n_168_,
    new_n_171_, new_n_172_, new_n_173_, new_n_178_, new_n_179_, new_n_180_,
    new_n_181_, new_n_182_, new_n_187_, new_n_188_, new_n_189_, new_n_190_,
    new_n_191_, new_n_192_, new_n_193_, new_n_197_, new_n_200_, new_n_203_,
    new_n_204_, new_n_205_, new_n_210_, new_n_211_, new_n_212_, new_n_213_,
    new_n_214_, new_n_219_, new_n_220_, new_n_221_, new_n_222_, new_n_223_,
    new_n_228_, new_n_229_, new_n_233_, new_n_234_, new_n_235_, new_n_236_,
    new_n_242_, new_n_243_, new_n_244_, new_n_245_, new_n_251_, new_n_252_,
    new_n_253_, new_n_254_, new_n_255_, new_n_256_, new_n_262_, new_n_263_,
    new_n_267_, new_n_268_, new_n_269_, new_n_270_, new_n_276_, new_n_277_,
    new_n_278_, new_n_279_, new_n_285_, new_n_286_, new_n_287_, new_n_288_,
    new_n_289_, new_n_290_, new_n_293_, new_n_296_, new_n_299_, new_n_300_,
    new_n_301_, new_n_306_, new_n_307_, new_n_308_, new_n_309_, new_n_310_,
    new_n_311_, new_n_316_, new_n_321_, new_n_322_, new_n_326_, new_n_327_,
    new_n_328_, new_n_329_, new_n_335_, new_n_336_, new_n_337_, new_n_338_,
    new_n_344_, new_n_345_, new_n_346_, new_n_347_, new_n_348_, new_n_349_,
    new_n_350_, new_n_351_, new_n_352_, new_n_353_, new_n_354_, new_n_355_,
    new_n_356_, new_n_357_, new_n_358_;
  assign A39 = ~new_n_358_;
  assign new_n_32_ = ~A202 & A203;
  assign new_n_33_ = A200 & new_n_32_;
  assign new_n_37_ = A202 & ~A203;
  assign new_n_38_ = ~A200 & new_n_37_;
  assign new_n_39_ = new_n_33_ | new_n_38_;
  assign new_n_40_ = ~A199 & new_n_39_;
  assign new_n_46_ = A202 & ~A203;
  assign new_n_47_ = A199 & new_n_46_;
  assign new_n_48_ = A201 | new_n_47_;
  assign new_n_49_ = A200 & new_n_48_;
  assign new_n_55_ = ~A202 & A203;
  assign new_n_56_ = ~A200 & new_n_55_;
  assign new_n_57_ = A201 | new_n_56_;
  assign new_n_58_ = A199 & new_n_57_;
  assign new_n_59_ = new_n_49_ | new_n_58_;
  assign new_n_60_ = new_n_40_ | new_n_59_;
  assign new_n_66_ = A169 | A170;
  assign new_n_67_ = A168 & new_n_66_;
  assign new_n_68_ = ~A167 & new_n_67_;
  assign new_n_69_ = A166 & new_n_68_;
  assign new_n_72_ = ~A166 & A167;
  assign new_n_73_ = new_n_69_ | new_n_72_;
  assign new_n_74_ = new_n_60_ & new_n_73_;
  assign new_n_81_ = ~A169 & ~A170;
  assign new_n_82_ = ~A168 | new_n_81_;
  assign new_n_83_ = ~A166 | new_n_82_;
  assign new_n_84_ = ~A167 & new_n_83_;
  assign new_n_87_ = A166 & A167;
  assign new_n_88_ = new_n_84_ | new_n_87_;
  assign new_n_91_ = A202 | ~A203;
  assign new_n_94_ = ~A199 & A200;
  assign new_n_97_ = A199 & ~A200;
  assign new_n_98_ = new_n_94_ | new_n_97_;
  assign new_n_99_ = new_n_91_ & new_n_98_;
  assign new_n_104_ = ~A202 | A203;
  assign new_n_105_ = A200 & new_n_104_;
  assign new_n_106_ = A199 & new_n_105_;
  assign new_n_107_ = new_n_99_ | new_n_106_;
  assign new_n_108_ = new_n_88_ & new_n_107_;
  assign new_n_109_ = ~A201 & new_n_108_;
  assign new_n_114_ = ~A202 | A203;
  assign new_n_120_ = ~A169 & ~A170;
  assign new_n_121_ = ~A168 | new_n_120_;
  assign new_n_122_ = ~A166 | new_n_121_;
  assign new_n_123_ = ~A167 & new_n_122_;
  assign new_n_126_ = A166 & A167;
  assign new_n_127_ = new_n_123_ | new_n_126_;
  assign new_n_128_ = new_n_114_ & new_n_127_;
  assign new_n_129_ = ~A200 & new_n_128_;
  assign new_n_130_ = ~A199 & new_n_129_;
  assign new_n_135_ = ~A268 & A269;
  assign new_n_136_ = A266 & new_n_135_;
  assign new_n_140_ = A268 & ~A269;
  assign new_n_141_ = ~A266 & new_n_140_;
  assign new_n_142_ = new_n_136_ | new_n_141_;
  assign new_n_143_ = ~A265 & new_n_142_;
  assign new_n_149_ = A268 & ~A269;
  assign new_n_150_ = A265 & new_n_149_;
  assign new_n_151_ = A267 | new_n_150_;
  assign new_n_152_ = A266 & new_n_151_;
  assign new_n_158_ = ~A268 & A269;
  assign new_n_159_ = ~A266 & new_n_158_;
  assign new_n_160_ = A267 | new_n_159_;
  assign new_n_161_ = A265 & new_n_160_;
  assign new_n_165_ = A301 | ~A302;
  assign new_n_168_ = ~A298 & A299;
  assign new_n_171_ = A298 & ~A299;
  assign new_n_172_ = new_n_168_ | new_n_171_;
  assign new_n_173_ = new_n_165_ & new_n_172_;
  assign new_n_178_ = ~A301 | A302;
  assign new_n_179_ = A299 & new_n_178_;
  assign new_n_180_ = A298 & new_n_179_;
  assign new_n_181_ = new_n_173_ | new_n_180_;
  assign new_n_182_ = ~A300 & new_n_181_;
  assign new_n_187_ = ~A301 | A302;
  assign new_n_188_ = ~A299 & new_n_187_;
  assign new_n_189_ = ~A298 & new_n_188_;
  assign new_n_190_ = new_n_182_ | new_n_189_;
  assign new_n_191_ = new_n_161_ | new_n_190_;
  assign new_n_192_ = new_n_152_ | new_n_191_;
  assign new_n_193_ = new_n_143_ | new_n_192_;
  assign new_n_197_ = A235 | ~A236;
  assign new_n_200_ = ~A232 & A233;
  assign new_n_203_ = A232 & ~A233;
  assign new_n_204_ = new_n_200_ | new_n_203_;
  assign new_n_205_ = new_n_197_ & new_n_204_;
  assign new_n_210_ = ~A235 | A236;
  assign new_n_211_ = A233 & new_n_210_;
  assign new_n_212_ = A232 & new_n_211_;
  assign new_n_213_ = new_n_205_ | new_n_212_;
  assign new_n_214_ = ~A234 & new_n_213_;
  assign new_n_219_ = ~A235 | A236;
  assign new_n_220_ = ~A233 & new_n_219_;
  assign new_n_221_ = ~A232 & new_n_220_;
  assign new_n_222_ = new_n_214_ | new_n_221_;
  assign new_n_223_ = new_n_193_ & new_n_222_;
  assign new_n_228_ = ~A301 & A302;
  assign new_n_229_ = A299 & new_n_228_;
  assign new_n_233_ = A301 & ~A302;
  assign new_n_234_ = ~A299 & new_n_233_;
  assign new_n_235_ = new_n_229_ | new_n_234_;
  assign new_n_236_ = ~A298 & new_n_235_;
  assign new_n_242_ = A301 & ~A302;
  assign new_n_243_ = A298 & new_n_242_;
  assign new_n_244_ = A300 | new_n_243_;
  assign new_n_245_ = A299 & new_n_244_;
  assign new_n_251_ = ~A301 & A302;
  assign new_n_252_ = ~A299 & new_n_251_;
  assign new_n_253_ = A300 | new_n_252_;
  assign new_n_254_ = A298 & new_n_253_;
  assign new_n_255_ = new_n_245_ | new_n_254_;
  assign new_n_256_ = new_n_236_ | new_n_255_;
  assign new_n_262_ = ~A235 & A236;
  assign new_n_263_ = A233 & new_n_262_;
  assign new_n_267_ = A235 & ~A236;
  assign new_n_268_ = ~A233 & new_n_267_;
  assign new_n_269_ = new_n_263_ | new_n_268_;
  assign new_n_270_ = ~A232 & new_n_269_;
  assign new_n_276_ = A235 & ~A236;
  assign new_n_277_ = A232 & new_n_276_;
  assign new_n_278_ = A234 | new_n_277_;
  assign new_n_279_ = A233 & new_n_278_;
  assign new_n_285_ = ~A235 & A236;
  assign new_n_286_ = ~A233 & new_n_285_;
  assign new_n_287_ = A234 | new_n_286_;
  assign new_n_288_ = A232 & new_n_287_;
  assign new_n_289_ = new_n_279_ | new_n_288_;
  assign new_n_290_ = new_n_270_ | new_n_289_;
  assign new_n_293_ = A268 | ~A269;
  assign new_n_296_ = ~A265 & A266;
  assign new_n_299_ = A265 & ~A266;
  assign new_n_300_ = new_n_296_ | new_n_299_;
  assign new_n_301_ = new_n_293_ & new_n_300_;
  assign new_n_306_ = ~A268 | A269;
  assign new_n_307_ = A266 & new_n_306_;
  assign new_n_308_ = A265 & new_n_307_;
  assign new_n_309_ = new_n_301_ | new_n_308_;
  assign new_n_310_ = new_n_290_ & new_n_309_;
  assign new_n_311_ = ~A267 & new_n_310_;
  assign new_n_316_ = ~A268 | A269;
  assign new_n_321_ = ~A235 & A236;
  assign new_n_322_ = A233 & new_n_321_;
  assign new_n_326_ = A235 & ~A236;
  assign new_n_327_ = ~A233 & new_n_326_;
  assign new_n_328_ = new_n_322_ | new_n_327_;
  assign new_n_329_ = ~A232 & new_n_328_;
  assign new_n_335_ = A235 & ~A236;
  assign new_n_336_ = A232 & new_n_335_;
  assign new_n_337_ = A234 | new_n_336_;
  assign new_n_338_ = A233 & new_n_337_;
  assign new_n_344_ = ~A235 & A236;
  assign new_n_345_ = ~A233 & new_n_344_;
  assign new_n_346_ = A234 | new_n_345_;
  assign new_n_347_ = A232 & new_n_346_;
  assign new_n_348_ = new_n_338_ | new_n_347_;
  assign new_n_349_ = new_n_329_ | new_n_348_;
  assign new_n_350_ = new_n_316_ & new_n_349_;
  assign new_n_351_ = ~A266 & new_n_350_;
  assign new_n_352_ = ~A265 & new_n_351_;
  assign new_n_353_ = new_n_311_ | new_n_352_;
  assign new_n_354_ = new_n_256_ & new_n_353_;
  assign new_n_355_ = new_n_223_ | new_n_354_;
  assign new_n_356_ = new_n_130_ | new_n_355_;
  assign new_n_357_ = new_n_109_ | new_n_356_;
  assign new_n_358_ = new_n_74_ | new_n_357_;
endmodule


