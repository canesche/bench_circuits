// Benchmark "tv80" written by ABC on Thu Oct  8 22:04:27 2020

module tv80 ( clock, 
    reset_n, clk, wait_n, int_n, nmi_n, busrq_n, \di[0] , \di[1] , \di[2] ,
    \di[3] , \di[4] , \di[5] , \di[6] , \di[7] ,
    m1_n, mreq_n, iorq_n, rd_n, wr_n, rfsh_n, halt_n, busak_n, \A[0] ,
    \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] , \A[9] ,
    \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \do[0] , \do[1] ,
    \do[2] , \do[3] , \do[4] , \do[5] , \do[6] , \do[7]   );
  input  clock;
  input  reset_n, clk, wait_n, int_n, nmi_n, busrq_n, \di[0] , \di[1] ,
    \di[2] , \di[3] , \di[4] , \di[5] , \di[6] , \di[7] ;
  output m1_n, mreq_n, iorq_n, rd_n, wr_n, rfsh_n, halt_n, busak_n, \A[0] ,
    \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] , \A[9] ,
    \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \do[0] , \do[1] ,
    \do[2] , \do[3] , \do[4] , \do[5] , \do[6] , \do[7] ;
  reg i_tv80_core_IncDecZ_reg, \\i_tv80_core_A_reg[1] ,
    \\i_tv80_core_A_reg[2] , \\i_tv80_core_A_reg[5] ,
    \\i_tv80_core_A_reg[6] , \\i_tv80_core_i_reg_RegsH_reg[0][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[0][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][4] ,
    \\i_tv80_core_i_reg_RegsH_reg[0][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][2] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][2] , \\i_tv80_core_A_reg[11] ,
    \\i_tv80_core_A_reg[12] , \\i_tv80_core_A_reg[13] ,
    \\i_tv80_core_A_reg[14] , \\i_tv80_core_A_reg[10] ,
    \\i_tv80_core_A_reg[4] , \\i_tv80_core_A_reg[0] ,
    \\i_tv80_core_A_reg[3] , \\i_tv80_core_A_reg[15] ,
    \\i_tv80_core_A_reg[8] , \\i_tv80_core_A_reg[7] ,
    \\i_tv80_core_A_reg[9] , \\i_tv80_core_i_reg_RegsH_reg[0][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[0][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][5] ,
    \\i_tv80_core_i_reg_RegsH_reg[0][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][3] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][6] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][6] ,
    \\i_tv80_core_i_reg_RegsH_reg[0][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][1] ,
    \\i_tv80_core_i_reg_RegsH_reg[4][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][7] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][7] ,
    \\i_tv80_core_i_reg_RegsH_reg[0][0] ,
    \\i_tv80_core_i_reg_RegsH_reg[1][0] ,
    \\i_tv80_core_i_reg_RegsH_reg[2][0] ,
    \\i_tv80_core_i_reg_RegsH_reg[3][0] ,
    \\i_tv80_core_i_reg_RegsH_reg[5][0] ,
    \\i_tv80_core_i_reg_RegsH_reg[6][0] ,
    \\i_tv80_core_i_reg_RegsH_reg[7][0] , \\i_tv80_core_tstate_reg[0] ,
    \\i_tv80_core_tstate_reg[1] , \\i_tv80_core_tstate_reg[2] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][5] , \\i_tv80_core_F_reg[2] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][5] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][4] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][4] , \\i_tv80_core_SP_reg[14] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][3] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][3] , \\i_tv80_core_ACC_reg[0] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][1] , \\i_tv80_core_do_reg[5] ,
    \\i_tv80_core_F_reg[1] , \\i_tv80_core_SP_reg[1] ,
    \\i_tv80_core_F_reg[6] , \\i_tv80_core_F_reg[0] ,
    \\i_tv80_core_ACC_reg[7] , \\i_tv80_core_do_reg[7] ,
    \\i_tv80_core_SP_reg[7] , \\i_tv80_core_do_reg[6] ,
    \\i_tv80_core_SP_reg[6] , \\i_tv80_core_ACC_reg[3] ,
    \\i_tv80_core_ACC_reg[5] , \\i_tv80_core_ACC_reg[6] ,
    \\i_tv80_core_ACC_reg[2] , \\i_tv80_core_ACC_reg[1] ,
    \\i_tv80_core_ACC_reg[4] , \\i_tv80_core_SP_reg[5] ,
    \\i_tv80_core_do_reg[4] , \\i_tv80_core_SP_reg[4] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[0][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][1] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][1] , \\i_tv80_core_do_reg[0] ,
    \\i_tv80_core_do_reg[1] , \\i_tv80_core_do_reg[2] ,
    \\i_tv80_core_do_reg[3] , \\i_tv80_core_i_reg_RegsL_reg[0][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[1][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[2][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[3][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[5][0] ,
    \\i_tv80_core_i_reg_RegsL_reg[7][0] , \\i_tv80_core_SP_reg[2] ,
    \\i_tv80_core_SP_reg[3] , \\i_tv80_core_SP_reg[0] ,
    \\i_tv80_core_i_reg_RegsL_reg[4][2] ,
    \\i_tv80_core_i_reg_RegsL_reg[6][0] , \\i_tv80_core_SP_reg[12] ,
    \\i_tv80_core_F_reg[7] , \\i_tv80_core_SP_reg[15] ,
    \\i_tv80_core_F_reg[3] , \\i_tv80_core_F_reg[5] ,
    \\i_tv80_core_SP_reg[10] , \\i_tv80_core_SP_reg[13] ,
    \\i_tv80_core_F_reg[4] , \\i_tv80_core_SP_reg[9] ,
    \\i_tv80_core_SP_reg[11] , \\i_tv80_core_SP_reg[8] ,
    \\i_tv80_core_mcycle_reg[1] , \\i_tv80_core_mcycle_reg[2] ,
    \\i_tv80_core_mcycle_reg[0] , \\i_tv80_core_TmpAddr_reg[14] ,
    i_tv80_core_IntE_FF1_reg, i_tv80_core_IntE_FF2_reg,
    i_tv80_core_m1_n_reg, i_tv80_core_IntCycle_reg,
    i_tv80_core_NMICycle_reg, \\i_tv80_core_BusA_reg[0] ,
    \\i_tv80_core_BusA_reg[5] , \\i_tv80_core_PC_reg[9] ,
    \\i_tv80_core_PC_reg[7] , \\i_tv80_core_Pre_XY_F_M_reg[2] ,
    \\i_tv80_core_BusA_reg[3] , \\i_tv80_core_PC_reg[11] ,
    \\i_tv80_core_PC_reg[12] , \\i_tv80_core_PC_reg[13] ,
    \\i_tv80_core_PC_reg[1] , \\i_tv80_core_PC_reg[2] ,
    \\i_tv80_core_PC_reg[3] , \\i_tv80_core_PC_reg[4] ,
    \\i_tv80_core_PC_reg[5] , \\i_tv80_core_PC_reg[6] ,
    \\i_tv80_core_PC_reg[8] , \\i_tv80_core_Pre_XY_F_M_reg[0] ,
    \\i_tv80_core_Pre_XY_F_M_reg[1] , \\i_tv80_core_BusA_reg[2] ,
    \\i_tv80_core_BusA_reg[4] , \\i_tv80_core_BusA_reg[6] ,
    \\i_tv80_core_PC_reg[15] , \\i_tv80_core_PC_reg[14] ,
    \\i_tv80_core_PC_reg[0] , \\i_tv80_core_PC_reg[10] ,
    \\i_tv80_core_TmpAddr_reg[10] , \\i_tv80_core_BusA_reg[7] ,
    \\i_tv80_core_TmpAddr_reg[15] , \\i_tv80_core_BusA_reg[1] ,
    \\i_tv80_core_TmpAddr_reg[12] , \\i_tv80_core_TmpAddr_reg[13] ,
    i_tv80_core_BTR_r_reg, \\i_tv80_core_TmpAddr_reg[11] ,
    i_tv80_core_Halt_FF_reg, \\i_tv80_core_Read_To_Reg_r_reg[4] ,
    \\i_tv80_core_TmpAddr_reg[9] , \\i_tv80_core_TmpAddr_reg[6] ,
    \\i_tv80_core_Read_To_Reg_r_reg[2] , \\i_tv80_core_RegBusA_r_reg[0] ,
    \\i_tv80_core_RegBusA_r_reg[13] , i_tv80_core_Auto_Wait_t2_reg,
    \\i_tv80_core_TmpAddr_reg[8] , \\i_tv80_core_Read_To_Reg_r_reg[0] ,
    \\i_tv80_core_Read_To_Reg_r_reg[1] , \\i_tv80_core_ALU_Op_r_reg[1] ,
    i_tv80_core_Save_ALU_r_reg, \\i_tv80_core_ALU_Op_r_reg[3] ,
    \\i_tv80_core_TmpAddr_reg[7] , \\i_tv80_core_RegBusA_r_reg[11] ,
    \\i_tv80_core_TmpAddr_reg[5] , i_tv80_core_BusAck_reg,
    \\i_tv80_core_RegBusA_r_reg[10] , \\i_tv80_core_RegBusA_r_reg[12] ,
    \\i_tv80_core_RegBusA_r_reg[14] , \\i_tv80_core_Read_To_Reg_r_reg[3] ,
    i_tv80_core_Auto_Wait_t1_reg, \\i_tv80_core_RegBusA_r_reg[15] ,
    \\i_tv80_core_RegBusA_r_reg[7] , \\i_tv80_core_RegBusA_r_reg[9] ,
    \\i_tv80_core_ALU_Op_r_reg[2] , \\i_tv80_core_ALU_Op_r_reg[0] ,
    \\i_tv80_core_RegBusA_r_reg[8] , \\i_tv80_core_TmpAddr_reg[4] ,
    \\i_tv80_core_RegBusA_r_reg[1] , \\i_tv80_core_RegBusA_r_reg[2] ,
    \\i_tv80_core_RegBusA_r_reg[5] , \\i_tv80_core_RegBusA_r_reg[6] ,
    \\i_tv80_core_BusB_reg[0] , \\i_tv80_core_TmpAddr_reg[3] ,
    \\i_tv80_core_RegBusA_r_reg[4] , \\i_tv80_core_RegBusA_r_reg[3] ,
    \\i_tv80_core_TmpAddr_reg[2] , \\i_tv80_core_BusB_reg[6] ,
    \\i_tv80_core_BusB_reg[4] , \\i_tv80_core_BusB_reg[1] ,
    \\i_tv80_core_BusB_reg[3] , \\i_tv80_core_BusB_reg[5] ,
    \\i_tv80_core_BusB_reg[2] , \\i_tv80_core_BusB_reg[7] ,
    \\i_tv80_core_TmpAddr_reg[1] , \\i_tv80_core_RegAddrC_reg[1] ,
    i_tv80_core_Z16_r_reg, iorq_n_reg, \\i_tv80_core_RegAddrB_r_reg[2] ,
    mreq_n_reg, \\i_tv80_core_TmpAddr_reg[0] ,
    \\i_tv80_core_RegAddrB_r_reg[0] , \\i_tv80_core_RegAddrB_r_reg[1] ,
    \\i_tv80_core_RegAddrC_reg[0] , \\i_tv80_core_R_reg[6] ,
    \\i_tv80_core_R_reg[5] , \\i_tv80_core_R_reg[3] ,
    \\i_tv80_core_R_reg[2] , \\i_tv80_core_R_reg[4] ,
    \\i_tv80_core_IR_reg[2] , \\i_tv80_core_R_reg[0] , rd_n_reg,
    \\i_tv80_core_ISet_reg[0] , \\i_tv80_core_R_reg[1] ,
    \\i_tv80_core_IR_reg[0] , \\i_tv80_core_IR_reg[1] ,
    \\i_tv80_core_IR_reg[5] , \\i_tv80_core_IR_reg[6] ,
    \\i_tv80_core_IR_reg[7] , \\i_tv80_core_ISet_reg[1] ,
    \\i_tv80_core_IR_reg[4] , \\i_tv80_core_IR_reg[3] ,
    i_tv80_core_Alternate_reg, i_tv80_core_XY_Ind_reg, wr_n_reg,
    \\i_tv80_core_mcycles_reg[0] , \\i_tv80_core_mcycles_reg[2] ,
    \\i_tv80_core_RegAddrA_r_reg[1] , \\i_tv80_core_mcycles_reg[1] ,
    \\i_tv80_core_RegAddrA_r_reg[2] , \\i_tv80_core_RegAddrA_r_reg[0] ,
    \\i_tv80_core_XY_State_reg[0] , \\i_tv80_core_XY_State_reg[1] ,
    \\i_tv80_core_Fp_reg[5] , \\i_tv80_core_Ap_reg[3] ,
    \\i_tv80_core_Ap_reg[5] , \\i_tv80_core_Fp_reg[7] ,
    \\i_tv80_core_Ap_reg[1] , \\i_tv80_core_Fp_reg[1] ,
    \\i_tv80_core_Fp_reg[3] , \\i_tv80_core_Fp_reg[0] ,
    \\i_tv80_core_Fp_reg[2] , \\i_tv80_core_Fp_reg[4] ,
    \\i_tv80_core_Fp_reg[6] , \\i_tv80_core_Ap_reg[0] ,
    \\i_tv80_core_Ap_reg[2] , \\i_tv80_core_Ap_reg[4] ,
    \\i_tv80_core_Ap_reg[6] , \\i_tv80_core_Ap_reg[7] ,
    \\i_tv80_core_IStatus_reg[1] , \\i_tv80_core_R_reg[7] ,
    \\i_tv80_core_IStatus_reg[0] , i_tv80_core_rfsh_n_reg,
    i_tv80_core_PreserveC_r_reg, \\i_tv80_core_I_reg[5] ,
    \\i_tv80_core_I_reg[2] , \\i_tv80_core_I_reg[4] ,
    \\i_tv80_core_I_reg[7] , \\i_tv80_core_I_reg[6] ,
    \\i_tv80_core_I_reg[0] , \\i_tv80_core_I_reg[1] ,
    \\i_tv80_core_I_reg[3] , i_tv80_core_Arith16_r_reg,
    i_tv80_core_No_BTR_reg, \\i_tv80_core_RegAddrC_reg[2] ,
    \\di_reg_reg[6] , \\di_reg_reg[3] , \\di_reg_reg[1] , \\di_reg_reg[7] ,
    \\di_reg_reg[2] , \\di_reg_reg[4] , \\di_reg_reg[5] , \\di_reg_reg[0] ,
    i_tv80_core_NMI_s_reg, i_tv80_core_BusReq_s_reg,
    i_tv80_core_Oldnmi_n_reg, i_tv80_core_INT_s_reg;
  wire \new_[407]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[464]_ , \new_[465]_ , \new_[466]_ , \new_[467]_ , \new_[468]_ ,
    \new_[469]_ , \new_[470]_ , \new_[471]_ , \new_[497]_ , \new_[498]_ ,
    \new_[499]_ , \new_[500]_ , \new_[501]_ , \new_[502]_ , \new_[503]_ ,
    \new_[504]_ , \new_[505]_ , \new_[506]_ , \new_[507]_ , \new_[508]_ ,
    \new_[509]_ , \new_[510]_ , \new_[511]_ , \new_[512]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ , \new_[571]_ ,
    \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ , \new_[576]_ ,
    \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[616]_ , \new_[617]_ , \new_[618]_ ,
    \new_[619]_ , \new_[620]_ , \new_[621]_ , \new_[622]_ , \new_[623]_ ,
    \new_[624]_ , \new_[625]_ , \new_[626]_ , \new_[627]_ , \new_[631]_ ,
    \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ , \new_[636]_ ,
    \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ , \new_[641]_ ,
    \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ , \new_[646]_ ,
    \new_[650]_ , \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ ,
    \new_[655]_ , \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ ,
    \new_[660]_ , \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ ,
    \new_[665]_ , \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ ,
    \new_[670]_ , \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ ,
    \new_[675]_ , \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ ,
    \new_[680]_ , \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ ,
    \new_[685]_ , \new_[686]_ , \new_[695]_ , \new_[696]_ , \new_[697]_ ,
    \new_[698]_ , \new_[699]_ , \new_[700]_ , \new_[701]_ , \new_[702]_ ,
    \new_[703]_ , \new_[704]_ , \new_[705]_ , \new_[709]_ , \new_[710]_ ,
    \new_[715]_ , \new_[716]_ , \new_[717]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ , \new_[731]_ ,
    \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ , \new_[736]_ ,
    \new_[737]_ , \new_[740]_ , \new_[741]_ , \new_[742]_ , \new_[743]_ ,
    \new_[744]_ , \new_[745]_ , \new_[746]_ , \new_[747]_ , \new_[748]_ ,
    \new_[749]_ , \new_[750]_ , \new_[751]_ , \new_[752]_ , \new_[753]_ ,
    \new_[755]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[766]_ ,
    \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ , \new_[771]_ ,
    \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ , \new_[776]_ ,
    \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[832]_ , \new_[833]_ ,
    \new_[834]_ , \new_[835]_ , \new_[836]_ , \new_[837]_ , \new_[838]_ ,
    \new_[839]_ , \new_[840]_ , \new_[841]_ , \new_[842]_ , \new_[843]_ ,
    \new_[844]_ , \new_[845]_ , \new_[846]_ , \new_[847]_ , \new_[848]_ ,
    \new_[849]_ , \new_[850]_ , \new_[851]_ , \new_[852]_ , \new_[853]_ ,
    \new_[854]_ , \new_[886]_ , \new_[887]_ , \new_[896]_ , \new_[898]_ ,
    \new_[899]_ , \new_[902]_ , \new_[904]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[921]_ , \new_[925]_ , \new_[926]_ ,
    \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ , \new_[931]_ ,
    \new_[932]_ , \new_[937]_ , \new_[939]_ , \new_[940]_ , \new_[941]_ ,
    \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ , \new_[946]_ ,
    \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ , \new_[951]_ ,
    \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ , \new_[956]_ ,
    \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ , \new_[961]_ ,
    \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ , \new_[966]_ ,
    \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ , \new_[971]_ ,
    \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ , \new_[976]_ ,
    \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ , \new_[981]_ ,
    \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ , \new_[986]_ ,
    \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ , \new_[991]_ ,
    \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ , \new_[996]_ ,
    \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ , \new_[1001]_ ,
    \new_[1002]_ , \new_[1003]_ , \new_[1004]_ , \new_[1005]_ ,
    \new_[1006]_ , \new_[1007]_ , \new_[1008]_ , \new_[1009]_ ,
    \new_[1010]_ , \new_[1011]_ , \new_[1012]_ , \new_[1013]_ ,
    \new_[1014]_ , \new_[1015]_ , \new_[1016]_ , \new_[1017]_ ,
    \new_[1018]_ , \new_[1019]_ , \new_[1020]_ , \new_[1021]_ ,
    \new_[1022]_ , \new_[1023]_ , \new_[1024]_ , \new_[1025]_ ,
    \new_[1026]_ , \new_[1027]_ , \new_[1028]_ , \new_[1029]_ ,
    \new_[1030]_ , \new_[1031]_ , \new_[1032]_ , \new_[1033]_ ,
    \new_[1034]_ , \new_[1035]_ , \new_[1036]_ , \new_[1037]_ ,
    \new_[1038]_ , \new_[1039]_ , \new_[1040]_ , \new_[1041]_ ,
    \new_[1042]_ , \new_[1043]_ , \new_[1044]_ , \new_[1045]_ ,
    \new_[1046]_ , \new_[1047]_ , \new_[1048]_ , \new_[1049]_ ,
    \new_[1050]_ , \new_[1051]_ , \new_[1052]_ , \new_[1053]_ ,
    \new_[1054]_ , \new_[1055]_ , \new_[1056]_ , \new_[1057]_ ,
    \new_[1058]_ , \new_[1059]_ , \new_[1060]_ , \new_[1061]_ ,
    \new_[1062]_ , \new_[1063]_ , \new_[1064]_ , \new_[1065]_ ,
    \new_[1066]_ , \new_[1067]_ , \new_[1068]_ , \new_[1069]_ ,
    \new_[1070]_ , \new_[1071]_ , \new_[1072]_ , \new_[1073]_ ,
    \new_[1074]_ , \new_[1075]_ , \new_[1076]_ , \new_[1077]_ ,
    \new_[1078]_ , \new_[1079]_ , \new_[1080]_ , \new_[1081]_ ,
    \new_[1082]_ , \new_[1083]_ , \new_[1084]_ , \new_[1085]_ ,
    \new_[1086]_ , \new_[1087]_ , \new_[1088]_ , \new_[1089]_ ,
    \new_[1090]_ , \new_[1091]_ , \new_[1092]_ , \new_[1093]_ ,
    \new_[1094]_ , \new_[1095]_ , \new_[1096]_ , \new_[1097]_ ,
    \new_[1098]_ , \new_[1099]_ , \new_[1100]_ , \new_[1101]_ ,
    \new_[1102]_ , \new_[1103]_ , \new_[1104]_ , \new_[1105]_ ,
    \new_[1106]_ , \new_[1107]_ , \new_[1108]_ , \new_[1109]_ ,
    \new_[1110]_ , \new_[1111]_ , \new_[1112]_ , \new_[1113]_ ,
    \new_[1114]_ , \new_[1116]_ , \new_[1117]_ , \new_[1118]_ ,
    \new_[1119]_ , \new_[1123]_ , \new_[1124]_ , \new_[1125]_ ,
    \new_[1126]_ , \new_[1127]_ , \new_[1128]_ , \new_[1129]_ ,
    \new_[1130]_ , \new_[1131]_ , \new_[1132]_ , \new_[1133]_ ,
    \new_[1134]_ , \new_[1135]_ , \new_[1136]_ , \new_[1137]_ ,
    \new_[1138]_ , \new_[1139]_ , \new_[1140]_ , \new_[1141]_ ,
    \new_[1142]_ , \new_[1143]_ , \new_[1144]_ , \new_[1145]_ ,
    \new_[1146]_ , \new_[1147]_ , \new_[1148]_ , \new_[1149]_ ,
    \new_[1150]_ , \new_[1151]_ , \new_[1152]_ , \new_[1153]_ ,
    \new_[1154]_ , \new_[1155]_ , \new_[1156]_ , \new_[1157]_ ,
    \new_[1158]_ , \new_[1160]_ , \new_[1161]_ , \new_[1162]_ ,
    \new_[1163]_ , \new_[1164]_ , \new_[1165]_ , \new_[1166]_ ,
    \new_[1167]_ , \new_[1168]_ , \new_[1169]_ , \new_[1170]_ ,
    \new_[1171]_ , \new_[1172]_ , \new_[1173]_ , \new_[1174]_ ,
    \new_[1175]_ , \new_[1176]_ , \new_[1177]_ , \new_[1178]_ ,
    \new_[1179]_ , \new_[1180]_ , \new_[1181]_ , \new_[1182]_ ,
    \new_[1183]_ , \new_[1184]_ , \new_[1185]_ , \new_[1186]_ ,
    \new_[1187]_ , \new_[1188]_ , \new_[1189]_ , \new_[1190]_ ,
    \new_[1191]_ , \new_[1192]_ , \new_[1193]_ , \new_[1194]_ ,
    \new_[1195]_ , \new_[1196]_ , \new_[1197]_ , \new_[1198]_ ,
    \new_[1199]_ , \new_[1200]_ , \new_[1201]_ , \new_[1202]_ ,
    \new_[1203]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1218]_ ,
    \new_[1219]_ , \new_[1220]_ , \new_[1221]_ , \new_[1222]_ ,
    \new_[1223]_ , \new_[1224]_ , \new_[1225]_ , \new_[1226]_ ,
    \new_[1227]_ , \new_[1228]_ , \new_[1229]_ , \new_[1230]_ ,
    \new_[1231]_ , \new_[1233]_ , \new_[1234]_ , \new_[1235]_ ,
    \new_[1236]_ , \new_[1237]_ , \new_[1238]_ , \new_[1239]_ ,
    \new_[1240]_ , \new_[1241]_ , \new_[1242]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1254]_ , \new_[1255]_ , \new_[1256]_ , \new_[1257]_ ,
    \new_[1258]_ , \new_[1259]_ , \new_[1260]_ , \new_[1261]_ ,
    \new_[1262]_ , \new_[1263]_ , \new_[1264]_ , \new_[1265]_ ,
    \new_[1266]_ , \new_[1267]_ , \new_[1268]_ , \new_[1269]_ ,
    \new_[1270]_ , \new_[1271]_ , \new_[1272]_ , \new_[1273]_ ,
    \new_[1274]_ , \new_[1275]_ , \new_[1276]_ , \new_[1277]_ ,
    \new_[1278]_ , \new_[1279]_ , \new_[1280]_ , \new_[1281]_ ,
    \new_[1282]_ , \new_[1283]_ , \new_[1284]_ , \new_[1285]_ ,
    \new_[1286]_ , \new_[1287]_ , \new_[1288]_ , \new_[1289]_ ,
    \new_[1290]_ , \new_[1291]_ , \new_[1292]_ , \new_[1293]_ ,
    \new_[1294]_ , \new_[1295]_ , \new_[1296]_ , \new_[1297]_ ,
    \new_[1298]_ , \new_[1299]_ , \new_[1300]_ , \new_[1301]_ ,
    \new_[1302]_ , \new_[1303]_ , \new_[1304]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1396]_ , \new_[1399]_ ,
    \new_[1400]_ , \new_[1401]_ , \new_[1402]_ , \new_[1403]_ ,
    \new_[1404]_ , \new_[1405]_ , \new_[1406]_ , \new_[1407]_ ,
    \new_[1408]_ , \new_[1409]_ , \new_[1410]_ , \new_[1411]_ ,
    \new_[1412]_ , \new_[1413]_ , \new_[1414]_ , \new_[1415]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1433]_ ,
    \new_[1434]_ , \new_[1435]_ , \new_[1436]_ , \new_[1437]_ ,
    \new_[1438]_ , \new_[1439]_ , \new_[1440]_ , \new_[1441]_ ,
    \new_[1442]_ , \new_[1443]_ , \new_[1444]_ , \new_[1445]_ ,
    \new_[1446]_ , \new_[1447]_ , \new_[1448]_ , \new_[1449]_ ,
    \new_[1450]_ , \new_[1451]_ , \new_[1452]_ , \new_[1453]_ ,
    \new_[1455]_ , \new_[1456]_ , \new_[1457]_ , \new_[1458]_ ,
    \new_[1459]_ , \new_[1460]_ , \new_[1461]_ , \new_[1462]_ ,
    \new_[1463]_ , \new_[1465]_ , \new_[1466]_ , \new_[1467]_ ,
    \new_[1468]_ , \new_[1469]_ , \new_[1470]_ , \new_[1471]_ ,
    \new_[1472]_ , \new_[1473]_ , \new_[1474]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1532]_ , \new_[1533]_ ,
    \new_[1534]_ , \new_[1535]_ , \new_[1536]_ , \new_[1537]_ ,
    \new_[1538]_ , \new_[1540]_ , \new_[1541]_ , \new_[1542]_ ,
    \new_[1543]_ , \new_[1544]_ , \new_[1545]_ , \new_[1546]_ ,
    \new_[1547]_ , \new_[1548]_ , \new_[1549]_ , \new_[1550]_ ,
    \new_[1551]_ , \new_[1552]_ , \new_[1553]_ , \new_[1554]_ ,
    \new_[1555]_ , \new_[1556]_ , \new_[1557]_ , \new_[1558]_ ,
    \new_[1559]_ , \new_[1560]_ , \new_[1561]_ , \new_[1562]_ ,
    \new_[1563]_ , \new_[1564]_ , \new_[1565]_ , \new_[1566]_ ,
    \new_[1567]_ , \new_[1568]_ , \new_[1569]_ , \new_[1570]_ ,
    \new_[1571]_ , \new_[1572]_ , \new_[1573]_ , \new_[1574]_ ,
    \new_[1575]_ , \new_[1576]_ , \new_[1577]_ , \new_[1578]_ ,
    \new_[1579]_ , \new_[1580]_ , \new_[1581]_ , \new_[1583]_ ,
    \new_[1584]_ , \new_[1585]_ , \new_[1586]_ , \new_[1587]_ ,
    \new_[1588]_ , \new_[1589]_ , \new_[1590]_ , \new_[1591]_ ,
    \new_[1592]_ , \new_[1593]_ , \new_[1594]_ , \new_[1595]_ ,
    \new_[1596]_ , \new_[1597]_ , \new_[1598]_ , \new_[1599]_ ,
    \new_[1600]_ , \new_[1601]_ , \new_[1602]_ , \new_[1603]_ ,
    \new_[1604]_ , \new_[1605]_ , \new_[1606]_ , \new_[1607]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1639]_ , \new_[1640]_ , \new_[1641]_ ,
    \new_[1642]_ , \new_[1643]_ , \new_[1646]_ , \new_[1647]_ ,
    \new_[1648]_ , \new_[1649]_ , \new_[1650]_ , \new_[1651]_ ,
    \new_[1652]_ , \new_[1653]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1703]_ , \new_[1704]_ , \new_[1705]_ ,
    \new_[1706]_ , \new_[1707]_ , \new_[1708]_ , \new_[1709]_ ,
    \new_[1710]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1724]_ , \new_[1725]_ ,
    \new_[1726]_ , \new_[1727]_ , \new_[1728]_ , \new_[1729]_ ,
    \new_[1730]_ , \new_[1731]_ , \new_[1732]_ , \new_[1733]_ ,
    \new_[1734]_ , \new_[1735]_ , \new_[1736]_ , \new_[1737]_ ,
    \new_[1738]_ , \new_[1739]_ , \new_[1740]_ , \new_[1741]_ ,
    \new_[1742]_ , \new_[1743]_ , \new_[1744]_ , \new_[1745]_ ,
    \new_[1746]_ , \new_[1747]_ , \new_[1748]_ , \new_[1749]_ ,
    \new_[1751]_ , \new_[1753]_ , \new_[1754]_ , \new_[1755]_ ,
    \new_[1756]_ , \new_[1757]_ , \new_[1758]_ , \new_[1759]_ ,
    \new_[1760]_ , \new_[1761]_ , \new_[1762]_ , \new_[1763]_ ,
    \new_[1764]_ , \new_[1765]_ , \new_[1770]_ , \new_[1771]_ ,
    \new_[1772]_ , \new_[1773]_ , \new_[1774]_ , \new_[1775]_ ,
    \new_[1776]_ , \new_[1777]_ , \new_[1778]_ , \new_[1779]_ ,
    \new_[1780]_ , \new_[1781]_ , \new_[1784]_ , \new_[1785]_ ,
    \new_[1786]_ , \new_[1787]_ , \new_[1788]_ , \new_[1789]_ ,
    \new_[1790]_ , \new_[1791]_ , \new_[1792]_ , \new_[1793]_ ,
    \new_[1794]_ , \new_[1795]_ , \new_[1796]_ , \new_[1797]_ ,
    \new_[1798]_ , \new_[1799]_ , \new_[1800]_ , \new_[1801]_ ,
    \new_[1802]_ , \new_[1803]_ , \new_[1804]_ , \new_[1805]_ ,
    \new_[1806]_ , \new_[1807]_ , \new_[1808]_ , \new_[1809]_ ,
    \new_[1810]_ , \new_[1811]_ , \new_[1812]_ , \new_[1813]_ ,
    \new_[1814]_ , \new_[1815]_ , \new_[1816]_ , \new_[1817]_ ,
    \new_[1818]_ , \new_[1819]_ , \new_[1820]_ , \new_[1821]_ ,
    \new_[1822]_ , \new_[1824]_ , \new_[1825]_ , \new_[1826]_ ,
    \new_[1827]_ , \new_[1828]_ , \new_[1829]_ , \new_[1830]_ ,
    \new_[1831]_ , \new_[1833]_ , \new_[1834]_ , \new_[1835]_ ,
    \new_[1836]_ , \new_[1837]_ , \new_[1838]_ , \new_[1839]_ ,
    \new_[1840]_ , \new_[1841]_ , \new_[1842]_ , \new_[1843]_ ,
    \new_[1844]_ , \new_[1845]_ , \new_[1846]_ , \new_[1847]_ ,
    \new_[1848]_ , \new_[1849]_ , \new_[1850]_ , \new_[1851]_ ,
    \new_[1852]_ , \new_[1853]_ , \new_[1854]_ , \new_[1855]_ ,
    \new_[1856]_ , \new_[1857]_ , \new_[1858]_ , \new_[1859]_ ,
    \new_[1860]_ , \new_[1861]_ , \new_[1862]_ , \new_[1863]_ ,
    \new_[1864]_ , \new_[1865]_ , \new_[1866]_ , \new_[1867]_ ,
    \new_[1868]_ , \new_[1869]_ , \new_[1870]_ , \new_[1871]_ ,
    \new_[1872]_ , \new_[1873]_ , \new_[1874]_ , \new_[1875]_ ,
    \new_[1876]_ , \new_[1877]_ , \new_[1878]_ , \new_[1879]_ ,
    \new_[1880]_ , \new_[1884]_ , \new_[1885]_ , \new_[1886]_ ,
    \new_[1887]_ , \new_[1888]_ , \new_[1889]_ , \new_[1892]_ ,
    \new_[1894]_ , \new_[1895]_ , \new_[1896]_ , \new_[1897]_ ,
    \new_[1898]_ , \new_[1899]_ , \new_[1900]_ , \new_[1901]_ ,
    \new_[1902]_ , \new_[1903]_ , \new_[1904]_ , \new_[1905]_ ,
    \new_[1906]_ , \new_[1907]_ , \new_[1908]_ , \new_[1909]_ ,
    \new_[1910]_ , \new_[1911]_ , \new_[1912]_ , \new_[1913]_ ,
    \new_[1914]_ , \new_[1915]_ , \new_[1916]_ , \new_[1917]_ ,
    \new_[1918]_ , \new_[1919]_ , \new_[1925]_ , \new_[1926]_ ,
    \new_[1927]_ , \new_[1928]_ , \new_[1929]_ , \new_[1930]_ ,
    \new_[1931]_ , \new_[1932]_ , \new_[1933]_ , \new_[1934]_ ,
    \new_[1935]_ , \new_[1936]_ , \new_[1937]_ , \new_[1938]_ ,
    \new_[1939]_ , \new_[1940]_ , \new_[1941]_ , \new_[1942]_ ,
    \new_[1943]_ , \new_[1944]_ , \new_[1945]_ , \new_[1947]_ ,
    \new_[1948]_ , \new_[1949]_ , \new_[1950]_ , \new_[1951]_ ,
    \new_[1952]_ , \new_[1953]_ , \new_[1954]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1986]_ ,
    \new_[1987]_ , \new_[1988]_ , \new_[1989]_ , \new_[1990]_ ,
    \new_[1991]_ , \new_[1992]_ , \new_[1993]_ , \new_[1994]_ ,
    \new_[1995]_ , \new_[1996]_ , \new_[1997]_ , \new_[1998]_ ,
    \new_[1999]_ , \new_[2000]_ , \new_[2001]_ , \new_[2002]_ ,
    \new_[2003]_ , \new_[2004]_ , \new_[2005]_ , \new_[2006]_ ,
    \new_[2007]_ , \new_[2009]_ , \new_[2010]_ , \new_[2011]_ ,
    \new_[2012]_ , \new_[2013]_ , \new_[2014]_ , \new_[2015]_ ,
    \new_[2016]_ , \new_[2017]_ , \new_[2018]_ , \new_[2019]_ ,
    \new_[2020]_ , \new_[2021]_ , \new_[2022]_ , \new_[2023]_ ,
    \new_[2024]_ , \new_[2025]_ , \new_[2026]_ , \new_[2027]_ ,
    \new_[2028]_ , \new_[2029]_ , \new_[2030]_ , \new_[2031]_ ,
    \new_[2032]_ , \new_[2033]_ , \new_[2034]_ , \new_[2035]_ ,
    \new_[2036]_ , \new_[2037]_ , \new_[2038]_ , \new_[2039]_ ,
    \new_[2040]_ , \new_[2041]_ , \new_[2042]_ , \new_[2043]_ ,
    \new_[2044]_ , \new_[2045]_ , \new_[2046]_ , \new_[2047]_ ,
    \new_[2048]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2076]_ , \new_[2077]_ , \new_[2078]_ , \new_[2079]_ ,
    \new_[2080]_ , \new_[2081]_ , \new_[2082]_ , \new_[2083]_ ,
    \new_[2084]_ , \new_[2085]_ , \new_[2086]_ , \new_[2087]_ ,
    \new_[2088]_ , \new_[2089]_ , \new_[2090]_ , \new_[2091]_ ,
    \new_[2092]_ , \new_[2093]_ , \new_[2094]_ , \new_[2095]_ ,
    \new_[2096]_ , \new_[2097]_ , \new_[2098]_ , \new_[2099]_ ,
    \new_[2100]_ , \new_[2101]_ , \new_[2102]_ , \new_[2103]_ ,
    \new_[2104]_ , \new_[2105]_ , \new_[2106]_ , \new_[2107]_ ,
    \new_[2108]_ , \new_[2109]_ , \new_[2110]_ , \new_[2111]_ ,
    \new_[2112]_ , \new_[2113]_ , \new_[2114]_ , \new_[2115]_ ,
    \new_[2116]_ , \new_[2117]_ , \new_[2118]_ , \new_[2119]_ ,
    \new_[2120]_ , \new_[2121]_ , \new_[2122]_ , \new_[2123]_ ,
    \new_[2124]_ , \new_[2125]_ , \new_[2126]_ , \new_[2127]_ ,
    \new_[2128]_ , \new_[2129]_ , \new_[2130]_ , \new_[2131]_ ,
    \new_[2132]_ , \new_[2133]_ , \new_[2134]_ , \new_[2135]_ ,
    \new_[2136]_ , \new_[2137]_ , \new_[2138]_ , \new_[2139]_ ,
    \new_[2140]_ , \new_[2141]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2168]_ , \new_[2169]_ ,
    \new_[2170]_ , \new_[2171]_ , \new_[2172]_ , \new_[2173]_ ,
    \new_[2174]_ , \new_[2175]_ , \new_[2176]_ , \new_[2177]_ ,
    \new_[2178]_ , \new_[2179]_ , \new_[2181]_ , \new_[2182]_ ,
    \new_[2183]_ , \new_[2184]_ , \new_[2185]_ , \new_[2186]_ ,
    \new_[2187]_ , \new_[2188]_ , \new_[2189]_ , \new_[2190]_ ,
    \new_[2191]_ , \new_[2192]_ , \new_[2193]_ , \new_[2194]_ ,
    \new_[2195]_ , \new_[2196]_ , \new_[2197]_ , \new_[2198]_ ,
    \new_[2199]_ , \new_[2200]_ , \new_[2201]_ , \new_[2202]_ ,
    \new_[2203]_ , \new_[2204]_ , \new_[2205]_ , \new_[2206]_ ,
    \new_[2207]_ , \new_[2208]_ , \new_[2209]_ , \new_[2210]_ ,
    \new_[2211]_ , \new_[2212]_ , \new_[2213]_ , \new_[2214]_ ,
    \new_[2215]_ , \new_[2216]_ , \new_[2217]_ , \new_[2218]_ ,
    \new_[2219]_ , \new_[2220]_ , \new_[2221]_ , \new_[2222]_ ,
    \new_[2223]_ , \new_[2224]_ , \new_[2225]_ , \new_[2226]_ ,
    \new_[2227]_ , \new_[2228]_ , \new_[2229]_ , \new_[2230]_ ,
    \new_[2231]_ , \new_[2232]_ , \new_[2233]_ , \new_[2234]_ ,
    \new_[2235]_ , \new_[2236]_ , \new_[2237]_ , \new_[2238]_ ,
    \new_[2239]_ , \new_[2240]_ , \new_[2241]_ , \new_[2242]_ ,
    \new_[2243]_ , \new_[2244]_ , \new_[2245]_ , \new_[2246]_ ,
    \new_[2247]_ , \new_[2248]_ , \new_[2249]_ , \new_[2250]_ ,
    \new_[2251]_ , \new_[2252]_ , \new_[2254]_ , \new_[2255]_ ,
    \new_[2256]_ , \new_[2257]_ , \new_[2258]_ , \new_[2259]_ ,
    \new_[2260]_ , \new_[2261]_ , \new_[2262]_ , \new_[2263]_ ,
    \new_[2264]_ , \new_[2265]_ , \new_[2266]_ , \new_[2267]_ ,
    \new_[2268]_ , \new_[2269]_ , \new_[2270]_ , \new_[2271]_ ,
    \new_[2272]_ , \new_[2273]_ , \new_[2274]_ , \new_[2275]_ ,
    \new_[2276]_ , \new_[2277]_ , \new_[2278]_ , \new_[2279]_ ,
    \new_[2280]_ , \new_[2281]_ , \new_[2282]_ , \new_[2283]_ ,
    \new_[2284]_ , \new_[2285]_ , \new_[2286]_ , \new_[2287]_ ,
    \new_[2288]_ , \new_[2289]_ , \new_[2290]_ , \new_[2291]_ ,
    \new_[2292]_ , \new_[2293]_ , \new_[2294]_ , \new_[2295]_ ,
    \new_[2296]_ , \new_[2297]_ , \new_[2298]_ , \new_[2299]_ ,
    \new_[2300]_ , \new_[2301]_ , \new_[2302]_ , \new_[2303]_ ,
    \new_[2304]_ , \new_[2305]_ , \new_[2306]_ , \new_[2307]_ ,
    \new_[2308]_ , \new_[2309]_ , \new_[2310]_ , \new_[2311]_ ,
    \new_[2312]_ , \new_[2313]_ , \new_[2314]_ , \new_[2315]_ ,
    \new_[2316]_ , \new_[2317]_ , \new_[2318]_ , \new_[2319]_ ,
    \new_[2320]_ , \new_[2321]_ , \new_[2322]_ , \new_[2323]_ ,
    \new_[2324]_ , \new_[2325]_ , \new_[2326]_ , \new_[2327]_ ,
    \new_[2328]_ , \new_[2329]_ , \new_[2330]_ , \new_[2331]_ ,
    \new_[2332]_ , \new_[2333]_ , \new_[2334]_ , \new_[2335]_ ,
    \new_[2336]_ , \new_[2337]_ , \new_[2338]_ , \new_[2339]_ ,
    \new_[2340]_ , \new_[2341]_ , \new_[2342]_ , \new_[2343]_ ,
    \new_[2344]_ , \new_[2345]_ , \new_[2346]_ , \new_[2347]_ ,
    \new_[2348]_ , \new_[2349]_ , \new_[2350]_ , \new_[2351]_ ,
    \new_[2352]_ , \new_[2353]_ , \new_[2354]_ , \new_[2355]_ ,
    \new_[2356]_ , \new_[2357]_ , \new_[2360]_ , \new_[2361]_ ,
    \new_[2362]_ , \new_[2363]_ , \new_[2364]_ , \new_[2365]_ ,
    \new_[2366]_ , \new_[2367]_ , \new_[2368]_ , \new_[2369]_ ,
    \new_[2370]_ , \new_[2371]_ , \new_[2372]_ , \new_[2373]_ ,
    \new_[2374]_ , \new_[2375]_ , \new_[2376]_ , \new_[2377]_ ,
    \new_[2378]_ , \new_[2379]_ , \new_[2380]_ , \new_[2381]_ ,
    \new_[2382]_ , \new_[2383]_ , \new_[2384]_ , \new_[2385]_ ,
    \new_[2386]_ , \new_[2387]_ , \new_[2388]_ , \new_[2389]_ ,
    \new_[2390]_ , \new_[2391]_ , \new_[2392]_ , \new_[2393]_ ,
    \new_[2394]_ , \new_[2395]_ , \new_[2396]_ , \new_[2397]_ ,
    \new_[2398]_ , \new_[2399]_ , \new_[2400]_ , \new_[2401]_ ,
    \new_[2402]_ , \new_[2403]_ , \new_[2404]_ , \new_[2405]_ ,
    \new_[2406]_ , \new_[2407]_ , \new_[2408]_ , \new_[2409]_ ,
    \new_[2410]_ , \new_[2411]_ , \new_[2412]_ , \new_[2413]_ ,
    \new_[2414]_ , \new_[2415]_ , \new_[2416]_ , \new_[2417]_ ,
    \new_[2418]_ , \new_[2419]_ , \new_[2420]_ , \new_[2421]_ ,
    \new_[2422]_ , \new_[2423]_ , \new_[2424]_ , \new_[2425]_ ,
    \new_[2426]_ , \new_[2428]_ , \new_[2429]_ , \new_[2430]_ ,
    \new_[2431]_ , \new_[2432]_ , \new_[2433]_ , \new_[2434]_ ,
    \new_[2435]_ , \new_[2436]_ , \new_[2437]_ , \new_[2438]_ ,
    \new_[2439]_ , \new_[2440]_ , \new_[2441]_ , \new_[2442]_ ,
    \new_[2443]_ , \new_[2444]_ , \new_[2445]_ , \new_[2446]_ ,
    \new_[2447]_ , \new_[2448]_ , \new_[2449]_ , \new_[2450]_ ,
    \new_[2451]_ , \new_[2452]_ , \new_[2453]_ , \new_[2454]_ ,
    \new_[2455]_ , \new_[2456]_ , \new_[2457]_ , \new_[2458]_ ,
    \new_[2459]_ , \new_[2460]_ , \new_[2461]_ , \new_[2462]_ ,
    \new_[2463]_ , \new_[2464]_ , \new_[2465]_ , \new_[2466]_ ,
    \new_[2467]_ , \new_[2468]_ , \new_[2469]_ , \new_[2470]_ ,
    \new_[2471]_ , \new_[2472]_ , \new_[2473]_ , \new_[2474]_ ,
    \new_[2475]_ , \new_[2476]_ , \new_[2477]_ , \new_[2478]_ ,
    \new_[2479]_ , \new_[2480]_ , \new_[2481]_ , \new_[2482]_ ,
    \new_[2483]_ , \new_[2484]_ , \new_[2485]_ , \new_[2486]_ ,
    \new_[2487]_ , \new_[2488]_ , \new_[2489]_ , \new_[2490]_ ,
    \new_[2491]_ , \new_[2492]_ , \new_[2493]_ , \new_[2494]_ ,
    \new_[2495]_ , \new_[2496]_ , \new_[2497]_ , \new_[2498]_ ,
    \new_[2499]_ , \new_[2500]_ , \new_[2501]_ , \new_[2502]_ ,
    \new_[2503]_ , \new_[2504]_ , \new_[2505]_ , \new_[2506]_ ,
    \new_[2507]_ , \new_[2508]_ , \new_[2509]_ , \new_[2510]_ ,
    \new_[2511]_ , \new_[2512]_ , \new_[2513]_ , \new_[2514]_ ,
    \new_[2515]_ , \new_[2516]_ , \new_[2517]_ , \new_[2518]_ ,
    \new_[2519]_ , \new_[2520]_ , \new_[2521]_ , \new_[2522]_ ,
    \new_[2523]_ , \new_[2524]_ , \new_[2525]_ , \new_[2526]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2549]_ ,
    \new_[2550]_ , \new_[2551]_ , \new_[2552]_ , \new_[2553]_ ,
    \new_[2554]_ , \new_[2555]_ , \new_[2556]_ , \new_[2557]_ ,
    \new_[2558]_ , \new_[2559]_ , \new_[2560]_ , \new_[2561]_ ,
    \new_[2562]_ , \new_[2563]_ , \new_[2564]_ , \new_[2565]_ ,
    \new_[2566]_ , \new_[2567]_ , \new_[2568]_ , \new_[2569]_ ,
    \new_[2570]_ , \new_[2571]_ , \new_[2572]_ , \new_[2573]_ ,
    \new_[2574]_ , \new_[2575]_ , \new_[2576]_ , \new_[2577]_ ,
    \new_[2578]_ , \new_[2579]_ , \new_[2580]_ , \new_[2581]_ ,
    \new_[2582]_ , \new_[2583]_ , \new_[2584]_ , \new_[2585]_ ,
    \new_[2586]_ , \new_[2587]_ , \new_[2588]_ , \new_[2589]_ ,
    \new_[2590]_ , \new_[2591]_ , \new_[2592]_ , \new_[2593]_ ,
    \new_[2594]_ , \new_[2595]_ , \new_[2596]_ , \new_[2597]_ ,
    \new_[2598]_ , \new_[2599]_ , \new_[2600]_ , \new_[2601]_ ,
    \new_[2602]_ , \new_[2603]_ , \new_[2604]_ , \new_[2605]_ ,
    \new_[2606]_ , \new_[2607]_ , \new_[2608]_ , \new_[2609]_ ,
    \new_[2610]_ , \new_[2611]_ , \new_[2612]_ , \new_[2613]_ ,
    \new_[2614]_ , \new_[2615]_ , \new_[2616]_ , \new_[2617]_ ,
    \new_[2618]_ , \new_[2619]_ , \new_[2620]_ , \new_[2621]_ ,
    \new_[2622]_ , \new_[2623]_ , \new_[2624]_ , \new_[2625]_ ,
    \new_[2626]_ , \new_[2627]_ , \new_[2628]_ , \new_[2629]_ ,
    \new_[2630]_ , \new_[2631]_ , \new_[2632]_ , \new_[2633]_ ,
    \new_[2634]_ , \new_[2635]_ , \new_[2636]_ , \new_[2637]_ ,
    \new_[2638]_ , \new_[2639]_ , \new_[2640]_ , \new_[2641]_ ,
    \new_[2642]_ , \new_[2643]_ , \new_[2644]_ , \new_[2645]_ ,
    \new_[2646]_ , \new_[2647]_ , \new_[2648]_ , \new_[2649]_ ,
    \new_[2650]_ , \new_[2651]_ , \new_[2652]_ , \new_[2653]_ ,
    \new_[2656]_ , \new_[2658]_ , \new_[2660]_ , \new_[2661]_ ,
    \new_[2662]_ , \new_[2663]_ , \new_[2664]_ , \new_[2665]_ ,
    \new_[2666]_ , \new_[2667]_ , \new_[2668]_ , \new_[2669]_ ,
    \new_[2670]_ , \new_[2671]_ , \new_[2672]_ , \new_[2673]_ ,
    \new_[2674]_ , \new_[2675]_ , \new_[2676]_ , \new_[2677]_ ,
    \new_[2678]_ , \new_[2679]_ , \new_[2680]_ , \new_[2681]_ ,
    \new_[2682]_ , \new_[2683]_ , \new_[2684]_ , \new_[2685]_ ,
    \new_[2686]_ , \new_[2687]_ , \new_[2688]_ , \new_[2689]_ ,
    \new_[2690]_ , \new_[2691]_ , \new_[2692]_ , \new_[2693]_ ,
    \new_[2694]_ , \new_[2695]_ , \new_[2696]_ , \new_[2697]_ ,
    \new_[2698]_ , \new_[2699]_ , \new_[2700]_ , \new_[2701]_ ,
    \new_[2702]_ , \new_[2703]_ , \new_[2704]_ , \new_[2706]_ ,
    \new_[2707]_ , \new_[2708]_ , \new_[2709]_ , \new_[2710]_ ,
    \new_[2711]_ , \new_[2712]_ , \new_[2713]_ , \new_[2714]_ ,
    \new_[2715]_ , \new_[2716]_ , \new_[2717]_ , \new_[2718]_ ,
    \new_[2719]_ , \new_[2720]_ , \new_[2723]_ , \new_[2727]_ ,
    \new_[2728]_ , \new_[2729]_ , \new_[2730]_ , \new_[2731]_ ,
    \new_[2732]_ , \new_[2733]_ , \new_[2734]_ , \new_[2735]_ ,
    \new_[2736]_ , \new_[2737]_ , \new_[2738]_ , \new_[2739]_ ,
    \new_[2740]_ , \new_[2741]_ , \new_[2742]_ , \new_[2743]_ ,
    \new_[2744]_ , \new_[2745]_ , \new_[2746]_ , \new_[2747]_ ,
    \new_[2748]_ , \new_[2749]_ , \new_[2750]_ , \new_[2751]_ ,
    \new_[2752]_ , \new_[2753]_ , \new_[2754]_ , \new_[2755]_ ,
    \new_[2756]_ , \new_[2757]_ , \new_[2758]_ , \new_[2759]_ ,
    \new_[2760]_ , \new_[2761]_ , \new_[2762]_ , \new_[2763]_ ,
    \new_[2764]_ , \new_[2765]_ , \new_[2766]_ , \new_[2767]_ ,
    \new_[2768]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2777]_ ,
    \new_[2779]_ , \new_[2780]_ , \new_[2787]_ , \new_[2789]_ ,
    \new_[2790]_ , \new_[2791]_ , \new_[2792]_ , \new_[2793]_ ,
    \new_[2794]_ , \new_[2795]_ , \new_[2796]_ , \new_[2797]_ ,
    \new_[2798]_ , \new_[2799]_ , \new_[2800]_ , \new_[2801]_ ,
    \new_[2802]_ , \new_[2803]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2806]_ , \new_[2807]_ , \new_[2808]_ , \new_[2809]_ ,
    \new_[2810]_ , \new_[2811]_ , \new_[2812]_ , \new_[2813]_ ,
    \new_[2814]_ , \new_[2815]_ , \new_[2816]_ , \new_[2817]_ ,
    \new_[2818]_ , \new_[2819]_ , \new_[2820]_ , \new_[2821]_ ,
    \new_[2822]_ , \new_[2823]_ , \new_[2824]_ , \new_[2825]_ ,
    \new_[2826]_ , \new_[2827]_ , \new_[2828]_ , \new_[2830]_ ,
    \new_[2831]_ , \new_[2833]_ , \new_[2834]_ , \new_[2835]_ ,
    \new_[2836]_ , \new_[2837]_ , \new_[2838]_ , \new_[2839]_ ,
    \new_[2840]_ , \new_[2841]_ , \new_[2842]_ , \new_[2843]_ ,
    \new_[2844]_ , \new_[2845]_ , \new_[2846]_ , \new_[2847]_ ,
    \new_[2848]_ , \new_[2849]_ , \new_[2850]_ , \new_[2851]_ ,
    \new_[2852]_ , \new_[2853]_ , \new_[2854]_ , \new_[2855]_ ,
    \new_[2856]_ , \new_[2857]_ , \new_[2858]_ , \new_[2859]_ ,
    \new_[2860]_ , \new_[2861]_ , \new_[2862]_ , \new_[2863]_ ,
    \new_[2864]_ , \new_[2865]_ , \new_[2866]_ , \new_[2867]_ ,
    \new_[2868]_ , \new_[2869]_ , \new_[2873]_ , \new_[2874]_ ,
    \new_[2875]_ , \new_[2876]_ , \new_[2877]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2880]_ , \new_[2881]_ , \new_[2882]_ ,
    \new_[2883]_ , \new_[2884]_ , \new_[2885]_ , \new_[2886]_ ,
    \new_[2887]_ , \new_[2888]_ , \new_[2889]_ , \new_[2890]_ ,
    \new_[2891]_ , \new_[2892]_ , \new_[2893]_ , \new_[2894]_ ,
    \new_[2895]_ , \new_[2896]_ , \new_[2897]_ , \new_[2898]_ ,
    \new_[2899]_ , \new_[2900]_ , \new_[2901]_ , \new_[2902]_ ,
    \new_[2903]_ , \new_[2904]_ , \new_[2905]_ , \new_[2906]_ ,
    \new_[2907]_ , \new_[2908]_ , \new_[2909]_ , \new_[2910]_ ,
    \new_[2911]_ , \new_[2912]_ , \new_[2913]_ , \new_[2914]_ ,
    \new_[2915]_ , \new_[2916]_ , \new_[2917]_ , \new_[2918]_ ,
    \new_[2919]_ , \new_[2920]_ , \new_[2921]_ , \new_[2922]_ ,
    \new_[2923]_ , \new_[2924]_ , \new_[2926]_ , \new_[2927]_ ,
    \new_[2928]_ , \new_[2929]_ , \new_[2930]_ , \new_[2931]_ ,
    \new_[2932]_ , \new_[2933]_ , \new_[2934]_ , \new_[2935]_ ,
    \new_[2936]_ , \new_[2937]_ , \new_[2938]_ , \new_[2939]_ ,
    \new_[2940]_ , \new_[2941]_ , \new_[2942]_ , \new_[2943]_ ,
    \new_[2944]_ , \new_[2945]_ , \new_[2946]_ , \new_[2947]_ ,
    \new_[2948]_ , \new_[2949]_ , \new_[2950]_ , \new_[2951]_ ,
    \new_[2952]_ , \new_[2953]_ , \new_[2954]_ , \new_[2955]_ ,
    \new_[2956]_ , \new_[2957]_ , \new_[2958]_ , \new_[2959]_ ,
    \new_[2960]_ , \new_[2961]_ , \new_[2962]_ , \new_[2963]_ ,
    \new_[2964]_ , \new_[2965]_ , \new_[2966]_ , \new_[2967]_ ,
    \new_[2968]_ , \new_[2969]_ , \new_[2970]_ , \new_[2971]_ ,
    \new_[2972]_ , \new_[2974]_ , \new_[2975]_ , \new_[2976]_ ,
    \new_[2977]_ , \new_[2979]_ , \new_[2980]_ , \new_[2981]_ ,
    \new_[2982]_ , \new_[2983]_ , \new_[2984]_ , \new_[2985]_ ,
    \new_[2986]_ , \new_[2987]_ , \new_[2988]_ , \new_[2989]_ ,
    \new_[2990]_ , \new_[2991]_ , \new_[2992]_ , \new_[2993]_ ,
    \new_[2994]_ , \new_[2995]_ , \new_[2996]_ , \new_[2997]_ ,
    \new_[2998]_ , \new_[2999]_ , \new_[3000]_ , \new_[3001]_ ,
    \new_[3002]_ , \new_[3003]_ , \new_[3004]_ , \new_[3005]_ ,
    \new_[3006]_ , \new_[3007]_ , \new_[3008]_ , \new_[3009]_ ,
    \new_[3010]_ , \new_[3014]_ , \new_[3015]_ , \new_[3016]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3019]_ , \new_[3020]_ ,
    \new_[3021]_ , \new_[3022]_ , \new_[3023]_ , \new_[3025]_ ,
    \new_[3026]_ , \new_[3027]_ , \new_[3028]_ , \new_[3029]_ ,
    \new_[3030]_ , \new_[3031]_ , \new_[3032]_ , \new_[3033]_ ,
    \new_[3034]_ , \new_[3035]_ , \new_[3036]_ , \new_[3037]_ ,
    \new_[3038]_ , \new_[3039]_ , \new_[3040]_ , \new_[3041]_ ,
    \new_[3042]_ , \new_[3043]_ , \new_[3044]_ , \new_[3045]_ ,
    \new_[3046]_ , \new_[3047]_ , \new_[3048]_ , \new_[3049]_ ,
    \new_[3051]_ , \new_[3052]_ , \new_[3053]_ , \new_[3054]_ ,
    \new_[3055]_ , \new_[3056]_ , \new_[3057]_ , \new_[3058]_ ,
    \new_[3059]_ , \new_[3060]_ , \new_[3061]_ , \new_[3062]_ ,
    \new_[3063]_ , \new_[3064]_ , \new_[3065]_ , \new_[3066]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3069]_ , \new_[3070]_ ,
    \new_[3071]_ , \new_[3072]_ , \new_[3073]_ , \new_[3074]_ ,
    \new_[3076]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3082]_ , \new_[3083]_ ,
    \new_[3084]_ , \new_[3085]_ , \new_[3086]_ , \new_[3087]_ ,
    \new_[3088]_ , \new_[3089]_ , \new_[3090]_ , \new_[3091]_ ,
    \new_[3092]_ , \new_[3093]_ , \new_[3094]_ , \new_[3095]_ ,
    \new_[3096]_ , \new_[3097]_ , \new_[3098]_ , \new_[3099]_ ,
    \new_[3100]_ , \new_[3101]_ , \new_[3102]_ , \new_[3103]_ ,
    \new_[3104]_ , \new_[3105]_ , \new_[3106]_ , \new_[3107]_ ,
    \new_[3108]_ , \new_[3109]_ , \new_[3110]_ , \new_[3111]_ ,
    \new_[3112]_ , \new_[3113]_ , \new_[3114]_ , \new_[3115]_ ,
    \new_[3117]_ , \new_[3118]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3124]_ ,
    \new_[3125]_ , \new_[3126]_ , \new_[3127]_ , \new_[3128]_ ,
    \new_[3129]_ , \new_[3130]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3135]_ , \new_[3136]_ ,
    \new_[3137]_ , \new_[3138]_ , \new_[3139]_ , \new_[3140]_ ,
    \new_[3141]_ , \new_[3142]_ , \new_[3143]_ , \new_[3144]_ ,
    \new_[3145]_ , \new_[3146]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3150]_ , \new_[3151]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3156]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3162]_ , \new_[3163]_ , \new_[3164]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3173]_ , \new_[3174]_ , \new_[3175]_ , \new_[3176]_ ,
    \new_[3177]_ , \new_[3178]_ , \new_[3179]_ , \new_[3180]_ ,
    \new_[3181]_ , \new_[3182]_ , \new_[3183]_ , \new_[3184]_ ,
    \new_[3185]_ , \new_[3186]_ , \new_[3187]_ , \new_[3188]_ ,
    \new_[3189]_ , \new_[3190]_ , \new_[3191]_ , \new_[3192]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3197]_ , \new_[3198]_ , \new_[3199]_ , \new_[3200]_ ,
    \new_[3201]_ , \new_[3202]_ , \new_[3203]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3222]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3226]_ , \new_[3227]_ , \new_[3228]_ ,
    \new_[3229]_ , \new_[3230]_ , \new_[3231]_ , \new_[3232]_ ,
    \new_[3233]_ , \new_[3234]_ , \new_[3235]_ , \new_[3236]_ ,
    \new_[3237]_ , \new_[3238]_ , \new_[3239]_ , \new_[3240]_ ,
    \new_[3241]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3246]_ , \new_[3247]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3251]_ , \new_[3252]_ ,
    \new_[3253]_ , \new_[3254]_ , \new_[3255]_ , \new_[3256]_ ,
    \new_[3257]_ , \new_[3258]_ , \new_[3259]_ , \new_[3260]_ ,
    \new_[3261]_ , \new_[3262]_ , \new_[3263]_ , \new_[3264]_ ,
    \new_[3265]_ , \new_[3266]_ , \new_[3267]_ , \new_[3268]_ ,
    \new_[3269]_ , \new_[3270]_ , \new_[3271]_ , \new_[3272]_ ,
    \new_[3273]_ , \new_[3274]_ , \new_[3275]_ , \new_[3276]_ ,
    \new_[3277]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3281]_ , \new_[3282]_ , \new_[3283]_ , \new_[3284]_ ,
    \new_[3285]_ , \new_[3286]_ , \new_[3287]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3294]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3298]_ , \new_[3299]_ , \new_[3300]_ ,
    \new_[3301]_ , \new_[3302]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3305]_ , \new_[3306]_ , \new_[3307]_ , \new_[3308]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3319]_ , \new_[3320]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3323]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3399]_ , \new_[3400]_ , \new_[3401]_ ,
    \new_[3402]_ , \new_[3403]_ , \new_[3404]_ , \new_[3405]_ ,
    \new_[3406]_ , \new_[3407]_ , \new_[3408]_ , \new_[3409]_ ,
    \new_[3410]_ , \new_[3411]_ , \new_[3412]_ , \new_[3413]_ ,
    \new_[3414]_ , \new_[3415]_ , \new_[3416]_ , \new_[3417]_ ,
    \new_[3418]_ , \new_[3419]_ , \new_[3420]_ , \new_[3421]_ ,
    \new_[3422]_ , \new_[3423]_ , \new_[3424]_ , \new_[3425]_ ,
    \new_[3426]_ , \new_[3427]_ , \new_[3428]_ , \new_[3429]_ ,
    \new_[3430]_ , \new_[3431]_ , \new_[3432]_ , \new_[3433]_ ,
    \new_[3434]_ , \new_[3435]_ , \new_[3436]_ , \new_[3437]_ ,
    \new_[3438]_ , \new_[3439]_ , \new_[3440]_ , \new_[3441]_ ,
    \new_[3442]_ , \new_[3443]_ , \new_[3444]_ , \new_[3445]_ ,
    \new_[3446]_ , \new_[3447]_ , \new_[3448]_ , \new_[3449]_ ,
    \new_[3450]_ , \new_[3451]_ , \new_[3452]_ , \new_[3453]_ ,
    \new_[3454]_ , \new_[3455]_ , \new_[3456]_ , \new_[3457]_ ,
    \new_[3458]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3493]_ ,
    \new_[3494]_ , \new_[3495]_ , \new_[3496]_ , \new_[3497]_ ,
    \new_[3498]_ , \new_[3499]_ , \new_[3500]_ , \new_[3501]_ ,
    \new_[3502]_ , \new_[3503]_ , \new_[3504]_ , \new_[3505]_ ,
    \new_[3506]_ , \new_[3507]_ , \new_[3508]_ , \new_[3509]_ ,
    \new_[3510]_ , \new_[3511]_ , \new_[3512]_ , \new_[3513]_ ,
    \new_[3514]_ , \new_[3515]_ , \new_[3516]_ , \new_[3517]_ ,
    \new_[3518]_ , \new_[3519]_ , \new_[3520]_ , \new_[3521]_ ,
    \new_[3522]_ , \new_[3523]_ , \new_[3524]_ , \new_[3525]_ ,
    \new_[3526]_ , \new_[3527]_ , \new_[3528]_ , \new_[3529]_ ,
    \new_[3530]_ , \new_[3531]_ , \new_[3532]_ , \new_[3533]_ ,
    \new_[3534]_ , \new_[3535]_ , \new_[3536]_ , \new_[3537]_ ,
    \new_[3538]_ , \new_[3539]_ , \new_[3540]_ , \new_[3541]_ ,
    \new_[3542]_ , \new_[3543]_ , \new_[3544]_ , \new_[3545]_ ,
    \new_[3546]_ , \new_[3547]_ , \new_[3548]_ , \new_[3549]_ ,
    \new_[3550]_ , \new_[3551]_ , \new_[3552]_ , \new_[3553]_ ,
    \new_[3554]_ , \new_[3555]_ , \new_[3556]_ , \new_[3557]_ ,
    \new_[3558]_ , \new_[3559]_ , \new_[3560]_ , \new_[3561]_ ,
    \new_[3562]_ , \new_[3563]_ , \new_[3564]_ , \new_[3565]_ ,
    \new_[3566]_ , \new_[3567]_ , \new_[3568]_ , \new_[3569]_ ,
    \new_[3570]_ , \new_[3571]_ , \new_[3572]_ , \new_[3573]_ ,
    \new_[3574]_ , \new_[3575]_ , \new_[3576]_ , \new_[3577]_ ,
    \new_[3578]_ , \new_[3579]_ , \new_[3580]_ , \new_[3581]_ ,
    \new_[3582]_ , \new_[3583]_ , \new_[3584]_ , \new_[3585]_ ,
    \new_[3586]_ , \new_[3587]_ , \new_[3588]_ , \new_[3589]_ ,
    \new_[3590]_ , \new_[3591]_ , \new_[3592]_ , \new_[3593]_ ,
    \new_[3594]_ , \new_[3595]_ , \new_[3596]_ , \new_[3597]_ ,
    \new_[3598]_ , \new_[3599]_ , \new_[3600]_ , \new_[3601]_ ,
    \new_[3602]_ , \new_[3603]_ , \new_[3604]_ , \new_[3605]_ ,
    \new_[3606]_ , \new_[3607]_ , \new_[3608]_ , \new_[3609]_ ,
    \new_[3610]_ , \new_[3611]_ , \new_[3612]_ , \new_[3613]_ ,
    \new_[3614]_ , \new_[3615]_ , \new_[3616]_ , \new_[3617]_ ,
    \new_[3618]_ , \new_[3619]_ , \new_[3620]_ , \new_[3621]_ ,
    \new_[3622]_ , \new_[3623]_ , \new_[3624]_ , \new_[3625]_ ,
    \new_[3626]_ , \new_[3627]_ , \new_[3628]_ , \new_[3629]_ ,
    \new_[3630]_ , \new_[3631]_ , \new_[3632]_ , \new_[3633]_ ,
    \new_[3634]_ , \new_[3635]_ , \new_[3636]_ , \new_[3637]_ ,
    \new_[3638]_ , \new_[3639]_ , \new_[3640]_ , \new_[3641]_ ,
    \new_[3642]_ , \new_[3643]_ , \new_[3644]_ , \new_[3645]_ ,
    \new_[3646]_ , \new_[3647]_ , \new_[3648]_ , \new_[3649]_ ,
    \new_[3650]_ , \new_[3651]_ , \new_[3652]_ , \new_[3653]_ ,
    \new_[3654]_ , \new_[3655]_ , \new_[3656]_ , \new_[3657]_ ,
    \new_[3658]_ , \new_[3659]_ , \new_[3660]_ , \new_[3661]_ ,
    \new_[3662]_ , \new_[3663]_ , \new_[3664]_ , \new_[3665]_ ,
    \new_[3666]_ , \new_[3667]_ , \new_[3668]_ , \new_[3669]_ ,
    \new_[3670]_ , \new_[3671]_ , \new_[3672]_ , \new_[3673]_ ,
    \new_[3674]_ , \new_[3675]_ , \new_[3676]_ , \new_[3677]_ ,
    \new_[3678]_ , \new_[3679]_ , \new_[3680]_ , \new_[3681]_ ,
    \new_[3682]_ , \new_[3683]_ , \new_[3684]_ , \new_[3685]_ ,
    \new_[3686]_ , \new_[3687]_ , \new_[3688]_ , \new_[3689]_ ,
    \new_[3690]_ , \new_[3691]_ , \new_[3692]_ , \new_[3693]_ ,
    \new_[3694]_ , \new_[3695]_ , \new_[3696]_ , \new_[3697]_ ,
    \new_[3698]_ , \new_[3699]_ , \new_[3700]_ , \new_[3701]_ ,
    \new_[3702]_ , \new_[3703]_ , \new_[3704]_ , \new_[3705]_ ,
    \new_[3706]_ , \new_[3707]_ , \new_[3708]_ , \new_[3709]_ ,
    \new_[3710]_ , \new_[3711]_ , \new_[3712]_ , \new_[3713]_ ,
    \new_[3714]_ , \new_[3715]_ , \new_[3717]_ , \new_[3718]_ ,
    \new_[3719]_ , \new_[3720]_ , \new_[3721]_ , \new_[3722]_ ,
    \new_[3723]_ , \new_[3724]_ , \new_[3725]_ , \new_[3726]_ ,
    \new_[3727]_ , \new_[3728]_ , \new_[3729]_ , \new_[3730]_ ,
    \new_[3731]_ , \new_[3732]_ , \new_[3733]_ , \new_[3734]_ ,
    \new_[3735]_ , \new_[3736]_ , \new_[3737]_ , \new_[3738]_ ,
    \new_[3739]_ , \new_[3740]_ , \new_[3741]_ , \new_[3742]_ ,
    \new_[3743]_ , \new_[3744]_ , \new_[3745]_ , \new_[3746]_ ,
    \new_[3747]_ , \new_[3748]_ , \new_[3749]_ , \new_[3750]_ ,
    \new_[3751]_ , \new_[3752]_ , \new_[3753]_ , \new_[3754]_ ,
    \new_[3755]_ , \new_[3756]_ , \new_[3757]_ , \new_[3758]_ ,
    \new_[3759]_ , \new_[3760]_ , \new_[3761]_ , \new_[3762]_ ,
    \new_[3763]_ , \new_[3764]_ , \new_[3765]_ , \new_[3766]_ ,
    \new_[3767]_ , \new_[3768]_ , \new_[3769]_ , \new_[3770]_ ,
    \new_[3771]_ , \new_[3772]_ , \new_[3773]_ , \new_[3774]_ ,
    \new_[3775]_ , \new_[3776]_ , \new_[3777]_ , \new_[3778]_ ,
    \new_[3779]_ , \new_[3780]_ , \new_[3781]_ , \new_[3782]_ ,
    \new_[3783]_ , \new_[3784]_ , \new_[3793]_ , \new_[3794]_ ,
    \new_[3795]_ , \new_[3796]_ , \new_[3797]_ , \new_[3798]_ ,
    \new_[3799]_ , \new_[3800]_ , \new_[3801]_ , \new_[3802]_ ,
    \new_[3803]_ , \new_[3804]_ , \new_[3805]_ , \new_[3806]_ ,
    \new_[3807]_ , \new_[3808]_ , \new_[3809]_ , \new_[3810]_ ,
    \new_[3811]_ , \new_[3812]_ , \new_[3813]_ , \new_[3814]_ ,
    \new_[3815]_ , \new_[3816]_ , \new_[3817]_ , \new_[3818]_ ,
    \new_[3819]_ , \new_[3820]_ , \new_[3821]_ , \new_[3822]_ ,
    \new_[3823]_ , \new_[3824]_ , \new_[3825]_ , \new_[3826]_ ,
    \new_[3827]_ , \new_[3828]_ , \new_[3829]_ , \new_[3830]_ ,
    \new_[3831]_ , \new_[3832]_ , \new_[3833]_ , \new_[3834]_ ,
    \new_[3835]_ , \new_[3836]_ , \new_[3837]_ , \new_[3838]_ ,
    \new_[3839]_ , \new_[3840]_ , \new_[3841]_ , \new_[3842]_ ,
    \new_[3843]_ , \new_[3844]_ , \new_[3845]_ , \new_[3846]_ ,
    \new_[3847]_ , \new_[3848]_ , \new_[3849]_ , \new_[3850]_ ,
    \new_[3851]_ , \new_[3852]_ , \new_[3853]_ , \new_[3854]_ ,
    \new_[3855]_ , \new_[3856]_ , \new_[3857]_ , \new_[3858]_ ,
    \new_[3859]_ , \new_[3860]_ , \new_[3861]_ , \new_[3862]_ ,
    \new_[3863]_ , \new_[3864]_ , \new_[3865]_ , \new_[3866]_ ,
    \new_[3867]_ , \new_[3868]_ , \new_[3869]_ , \new_[3870]_ ,
    \new_[3871]_ , \new_[3872]_ , \new_[3873]_ , \new_[3874]_ ,
    \new_[3875]_ , \new_[3876]_ , \new_[3877]_ , \new_[3878]_ ,
    \new_[3879]_ , \new_[3880]_ , \new_[3881]_ , \new_[3882]_ ,
    \new_[3883]_ , \new_[3884]_ , \new_[3885]_ , \new_[3886]_ ,
    \new_[3887]_ , \new_[3888]_ , \new_[3889]_ , \new_[3890]_ ,
    \new_[3891]_ , \new_[3892]_ , \new_[3893]_ , \new_[3894]_ ,
    \new_[3895]_ , \new_[3896]_ , \new_[3897]_ , \new_[3898]_ ,
    \new_[3899]_ , \new_[3900]_ , \new_[3901]_ , \new_[3902]_ ,
    \new_[3903]_ , \new_[3904]_ , \new_[3905]_ , \new_[3906]_ ,
    \new_[3907]_ , \new_[3908]_ , \new_[3909]_ , \new_[3910]_ ,
    \new_[3911]_ , \new_[3912]_ , \new_[3913]_ , \new_[3914]_ ,
    \new_[3915]_ , \new_[3916]_ , \new_[3917]_ , \new_[3918]_ ,
    \new_[3919]_ , \new_[3920]_ , \new_[3921]_ , \new_[3922]_ ,
    \new_[3923]_ , \new_[3924]_ , \new_[3925]_ , \new_[3926]_ ,
    \new_[3927]_ , \new_[3928]_ , \new_[3929]_ , \new_[3930]_ ,
    \new_[3931]_ , \new_[3932]_ , \new_[3933]_ , \new_[3934]_ ,
    \new_[3935]_ , \new_[3936]_ , \new_[3937]_ , \new_[3938]_ ,
    \new_[3939]_ , \new_[3940]_ , \new_[3941]_ , \new_[3942]_ ,
    \new_[3943]_ , \new_[3944]_ , \new_[3945]_ , \new_[3946]_ ,
    \new_[3947]_ , \new_[3948]_ , \new_[3949]_ , \new_[3950]_ ,
    \new_[3951]_ , \new_[3952]_ , \new_[3953]_ , \new_[3954]_ ,
    \new_[3955]_ , \new_[3956]_ , \new_[3957]_ , \new_[3958]_ ,
    \new_[3959]_ , \new_[3960]_ , \new_[3961]_ , \new_[3962]_ ,
    \new_[3963]_ , \new_[3964]_ , \new_[3965]_ , \new_[3967]_ ,
    \new_[3968]_ , \new_[3969]_ , \new_[3970]_ , \new_[3971]_ ,
    \new_[3972]_ , \new_[3973]_ , \new_[3974]_ , \new_[3975]_ ,
    \new_[3976]_ , \new_[3977]_ , \new_[3978]_ , \new_[3980]_ ,
    \new_[3981]_ , \new_[3982]_ , \new_[3983]_ , \new_[3984]_ ,
    \new_[3985]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3989]_ , \new_[3990]_ , \new_[3991]_ , \new_[3992]_ ,
    \new_[3993]_ , \new_[3994]_ , \new_[3995]_ , \new_[3996]_ ,
    \new_[3997]_ , \new_[3998]_ , \new_[3999]_ , \new_[4000]_ ,
    \new_[4001]_ , \new_[4002]_ , \new_[4003]_ , \new_[4004]_ ,
    \new_[4005]_ , \new_[4006]_ , \new_[4007]_ , \new_[4008]_ ,
    \new_[4009]_ , \new_[4010]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4013]_ , \new_[4014]_ , \new_[4015]_ , \new_[4016]_ ,
    \new_[4017]_ , \new_[4018]_ , \new_[4019]_ , \new_[4020]_ ,
    \new_[4021]_ , \new_[4022]_ , \new_[4023]_ , \new_[4024]_ ,
    \new_[4025]_ , \new_[4026]_ , \new_[4027]_ , \new_[4028]_ ,
    \new_[4029]_ , \new_[4030]_ , \new_[4031]_ , \new_[4032]_ ,
    \new_[4033]_ , \new_[4034]_ , \new_[4035]_ , \new_[4036]_ ,
    \new_[4037]_ , \new_[4038]_ , \new_[4039]_ , \new_[4040]_ ,
    \new_[4041]_ , \new_[4042]_ , \new_[4043]_ , \new_[4044]_ ,
    \new_[4045]_ , \new_[4046]_ , \new_[4047]_ , \new_[4048]_ ,
    \new_[4049]_ , \new_[4050]_ , \new_[4051]_ , \new_[4052]_ ,
    \new_[4053]_ , \new_[4054]_ , \new_[4055]_ , \new_[4056]_ ,
    \new_[4057]_ , \new_[4058]_ , \new_[4059]_ , \new_[4060]_ ,
    \new_[4061]_ , \new_[4062]_ , \new_[4063]_ , \new_[4064]_ ,
    \new_[4065]_ , \new_[4066]_ , \new_[4067]_ , \new_[4068]_ ,
    \new_[4069]_ , \new_[4070]_ , \new_[4071]_ , \new_[4072]_ ,
    \new_[4073]_ , \new_[4074]_ , \new_[4075]_ , \new_[4076]_ ,
    \new_[4077]_ , \new_[4078]_ , \new_[4079]_ , \new_[4080]_ ,
    \new_[4081]_ , \new_[4082]_ , \new_[4083]_ , \new_[4084]_ ,
    \new_[4085]_ , \new_[4086]_ , \new_[4087]_ , \new_[4088]_ ,
    \new_[4089]_ , \new_[4090]_ , \new_[4091]_ , \new_[4092]_ ,
    \new_[4093]_ , \new_[4094]_ , \new_[4095]_ , \new_[4096]_ ,
    \new_[4097]_ , \new_[4098]_ , \new_[4099]_ , \new_[4100]_ ,
    \new_[4101]_ , \new_[4102]_ , \new_[4103]_ , \new_[4104]_ ,
    \new_[4105]_ , \new_[4106]_ , \new_[4107]_ , \new_[4108]_ ,
    \new_[4109]_ , \new_[4110]_ , \new_[4111]_ , \new_[4112]_ ,
    \new_[4113]_ , \new_[4114]_ , \new_[4115]_ , \new_[4116]_ ,
    \new_[4117]_ , \new_[4118]_ , \new_[4119]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4122]_ , \new_[4123]_ , \new_[4124]_ ,
    \new_[4125]_ , \new_[4126]_ , \new_[4127]_ , \new_[4128]_ ,
    \new_[4129]_ , \new_[4130]_ , \new_[4131]_ , \new_[4132]_ ,
    \new_[4133]_ , \new_[4134]_ , \new_[4135]_ , \new_[4136]_ ,
    \new_[4137]_ , \new_[4138]_ , \new_[4139]_ , \new_[4140]_ ,
    \new_[4141]_ , \new_[4142]_ , \new_[4143]_ , \new_[4144]_ ,
    \new_[4145]_ , \new_[4146]_ , \new_[4147]_ , \new_[4148]_ ,
    \new_[4149]_ , \new_[4150]_ , \new_[4151]_ , \new_[4152]_ ,
    \new_[4153]_ , \new_[4154]_ , \new_[4155]_ , \new_[4156]_ ,
    \new_[4157]_ , \new_[4158]_ , \new_[4159]_ , \new_[4160]_ ,
    \new_[4161]_ , \new_[4162]_ , \new_[4163]_ , \new_[4164]_ ,
    \new_[4165]_ , \new_[4166]_ , \new_[4167]_ , \new_[4168]_ ,
    \new_[4169]_ , \new_[4170]_ , \new_[4171]_ , \new_[4172]_ ,
    \new_[4173]_ , \new_[4174]_ , \new_[4175]_ , \new_[4176]_ ,
    \new_[4177]_ , \new_[4178]_ , \new_[4179]_ , \new_[4180]_ ,
    \new_[4181]_ , \new_[4182]_ , \new_[4183]_ , \new_[4184]_ ,
    \new_[4185]_ , \new_[4186]_ , \new_[4187]_ , \new_[4188]_ ,
    \new_[4189]_ , \new_[4190]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4193]_ , \new_[4194]_ , \new_[4195]_ , \new_[4196]_ ,
    \new_[4197]_ , \new_[4198]_ , \new_[4199]_ , \new_[4200]_ ,
    \new_[4201]_ , \new_[4202]_ , \new_[4203]_ , \new_[4204]_ ,
    \new_[4205]_ , \new_[4206]_ , \new_[4207]_ , \new_[4208]_ ,
    \new_[4209]_ , \new_[4210]_ , \new_[4211]_ , \new_[4212]_ ,
    \new_[4213]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4219]_ , \new_[4220]_ , \new_[4221]_ ,
    \new_[4222]_ , \new_[4223]_ , \new_[4224]_ , \new_[4225]_ ,
    \new_[4226]_ , \new_[4227]_ , \new_[4228]_ , \new_[4229]_ ,
    \new_[4230]_ , \new_[4231]_ , \new_[4232]_ , \new_[4233]_ ,
    \new_[4234]_ , \new_[4235]_ , \new_[4236]_ , \new_[4237]_ ,
    \new_[4238]_ , \new_[4239]_ , \new_[4240]_ , \new_[4241]_ ,
    \new_[4242]_ , \new_[4243]_ , \new_[4244]_ , \new_[4245]_ ,
    \new_[4246]_ , \new_[4247]_ , \new_[4248]_ , \new_[4249]_ ,
    \new_[4250]_ , \new_[4251]_ , \new_[4252]_ , \new_[4253]_ ,
    \new_[4254]_ , \new_[4255]_ , \new_[4256]_ , \new_[4257]_ ,
    \new_[4258]_ , \new_[4259]_ , \new_[4260]_ , \new_[4261]_ ,
    \new_[4262]_ , \new_[4263]_ , \new_[4264]_ , \new_[4265]_ ,
    \new_[4266]_ , \new_[4267]_ , \new_[4268]_ , \new_[4269]_ ,
    \new_[4270]_ , \new_[4271]_ , \new_[4272]_ , \new_[4273]_ ,
    \new_[4274]_ , \new_[4275]_ , \new_[4276]_ , \new_[4277]_ ,
    \new_[4278]_ , \new_[4279]_ , \new_[4280]_ , \new_[4281]_ ,
    \new_[4282]_ , \new_[4283]_ , \new_[4284]_ , \new_[4285]_ ,
    \new_[4286]_ , \new_[4287]_ , \new_[4288]_ , \new_[4289]_ ,
    \new_[4290]_ , \new_[4291]_ , \new_[4292]_ , \new_[4293]_ ,
    \new_[4294]_ , \new_[4295]_ , \new_[4296]_ , \new_[4297]_ ,
    \new_[4298]_ , \new_[4299]_ , \new_[4300]_ , \new_[4301]_ ,
    \new_[4302]_ , \new_[4303]_ , \new_[4304]_ , \new_[4305]_ ,
    \new_[4306]_ , \new_[4307]_ , \new_[4308]_ , \new_[4309]_ ,
    \new_[4310]_ , \new_[4311]_ , \new_[4312]_ , \new_[4313]_ ,
    \new_[4314]_ , \new_[4315]_ , \new_[4316]_ , \new_[4317]_ ,
    \new_[4318]_ , \new_[4319]_ , \new_[4320]_ , \new_[4321]_ ,
    \new_[4322]_ , \new_[4323]_ , \new_[4324]_ , \new_[4325]_ ,
    \new_[4326]_ , \new_[4327]_ , \new_[4328]_ , \new_[4329]_ ,
    \new_[4330]_ , \new_[4331]_ , \new_[4332]_ , \new_[4333]_ ,
    \new_[4334]_ , \new_[4335]_ , \new_[4336]_ , \new_[4337]_ ,
    \new_[4338]_ , \new_[4339]_ , \new_[4340]_ , \new_[4341]_ ,
    \new_[4342]_ , \new_[4343]_ , \new_[4344]_ , \new_[4345]_ ,
    \new_[4346]_ , \new_[4347]_ , \new_[4348]_ , \new_[4349]_ ,
    \new_[4350]_ , \new_[4351]_ , \new_[4352]_ , \new_[4353]_ ,
    \new_[4354]_ , \new_[4355]_ , \new_[4356]_ , \new_[4357]_ ,
    \new_[4358]_ , \new_[4359]_ , \new_[4360]_ , \new_[4361]_ ,
    \new_[4362]_ , \new_[4363]_ , \new_[4364]_ , \new_[4365]_ ,
    \new_[4366]_ , \new_[4367]_ , \new_[4368]_ , \new_[4369]_ ,
    \new_[4370]_ , \new_[4371]_ , \new_[4372]_ , \new_[4373]_ ,
    \new_[4374]_ , \new_[4375]_ , \new_[4376]_ , \new_[4377]_ ,
    \new_[4378]_ , \new_[4379]_ , \new_[4380]_ , \new_[4381]_ ,
    \new_[4382]_ , \new_[4383]_ , \new_[4384]_ , \new_[4385]_ ,
    \new_[4386]_ , \new_[4387]_ , \new_[4388]_ , \new_[4389]_ ,
    \new_[4390]_ , \new_[4391]_ , \new_[4392]_ , \new_[4393]_ ,
    \new_[4394]_ , \new_[4395]_ , \new_[4396]_ , \new_[4397]_ ,
    \new_[4398]_ , \new_[4399]_ , \new_[4400]_ , \new_[4401]_ ,
    \new_[4402]_ , \new_[4403]_ , \new_[4404]_ , \new_[4405]_ ,
    \new_[4406]_ , \new_[4407]_ , \new_[4408]_ , \new_[4409]_ ,
    \new_[4410]_ , \new_[4411]_ , \new_[4412]_ , \new_[4413]_ ,
    \new_[4414]_ , \new_[4415]_ , \new_[4416]_ , \new_[4417]_ ,
    \new_[4418]_ , \new_[4419]_ , \new_[4420]_ , \new_[4421]_ ,
    \new_[4422]_ , \new_[4423]_ , \new_[4424]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4429]_ , \new_[4430]_ ,
    \new_[4431]_ , \new_[4432]_ , \new_[4433]_ , \new_[4434]_ ,
    \new_[4435]_ , \new_[4436]_ , \new_[4437]_ , \new_[4438]_ ,
    \new_[4439]_ , \new_[4440]_ , \new_[4441]_ , \new_[4442]_ ,
    \new_[4443]_ , \new_[4444]_ , \new_[4445]_ , \new_[4446]_ ,
    \new_[4447]_ , \new_[4448]_ , \new_[4449]_ , \new_[4450]_ ,
    \new_[4451]_ , \new_[4452]_ , \new_[4453]_ , \new_[4454]_ ,
    \new_[4455]_ , \new_[4456]_ , \new_[4457]_ , \new_[4458]_ ,
    \new_[4459]_ , \new_[4460]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4463]_ , \new_[4464]_ , \new_[4465]_ , \new_[4466]_ ,
    \new_[4467]_ , \new_[4468]_ , \new_[4469]_ , \new_[4470]_ ,
    \new_[4471]_ , \new_[4472]_ , \new_[4473]_ , \new_[4474]_ ,
    \new_[4475]_ , \new_[4476]_ , \new_[4477]_ , \new_[4478]_ ,
    \new_[4479]_ , \new_[4480]_ , \new_[4481]_ , \new_[4482]_ ,
    \new_[4483]_ , \new_[4484]_ , \new_[4485]_ , \new_[4486]_ ,
    \new_[4487]_ , \new_[4488]_ , \new_[4489]_ , \new_[4490]_ ,
    \new_[4491]_ , \new_[4492]_ , \new_[4493]_ , \new_[4494]_ ,
    \new_[4495]_ , \new_[4496]_ , \new_[4497]_ , \new_[4498]_ ,
    \new_[4499]_ , \new_[4500]_ , \new_[4501]_ , \new_[4502]_ ,
    \new_[4503]_ , \new_[4504]_ , \new_[4505]_ , \new_[4506]_ ,
    \new_[4507]_ , \new_[4508]_ , \new_[4509]_ , \new_[4510]_ ,
    \new_[4511]_ , \new_[4512]_ , \new_[4513]_ , \new_[4514]_ ,
    \new_[4515]_ , \new_[4516]_ , \new_[4517]_ , \new_[4518]_ ,
    \new_[4519]_ , \new_[4520]_ , \new_[4521]_ , \new_[4522]_ ,
    \new_[4523]_ , \new_[4524]_ , \new_[4525]_ , \new_[4526]_ ,
    \new_[4527]_ , \new_[4528]_ , \new_[4529]_ , \new_[4530]_ ,
    \new_[4531]_ , \new_[4532]_ , \new_[4533]_ , \new_[4534]_ ,
    \new_[4535]_ , \new_[4536]_ , \new_[4537]_ , \new_[4538]_ ,
    \new_[4539]_ , \new_[4540]_ , \new_[4541]_ , \new_[4542]_ ,
    \new_[4543]_ , \new_[4544]_ , \new_[4545]_ , \new_[4546]_ ,
    \new_[4547]_ , \new_[4548]_ , \new_[4549]_ , \new_[4550]_ ,
    \new_[4551]_ , \new_[4552]_ , \new_[4553]_ , \new_[4554]_ ,
    \new_[4555]_ , \new_[4556]_ , \new_[4557]_ , \new_[4558]_ ,
    \new_[4559]_ , \new_[4560]_ , \new_[4561]_ , \new_[4562]_ ,
    \new_[4563]_ , \new_[4564]_ , \new_[4565]_ , \new_[4566]_ ,
    \new_[4567]_ , \new_[4568]_ , \new_[4569]_ , \new_[4570]_ ,
    \new_[4571]_ , \new_[4572]_ , \new_[4573]_ , \new_[4574]_ ,
    \new_[4575]_ , \new_[4576]_ , \new_[4577]_ , \new_[4578]_ ,
    \new_[4579]_ , \new_[4580]_ , \new_[4581]_ , \new_[4582]_ ,
    \new_[4583]_ , \new_[4584]_ , \new_[4585]_ , \new_[4586]_ ,
    \new_[4587]_ , \new_[4588]_ , \new_[4589]_ , \new_[4590]_ ,
    \new_[4591]_ , \new_[4592]_ , \new_[4593]_ , \new_[4594]_ ,
    \new_[4595]_ , \new_[4596]_ , \new_[4597]_ , \new_[4598]_ ,
    \new_[4599]_ , \new_[4600]_ , \new_[4601]_ , \new_[4602]_ ,
    \new_[4603]_ , \new_[4604]_ , \new_[4605]_ , \new_[4606]_ ,
    \new_[4607]_ , \new_[4608]_ , \new_[4609]_ , \new_[4610]_ ,
    \new_[4611]_ , \new_[4612]_ , \new_[4613]_ , \new_[4614]_ ,
    \new_[4615]_ , \new_[4616]_ , \new_[4617]_ , \new_[4618]_ ,
    \new_[4619]_ , \new_[4620]_ , \new_[4621]_ , \new_[4622]_ ,
    \new_[4623]_ , \new_[4624]_ , \new_[4625]_ , \new_[4626]_ ,
    \new_[4627]_ , \new_[4628]_ , \new_[4629]_ , \new_[4630]_ ,
    \new_[4631]_ , \new_[4632]_ , \new_[4633]_ , \new_[4634]_ ,
    \new_[4635]_ , \new_[4636]_ , \new_[4637]_ , \new_[4638]_ ,
    \new_[4639]_ , \new_[4640]_ , \new_[4641]_ , \new_[4642]_ ,
    \new_[4643]_ , \new_[4644]_ , \new_[4645]_ , \new_[4646]_ ,
    \new_[4647]_ , \new_[4648]_ , \new_[4649]_ , \new_[4650]_ ,
    \new_[4651]_ , \new_[4652]_ , \new_[4653]_ , \new_[4654]_ ,
    \new_[4655]_ , \new_[4656]_ , \new_[4657]_ , \new_[4658]_ ,
    \new_[4659]_ , \new_[4660]_ , \new_[4661]_ , \new_[4662]_ ,
    \new_[4663]_ , \new_[4664]_ , \new_[4665]_ , \new_[4666]_ ,
    \new_[4667]_ , \new_[4668]_ , \new_[4669]_ , \new_[4670]_ ,
    \new_[4671]_ , \new_[4672]_ , \new_[4673]_ , \new_[4674]_ ,
    \new_[4675]_ , \new_[4676]_ , \new_[4677]_ , \new_[4678]_ ,
    \new_[4679]_ , \new_[4680]_ , \new_[4681]_ , \new_[4682]_ ,
    \new_[4683]_ , \new_[4684]_ , \new_[4685]_ , \new_[4686]_ ,
    \new_[4687]_ , \new_[4688]_ , \new_[4689]_ , \new_[4690]_ ,
    \new_[4691]_ , \new_[4692]_ , \new_[4693]_ , \new_[4694]_ ,
    \new_[4695]_ , \new_[4704]_ , \new_[4705]_ , \new_[4706]_ ,
    \new_[4707]_ , \new_[4708]_ , \new_[4709]_ , \new_[4710]_ ,
    \new_[4711]_ , \new_[4712]_ , \new_[4713]_ , \new_[4714]_ ,
    \new_[4715]_ , \new_[4716]_ , \new_[4717]_ , \new_[4718]_ ,
    \new_[4719]_ , \new_[4720]_ , \new_[4721]_ , \new_[4722]_ ,
    \new_[4723]_ , \new_[4724]_ , \new_[4725]_ , \new_[4726]_ ,
    \new_[4727]_ , \new_[4728]_ , \new_[4729]_ , \new_[4730]_ ,
    \new_[4731]_ , \new_[4732]_ , \new_[4733]_ , \new_[4734]_ ,
    \new_[4735]_ , \new_[4736]_ , \new_[4737]_ , \new_[4738]_ ,
    \new_[4739]_ , \new_[4740]_ , \new_[4741]_ , \new_[4742]_ ,
    \new_[4743]_ , \new_[4744]_ , \new_[4745]_ , \new_[4746]_ ,
    \new_[4747]_ , \new_[4748]_ , \new_[4749]_ , \new_[4750]_ ,
    \new_[4751]_ , \new_[4752]_ , \new_[4753]_ , \new_[4754]_ ,
    \new_[4755]_ , \new_[4756]_ , \new_[4757]_ , \new_[4758]_ ,
    \new_[4759]_ , \new_[4760]_ , \new_[4761]_ , \new_[4762]_ ,
    \new_[4763]_ , \new_[4764]_ , \new_[4765]_ , \new_[4766]_ ,
    \new_[4767]_ , \new_[4768]_ , \new_[4769]_ , \new_[4770]_ ,
    \new_[4771]_ , \new_[4772]_ , \new_[4773]_ , \new_[4774]_ ,
    \new_[4775]_ , \new_[4776]_ , \new_[4777]_ , \new_[4778]_ ,
    \new_[4779]_ , \new_[4780]_ , \new_[4781]_ , \new_[4782]_ ,
    \new_[4783]_ , \new_[4784]_ , \new_[4785]_ , \new_[4786]_ ,
    \new_[4787]_ , \new_[4788]_ , \new_[4789]_ , \new_[4790]_ ,
    \new_[4791]_ , \new_[4792]_ , \new_[4793]_ , \new_[4794]_ ,
    \new_[4795]_ , \new_[4796]_ , \new_[4797]_ , \new_[4798]_ ,
    \new_[4799]_ , \new_[4800]_ , \new_[4801]_ , \new_[4802]_ ,
    \new_[4803]_ , \new_[4804]_ , \new_[4805]_ , \new_[4806]_ ,
    \new_[4807]_ , \new_[4808]_ , \new_[4809]_ , \new_[4810]_ ,
    \new_[4811]_ , \new_[4812]_ , \new_[4813]_ , \new_[4814]_ ,
    \new_[4815]_ , \new_[4816]_ , \new_[4817]_ , \new_[4818]_ ,
    \new_[4819]_ , \new_[4820]_ , \new_[4821]_ , \new_[4822]_ ,
    \new_[4823]_ , \new_[4824]_ , \new_[4825]_ , \new_[4826]_ ,
    \new_[4827]_ , \new_[4828]_ , \new_[4829]_ , \new_[4830]_ ,
    \new_[4831]_ , \new_[4832]_ , \new_[4833]_ , \new_[4834]_ ,
    \new_[4835]_ , \new_[4836]_ , \new_[4837]_ , \new_[4838]_ ,
    \new_[4839]_ , \new_[4840]_ , \new_[4841]_ , \new_[4842]_ ,
    \new_[4843]_ , \new_[4844]_ , \new_[4845]_ , \new_[4846]_ ,
    \new_[4847]_ , \new_[4848]_ , \new_[4849]_ , \new_[4850]_ ,
    \new_[4851]_ , \new_[4852]_ , \new_[4853]_ , \new_[4854]_ ,
    \new_[4855]_ , \new_[4856]_ , \new_[4857]_ , \new_[4858]_ ,
    \new_[4859]_ , \new_[4860]_ , \new_[4861]_ , \new_[4862]_ ,
    \new_[4863]_ , \new_[4864]_ , \new_[4865]_ , \new_[4866]_ ,
    \new_[4867]_ , \new_[4868]_ , \new_[4869]_ , \new_[4870]_ ,
    \new_[4871]_ , \new_[4872]_ , \new_[4873]_ , \new_[4874]_ ,
    \new_[4875]_ , \new_[4876]_ , \new_[4877]_ , \new_[4878]_ ,
    \new_[4879]_ , \new_[4880]_ , \new_[4881]_ , \new_[4882]_ ,
    \new_[4883]_ , \new_[4884]_ , \new_[4885]_ , \new_[4886]_ ,
    \new_[4887]_ , \new_[4888]_ , \new_[4889]_ , \new_[4890]_ ,
    \new_[4891]_ , \new_[4892]_ , \new_[4893]_ , \new_[4894]_ ,
    \new_[4895]_ , \new_[4896]_ , \new_[4897]_ , \new_[4898]_ ,
    \new_[4899]_ , \new_[4900]_ , \new_[4901]_ , \new_[4902]_ ,
    \new_[4903]_ , \new_[4904]_ , \new_[4905]_ , \new_[4906]_ ,
    \new_[4907]_ , \new_[4908]_ , \new_[4909]_ , \new_[4910]_ ,
    \new_[4911]_ , \new_[4912]_ , \new_[4913]_ , \new_[4914]_ ,
    \new_[4915]_ , \new_[4916]_ , \new_[4917]_ , \new_[4918]_ ,
    \new_[4919]_ , \new_[4920]_ , \new_[4921]_ , \new_[4922]_ ,
    \new_[4923]_ , \new_[4924]_ , \new_[4925]_ , \new_[4926]_ ,
    \new_[4927]_ , \new_[4928]_ , \new_[4929]_ , \new_[4930]_ ,
    \new_[4931]_ , \new_[4932]_ , \new_[4933]_ , \new_[4934]_ ,
    \new_[4935]_ , \new_[4936]_ , \new_[4937]_ , \new_[4938]_ ,
    \new_[4939]_ , \new_[4940]_ , \new_[4941]_ , \new_[4942]_ ,
    \new_[4943]_ , \new_[4944]_ , \new_[4945]_ , \new_[4946]_ ,
    \new_[4947]_ , \new_[4948]_ , \new_[4949]_ , \new_[4950]_ ,
    \new_[4951]_ , \new_[4952]_ , \new_[4953]_ , \new_[4954]_ ,
    \new_[4955]_ , \new_[4956]_ , \new_[4957]_ , \new_[4958]_ ,
    \new_[4959]_ , \new_[4960]_ , \new_[4961]_ , \new_[4962]_ ,
    \new_[4963]_ , \new_[4964]_ , \new_[4965]_ , \new_[4966]_ ,
    \new_[4967]_ , \new_[4968]_ , \new_[4969]_ , \new_[4970]_ ,
    \new_[4971]_ , \new_[4972]_ , \new_[4973]_ , \new_[4974]_ ,
    \new_[4975]_ , \new_[4976]_ , \new_[4977]_ , \new_[4978]_ ,
    \new_[4979]_ , \new_[4980]_ , \new_[4981]_ , \new_[4982]_ ,
    \new_[4983]_ , \new_[4984]_ , \new_[4985]_ , \new_[4986]_ ,
    \new_[4987]_ , \new_[4988]_ , \new_[4989]_ , \new_[4990]_ ,
    \new_[4991]_ , \new_[4992]_ , \new_[4993]_ , \new_[4994]_ ,
    \new_[4995]_ , \new_[4996]_ , \new_[4997]_ , \new_[4998]_ ,
    \new_[4999]_ , \new_[5000]_ , \new_[5001]_ , \new_[5002]_ ,
    \new_[5003]_ , \new_[5004]_ , \new_[5005]_ , \new_[5006]_ ,
    \new_[5007]_ , \new_[5008]_ , \new_[5009]_ , \new_[5010]_ ,
    \new_[5011]_ , \new_[5012]_ , \new_[5013]_ , \new_[5014]_ ,
    \new_[5015]_ , \new_[5016]_ , \new_[5017]_ , \new_[5018]_ ,
    \new_[5019]_ , \new_[5020]_ , \new_[5021]_ , \new_[5022]_ ,
    \new_[5023]_ , \new_[5024]_ , \new_[5025]_ , \new_[5026]_ ,
    \new_[5027]_ , \new_[5028]_ , \new_[5029]_ , \new_[5030]_ ,
    \new_[5031]_ , \new_[5032]_ , \new_[5033]_ , \new_[5034]_ ,
    \new_[5035]_ , \new_[5036]_ , \new_[5037]_ , \new_[5038]_ ,
    \new_[5039]_ , \new_[5040]_ , \new_[5041]_ , \new_[5042]_ ,
    \new_[5043]_ , \new_[5044]_ , \new_[5045]_ , \new_[5046]_ ,
    \new_[5047]_ , \new_[5048]_ , \new_[5049]_ , \new_[5050]_ ,
    \new_[5051]_ , \new_[5052]_ , \new_[5053]_ , \new_[5054]_ ,
    \new_[5055]_ , \new_[5056]_ , \new_[5057]_ , \new_[5058]_ ,
    \new_[5059]_ , \new_[5060]_ , \new_[5061]_ , \new_[5062]_ ,
    \new_[5063]_ , \new_[5064]_ , \new_[5065]_ , \new_[5066]_ ,
    \new_[5067]_ , \new_[5068]_ , \new_[5069]_ , \new_[5070]_ ,
    \new_[5071]_ , \new_[5072]_ , \new_[5073]_ , \new_[5074]_ ,
    \new_[5075]_ , \new_[5076]_ , \new_[5077]_ , \new_[5078]_ ,
    \new_[5079]_ , \new_[5080]_ , \new_[5081]_ , \new_[5082]_ ,
    \new_[5083]_ , \new_[5084]_ , \new_[5085]_ , \new_[5086]_ ,
    \new_[5087]_ , \new_[5088]_ , \new_[5089]_ , \new_[5090]_ ,
    \new_[5091]_ , \new_[5092]_ , \new_[5093]_ , \new_[5094]_ ,
    \new_[5095]_ , \new_[5096]_ , \new_[5097]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5100]_ , \new_[5101]_ , \new_[5102]_ ,
    \new_[5103]_ , \new_[5104]_ , \new_[5105]_ , \new_[5106]_ ,
    \new_[5107]_ , \new_[5108]_ , \new_[5109]_ , \new_[5110]_ ,
    \new_[5111]_ , \new_[5112]_ , \new_[5113]_ , \new_[5114]_ ,
    \new_[5115]_ , \new_[5116]_ , \new_[5117]_ , \new_[5118]_ ,
    \new_[5119]_ , \new_[5120]_ , \new_[5121]_ , \new_[5122]_ ,
    \new_[5123]_ , \new_[5124]_ , \new_[5125]_ , \new_[5126]_ ,
    \new_[5127]_ , \new_[5128]_ , \new_[5129]_ , \new_[5130]_ ,
    \new_[5131]_ , \new_[5132]_ , \new_[5133]_ , \new_[5134]_ ,
    \new_[5135]_ , \new_[5136]_ , \new_[5137]_ , \new_[5138]_ ,
    \new_[5139]_ , \new_[5140]_ , \new_[5141]_ , \new_[5142]_ ,
    \new_[5143]_ , \new_[5144]_ , \new_[5145]_ , \new_[5146]_ ,
    \new_[5147]_ , \new_[5148]_ , \new_[5149]_ , \new_[5150]_ ,
    \new_[5151]_ , \new_[5152]_ , \new_[5153]_ , \new_[5154]_ ,
    \new_[5155]_ , \new_[5156]_ , \new_[5157]_ , \new_[5158]_ ,
    \new_[5159]_ , \new_[5160]_ , \new_[5161]_ , \new_[5162]_ ,
    \new_[5163]_ , \new_[5164]_ , \new_[5165]_ , \new_[5166]_ ,
    \new_[5167]_ , \new_[5168]_ , \new_[5169]_ , \new_[5170]_ ,
    \new_[5171]_ , \new_[5172]_ , \new_[5173]_ , \new_[5174]_ ,
    \new_[5175]_ , \new_[5176]_ , \new_[5177]_ , \new_[5178]_ ,
    \new_[5179]_ , \new_[5180]_ , \new_[5181]_ , \new_[5182]_ ,
    \new_[5183]_ , \new_[5184]_ , \new_[5185]_ , \new_[5186]_ ,
    \new_[5187]_ , \new_[5188]_ , \new_[5189]_ , \new_[5190]_ ,
    \new_[5191]_ , \new_[5192]_ , \new_[5193]_ , \new_[5194]_ ,
    \new_[5195]_ , \new_[5196]_ , \new_[5197]_ , \new_[5198]_ ,
    \new_[5199]_ , \new_[5200]_ , \new_[5201]_ , \new_[5202]_ ,
    \new_[5203]_ , \new_[5204]_ , \new_[5205]_ , \new_[5206]_ ,
    \new_[5207]_ , \new_[5208]_ , \new_[5209]_ , \new_[5210]_ ,
    \new_[5211]_ , \new_[5212]_ , \new_[5213]_ , \new_[5214]_ ,
    \new_[5215]_ , \new_[5216]_ , \new_[5217]_ , \new_[5218]_ ,
    \new_[5219]_ , \new_[5220]_ , \new_[5221]_ , \new_[5222]_ ,
    \new_[5223]_ , \new_[5224]_ , \new_[5225]_ , \new_[5226]_ ,
    \new_[5227]_ , \new_[5228]_ , \new_[5229]_ , \new_[5230]_ ,
    \new_[5231]_ , \new_[5232]_ , \new_[5233]_ , \new_[5234]_ ,
    \new_[5235]_ , \new_[5236]_ , \new_[5237]_ , \new_[5238]_ ,
    \new_[5239]_ , \new_[5240]_ , \new_[5241]_ , \new_[5242]_ ,
    \new_[5243]_ , \new_[5244]_ , \new_[5245]_ , \new_[5246]_ ,
    \new_[5247]_ , \new_[5248]_ , \new_[5249]_ , \new_[5250]_ ,
    \new_[5251]_ , \new_[5252]_ , \new_[5253]_ , \new_[5254]_ ,
    \new_[5255]_ , \new_[5256]_ , \new_[5257]_ , \new_[5258]_ ,
    \new_[5259]_ , \new_[5260]_ , \new_[5261]_ , \new_[5262]_ ,
    \new_[5263]_ , \new_[5264]_ , \new_[5265]_ , \new_[5266]_ ,
    \new_[5267]_ , \new_[5268]_ , \new_[5269]_ , \new_[5270]_ ,
    \new_[5271]_ , \new_[5272]_ , \new_[5273]_ , \new_[5274]_ ,
    \new_[5275]_ , \new_[5276]_ , \new_[5277]_ , \new_[5278]_ ,
    \new_[5279]_ , \new_[5280]_ , \new_[5281]_ , \new_[5282]_ ,
    \new_[5283]_ , \new_[5284]_ , \new_[5285]_ , \new_[5286]_ ,
    \new_[5287]_ , \new_[5288]_ , \new_[5289]_ , \new_[5290]_ ,
    \new_[5291]_ , \new_[5292]_ , \new_[5293]_ , \new_[5294]_ ,
    \new_[5295]_ , \new_[5296]_ , \new_[5297]_ , \new_[5298]_ ,
    \new_[5299]_ , \new_[5300]_ , \new_[5301]_ , \new_[5302]_ ,
    \new_[5303]_ , \new_[5304]_ , \new_[5305]_ , \new_[5306]_ ,
    \new_[5307]_ , \new_[5308]_ , \new_[5310]_ , \new_[5311]_ ,
    \new_[5312]_ , \new_[5313]_ , \new_[5314]_ , \new_[5315]_ ,
    \new_[5316]_ , \new_[5317]_ , \new_[5318]_ , \new_[5319]_ ,
    \new_[5320]_ , \new_[5321]_ , \new_[5322]_ , \new_[5323]_ ,
    \new_[5324]_ , \new_[5325]_ , \new_[5326]_ , \new_[5327]_ ,
    \new_[5328]_ , \new_[5329]_ , \new_[5330]_ , \new_[5331]_ ,
    \new_[5332]_ , \new_[5333]_ , \new_[5334]_ , \new_[5335]_ ,
    \new_[5336]_ , \new_[5337]_ , \new_[5338]_ , \new_[5339]_ ,
    \new_[5340]_ , \new_[5341]_ , \new_[5342]_ , \new_[5343]_ ,
    \new_[5344]_ , \new_[5345]_ , \new_[5346]_ , \new_[5347]_ ,
    \new_[5348]_ , \new_[5349]_ , \new_[5350]_ , \new_[5351]_ ,
    \new_[5352]_ , \new_[5353]_ , \new_[5354]_ , \new_[5355]_ ,
    \new_[5356]_ , \new_[5357]_ , \new_[5358]_ , \new_[5359]_ ,
    \new_[5360]_ , \new_[5361]_ , \new_[5362]_ , \new_[5363]_ ,
    \new_[5364]_ , \new_[5365]_ , \new_[5366]_ , \new_[5367]_ ,
    \new_[5368]_ , \new_[5369]_ , \new_[5370]_ , \new_[5371]_ ,
    \new_[5372]_ , \new_[5373]_ , \new_[5374]_ , \new_[5375]_ ,
    \new_[5376]_ , \new_[5377]_ , \new_[5378]_ , \new_[5379]_ ,
    \new_[5380]_ , \new_[5381]_ , \new_[5382]_ , \new_[5383]_ ,
    \new_[5384]_ , \new_[5385]_ , \new_[5386]_ , \new_[5387]_ ,
    \new_[5388]_ , \new_[5389]_ , \new_[5390]_ , \new_[5391]_ ,
    \new_[5392]_ , \new_[5393]_ , \new_[5394]_ , \new_[5395]_ ,
    \new_[5396]_ , \new_[5397]_ , \new_[5398]_ , \new_[5399]_ ,
    \new_[5400]_ , \new_[5401]_ , \new_[5402]_ , \new_[5403]_ ,
    \new_[5404]_ , \new_[5405]_ , \new_[5406]_ , \new_[5407]_ ,
    \new_[5408]_ , \new_[5409]_ , \new_[5410]_ , \new_[5411]_ ,
    \new_[5412]_ , \new_[5413]_ , \new_[5414]_ , \new_[5415]_ ,
    \new_[5416]_ , \new_[5417]_ , \new_[5418]_ , \new_[5419]_ ,
    \new_[5420]_ , \new_[5421]_ , \new_[5422]_ , \new_[5423]_ ,
    \new_[5424]_ , \new_[5425]_ , \new_[5426]_ , \new_[5427]_ ,
    \new_[5428]_ , \new_[5429]_ , \new_[5430]_ , \new_[5431]_ ,
    \new_[5432]_ , \new_[5433]_ , \new_[5434]_ , \new_[5435]_ ,
    \new_[5436]_ , \new_[5437]_ , \new_[5438]_ , \new_[5439]_ ,
    \new_[5440]_ , \new_[5441]_ , \new_[5442]_ , \new_[5443]_ ,
    \new_[5444]_ , \new_[5445]_ , \new_[5446]_ , \new_[5447]_ ,
    \new_[5448]_ , \new_[5449]_ , \new_[5450]_ , \new_[5451]_ ,
    \new_[5452]_ , \new_[5453]_ , \new_[5454]_ , \new_[5455]_ ,
    \new_[5456]_ , \new_[5457]_ , \new_[5458]_ , \new_[5459]_ ,
    \new_[5460]_ , \new_[5461]_ , \new_[5462]_ , \new_[5463]_ ,
    \new_[5464]_ , \new_[5465]_ , \new_[5466]_ , \new_[5467]_ ,
    \new_[5468]_ , \new_[5469]_ , \new_[5470]_ , \new_[5471]_ ,
    \new_[5472]_ , \new_[5473]_ , \new_[5474]_ , \new_[5475]_ ,
    \new_[5476]_ , \new_[5477]_ , \new_[5478]_ , \new_[5479]_ ,
    \new_[5480]_ , \new_[5481]_ , \new_[5482]_ , \new_[5483]_ ,
    \new_[5484]_ , \new_[5485]_ , \new_[5486]_ , \new_[5487]_ ,
    \new_[5488]_ , \new_[5489]_ , \new_[5490]_ , \new_[5491]_ ,
    \new_[5492]_ , \new_[5493]_ , \new_[5494]_ , \new_[5495]_ ,
    \new_[5496]_ , \new_[5497]_ , \new_[5498]_ , \new_[5499]_ ,
    \new_[5500]_ , \new_[5501]_ , \new_[5502]_ , \new_[5503]_ ,
    \new_[5504]_ , \new_[5505]_ , \new_[5506]_ , \new_[5507]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5510]_ , \new_[5511]_ ,
    \new_[5512]_ , \new_[5513]_ , \new_[5514]_ , \new_[5515]_ ,
    \new_[5516]_ , \new_[5517]_ , \new_[5518]_ , \new_[5519]_ ,
    \new_[5520]_ , \new_[5521]_ , \new_[5522]_ , \new_[5523]_ ,
    \new_[5524]_ , \new_[5525]_ , \new_[5526]_ , \new_[5527]_ ,
    \new_[5528]_ , \new_[5529]_ , \new_[5530]_ , \new_[5531]_ ,
    \new_[5532]_ , \new_[5533]_ , \new_[5534]_ , \new_[5535]_ ,
    \new_[5536]_ , \new_[5537]_ , \new_[5538]_ , \new_[5539]_ ,
    \new_[5540]_ , \new_[5541]_ , \new_[5542]_ , \new_[5543]_ ,
    \new_[5544]_ , \new_[5545]_ , \new_[5546]_ , \new_[5547]_ ,
    \new_[5548]_ , \new_[5549]_ , \new_[5550]_ , \new_[5551]_ ,
    \new_[5552]_ , \new_[5553]_ , \new_[5554]_ , \new_[5555]_ ,
    \new_[5556]_ , \new_[5557]_ , \new_[5558]_ , \new_[5559]_ ,
    \new_[5560]_ , \new_[5561]_ , \new_[5562]_ , \new_[5563]_ ,
    \new_[5564]_ , \new_[5565]_ , \new_[5566]_ , \new_[5567]_ ,
    \new_[5568]_ , \new_[5569]_ , \new_[5570]_ , \new_[5571]_ ,
    \new_[5572]_ , \new_[5573]_ , \new_[5574]_ , \new_[5575]_ ,
    \new_[5576]_ , \new_[5577]_ , \new_[5578]_ , \new_[5579]_ ,
    \new_[5580]_ , \new_[5581]_ , \new_[5582]_ , \new_[5583]_ ,
    \new_[5584]_ , \new_[5585]_ , \new_[5586]_ , \new_[5587]_ ,
    \new_[5588]_ , \new_[5589]_ , \new_[5590]_ , \new_[5591]_ ,
    \new_[5592]_ , \new_[5593]_ , \new_[5594]_ , \new_[5595]_ ,
    \new_[5596]_ , \new_[5597]_ , \new_[5598]_ , \new_[5599]_ ,
    \new_[5600]_ , \new_[5601]_ , \new_[5602]_ , \new_[5603]_ ,
    \new_[5604]_ , \new_[5605]_ , \new_[5606]_ , \new_[5607]_ ,
    \new_[5608]_ , \new_[5609]_ , \new_[5610]_ , \new_[5611]_ ,
    \new_[5612]_ , \new_[5613]_ , \new_[5614]_ , \new_[5615]_ ,
    \new_[5616]_ , \new_[5617]_ , \new_[5618]_ , \new_[5619]_ ,
    \new_[5620]_ , \new_[5621]_ , \new_[5622]_ , \new_[5623]_ ,
    \new_[5624]_ , \new_[5625]_ , \new_[5626]_ , \new_[5627]_ ,
    \new_[5628]_ , \new_[5629]_ , \new_[5630]_ , \new_[5631]_ ,
    \new_[5632]_ , \new_[5633]_ , \new_[5634]_ , \new_[5635]_ ,
    \new_[5636]_ , \new_[5637]_ , \new_[5638]_ , \new_[5639]_ ,
    \new_[5640]_ , \new_[5641]_ , \new_[5642]_ , \new_[5643]_ ,
    \new_[5644]_ , \new_[5645]_ , \new_[5646]_ , \new_[5647]_ ,
    \new_[5648]_ , \new_[5649]_ , \new_[5650]_ , \new_[5651]_ ,
    \new_[5652]_ , \new_[5653]_ , \new_[5654]_ , \new_[5655]_ ,
    \new_[5656]_ , \new_[5657]_ , \new_[5658]_ , \new_[5659]_ ,
    \new_[5660]_ , \new_[5661]_ , \new_[5662]_ , \new_[5663]_ ,
    \new_[5664]_ , \new_[5665]_ , \new_[5666]_ , \new_[5667]_ ,
    \new_[5668]_ , \new_[5669]_ , \new_[5670]_ , \new_[5671]_ ,
    \new_[5672]_ , \new_[5673]_ , \new_[5674]_ , \new_[5675]_ ,
    \new_[5676]_ , \new_[5677]_ , \new_[5678]_ , \new_[5679]_ ,
    \new_[5680]_ , \new_[5681]_ , \new_[5682]_ , \new_[5683]_ ,
    \new_[5684]_ , \new_[5685]_ , \new_[5686]_ , \new_[5687]_ ,
    \new_[5688]_ , \new_[5689]_ , \new_[5690]_ , \new_[5691]_ ,
    \new_[5692]_ , \new_[5693]_ , \new_[5694]_ , \new_[5695]_ ,
    \new_[5696]_ , \new_[5697]_ , \new_[5698]_ , \new_[5699]_ ,
    \new_[5700]_ , \new_[5701]_ , \new_[5702]_ , \new_[5703]_ ,
    \new_[5704]_ , \new_[5705]_ , \new_[5706]_ , \new_[5707]_ ,
    \new_[5708]_ , \new_[5709]_ , \new_[5710]_ , \new_[5711]_ ,
    \new_[5712]_ , \new_[5713]_ , \new_[5714]_ , \new_[5715]_ ,
    \new_[5716]_ , \new_[5717]_ , \new_[5718]_ , \new_[5719]_ ,
    \new_[5720]_ , \new_[5721]_ , \new_[5722]_ , \new_[5723]_ ,
    \new_[5724]_ , \new_[5725]_ , \new_[5726]_ , \new_[5727]_ ,
    \new_[5728]_ , \new_[5729]_ , \new_[5730]_ , \new_[5731]_ ,
    \new_[5732]_ , \new_[5733]_ , \new_[5734]_ , \new_[5735]_ ,
    \new_[5736]_ , \new_[5737]_ , \new_[5738]_ , \new_[5739]_ ,
    \new_[5740]_ , \new_[5741]_ , \new_[5742]_ , \new_[5743]_ ,
    \new_[5744]_ , \new_[5745]_ , \new_[5746]_ , \new_[5747]_ ,
    \new_[5748]_ , \new_[5749]_ , \new_[5750]_ , \new_[5751]_ ,
    \new_[5752]_ , \new_[5753]_ , \new_[5754]_ , \new_[5755]_ ,
    \new_[5756]_ , \new_[5757]_ , \new_[5758]_ , \new_[5759]_ ,
    \new_[5760]_ , \new_[5761]_ , \new_[5762]_ , \new_[5763]_ ,
    \new_[5764]_ , \new_[5765]_ , \new_[5766]_ , \new_[5767]_ ,
    \new_[5768]_ , \new_[5769]_ , \new_[5770]_ , \new_[5771]_ ,
    \new_[5772]_ , \new_[5773]_ , \new_[5774]_ , \new_[5775]_ ,
    \new_[5776]_ , \new_[5777]_ , \new_[5778]_ , \new_[5779]_ ,
    \new_[5780]_ , \new_[5781]_ , \new_[5782]_ , \new_[5783]_ ,
    \new_[5784]_ , \new_[5785]_ , \new_[5786]_ , \new_[5787]_ ,
    \new_[5788]_ , \new_[5789]_ , \new_[5790]_ , \new_[5791]_ ,
    \new_[5792]_ , \new_[5793]_ , \new_[5794]_ , \new_[5795]_ ,
    \new_[5796]_ , \new_[5797]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5800]_ , \new_[5801]_ , \new_[5802]_ , \new_[5803]_ ,
    \new_[5804]_ , \new_[5805]_ , \new_[5806]_ , \new_[5807]_ ,
    \new_[5808]_ , \new_[5809]_ , \new_[5810]_ , \new_[5811]_ ,
    \new_[5812]_ , \new_[5813]_ , \new_[5814]_ , \new_[5815]_ ,
    \new_[5816]_ , \new_[5817]_ , \new_[5818]_ , \new_[5819]_ ,
    \new_[5820]_ , \new_[5821]_ , \new_[5822]_ , \new_[5823]_ ,
    \new_[5824]_ , \new_[5825]_ , \new_[5826]_ , \new_[5827]_ ,
    \new_[5828]_ , \new_[5829]_ , \new_[5830]_ , \new_[5831]_ ,
    \new_[5832]_ , \new_[5833]_ , \new_[5834]_ , \new_[5835]_ ,
    \new_[5836]_ , \new_[5837]_ , \new_[5838]_ , \new_[5839]_ ,
    \new_[5840]_ , \new_[5841]_ , \new_[5842]_ , \new_[5843]_ ,
    \new_[5844]_ , \new_[5845]_ , \new_[5846]_ , \new_[5847]_ ,
    \new_[5848]_ , \new_[5849]_ , \new_[5850]_ , \new_[5851]_ ,
    \new_[5852]_ , \new_[5853]_ , \new_[5854]_ , \new_[5855]_ ,
    \new_[5856]_ , \new_[5857]_ , \new_[5858]_ , \new_[5859]_ ,
    \new_[5860]_ , \new_[5861]_ , \new_[5862]_ , \new_[5863]_ ,
    \new_[5864]_ , \new_[5865]_ , \new_[5866]_ , \new_[5867]_ ,
    \new_[5868]_ , \new_[5869]_ , \new_[5870]_ , \new_[5871]_ ,
    \new_[5872]_ , \new_[5873]_ , \new_[5874]_ , \new_[5875]_ ,
    \new_[5876]_ , \new_[5877]_ , \new_[5878]_ , \new_[5879]_ ,
    \new_[5880]_ , \new_[5881]_ , \new_[5882]_ , \new_[5883]_ ,
    \new_[5884]_ , \new_[5885]_ , \new_[5886]_ , \new_[5887]_ ,
    \new_[5888]_ , \new_[5889]_ , \new_[5890]_ , \new_[5891]_ ,
    \new_[5892]_ , \new_[5893]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5896]_ , \new_[5897]_ , \new_[5898]_ , \new_[5899]_ ,
    \new_[5900]_ , \new_[5901]_ , \new_[5902]_ , \new_[5903]_ ,
    \new_[5904]_ , \new_[5905]_ , \new_[5906]_ , \new_[5907]_ ,
    \new_[5908]_ , \new_[5909]_ , \new_[5910]_ , \new_[5911]_ ,
    \new_[5912]_ , \new_[5913]_ , \new_[5914]_ , \new_[5915]_ ,
    \new_[5916]_ , \new_[5917]_ , \new_[5918]_ , \new_[5919]_ ,
    \new_[5920]_ , \new_[5921]_ , \new_[5922]_ , \new_[5923]_ ,
    \new_[5924]_ , \new_[5925]_ , \new_[5926]_ , \new_[5927]_ ,
    \new_[5928]_ , \new_[5929]_ , \new_[5930]_ , \new_[5931]_ ,
    \new_[5932]_ , \new_[5933]_ , \new_[5934]_ , \new_[5935]_ ,
    \new_[5936]_ , \new_[5937]_ , \new_[5938]_ , \new_[5939]_ ,
    \new_[5940]_ , \new_[5941]_ , \new_[5942]_ , \new_[5943]_ ,
    \new_[5944]_ , \new_[5945]_ , \new_[5946]_ , \new_[5947]_ ,
    \new_[5948]_ , \new_[5949]_ , \new_[5950]_ , \new_[5951]_ ,
    \new_[5952]_ , \new_[5953]_ , \new_[5954]_ , \new_[5955]_ ,
    \new_[5956]_ , \new_[5957]_ , \new_[5958]_ , \new_[5959]_ ,
    \new_[5960]_ , \new_[5961]_ , \new_[5962]_ , \new_[5963]_ ,
    \new_[5964]_ , \new_[5965]_ , \new_[5966]_ , \new_[5967]_ ,
    \new_[5968]_ , \new_[5969]_ , \new_[5970]_ , \new_[5971]_ ,
    \new_[5972]_ , \new_[5973]_ , \new_[5974]_ , \new_[5975]_ ,
    \new_[5976]_ , \new_[5977]_ , \new_[5978]_ , \new_[5979]_ ,
    \new_[5980]_ , \new_[5981]_ , \new_[5982]_ , \new_[5983]_ ,
    \new_[5984]_ , \new_[5985]_ , \new_[5986]_ , \new_[5987]_ ,
    \new_[5988]_ , \new_[5989]_ , \new_[5990]_ , \new_[5991]_ ,
    \new_[5992]_ , \new_[5993]_ , \new_[5994]_ , \new_[5995]_ ,
    \new_[5996]_ , \new_[5997]_ , \new_[5998]_ , \new_[5999]_ ,
    \new_[6000]_ , \new_[6001]_ , \new_[6002]_ , \new_[6003]_ ,
    \new_[6004]_ , \new_[6005]_ , \new_[6006]_ , \new_[6007]_ ,
    \new_[6008]_ , \new_[6009]_ , \new_[6010]_ , \new_[6011]_ ,
    \new_[6012]_ , \new_[6013]_ , \new_[6014]_ , \new_[6015]_ ,
    \new_[6016]_ , \new_[6017]_ , \new_[6018]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6021]_ , \new_[6022]_ , \new_[6023]_ ,
    \new_[6024]_ , \new_[6025]_ , \new_[6026]_ , \new_[6027]_ ,
    \new_[6028]_ , \new_[6029]_ , \new_[6030]_ , \new_[6031]_ ,
    \new_[6032]_ , \new_[6033]_ , \new_[6034]_ , \new_[6035]_ ,
    \new_[6036]_ , \new_[6037]_ , \new_[6038]_ , \new_[6039]_ ,
    \new_[6040]_ , \new_[6041]_ , \new_[6042]_ , \new_[6043]_ ,
    \new_[6044]_ , \new_[6045]_ , \new_[6046]_ , \new_[6047]_ ,
    \new_[6048]_ , \new_[6049]_ , \new_[6050]_ , \new_[6051]_ ,
    \new_[6052]_ , \new_[6053]_ , \new_[6054]_ , \new_[6055]_ ,
    \new_[6056]_ , \new_[6057]_ , \new_[6058]_ , \new_[6059]_ ,
    \new_[6060]_ , \new_[6061]_ , \new_[6062]_ , \new_[6063]_ ,
    \new_[6064]_ , \new_[6065]_ , \new_[6066]_ , \new_[6067]_ ,
    \new_[6068]_ , \new_[6069]_ , \new_[6070]_ , \new_[6071]_ ,
    \new_[6072]_ , \new_[6073]_ , \new_[6074]_ , \new_[6075]_ ,
    \new_[6076]_ , \new_[6077]_ , \new_[6078]_ , \new_[6079]_ ,
    \new_[6080]_ , \new_[6081]_ , \new_[6082]_ , \new_[6083]_ ,
    \new_[6084]_ , \new_[6085]_ , \new_[6086]_ , \new_[6087]_ ,
    \new_[6088]_ , \new_[6089]_ , \new_[6090]_ , \new_[6091]_ ,
    \new_[6092]_ , \new_[6093]_ , \new_[6094]_ , \new_[6095]_ ,
    \new_[6096]_ , \new_[6097]_ , \new_[6098]_ , \new_[6099]_ ,
    \new_[6100]_ , \new_[6101]_ , \new_[6102]_ , \new_[6103]_ ,
    \new_[6104]_ , \new_[6105]_ , \new_[6106]_ , \new_[6107]_ ,
    \new_[6108]_ , \new_[6109]_ , \new_[6110]_ , \new_[6111]_ ,
    \new_[6112]_ , \new_[6113]_ , \new_[6114]_ , \new_[6115]_ ,
    \new_[6116]_ , \new_[6117]_ , \new_[6118]_ , \new_[6119]_ ,
    \new_[6120]_ , \new_[6121]_ , \new_[6122]_ , \new_[6123]_ ,
    \new_[6124]_ , \new_[6125]_ , \new_[6126]_ , \new_[6127]_ ,
    \new_[6128]_ , \new_[6129]_ , \new_[6130]_ , \new_[6131]_ ,
    \new_[6132]_ , \new_[6133]_ , \new_[6134]_ , \new_[6135]_ ,
    \new_[6136]_ , \new_[6137]_ , \new_[6138]_ , \new_[6139]_ ,
    \new_[6140]_ , \new_[6141]_ , \new_[6142]_ , \new_[6143]_ ,
    \new_[6144]_ , \new_[6145]_ , \new_[6146]_ , \new_[6147]_ ,
    \new_[6148]_ , \new_[6149]_ , \new_[6150]_ , \new_[6151]_ ,
    \new_[6152]_ , \new_[6153]_ , \new_[6155]_ , \new_[6156]_ ,
    \new_[6157]_ , \new_[6158]_ , \new_[6159]_ , \new_[6160]_ ,
    \new_[6161]_ , \new_[6162]_ , \new_[6163]_ , \new_[6164]_ ,
    \new_[6165]_ , \new_[6166]_ , \new_[6167]_ , \new_[6168]_ ,
    \new_[6169]_ , \new_[6170]_ , \new_[6171]_ , \new_[6172]_ ,
    \new_[6173]_ , \new_[6174]_ , \new_[6175]_ , \new_[6176]_ ,
    \new_[6177]_ , \new_[6178]_ , \new_[6179]_ , \new_[6180]_ ,
    \new_[6181]_ , \new_[6182]_ , \new_[6183]_ , \new_[6184]_ ,
    \new_[6185]_ , \new_[6186]_ , \new_[6187]_ , \new_[6188]_ ,
    \new_[6189]_ , \new_[6190]_ , \new_[6191]_ , \new_[6192]_ ,
    \new_[6193]_ , \new_[6194]_ , \new_[6195]_ , \new_[6196]_ ,
    \new_[6197]_ , \new_[6198]_ , \new_[6199]_ , \new_[6200]_ ,
    \new_[6201]_ , \new_[6202]_ , \new_[6203]_ , \new_[6204]_ ,
    \new_[6205]_ , \new_[6206]_ , \new_[6207]_ , \new_[6208]_ ,
    \new_[6209]_ , \new_[6210]_ , \new_[6211]_ , \new_[6212]_ ,
    \new_[6213]_ , \new_[6214]_ , \new_[6215]_ , \new_[6216]_ ,
    \new_[6217]_ , \new_[6218]_ , \new_[6219]_ , \new_[6220]_ ,
    \new_[6221]_ , \new_[6222]_ , \new_[6223]_ , \new_[6224]_ ,
    \new_[6225]_ , \new_[6226]_ , \new_[6227]_ , \new_[6228]_ ,
    \new_[6229]_ , \new_[6231]_ , \new_[6232]_ , \new_[6233]_ ,
    \new_[6234]_ , \new_[6235]_ , \new_[6236]_ , \new_[6237]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6240]_ , \new_[6241]_ ,
    \new_[6242]_ , \new_[6243]_ , \new_[6244]_ , \new_[6245]_ ,
    \new_[6246]_ , \new_[6247]_ , \new_[6248]_ , \new_[6249]_ ,
    \new_[6250]_ , \new_[6251]_ , \new_[6252]_ , \new_[6254]_ ,
    \new_[6255]_ , \new_[6256]_ , \new_[6257]_ , \new_[6258]_ ,
    \new_[6259]_ , \new_[6260]_ , \new_[6261]_ , \new_[6262]_ ,
    \new_[6263]_ , \new_[6264]_ , \new_[6265]_ , \new_[6266]_ ,
    \new_[6267]_ , \new_[6268]_ , \new_[6269]_ , \new_[6270]_ ,
    \new_[6271]_ , \new_[6272]_ , \new_[6273]_ , \new_[6274]_ ,
    \new_[6275]_ , \new_[6276]_ , \new_[6277]_ , \new_[6278]_ ,
    \new_[6279]_ , \new_[6280]_ , \new_[6281]_ , \new_[6282]_ ,
    \new_[6283]_ , \new_[6284]_ , \new_[6285]_ , \new_[6286]_ ,
    \new_[6287]_ , \new_[6288]_ , \new_[6289]_ , \new_[6290]_ ,
    \new_[6291]_ , \new_[6292]_ , \new_[6293]_ , \new_[6294]_ ,
    \new_[6295]_ , \new_[6296]_ , \new_[6297]_ , \new_[6298]_ ,
    \new_[6299]_ , \new_[6300]_ , \new_[6301]_ , \new_[6302]_ ,
    \new_[6303]_ , \new_[6304]_ , \new_[6305]_ , \new_[6306]_ ,
    \new_[6307]_ , \new_[6308]_ , \new_[6309]_ , \new_[6310]_ ,
    \new_[6311]_ , \new_[6312]_ , \new_[6313]_ , \new_[6314]_ ,
    \new_[6315]_ , \new_[6316]_ , \new_[6317]_ , \new_[6318]_ ,
    \new_[6319]_ , \new_[6320]_ , \new_[6321]_ , \new_[6322]_ ,
    \new_[6323]_ , \new_[6324]_ , \new_[6325]_ , \new_[6326]_ ,
    \new_[6327]_ , \new_[6328]_ , \new_[6329]_ , \new_[6330]_ ,
    \new_[6331]_ , \new_[6332]_ , \new_[6333]_ , \new_[6334]_ ,
    \new_[6335]_ , \new_[6336]_ , \new_[6337]_ , \new_[6338]_ ,
    \new_[6339]_ , \new_[6340]_ , \new_[6341]_ , \new_[6342]_ ,
    \new_[6343]_ , \new_[6344]_ , \new_[6345]_ , \new_[6346]_ ,
    \new_[6347]_ , \new_[6348]_ , \new_[6349]_ , \new_[6350]_ ,
    \new_[6351]_ , \new_[6352]_ , \new_[6353]_ , \new_[6354]_ ,
    \new_[6355]_ , \new_[6356]_ , \new_[6357]_ , \new_[6358]_ ,
    \new_[6359]_ , \new_[6360]_ , \new_[6361]_ , \new_[6362]_ ,
    \new_[6363]_ , \new_[6364]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6367]_ , \new_[6368]_ , \new_[6369]_ , \new_[6370]_ ,
    \new_[6371]_ , \new_[6372]_ , \new_[6373]_ , \new_[6374]_ ,
    \new_[6375]_ , \new_[6376]_ , \new_[6377]_ , \new_[6378]_ ,
    \new_[6379]_ , \new_[6380]_ , \new_[6381]_ , \new_[6382]_ ,
    \new_[6384]_ , \new_[6385]_ , \new_[6386]_ , \new_[6387]_ ,
    \new_[6388]_ , \new_[6389]_ , \new_[6390]_ , \new_[6391]_ ,
    \new_[6392]_ , \new_[6393]_ , \new_[6394]_ , \new_[6395]_ ,
    \new_[6396]_ , \new_[6397]_ , \new_[6398]_ , \new_[6399]_ ,
    \new_[6400]_ , \new_[6401]_ , \new_[6402]_ , \new_[6403]_ ,
    \new_[6404]_ , \new_[6405]_ , \new_[6406]_ , \new_[6407]_ ,
    \new_[6408]_ , \new_[6409]_ , \new_[6410]_ , \new_[6411]_ ,
    \new_[6412]_ , \new_[6413]_ , \new_[6414]_ , \new_[6415]_ ,
    \new_[6416]_ , \new_[6417]_ , \new_[6418]_ , \new_[6419]_ ,
    \new_[6420]_ , \new_[6421]_ , \new_[6422]_ , \new_[6423]_ ,
    \new_[6424]_ , \new_[6425]_ , \new_[6426]_ , \new_[6427]_ ,
    \new_[6428]_ , \new_[6429]_ , \new_[6430]_ , \new_[6431]_ ,
    \new_[6432]_ , \new_[6433]_ , \new_[6434]_ , \new_[6435]_ ,
    \new_[6436]_ , \new_[6437]_ , \new_[6438]_ , \new_[6439]_ ,
    \new_[6440]_ , \new_[6441]_ , \new_[6442]_ , \new_[6443]_ ,
    \new_[6444]_ , \new_[6445]_ , \new_[6446]_ , \new_[6447]_ ,
    \new_[6448]_ , \new_[6449]_ , \new_[6450]_ , \new_[6451]_ ,
    \new_[6452]_ , \new_[6453]_ , \new_[6454]_ , \new_[6455]_ ,
    \new_[6456]_ , \new_[6457]_ , \new_[6458]_ , \new_[6459]_ ,
    \new_[6460]_ , \new_[6461]_ , \new_[6462]_ , \new_[6463]_ ,
    \new_[6464]_ , \new_[6465]_ , \new_[6466]_ , \new_[6467]_ ,
    \new_[6468]_ , \new_[6469]_ , \new_[6470]_ , \new_[6471]_ ,
    \new_[6472]_ , \new_[6473]_ , \new_[6474]_ , \new_[6475]_ ,
    \new_[6476]_ , \new_[6477]_ , \new_[6478]_ , \new_[6479]_ ,
    \new_[6480]_ , \new_[6481]_ , \new_[6482]_ , \new_[6483]_ ,
    \new_[6484]_ , \new_[6485]_ , \new_[6486]_ , \new_[6487]_ ,
    \new_[6488]_ , \new_[6489]_ , \new_[6490]_ , \new_[6491]_ ,
    \new_[6492]_ , \new_[6493]_ , \new_[6494]_ , \new_[6495]_ ,
    \new_[6496]_ , \new_[6497]_ , \new_[6498]_ , \new_[6499]_ ,
    \new_[6500]_ , \new_[6501]_ , \new_[6502]_ , \new_[6503]_ ,
    \new_[6504]_ , \new_[6505]_ , \new_[6506]_ , \new_[6507]_ ,
    \new_[6508]_ , \new_[6509]_ , \new_[6510]_ , \new_[6511]_ ,
    \new_[6512]_ , \new_[6513]_ , \new_[6514]_ , \new_[6515]_ ,
    \new_[6516]_ , \new_[6517]_ , \new_[6518]_ , \new_[6519]_ ,
    \new_[6520]_ , \new_[6521]_ , \new_[6522]_ , \new_[6523]_ ,
    \new_[6524]_ , \new_[6525]_ , \new_[6526]_ , \new_[6527]_ ,
    \new_[6528]_ , \new_[6529]_ , \new_[6530]_ , \new_[6531]_ ,
    \new_[6532]_ , \new_[6533]_ , \new_[6534]_ , \new_[6535]_ ,
    \new_[6536]_ , \new_[6537]_ , \new_[6538]_ , \new_[6539]_ ,
    \new_[6540]_ , \new_[6541]_ , \new_[6542]_ , \new_[6543]_ ,
    \new_[6544]_ , \new_[6545]_ , \new_[6546]_ , \new_[6547]_ ,
    \new_[6548]_ , \new_[6549]_ , \new_[6550]_ , \new_[6551]_ ,
    \new_[6552]_ , \new_[6553]_ , \new_[6554]_ , \new_[6555]_ ,
    \new_[6556]_ , \new_[6557]_ , \new_[6558]_ , \new_[6559]_ ,
    \new_[6560]_ , \new_[6561]_ , \new_[6563]_ , \new_[6564]_ ,
    \new_[6565]_ , \new_[6566]_ , \new_[6567]_ , \new_[6568]_ ,
    \new_[6569]_ , \new_[6570]_ , \new_[6571]_ , \new_[6572]_ ,
    \new_[6573]_ , \new_[6574]_ , \new_[6575]_ , \new_[6576]_ ,
    \new_[6577]_ , \new_[6578]_ , \new_[6580]_ , \new_[6581]_ ,
    \new_[6582]_ , \new_[6583]_ , \new_[6584]_ , \new_[6586]_ ,
    \new_[6587]_ , \new_[6588]_ , \new_[6589]_ , \new_[6590]_ ,
    \new_[6591]_ , \new_[6592]_ , \new_[6593]_ , \new_[6595]_ ,
    \new_[6596]_ , \new_[6597]_ , \new_[6598]_ , \new_[6599]_ ,
    \new_[6600]_ , \new_[6601]_ , \new_[6602]_ , \new_[6603]_ ,
    \new_[6604]_ , \new_[6605]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6608]_ , \new_[6609]_ , \new_[6610]_ , \new_[6611]_ ,
    \new_[6612]_ , \new_[6613]_ , \new_[6614]_ , \new_[6615]_ ,
    \new_[6616]_ , \new_[6617]_ , \new_[6618]_ , \new_[6619]_ ,
    \new_[6620]_ , \new_[6621]_ , \new_[6622]_ , \new_[6623]_ ,
    \new_[6624]_ , \new_[6625]_ , \new_[6626]_ , \new_[6627]_ ,
    \new_[6629]_ , \new_[6630]_ , \new_[6631]_ , \new_[6632]_ ,
    \new_[6633]_ , \new_[6634]_ , \new_[6635]_ , \new_[6637]_ ,
    \new_[6638]_ , \new_[6639]_ , \new_[6640]_ , \new_[6641]_ ,
    \new_[6642]_ , \new_[6643]_ , \new_[6644]_ , \new_[6645]_ ,
    \new_[6646]_ , \new_[6647]_ , \new_[6648]_ , \new_[6649]_ ,
    \new_[6651]_ , \new_[6652]_ , \new_[6653]_ , \new_[6654]_ ,
    \new_[6655]_ , \new_[6656]_ , \new_[6657]_ , \new_[6658]_ ,
    \new_[6659]_ , \new_[6660]_ , \new_[6661]_ , \new_[6662]_ ,
    \new_[6663]_ , \new_[6664]_ , \new_[6665]_ , \new_[6666]_ ,
    \new_[6667]_ , \new_[6668]_ , \new_[6669]_ , \new_[6670]_ ,
    \new_[6671]_ , \new_[6672]_ , \new_[6673]_ , \new_[6674]_ ,
    \new_[6675]_ , \new_[6676]_ , \new_[6677]_ , \new_[6678]_ ,
    \new_[6679]_ , \new_[6680]_ , \new_[6681]_ , \new_[6682]_ ,
    \new_[6683]_ , \new_[6684]_ , \new_[6685]_ , \new_[6686]_ ,
    \new_[6687]_ , \new_[6688]_ , \new_[6689]_ , \new_[6690]_ ,
    \new_[6691]_ , \new_[6692]_ , \new_[6693]_ , \new_[6694]_ ,
    \new_[6695]_ , \new_[6696]_ , \new_[6697]_ , \new_[6698]_ ,
    \new_[6699]_ , \new_[6700]_ , \new_[6701]_ , \new_[6702]_ ,
    \new_[6703]_ , \new_[6704]_ , \new_[6705]_ , \new_[6706]_ ,
    \new_[6707]_ , \new_[6708]_ , \new_[6709]_ , \new_[6710]_ ,
    \new_[6711]_ , \new_[6712]_ , \new_[6713]_ , \new_[6714]_ ,
    \new_[6715]_ , \new_[6716]_ , \new_[6717]_ , \new_[6718]_ ,
    \new_[6719]_ , \new_[6720]_ , \new_[6721]_ , \new_[6722]_ ,
    \new_[6723]_ , \new_[6724]_ , \new_[6725]_ , \new_[6726]_ ,
    \new_[6727]_ , \new_[6728]_ , \new_[6729]_ , \new_[6730]_ ,
    \new_[6731]_ , \new_[6732]_ , \new_[6733]_ , \new_[6734]_ ,
    \new_[6735]_ , \new_[6736]_ , \new_[6737]_ , \new_[6738]_ ,
    \new_[6739]_ , \new_[6745]_ , \new_[6747]_ , \new_[6753]_ ,
    \new_[6754]_ , \new_[6756]_ , \new_[6757]_ , \new_[6758]_ ,
    \new_[6760]_ , \new_[6761]_ , \new_[6762]_ , \new_[6764]_ ,
    \new_[6765]_ , \new_[6766]_ , \new_[6768]_ , \new_[6769]_ ,
    \new_[6770]_ , \new_[6771]_ , \new_[6772]_ , \new_[6773]_ ,
    \new_[6774]_ , \new_[6775]_ , \new_[6776]_ , \new_[6777]_ ,
    \new_[6778]_ , \new_[6779]_ , \new_[6780]_ , \new_[6781]_ ,
    \new_[6782]_ , \new_[6783]_ , \new_[6784]_ , \new_[6785]_ ,
    \new_[6786]_ , \new_[6787]_ , \new_[6788]_ , \new_[6789]_ ,
    \new_[6790]_ , \new_[6791]_ , \new_[6792]_ , \new_[6793]_ ,
    \new_[6794]_ , \new_[6795]_ , \new_[6796]_ , \new_[6797]_ ,
    \new_[6798]_ , \new_[6799]_ , \new_[6800]_ , \new_[6801]_ ,
    \new_[6802]_ , \new_[6803]_ , \new_[6804]_ , \new_[6805]_ ,
    \new_[6806]_ , \new_[6807]_ , \new_[6808]_ , \new_[6809]_ ,
    \new_[6810]_ , \new_[6811]_ , \new_[6812]_ , \new_[6813]_ ,
    \new_[6814]_ , \new_[6815]_ , \new_[6816]_ , \new_[6817]_ ,
    \new_[6818]_ , \new_[6819]_ , \new_[6820]_ , \new_[6821]_ ,
    \new_[6822]_ , \new_[6823]_ , \new_[6824]_ , \new_[6825]_ ,
    \new_[6826]_ , \new_[6827]_ , \new_[6829]_ , \new_[6830]_ ,
    \new_[6831]_ , \new_[6832]_ , \new_[6834]_ , \new_[6835]_ ,
    \new_[6836]_ , \new_[6837]_ , \new_[6838]_ , \new_[6839]_ ,
    \new_[6840]_ , \new_[6841]_ , \new_[6842]_ , \new_[6843]_ ,
    \new_[6845]_ , \new_[6846]_ , \new_[6847]_ , \new_[6848]_ ,
    \new_[6849]_ , \new_[6851]_ , \new_[6852]_ , \new_[6853]_ ,
    \new_[6854]_ , \new_[6855]_ , \new_[6856]_ , \new_[6858]_ ,
    \new_[6859]_ , \new_[6860]_ , \new_[6862]_ , \new_[6863]_ ,
    \new_[6864]_ , \new_[6865]_ , \new_[6866]_ , \new_[6867]_ ,
    \new_[6868]_ , \new_[6870]_ , \new_[6871]_ , \new_[6872]_ ,
    \new_[6873]_ , \new_[6874]_ , \new_[6875]_ , \new_[6876]_ ,
    \new_[6877]_ , \new_[6879]_ , \new_[6880]_ , \new_[6881]_ ,
    \new_[6882]_ , \new_[6883]_ , \new_[6884]_ , \new_[6885]_ ,
    \new_[6886]_ , \new_[6887]_ , \new_[6888]_ , \new_[6889]_ ,
    \new_[6890]_ , \new_[6891]_ , \new_[6892]_ , \new_[6893]_ ,
    \new_[6894]_ , \new_[6895]_ , \new_[6897]_ , \new_[6898]_ ,
    \new_[6899]_ , \new_[6900]_ , \new_[6901]_ , \new_[6902]_ ,
    \new_[6903]_ , \new_[6904]_ , \new_[6906]_ , \new_[6907]_ ,
    \new_[6908]_ , \new_[6909]_ , \new_[6910]_ , \new_[6911]_ ,
    \new_[6912]_ , \new_[6913]_ , \new_[6914]_ , \new_[6915]_ ,
    \new_[6916]_ , \new_[6917]_ , \new_[6918]_ , \new_[6919]_ ,
    \new_[6920]_ , \new_[6921]_ , \new_[6922]_ , \new_[6923]_ ,
    \new_[6924]_ , \new_[6925]_ , \new_[6926]_ , \new_[6927]_ ,
    \new_[6928]_ , \new_[6929]_ , \new_[6930]_ , \new_[6931]_ ,
    \new_[6932]_ , \new_[6933]_ , \new_[6934]_ , \new_[6935]_ ,
    \new_[6936]_ , \new_[6937]_ , \new_[6938]_ , \new_[6939]_ ,
    \new_[6940]_ , \new_[6941]_ , \new_[6942]_ , \new_[6943]_ ,
    \new_[6944]_ , \new_[6945]_ , \new_[6946]_ , \new_[6947]_ ,
    \new_[6948]_ , \new_[6949]_ , \new_[6950]_ , \new_[6951]_ ,
    \new_[6952]_ , \new_[6953]_ , \new_[6954]_ , \new_[6955]_ ,
    \new_[6956]_ , \new_[6957]_ , \new_[6958]_ , \new_[6959]_ ,
    \new_[6960]_ , \new_[6961]_ , \new_[6962]_ , \new_[6963]_ ,
    \new_[6964]_ , \new_[6965]_ , \new_[6966]_ , \new_[6967]_ ,
    \new_[6968]_ , \new_[6969]_ , \new_[6970]_ , \new_[6971]_ ,
    \new_[6972]_ , \new_[6973]_ , \new_[6974]_ , \new_[6975]_ ,
    \new_[6976]_ , \new_[6977]_ , \new_[6978]_ , \new_[6979]_ ,
    \new_[6980]_ , \new_[6981]_ , \new_[6982]_ , \new_[6983]_ ,
    \new_[6984]_ , \new_[6985]_ , \new_[6986]_ , \new_[6987]_ ,
    \new_[6988]_ , \new_[6989]_ , \new_[6990]_ , \new_[6991]_ ,
    \new_[6992]_ , \new_[6993]_ , \new_[6994]_ , \new_[6995]_ ,
    \new_[6996]_ , \new_[6997]_ , \new_[6998]_ , \new_[6999]_ ,
    \new_[7000]_ , \new_[7001]_ , \new_[7002]_ , \new_[7003]_ ,
    \new_[7004]_ , \new_[7005]_ , \new_[7006]_ , \new_[7007]_ ,
    \new_[7008]_ , \new_[7009]_ , \new_[7010]_ , \new_[7011]_ ,
    \new_[7012]_ , \new_[7013]_ , \new_[7014]_ , \new_[7015]_ ,
    \new_[7016]_ , \new_[7017]_ , \new_[7018]_ , \new_[7019]_ ,
    \new_[7020]_ , \new_[7021]_ , \new_[7022]_ , \new_[7023]_ ,
    \new_[7024]_ , \new_[7025]_ , \new_[7026]_ , \new_[7027]_ ,
    \new_[7028]_ , \new_[7029]_ , \new_[7030]_ , \new_[7031]_ ,
    \new_[7032]_ , \new_[7033]_ , \new_[7034]_ , \new_[7035]_ ,
    \new_[7036]_ , \new_[7037]_ , \new_[7038]_ , \new_[7039]_ ,
    \new_[7040]_ , \new_[7041]_ , \new_[7042]_ , \new_[7043]_ ,
    \new_[7044]_ , \new_[7045]_ , \new_[7046]_ , \new_[7047]_ ,
    \new_[7048]_ , \new_[7049]_ , \new_[7050]_ , \new_[7051]_ ,
    \new_[7052]_ , \new_[7053]_ , \new_[7054]_ , \new_[7055]_ ,
    \new_[7056]_ , \new_[7057]_ , \new_[7058]_ , \new_[7059]_ ,
    \new_[7060]_ , \new_[7061]_ , \new_[7062]_ , \new_[7063]_ ,
    \new_[7064]_ , \new_[7065]_ , \new_[7066]_ , \new_[7067]_ ,
    \new_[7068]_ , \new_[7069]_ , \new_[7070]_ , \new_[7071]_ ,
    \new_[7072]_ , \new_[7073]_ , \new_[7074]_ , \new_[7075]_ ,
    \new_[7076]_ , \new_[7077]_ , \new_[7078]_ , \new_[7079]_ ,
    \new_[7080]_ , \new_[7081]_ , \new_[7082]_ , \new_[7083]_ ,
    \new_[7084]_ , \new_[7085]_ , \new_[7086]_ , \new_[7087]_ ,
    \new_[7088]_ , \new_[7089]_ , \new_[7090]_ , \new_[7091]_ ,
    \new_[7092]_ , \new_[7093]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7096]_ , \new_[7097]_ , \new_[7098]_ , \new_[7099]_ ,
    \new_[7100]_ , \new_[7101]_ , \new_[7102]_ , \new_[7103]_ ,
    \new_[7104]_ , \new_[7105]_ , \new_[7106]_ , \new_[7107]_ ,
    \new_[7108]_ , \new_[7109]_ , \new_[7110]_ , \new_[7111]_ ,
    \new_[7112]_ , \new_[7113]_ , \new_[7114]_ , \new_[7115]_ ,
    \new_[7116]_ , \new_[7117]_ , \new_[7118]_ , \new_[7119]_ ,
    \new_[7120]_ , \new_[7121]_ , \new_[7122]_ , \new_[7123]_ ,
    \new_[7124]_ , \new_[7125]_ , \new_[7126]_ , \new_[7127]_ ,
    \new_[7128]_ , \new_[7129]_ , \new_[7130]_ , \new_[7131]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7134]_ , \new_[7135]_ ,
    \new_[7136]_ , \new_[7137]_ , \new_[7138]_ , \new_[7139]_ ,
    \new_[7140]_ , \new_[7141]_ , \new_[7142]_ , \new_[7143]_ ,
    \new_[7144]_ , \new_[7145]_ , \new_[7146]_ , \new_[7147]_ ,
    \new_[7148]_ , \new_[7149]_ , \new_[7150]_ , \new_[7151]_ ,
    \new_[7152]_ , \new_[7153]_ , \new_[7154]_ , \new_[7155]_ ,
    \new_[7156]_ , \new_[7157]_ , \new_[7158]_ , \new_[7159]_ ,
    \new_[7160]_ , \new_[7161]_ , \new_[7162]_ , \new_[7163]_ ,
    \new_[7164]_ , \new_[7165]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7168]_ , \new_[7169]_ , \new_[7170]_ , \new_[7171]_ ,
    \new_[7172]_ , \new_[7173]_ , \new_[7174]_ , \new_[7175]_ ,
    \new_[7176]_ , \new_[7177]_ , \new_[7178]_ , \new_[7179]_ ,
    \new_[7180]_ , \new_[7181]_ , \new_[7182]_ , \new_[7183]_ ,
    \new_[7184]_ , \new_[7185]_ , \new_[7186]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7189]_ , \new_[7190]_ , \new_[7191]_ ,
    \new_[7192]_ , \new_[7193]_ , \new_[7194]_ , \new_[7195]_ ,
    \new_[7196]_ , \new_[7197]_ , \new_[7198]_ , \new_[7199]_ ,
    \new_[7200]_ , \new_[7201]_ , \new_[7202]_ , \new_[7203]_ ,
    \new_[7204]_ , \new_[7205]_ , \new_[7206]_ , \new_[7207]_ ,
    \new_[7208]_ , \new_[7209]_ , \new_[7210]_ , \new_[7211]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7214]_ , \new_[7215]_ ,
    \new_[7216]_ , \new_[7217]_ , \new_[7218]_ , \new_[7219]_ ,
    \new_[7220]_ , \new_[7221]_ , \new_[7222]_ , \new_[7223]_ ,
    \new_[7224]_ , \new_[7225]_ , \new_[7226]_ , \new_[7227]_ ,
    \new_[7228]_ , \new_[7229]_ , \new_[7230]_ , \new_[7231]_ ,
    \new_[7232]_ , \new_[7233]_ , \new_[7234]_ , \new_[7235]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7241]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7244]_ , \new_[7245]_ , \new_[7246]_ , \new_[7247]_ ,
    \new_[7248]_ , \new_[7249]_ , \new_[7250]_ , \new_[7251]_ ,
    \new_[7252]_ , \new_[7253]_ , \new_[7254]_ , \new_[7255]_ ,
    \new_[7256]_ , \new_[7257]_ , \new_[7258]_ , \new_[7259]_ ,
    \new_[7260]_ , \new_[7261]_ , \new_[7262]_ , \new_[7263]_ ,
    \new_[7264]_ , \new_[7265]_ , \new_[7266]_ , \new_[7267]_ ,
    \new_[7268]_ , \new_[7269]_ , \new_[7270]_ , \new_[7271]_ ,
    \new_[7272]_ , \new_[7273]_ , \new_[7274]_ , \new_[7275]_ ,
    \new_[7276]_ , \new_[7277]_ , \new_[7278]_ , \new_[7279]_ ,
    \new_[7280]_ , \new_[7281]_ , \new_[7282]_ , \new_[7283]_ ,
    \new_[7284]_ , \new_[7285]_ , \new_[7286]_ , \new_[7287]_ ,
    \new_[7288]_ , \new_[7289]_ , \new_[7290]_ , \new_[7291]_ ,
    \new_[7292]_ , \new_[7293]_ , \new_[7294]_ , \new_[7295]_ ,
    \new_[7296]_ , \new_[7297]_ , \new_[7298]_ , \new_[7299]_ ,
    \new_[7300]_ , \new_[7301]_ , \new_[7302]_ , \new_[7303]_ ,
    \new_[7304]_ , \new_[7305]_ , \new_[7306]_ , \new_[7307]_ ,
    \new_[7308]_ , \new_[7309]_ , \new_[7310]_ , \new_[7311]_ ,
    \new_[7312]_ , \new_[7313]_ , \new_[7314]_ , \new_[7315]_ ,
    \new_[7316]_ , \new_[7317]_ , \new_[7318]_ , \new_[7319]_ ,
    \new_[7320]_ , \new_[7321]_ , \new_[7322]_ , \new_[7323]_ ,
    \new_[7324]_ , \new_[7325]_ , \new_[7326]_ , \new_[7327]_ ,
    \new_[7328]_ , \new_[7329]_ , \new_[7330]_ , \new_[7331]_ ,
    \new_[7332]_ , \new_[7333]_ , \new_[7334]_ , \new_[7335]_ ,
    \new_[7336]_ , \new_[7337]_ , \new_[7338]_ , \new_[7339]_ ,
    \new_[7340]_ , \new_[7341]_ , \new_[7342]_ , \new_[7343]_ ,
    \new_[7344]_ , \new_[7345]_ , \new_[7346]_ , \new_[7347]_ ,
    \new_[7348]_ , \new_[7349]_ , \new_[7350]_ , \new_[7351]_ ,
    \new_[7352]_ , \new_[7353]_ , \new_[7354]_ , \new_[7355]_ ,
    \new_[7356]_ , \new_[7357]_ , \new_[7358]_ , \new_[7359]_ ,
    \new_[7360]_ , \new_[7361]_ , \new_[7362]_ , \new_[7363]_ ,
    \new_[7364]_ , \new_[7365]_ , \new_[7366]_ , \new_[7367]_ ,
    \new_[7368]_ , \new_[7369]_ , \new_[7370]_ , \new_[7371]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7374]_ , \new_[7375]_ ,
    \new_[7376]_ , \new_[7377]_ , \new_[7378]_ , \new_[7379]_ ,
    \new_[7381]_ , \new_[7382]_ , \new_[7383]_ , \new_[7384]_ ,
    \new_[7385]_ , \new_[7387]_ , \new_[7388]_ , \new_[7389]_ ,
    \new_[7390]_ , \new_[7391]_ , \new_[7392]_ , \new_[7393]_ ,
    \new_[7394]_ , \new_[7396]_ , \new_[7397]_ , \new_[7398]_ ,
    \new_[7399]_ , \new_[7400]_ , \new_[7401]_ , \new_[7402]_ ,
    \new_[7403]_ , \new_[7404]_ , \new_[7405]_ , \new_[7406]_ ,
    \new_[7407]_ , \new_[7408]_ , \new_[7409]_ , \new_[7410]_ ,
    \new_[7411]_ , \new_[7412]_ , \new_[7413]_ , \new_[7414]_ ,
    \new_[7415]_ , \new_[7416]_ , \new_[7418]_ , \new_[7419]_ ,
    \new_[7420]_ , \new_[7421]_ , \new_[7423]_ , \new_[7424]_ ,
    \new_[7425]_ , \new_[7426]_ , \new_[7427]_ , \new_[7428]_ ,
    \new_[7429]_ , \new_[7430]_ , \new_[7431]_ , \new_[7432]_ ,
    \new_[7433]_ , \new_[7434]_ , \new_[7435]_ , \new_[7436]_ ,
    \new_[7437]_ , \new_[7438]_ , \new_[7439]_ , \new_[7440]_ ,
    \new_[7441]_ , \new_[7442]_ , \new_[7443]_ , \new_[7444]_ ,
    \new_[7445]_ , \new_[7446]_ , \new_[7447]_ , \new_[7448]_ ,
    \new_[7449]_ , \new_[7450]_ , \new_[7451]_ , \new_[7452]_ ,
    \new_[7453]_ , \new_[7454]_ , \new_[7455]_ , \new_[7456]_ ,
    \new_[7457]_ , \new_[7458]_ , \new_[7459]_ , \new_[7460]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7464]_ ,
    \new_[7465]_ , \new_[7466]_ , \new_[7467]_ , \new_[7468]_ ,
    \new_[7469]_ , \new_[7470]_ , \new_[7471]_ , \new_[7472]_ ,
    \new_[7473]_ , \new_[7474]_ , \new_[7475]_ , \new_[7476]_ ,
    \new_[7477]_ , \new_[7478]_ , \new_[7479]_ , \new_[7480]_ ,
    \new_[7481]_ , \new_[7482]_ , \new_[7483]_ , \new_[7484]_ ,
    \new_[7485]_ , \new_[7486]_ , \new_[7487]_ , \new_[7488]_ ,
    \new_[7489]_ , \new_[7490]_ , \new_[7491]_ , \new_[7492]_ ,
    \new_[7493]_ , \new_[7494]_ , \new_[7495]_ , \new_[7496]_ ,
    \new_[7497]_ , \new_[7498]_ , \new_[7499]_ , \new_[7500]_ ,
    \new_[7501]_ , \new_[7502]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7505]_ , \new_[7507]_ , \new_[7508]_ , \new_[7509]_ ,
    \new_[7510]_ , \new_[7511]_ , \new_[7512]_ , \new_[7513]_ ,
    \new_[7514]_ , \new_[7515]_ , \new_[7516]_ , \new_[7517]_ ,
    \new_[7518]_ , \new_[7519]_ , \new_[7520]_ , \new_[7521]_ ,
    \new_[7522]_ , \new_[7523]_ , \new_[7524]_ , \new_[7525]_ ,
    \new_[7526]_ , \new_[7527]_ , \new_[7528]_ , \new_[7529]_ ,
    \new_[7530]_ , \new_[7531]_ , \new_[7532]_ , \new_[7533]_ ,
    \new_[7534]_ , \new_[7535]_ , \new_[7536]_ , \new_[7537]_ ,
    \new_[7538]_ , \new_[7539]_ , \new_[7540]_ , \new_[7541]_ ,
    \new_[7542]_ , \new_[7543]_ , \new_[7544]_ , \new_[7545]_ ,
    \new_[7546]_ , \new_[7547]_ , \new_[7548]_ , \new_[7549]_ ,
    \new_[7550]_ , \new_[7551]_ , \new_[7552]_ , \new_[7553]_ ,
    \new_[7554]_ , \new_[7555]_ , \new_[7556]_ , \new_[7557]_ ,
    \new_[7558]_ , \new_[7559]_ , \new_[7560]_ , \new_[7561]_ ,
    \new_[7562]_ , \new_[7563]_ , \new_[7564]_ , \new_[7565]_ ,
    \new_[7566]_ , \new_[7567]_ , \new_[7568]_ , \new_[7569]_ ,
    \new_[7570]_ , n94, n99, n104, n109, n114, n119, n124, n129, n134,
    n139, n144, n149, n154, n159, n164, n169, n174, n179, n184, n189, n194,
    n199, n204, n209, n214, n219, n224, n229, n234, n239, n244, n249, n254,
    n259, n264, n269, n274, n279, n284, n289, n294, n299, n304, n309, n314,
    n319, n324, n329, n334, n339, n344, n349, n354, n359, n364, n369, n374,
    n379, n384, n389, n394, n399, n404, n409, n414, n419, n424, n429, n434,
    n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489, n494,
    n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549, n554,
    n559, n564, n569, n574, n579, n584, n589, n594, n599, n604, n609, n614,
    n619, n624, n629, n634, n639, n644, n649, n654, n659, n664, n669, n674,
    n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729, n734,
    n739, n744, n749, n754, n759, n764, n769, n774, n779, n784, n789, n794,
    n799, n804, n809, n814, n819, n824, n829, n834, n839, n844, n849, n854,
    n859, n864, n869, n874, n879, n884, n889, n894, n899, n904, n909, n914,
    n919, n924, n929, n934, n939, n944, n949, n954, n959, n964, n969, n974,
    n979, n984, n989, n994, n999, n1004, n1009, n1014, n1019, n1024, n1029,
    n1034, n1039, n1044, n1049, n1054, n1059, n1064, n1069, n1074, n1079,
    n1084, n1089, n1094, n1099, n1104, n1109, n1114, n1119, n1124, n1129,
    n1134, n1139, n1144, n1149, n1154, n1159, n1164, n1169, n1174, n1179,
    n1184, n1189, n1194, n1199, n1204, n1209, n1214, n1219, n1224, n1229,
    n1234, n1239, n1244, n1249, n1254, n1259, n1264, n1269, n1274, n1279,
    n1284, n1289, n1294, n1299, n1304, n1309, n1314, n1319, n1324, n1329,
    n1334, n1339, n1344, n1349, n1354, n1359, n1364, n1369, n1374, n1379,
    n1384, n1389, n1394, n1399, n1404, n1409, n1414, n1419, n1424, n1429,
    n1434, n1439, n1444, n1449, n1454, n1459, n1464, n1469, n1474, n1479,
    n1484, n1489, n1494, n1499, n1504, n1509, n1514, n1519, n1524, n1529,
    n1534, n1539, n1544, n1549, n1554, n1559, n1564, n1569, n1574, n1579,
    n1584, n1589, n1594, n1599, n1604, n1609, n1614, n1619, n1624, n1629,
    n1634, n1639, n1644, n1649, n1654, n1659, n1664, n1669, n1674, n1679,
    n1684, n1689, n1694, n1699, n1704, n1709, n1714, n1719, n1724, n1729,
    n1734, n1739, n1744, n1749, n1754, n1759, n1764, n1769, n1774, n1779,
    n1784, n1789, n1794, n1799, n1804, n1809, n1814, n1819, n1824, n1829,
    n1834, n1839, n1844, n1849, n1854, n1859, n1864, n1869, n1874, n1879,
    n1884;
  assign \new_[407]_  = i_tv80_core_IncDecZ_reg;
  assign \A[1]  = \\i_tv80_core_A_reg[1] ;
  assign \A[2]  = \\i_tv80_core_A_reg[2] ;
  assign \A[5]  = \\i_tv80_core_A_reg[5] ;
  assign \A[6]  = \\i_tv80_core_A_reg[6] ;
  assign \new_[412]_  = ~\\i_tv80_core_i_reg_RegsH_reg[0][6] ;
  assign \new_[413]_  = ~\\i_tv80_core_i_reg_RegsH_reg[1][6] ;
  assign \new_[414]_  = ~\\i_tv80_core_i_reg_RegsH_reg[2][6] ;
  assign \new_[415]_  = ~\\i_tv80_core_i_reg_RegsH_reg[3][6] ;
  assign \new_[416]_  = ~\\i_tv80_core_i_reg_RegsH_reg[4][6] ;
  assign \new_[417]_  = ~\\i_tv80_core_i_reg_RegsH_reg[5][6] ;
  assign \new_[418]_  = ~\\i_tv80_core_i_reg_RegsH_reg[6][6] ;
  assign \new_[419]_  = ~\\i_tv80_core_i_reg_RegsH_reg[7][6] ;
  assign \new_[420]_  = ~\\i_tv80_core_i_reg_RegsH_reg[0][4] ;
  assign \new_[421]_  = ~\\i_tv80_core_i_reg_RegsH_reg[1][4] ;
  assign \new_[422]_  = ~\\i_tv80_core_i_reg_RegsH_reg[2][4] ;
  assign \new_[423]_  = ~\\i_tv80_core_i_reg_RegsH_reg[3][4] ;
  assign \new_[424]_  = ~\\i_tv80_core_i_reg_RegsH_reg[4][4] ;
  assign \new_[425]_  = ~\\i_tv80_core_i_reg_RegsH_reg[5][4] ;
  assign \new_[426]_  = ~\\i_tv80_core_i_reg_RegsH_reg[6][4] ;
  assign \new_[427]_  = ~\\i_tv80_core_i_reg_RegsH_reg[7][4] ;
  assign \new_[428]_  = \\i_tv80_core_i_reg_RegsH_reg[0][2] ;
  assign \new_[429]_  = \\i_tv80_core_i_reg_RegsH_reg[1][2] ;
  assign \new_[430]_  = \\i_tv80_core_i_reg_RegsH_reg[2][2] ;
  assign \new_[431]_  = \\i_tv80_core_i_reg_RegsH_reg[3][2] ;
  assign \new_[432]_  = \\i_tv80_core_i_reg_RegsH_reg[4][2] ;
  assign \new_[433]_  = \\i_tv80_core_i_reg_RegsH_reg[5][2] ;
  assign \new_[434]_  = \\i_tv80_core_i_reg_RegsH_reg[6][2] ;
  assign \new_[435]_  = \\i_tv80_core_i_reg_RegsH_reg[7][2] ;
  assign n94 = ~\new_[7401]_ ;
  assign n119 = ~\new_[1068]_  | (~\new_[497]_  & ~\new_[6903]_ );
  assign n134 = ~\new_[1081]_  | (~\new_[499]_  & ~\new_[1185]_ );
  assign n104 = ~\new_[6623]_  & (~\new_[6033]_  | ~\new_[502]_ );
  assign n139 = ~\new_[1088]_  | (~\new_[500]_  & ~\new_[1189]_ );
  assign n154 = ~\new_[1100]_  | (~\new_[498]_  & ~\new_[1189]_ );
  assign n99 = ~\new_[6623]_  & (~\new_[6063]_  | ~\new_[501]_ );
  assign n109 = ~\new_[6623]_  & (~\new_[6052]_  | ~\new_[503]_ );
  assign \A[11]  = \\i_tv80_core_A_reg[11] ;
  assign \A[12]  = \\i_tv80_core_A_reg[12] ;
  assign \A[13]  = \\i_tv80_core_A_reg[13] ;
  assign \A[14]  = \\i_tv80_core_A_reg[14] ;
  assign \A[10]  = \\i_tv80_core_A_reg[10] ;
  assign \A[4]  = \\i_tv80_core_A_reg[4] ;
  assign \A[0]  = \\i_tv80_core_A_reg[0] ;
  assign \A[3]  = \\i_tv80_core_A_reg[3] ;
  assign \A[15]  = \\i_tv80_core_A_reg[15] ;
  assign \A[8]  = \\i_tv80_core_A_reg[8] ;
  assign \A[7]  = \\i_tv80_core_A_reg[7] ;
  assign \A[9]  = \\i_tv80_core_A_reg[9] ;
  assign n299 = \\i_tv80_core_i_reg_RegsH_reg[0][7] ;
  assign n304 = \\i_tv80_core_i_reg_RegsH_reg[1][7] ;
  assign n309 = \\i_tv80_core_i_reg_RegsH_reg[2][7] ;
  assign n314 = \\i_tv80_core_i_reg_RegsH_reg[3][7] ;
  assign n319 = \\i_tv80_core_i_reg_RegsH_reg[4][7] ;
  assign n324 = \\i_tv80_core_i_reg_RegsH_reg[5][7] ;
  assign n329 = \\i_tv80_core_i_reg_RegsH_reg[6][7] ;
  assign n334 = \\i_tv80_core_i_reg_RegsH_reg[7][7] ;
  assign \new_[464]_  = ~\\i_tv80_core_i_reg_RegsH_reg[0][5] ;
  assign \new_[465]_  = ~\\i_tv80_core_i_reg_RegsH_reg[1][5] ;
  assign \new_[466]_  = ~\\i_tv80_core_i_reg_RegsH_reg[2][5] ;
  assign \new_[467]_  = ~\\i_tv80_core_i_reg_RegsH_reg[3][5] ;
  assign \new_[468]_  = ~\\i_tv80_core_i_reg_RegsH_reg[4][5] ;
  assign \new_[469]_  = ~\\i_tv80_core_i_reg_RegsH_reg[7][5] ;
  assign \new_[470]_  = ~\\i_tv80_core_i_reg_RegsH_reg[5][5] ;
  assign \new_[471]_  = ~\\i_tv80_core_i_reg_RegsH_reg[6][5] ;
  assign n114 = ~\new_[6623]_  & (~\new_[6051]_  | ~\new_[504]_ );
  assign n164 = ~\new_[1071]_  | (~\new_[521]_  & ~\new_[1185]_ );
  assign n174 = ~\new_[1079]_  | (~\new_[522]_  & ~\new_[1190]_ );
  assign n179 = ~\new_[1086]_  | (~\new_[523]_  & ~\new_[1189]_ );
  assign n194 = ~\new_[1098]_  | (~\new_[525]_  & ~\new_[1186]_ );
  assign n199 = ~\new_[1065]_  | (~\new_[550]_  & ~\new_[1191]_ );
  assign n214 = ~\new_[1077]_  | (~\new_[552]_  & ~\new_[1185]_ );
  assign n219 = ~\new_[1084]_  | (~\new_[553]_  & ~\new_[1185]_ );
  assign n234 = ~\new_[1096]_  | (~\new_[555]_  & ~\new_[6903]_ );
  assign n279 = ~\new_[546]_  & ~\new_[6329]_ ;
  assign n264 = ~\new_[548]_  & ~\new_[6402]_ ;
  assign n274 = ~\new_[547]_  & ~\new_[6413]_ ;
  assign n289 = ~\new_[549]_  & ~\new_[6382]_ ;
  assign n339 = ~\new_[1067]_  | (~\new_[561]_  & ~\new_[1191]_ );
  assign n284 = ~\new_[551]_  & ~\new_[6403]_ ;
  assign n294 = ~\new_[554]_  & ~\new_[6370]_ ;
  assign n354 = ~\new_[1080]_  | (~\new_[563]_  & ~\new_[1185]_ );
  assign n359 = ~\new_[1087]_  | (~\new_[564]_  & ~\new_[1189]_ );
  assign n364 = ~\new_[1099]_  | (~\new_[565]_  & ~\new_[1186]_ );
  assign n269 = ~\new_[524]_  & ~\new_[6424]_ ;
  assign n259 = ~\new_[526]_  & ~\new_[6382]_ ;
  assign n239 = ~\new_[527]_  & ~\new_[6426]_ ;
  assign n244 = ~\new_[541]_  & ~\new_[6329]_ ;
  assign n249 = ~\new_[544]_  & ~\new_[6370]_ ;
  assign n254 = ~\new_[545]_  & ~\new_[6424]_ ;
  assign \new_[497]_  = ~\new_[2413]_  | (~\new_[6847]_  & ~\new_[7397]_ );
  assign \new_[498]_  = ~\new_[2507]_  | (~\new_[6847]_  & ~\new_[2625]_ );
  assign \new_[499]_  = ~\new_[2336]_  | (~\new_[6847]_  & ~\new_[2622]_ );
  assign \new_[500]_  = ~\new_[2343]_  | (~\new_[6847]_  & ~\new_[2423]_ );
  assign \new_[501]_  = ~\new_[556]_  | ~busak_n;
  assign \new_[502]_  = ~\new_[557]_  | ~busak_n;
  assign \new_[503]_  = ~\new_[558]_  | ~busak_n;
  assign \new_[504]_  = ~\new_[559]_  | ~busak_n;
  assign \new_[505]_  = ~\\i_tv80_core_i_reg_RegsH_reg[0][3] ;
  assign \new_[506]_  = ~\\i_tv80_core_i_reg_RegsH_reg[1][3] ;
  assign \new_[507]_  = ~\\i_tv80_core_i_reg_RegsH_reg[2][3] ;
  assign \new_[508]_  = ~\\i_tv80_core_i_reg_RegsH_reg[3][3] ;
  assign \new_[509]_  = ~\\i_tv80_core_i_reg_RegsH_reg[4][3] ;
  assign \new_[510]_  = ~\\i_tv80_core_i_reg_RegsH_reg[5][3] ;
  assign \new_[511]_  = ~\\i_tv80_core_i_reg_RegsH_reg[6][3] ;
  assign \new_[512]_  = ~\\i_tv80_core_i_reg_RegsH_reg[7][3] ;
  assign \new_[520]_  = \\i_tv80_core_i_reg_RegsH_reg[5][1] ;
  assign \new_[521]_  = ~\new_[2482]_  | (~\new_[6769]_  & ~\new_[6846]_ );
  assign \new_[522]_  = ~\new_[2334]_  | (~\new_[6769]_  & ~\new_[2622]_ );
  assign \new_[523]_  = ~\new_[2341]_  | (~\new_[6769]_  & ~\new_[2423]_ );
  assign \new_[524]_  = (~\new_[616]_  | ~\new_[6126]_ ) & (~\A[0]  | ~\new_[6239]_ );
  assign \new_[525]_  = ~\new_[2503]_  | (~\new_[6769]_  & ~\new_[2626]_ );
  assign \new_[526]_  = (~\new_[6132]_  | ~\new_[617]_ ) & (~\A[10]  | ~\new_[6149]_ );
  assign \new_[527]_  = (~\new_[618]_  | ~\new_[6126]_ ) & (~\A[11]  | ~\new_[6149]_ );
  assign \new_[528]_  = \\i_tv80_core_i_reg_RegsL_reg[0][6] ;
  assign \new_[529]_  = \\i_tv80_core_i_reg_RegsL_reg[1][6] ;
  assign \new_[530]_  = \\i_tv80_core_i_reg_RegsL_reg[2][6] ;
  assign \new_[531]_  = \\i_tv80_core_i_reg_RegsL_reg[5][6] ;
  assign \new_[532]_  = \\i_tv80_core_i_reg_RegsL_reg[6][6] ;
  assign \new_[533]_  = \\i_tv80_core_i_reg_RegsL_reg[7][6] ;
  assign \new_[534]_  = \\i_tv80_core_i_reg_RegsL_reg[3][6] ;
  assign \new_[535]_  = \\i_tv80_core_i_reg_RegsL_reg[4][6] ;
  assign \new_[536]_  = \\i_tv80_core_i_reg_RegsH_reg[0][1] ;
  assign \new_[537]_  = \\i_tv80_core_i_reg_RegsH_reg[1][1] ;
  assign \new_[538]_  = \\i_tv80_core_i_reg_RegsH_reg[2][1] ;
  assign \new_[539]_  = \\i_tv80_core_i_reg_RegsH_reg[3][1] ;
  assign \new_[540]_  = \\i_tv80_core_i_reg_RegsH_reg[4][1] ;
  assign \new_[541]_  = (~\new_[619]_  | ~\new_[6126]_ ) & (~\A[12]  | ~\new_[6149]_ );
  assign \new_[542]_  = \\i_tv80_core_i_reg_RegsH_reg[6][1] ;
  assign \new_[543]_  = \\i_tv80_core_i_reg_RegsH_reg[7][1] ;
  assign \new_[544]_  = (~\new_[620]_  | ~\new_[6314]_ ) & (~\A[13]  | ~\new_[6165]_ );
  assign \new_[545]_  = (~\new_[621]_  | ~\new_[6314]_ ) & (~\A[14]  | ~\new_[6322]_ );
  assign \new_[546]_  = (~\new_[622]_  | ~\new_[6263]_ ) & (~\A[15]  | ~\new_[6239]_ );
  assign \new_[547]_  = (~\new_[6263]_  | ~\new_[623]_ ) & (~\A[3]  | ~\new_[6322]_ );
  assign \new_[548]_  = (~\new_[624]_  | ~\new_[6263]_ ) & (~\A[4]  | ~\new_[6322]_ );
  assign \new_[549]_  = (~\new_[625]_  | ~\new_[6314]_ ) & (~\A[7]  | ~\new_[6438]_ );
  assign \new_[550]_  = ~\new_[2407]_  | (~\new_[6910]_  & ~\new_[7397]_ );
  assign \new_[551]_  = (~\new_[626]_  | ~\new_[6132]_ ) & (~\A[8]  | ~\new_[6438]_ );
  assign \new_[552]_  = ~\new_[2332]_  | (~\new_[6910]_  & ~\new_[2422]_ );
  assign \new_[553]_  = ~\new_[2339]_  | (~\new_[6910]_  & ~\new_[2623]_ );
  assign \new_[554]_  = (~\new_[627]_  | ~\new_[6132]_ ) & (~\A[9]  | ~\new_[6149]_ );
  assign \new_[555]_  = ~\new_[2501]_  | (~\new_[6910]_  & ~\new_[2625]_ );
  assign \new_[556]_  = ~\new_[3137]_  | (~\new_[634]_  & ~\new_[6712]_ );
  assign \new_[557]_  = ~\new_[3138]_  | (~\new_[635]_  & ~\new_[3234]_ );
  assign \new_[558]_  = ~\new_[3136]_  | (~\new_[636]_  & ~\new_[6712]_ );
  assign \new_[559]_  = ~\new_[3140]_  | (~\new_[637]_  & ~\new_[6712]_ );
  assign \new_[560]_  = \\i_tv80_core_i_reg_RegsH_reg[4][0] ;
  assign \new_[561]_  = ~\new_[2406]_  | (~\new_[7392]_  & ~\new_[2529]_ );
  assign \new_[562]_  = \\i_tv80_core_i_reg_RegsL_reg[7][7] ;
  assign \new_[563]_  = ~\new_[2335]_  | (~\new_[7431]_  & ~\new_[2622]_ );
  assign \new_[564]_  = ~\new_[2342]_  | (~\new_[7392]_  & ~\new_[2423]_ );
  assign \new_[565]_  = ~\new_[2506]_  | (~\new_[7392]_  & ~\new_[2626]_ );
  assign n379 = ~\new_[1066]_  | (~\new_[638]_  & ~\new_[6903]_ );
  assign \new_[567]_  = \\i_tv80_core_i_reg_RegsL_reg[0][7] ;
  assign \new_[568]_  = \\i_tv80_core_i_reg_RegsL_reg[1][7] ;
  assign \new_[569]_  = \\i_tv80_core_i_reg_RegsL_reg[2][7] ;
  assign \new_[570]_  = \\i_tv80_core_i_reg_RegsL_reg[3][7] ;
  assign \new_[571]_  = \\i_tv80_core_i_reg_RegsL_reg[4][7] ;
  assign \new_[572]_  = \\i_tv80_core_i_reg_RegsL_reg[5][7] ;
  assign \new_[573]_  = \\i_tv80_core_i_reg_RegsL_reg[6][7] ;
  assign \new_[574]_  = \\i_tv80_core_i_reg_RegsH_reg[0][0] ;
  assign \new_[575]_  = \\i_tv80_core_i_reg_RegsH_reg[1][0] ;
  assign \new_[576]_  = \\i_tv80_core_i_reg_RegsH_reg[2][0] ;
  assign \new_[577]_  = \\i_tv80_core_i_reg_RegsH_reg[3][0] ;
  assign \new_[578]_  = \\i_tv80_core_i_reg_RegsH_reg[5][0] ;
  assign \new_[579]_  = \\i_tv80_core_i_reg_RegsH_reg[6][0] ;
  assign \new_[580]_  = \\i_tv80_core_i_reg_RegsH_reg[7][0] ;
  assign n384 = ~\new_[1070]_  | (~\new_[639]_  & ~\new_[6856]_ );
  assign n389 = ~\new_[1074]_  | (~\new_[640]_  & ~\new_[1190]_ );
  assign n394 = ~\new_[1078]_  | (~\new_[641]_  & ~\new_[1190]_ );
  assign n399 = ~\new_[1085]_  | (~\new_[642]_  & ~\new_[1190]_ );
  assign n404 = ~\new_[1091]_  | (~\new_[643]_  & ~\new_[7430]_ );
  assign n409 = ~\new_[1093]_  | (~\new_[644]_  & ~\new_[7430]_ );
  assign n414 = ~\new_[1097]_  | (~\new_[645]_  & ~\new_[6856]_ );
  assign n424 = ~\new_[966]_  | ~\new_[666]_ ;
  assign n429 = ~\new_[973]_  | ~\new_[667]_ ;
  assign n434 = ~\new_[979]_  | ~\new_[668]_ ;
  assign n454 = ~\new_[984]_  | ~\new_[669]_ ;
  assign n459 = ~\new_[989]_  | ~\new_[670]_ ;
  assign n439 = ~\new_[996]_  | ~\new_[631]_ ;
  assign n444 = ~\new_[1000]_  | ~\new_[632]_ ;
  assign \new_[595]_  = \\i_tv80_core_tstate_reg[0] ;
  assign \new_[596]_  = \\i_tv80_core_tstate_reg[1] ;
  assign \new_[597]_  = \\i_tv80_core_tstate_reg[2] ;
  assign n449 = ~\new_[961]_  | ~\new_[633]_ ;
  assign n474 = ~\new_[1073]_  | (~\new_[671]_  & ~\new_[1190]_ );
  assign n479 = ~\new_[1076]_  | (~\new_[672]_  & ~\new_[1190]_ );
  assign n484 = ~\new_[1083]_  | (~\new_[673]_  & ~\new_[1190]_ );
  assign n419 = ~\new_[1090]_  | (~\new_[674]_  & ~\new_[1190]_ );
  assign n494 = ~\new_[1095]_  | (~\new_[675]_  & ~\new_[1185]_ );
  assign n564 = ~\new_[1089]_  | (~\new_[700]_  & ~\new_[1186]_ );
  assign n499 = ~\new_[1082]_  | (~\new_[698]_  & ~\new_[6856]_ );
  assign n569 = ~\new_[1092]_  | (~\new_[701]_  & ~\new_[1186]_ );
  assign n574 = ~\new_[1094]_  | (~\new_[702]_  & ~\new_[1191]_ );
  assign n509 = ~\new_[967]_  | ~\new_[676]_ ;
  assign n514 = ~\new_[974]_  | ~\new_[677]_ ;
  assign n519 = ~\new_[980]_  | ~\new_[678]_ ;
  assign n524 = ~\new_[985]_  | ~\new_[682]_ ;
  assign n529 = ~\new_[990]_  | ~\new_[679]_ ;
  assign n534 = ~\new_[997]_  | ~\new_[680]_ ;
  assign n504 = ~\new_[1005]_  | ~\new_[681]_ ;
  assign n539 = ~\new_[1001]_  | ~\new_[683]_ ;
  assign \new_[616]_  = ~\new_[3124]_  | (~\new_[709]_  & ~\new_[3360]_ );
  assign \new_[617]_  = ~\new_[3133]_  | (~\new_[710]_  & ~\new_[6712]_ );
  assign \new_[618]_  = ~\new_[3134]_  | (~\new_[715]_  & ~\new_[3288]_ );
  assign \new_[619]_  = ~\new_[3135]_  | (~\new_[716]_  & ~\new_[3360]_ );
  assign \new_[620]_  = ~\new_[3128]_  | (~\new_[717]_  & ~\new_[3234]_ );
  assign \new_[621]_  = ~\new_[3131]_  | (~\new_[719]_  & ~\new_[3287]_ );
  assign \new_[622]_  = ~\new_[3127]_  | (~\new_[720]_  & ~\new_[6712]_ );
  assign \new_[623]_  = ~\new_[3139]_  | (~\new_[721]_  & ~\new_[6712]_ );
  assign \new_[624]_  = ~\new_[3132]_  | (~\new_[722]_  & ~\new_[3360]_ );
  assign \new_[625]_  = ~\new_[3130]_  | (~\new_[723]_  & ~\new_[3288]_ );
  assign \new_[626]_  = ~\new_[3129]_  | (~\new_[724]_  & ~\new_[3287]_ );
  assign \new_[627]_  = ~\new_[3141]_  | (~\new_[725]_  & ~\new_[3234]_ );
  assign n549 = ~\new_[1069]_  | (~\new_[695]_  & ~\new_[1191]_ );
  assign n554 = ~\new_[1072]_  | (~\new_[696]_  & ~\new_[6903]_ );
  assign n559 = ~\new_[1075]_  | (~\new_[697]_  & ~\new_[6856]_ );
  assign \new_[631]_  = ~\new_[748]_  | ~\new_[1105]_  | ~\new_[2511]_ ;
  assign \new_[632]_  = ~\new_[749]_  | ~\new_[1105]_  | ~\new_[2514]_ ;
  assign \new_[633]_  = ~\new_[750]_  | ~\new_[1105]_  | ~\new_[2519]_ ;
  assign \new_[634]_  = ~\new_[699]_  & (~\new_[2127]_  | ~\A[1] );
  assign \new_[635]_  = ~\new_[703]_  & (~\new_[2127]_  | ~\A[2] );
  assign \new_[636]_  = ~\new_[704]_  & (~\new_[2127]_  | ~\A[5] );
  assign \new_[637]_  = ~\new_[705]_  & (~\new_[2127]_  | ~\A[6] );
  assign \new_[638]_  = ~\new_[2408]_  | (~\new_[741]_  & ~\new_[7397]_ );
  assign \new_[639]_  = ~\new_[2488]_  | (~\new_[741]_  & ~\new_[6846]_ );
  assign \new_[640]_  = ~\new_[2615]_  | (~\new_[741]_  & ~\new_[2711]_ );
  assign \new_[641]_  = ~\new_[2333]_  | (~\new_[741]_  & ~\new_[2422]_ );
  assign \new_[642]_  = ~\new_[2340]_  | (~\new_[741]_  & ~\new_[2623]_ );
  assign \new_[643]_  = ~\new_[2496]_  | (~\new_[741]_  & ~\new_[6907]_ );
  assign \new_[644]_  = ~\new_[2419]_  | (~\new_[741]_  & ~\new_[6853]_ );
  assign \new_[645]_  = ~\new_[2502]_  | (~\new_[741]_  & ~\new_[2625]_ );
  assign \new_[646]_  = \\i_tv80_core_i_reg_RegsL_reg[4][4] ;
  assign n584 = ~\new_[6441]_  & (~\new_[5400]_  | ~\new_[795]_ );
  assign n579 = ~\new_[727]_  & ~\new_[6371]_ ;
  assign n589 = ~\new_[728]_  & ~\new_[6441]_ ;
  assign \new_[650]_  = \\i_tv80_core_i_reg_RegsL_reg[0][5] ;
  assign \new_[651]_  = \\i_tv80_core_F_reg[2] ;
  assign \new_[652]_  = \\i_tv80_core_i_reg_RegsL_reg[1][5] ;
  assign \new_[653]_  = \\i_tv80_core_i_reg_RegsL_reg[2][5] ;
  assign \new_[654]_  = \\i_tv80_core_i_reg_RegsL_reg[3][5] ;
  assign \new_[655]_  = \\i_tv80_core_i_reg_RegsL_reg[4][5] ;
  assign \new_[656]_  = \\i_tv80_core_i_reg_RegsL_reg[5][5] ;
  assign \new_[657]_  = \\i_tv80_core_i_reg_RegsL_reg[6][5] ;
  assign \new_[658]_  = \\i_tv80_core_i_reg_RegsL_reg[7][5] ;
  assign \new_[659]_  = \\i_tv80_core_i_reg_RegsL_reg[0][4] ;
  assign \new_[660]_  = \\i_tv80_core_i_reg_RegsL_reg[1][4] ;
  assign \new_[661]_  = \\i_tv80_core_i_reg_RegsL_reg[2][4] ;
  assign \new_[662]_  = \\i_tv80_core_i_reg_RegsL_reg[3][4] ;
  assign \new_[663]_  = \\i_tv80_core_i_reg_RegsL_reg[6][4] ;
  assign \new_[664]_  = \\i_tv80_core_i_reg_RegsL_reg[7][4] ;
  assign \new_[665]_  = \\i_tv80_core_i_reg_RegsL_reg[5][4] ;
  assign \new_[666]_  = ~\new_[743]_  | ~\new_[1105]_  | ~\new_[2415]_ ;
  assign \new_[667]_  = ~\new_[744]_  | ~\new_[1105]_  | ~\new_[2486]_ ;
  assign \new_[668]_  = ~\new_[745]_  | ~\new_[1105]_  | ~\new_[2618]_ ;
  assign \new_[669]_  = ~\new_[746]_  | ~\new_[1105]_  | ~\new_[2347]_ ;
  assign \new_[670]_  = ~\new_[747]_  | ~\new_[1105]_  | ~\new_[2350]_ ;
  assign \new_[671]_  = ~\new_[2613]_  | (~\new_[7474]_  & ~\new_[6830]_ );
  assign \new_[672]_  = ~\new_[2331]_  | (~\new_[7474]_  & ~\new_[2622]_ );
  assign \new_[673]_  = ~\new_[2338]_  | (~\new_[7474]_  & ~\new_[2423]_ );
  assign \new_[674]_  = ~\new_[2495]_  | (~\new_[7474]_  & ~\new_[7432]_ );
  assign \new_[675]_  = ~\new_[2498]_  | (~\new_[7474]_  & ~\new_[2625]_ );
  assign \new_[676]_  = ~\new_[808]_  | ~\new_[1105]_  | ~\new_[2416]_ ;
  assign \new_[677]_  = ~\new_[818]_  | ~\new_[1105]_  | ~\new_[2487]_ ;
  assign \new_[678]_  = ~\new_[817]_  | ~\new_[1180]_  | ~\new_[2619]_ ;
  assign \new_[679]_  = ~\new_[820]_  | ~\new_[1105]_  | ~\new_[2351]_ ;
  assign \new_[680]_  = ~\new_[819]_  | ~\new_[1180]_  | ~\new_[2512]_ ;
  assign \new_[681]_  = ~\new_[7497]_  | ~\new_[1105]_  | ~\new_[2520]_ ;
  assign \new_[682]_  = ~\new_[822]_  | ~\new_[1105]_  | ~\new_[2348]_ ;
  assign \new_[683]_  = ~\new_[821]_  | ~\new_[1180]_  | ~\new_[2516]_ ;
  assign \new_[684]_  = \\i_tv80_core_SP_reg[14] ;
  assign \new_[685]_  = \\i_tv80_core_i_reg_RegsL_reg[5][3] ;
  assign \new_[686]_  = \\i_tv80_core_i_reg_RegsL_reg[6][3] ;
  assign n599 = ~\new_[965]_  | ~\new_[800]_ ;
  assign n609 = ~\new_[971]_  | ~\new_[801]_ ;
  assign n614 = ~\new_[978]_  | ~\new_[802]_ ;
  assign n619 = ~\new_[983]_  | ~\new_[803]_ ;
  assign n624 = ~\new_[1006]_  | ~\new_[804]_ ;
  assign n629 = ~\new_[995]_  | ~\new_[805]_ ;
  assign n634 = ~\new_[1007]_  | ~\new_[806]_ ;
  assign n639 = ~\new_[1004]_  | ~\new_[807]_ ;
  assign \new_[695]_  = ~\new_[2409]_  | (~\new_[6868]_  & ~\new_[7382]_ );
  assign \new_[696]_  = ~\new_[2612]_  | (~\new_[6868]_  & ~\new_[6830]_ );
  assign \new_[697]_  = ~\new_[2241]_  | (~\new_[6868]_  & ~\new_[2422]_ );
  assign \new_[698]_  = ~\new_[2242]_  | (~\new_[6868]_  & ~\new_[2623]_ );
  assign \new_[699]_  = ~\new_[2128]_  & (~\new_[898]_  | ~\new_[3862]_ );
  assign \new_[700]_  = ~\new_[2494]_  | (~\new_[6868]_  & ~\new_[6907]_ );
  assign \new_[701]_  = ~\new_[2418]_  | (~\new_[6868]_  & ~\new_[7419]_ );
  assign \new_[702]_  = ~\new_[2497]_  | (~\new_[6868]_  & ~\new_[2626]_ );
  assign \new_[703]_  = ~\new_[2128]_  & (~\new_[899]_  | ~\new_[3863]_ );
  assign \new_[704]_  = ~\new_[2128]_  & (~\new_[902]_  | ~\new_[3855]_ );
  assign \new_[705]_  = ~\new_[2128]_  & (~\new_[904]_  | ~\new_[3856]_ );
  assign n644 = ~\new_[964]_  | ~\new_[809]_ ;
  assign n649 = ~\new_[970]_  | ~\new_[810]_ ;
  assign n654 = ~\new_[977]_  | ~\new_[811]_ ;
  assign \new_[709]_  = ~\new_[832]_  & (~\new_[2127]_  | ~\A[0] );
  assign \new_[710]_  = ~\new_[833]_  & (~\new_[2127]_  | ~\A[10] );
  assign n659 = ~\new_[982]_  | ~\new_[812]_ ;
  assign n594 = ~\new_[988]_  | ~\new_[813]_ ;
  assign n674 = ~\new_[994]_  | ~\new_[814]_ ;
  assign n664 = ~\new_[999]_  | ~\new_[815]_ ;
  assign \new_[715]_  = ~\new_[834]_  & (~\new_[2129]_  | ~\A[11] );
  assign \new_[716]_  = ~\new_[835]_  & (~\new_[2127]_  | ~\A[12] );
  assign \new_[717]_  = ~\new_[836]_  & (~\new_[2127]_  | ~\A[13] );
  assign n669 = ~\new_[1003]_  | ~\new_[816]_ ;
  assign \new_[719]_  = ~\new_[837]_  & (~\new_[2129]_  | ~\A[14] );
  assign \new_[720]_  = ~\new_[838]_  & (~\new_[2129]_  | ~\A[15] );
  assign \new_[721]_  = ~\new_[839]_  & (~\new_[2127]_  | ~\A[3] );
  assign \new_[722]_  = ~\new_[840]_  & (~\new_[2127]_  | ~\A[4] );
  assign \new_[723]_  = ~\new_[841]_  & (~\new_[2127]_  | ~\A[7] );
  assign \new_[724]_  = ~\new_[842]_  & (~\new_[2127]_  | ~\A[8] );
  assign \new_[725]_  = ~\new_[843]_  & (~\new_[2127]_  | ~\A[9] );
  assign n604 = ~\new_[798]_  | ~\new_[6376]_ ;
  assign \new_[727]_  = (~\new_[915]_  | ~\new_[5847]_ ) & (~\new_[5614]_  | ~\new_[595]_ );
  assign \new_[728]_  = (~\new_[914]_  | ~\new_[6055]_ ) & (~\new_[5614]_  | ~\new_[597]_ );
  assign \new_[729]_  = ~\new_[1059]_  & ~\new_[854]_ ;
  assign \new_[730]_  = \\i_tv80_core_i_reg_RegsL_reg[0][3] ;
  assign \new_[731]_  = \\i_tv80_core_i_reg_RegsL_reg[1][3] ;
  assign \new_[732]_  = \\i_tv80_core_i_reg_RegsL_reg[3][3] ;
  assign \new_[733]_  = \\i_tv80_core_i_reg_RegsL_reg[4][3] ;
  assign \new_[734]_  = \\i_tv80_core_i_reg_RegsL_reg[7][3] ;
  assign \new_[735]_  = \\i_tv80_core_i_reg_RegsL_reg[2][3] ;
  assign \new_[736]_  = \\i_tv80_core_ACC_reg[0] ;
  assign \new_[737]_  = \\i_tv80_core_i_reg_RegsL_reg[4][1] ;
  assign \do[5]  = \\i_tv80_core_do_reg[5] ;
  assign n679 = ~\new_[896]_  | ~\new_[6304]_ ;
  assign \new_[740]_  = \\i_tv80_core_F_reg[1] ;
  assign \new_[741]_  = \new_[823]_ ;
  assign \new_[742]_  = \\i_tv80_core_SP_reg[1] ;
  assign \new_[743]_  = ~\new_[916]_  | ~\new_[7398]_ ;
  assign \new_[744]_  = ~\new_[916]_  | ~\new_[7383]_ ;
  assign \new_[745]_  = ~\new_[916]_  | ~\new_[7389]_ ;
  assign \new_[746]_  = ~\new_[916]_  | ~\new_[2524]_ ;
  assign \new_[747]_  = ~\new_[916]_  | ~\new_[2526]_ ;
  assign \new_[748]_  = ~\new_[916]_  | ~\new_[7426]_ ;
  assign \new_[749]_  = ~\new_[916]_  | ~\new_[7514]_ ;
  assign \new_[750]_  = ~\new_[916]_  | ~\new_[7498]_ ;
  assign \new_[751]_  = \\i_tv80_core_F_reg[6] ;
  assign \new_[752]_  = \\i_tv80_core_F_reg[0] ;
  assign \new_[753]_  = \\i_tv80_core_ACC_reg[7] ;
  assign \do[7]  = \\i_tv80_core_do_reg[7] ;
  assign \new_[755]_  = \\i_tv80_core_SP_reg[7] ;
  assign \do[6]  = \\i_tv80_core_do_reg[6] ;
  assign \new_[757]_  = \\i_tv80_core_SP_reg[6] ;
  assign \new_[758]_  = \\i_tv80_core_ACC_reg[3] ;
  assign \new_[759]_  = \\i_tv80_core_ACC_reg[5] ;
  assign \new_[760]_  = \\i_tv80_core_ACC_reg[6] ;
  assign \new_[761]_  = \\i_tv80_core_ACC_reg[2] ;
  assign \new_[762]_  = \\i_tv80_core_ACC_reg[1] ;
  assign \new_[763]_  = \\i_tv80_core_ACC_reg[4] ;
  assign \new_[764]_  = \\i_tv80_core_SP_reg[5] ;
  assign \do[4]  = \\i_tv80_core_do_reg[4] ;
  assign \new_[766]_  = \\i_tv80_core_SP_reg[4] ;
  assign \new_[767]_  = \\i_tv80_core_i_reg_RegsL_reg[0][2] ;
  assign \new_[768]_  = \\i_tv80_core_i_reg_RegsL_reg[1][2] ;
  assign \new_[769]_  = \\i_tv80_core_i_reg_RegsL_reg[2][2] ;
  assign \new_[770]_  = \\i_tv80_core_i_reg_RegsL_reg[3][2] ;
  assign \new_[771]_  = \\i_tv80_core_i_reg_RegsL_reg[5][2] ;
  assign \new_[772]_  = \\i_tv80_core_i_reg_RegsL_reg[6][2] ;
  assign \new_[773]_  = \\i_tv80_core_i_reg_RegsL_reg[7][2] ;
  assign \new_[774]_  = \\i_tv80_core_i_reg_RegsL_reg[0][1] ;
  assign \new_[775]_  = \\i_tv80_core_i_reg_RegsL_reg[1][1] ;
  assign \new_[776]_  = \\i_tv80_core_i_reg_RegsL_reg[2][1] ;
  assign \new_[777]_  = \\i_tv80_core_i_reg_RegsL_reg[3][1] ;
  assign \new_[778]_  = \\i_tv80_core_i_reg_RegsL_reg[5][1] ;
  assign \new_[779]_  = \\i_tv80_core_i_reg_RegsL_reg[6][1] ;
  assign \new_[780]_  = \\i_tv80_core_i_reg_RegsL_reg[7][1] ;
  assign \do[0]  = \\i_tv80_core_do_reg[0] ;
  assign \do[1]  = \\i_tv80_core_do_reg[1] ;
  assign \do[2]  = \\i_tv80_core_do_reg[2] ;
  assign \do[3]  = \\i_tv80_core_do_reg[3] ;
  assign \new_[785]_  = \\i_tv80_core_i_reg_RegsL_reg[0][0] ;
  assign \new_[786]_  = \\i_tv80_core_i_reg_RegsL_reg[1][0] ;
  assign \new_[787]_  = \\i_tv80_core_i_reg_RegsL_reg[2][0] ;
  assign \new_[788]_  = \\i_tv80_core_i_reg_RegsL_reg[3][0] ;
  assign \new_[789]_  = \\i_tv80_core_i_reg_RegsL_reg[4][0] ;
  assign \new_[790]_  = \\i_tv80_core_i_reg_RegsL_reg[5][0] ;
  assign \new_[791]_  = \\i_tv80_core_i_reg_RegsL_reg[7][0] ;
  assign \new_[792]_  = \\i_tv80_core_SP_reg[2] ;
  assign \new_[793]_  = \\i_tv80_core_SP_reg[3] ;
  assign \new_[794]_  = \\i_tv80_core_SP_reg[0] ;
  assign \new_[795]_  = ~\new_[5847]_  | ~\new_[6055]_  | ~\new_[921]_ ;
  assign \new_[796]_  = \\i_tv80_core_i_reg_RegsL_reg[4][2] ;
  assign \new_[797]_  = \\i_tv80_core_i_reg_RegsL_reg[6][0] ;
  assign \new_[798]_  = (~\new_[1055]_  | ~\new_[6326]_ ) & (~\new_[6521]_  | ~\new_[6226]_ );
  assign \new_[799]_  = \\i_tv80_core_SP_reg[12] ;
  assign \new_[800]_  = ~\new_[1180]_  | ~\new_[1017]_  | ~\new_[2414]_ ;
  assign \new_[801]_  = ~\new_[1018]_  | ~\new_[1105]_  | ~\new_[2485]_ ;
  assign \new_[802]_  = ~\new_[1180]_  | ~\new_[1019]_  | ~\new_[2614]_ ;
  assign \new_[803]_  = ~\new_[1020]_  | ~\new_[1105]_  | ~\new_[2337]_ ;
  assign \new_[804]_  = ~\new_[1021]_  | ~\new_[1105]_  | ~\new_[2353]_ ;
  assign \new_[805]_  = ~\new_[1022]_  | ~\new_[1180]_  | ~\new_[2499]_ ;
  assign \new_[806]_  = ~\new_[1180]_  | ~\new_[1023]_  | ~\new_[2489]_ ;
  assign \new_[807]_  = ~\new_[1024]_  | ~\new_[1105]_  | ~\new_[2505]_ ;
  assign \new_[808]_  = ~\new_[7499]_  | ~\new_[2530]_ ;
  assign \new_[809]_  = ~\new_[1033]_  | ~\new_[1105]_  | ~\new_[2412]_ ;
  assign \new_[810]_  = ~\new_[1034]_  | ~\new_[1105]_  | ~\new_[2484]_ ;
  assign \new_[811]_  = ~\new_[1035]_  | ~\new_[1180]_  | ~\new_[2616]_ ;
  assign \new_[812]_  = ~\new_[1040]_  | ~\new_[1105]_  | ~\new_[2354]_ ;
  assign \new_[813]_  = ~\new_[1042]_  | ~\new_[1105]_  | ~\new_[2352]_ ;
  assign \new_[814]_  = ~\new_[1044]_  | ~\new_[1105]_  | ~\new_[2515]_ ;
  assign \new_[815]_  = ~\new_[1046]_  | ~\new_[1105]_  | ~\new_[2521]_ ;
  assign \new_[816]_  = ~\new_[1048]_  | ~\new_[1105]_  | ~\new_[2490]_ ;
  assign \new_[817]_  = ~\new_[7499]_  | ~\new_[2710]_ ;
  assign \new_[818]_  = ~\new_[7499]_  | ~\new_[7383]_ ;
  assign \new_[819]_  = ~\new_[7499]_  | ~\new_[7426]_ ;
  assign \new_[820]_  = ~\new_[7499]_  | ~\new_[2526]_ ;
  assign \new_[821]_  = ~\new_[7499]_  | ~\new_[2624]_ ;
  assign \new_[822]_  = ~\new_[7499]_  | ~\new_[2524]_ ;
  assign \new_[823]_  = ~\new_[3771]_  | (~\new_[1049]_  & ~\new_[7466]_ );
  assign n694 = ~\new_[963]_  | ~\new_[925]_ ;
  assign n699 = ~\new_[969]_  | ~\new_[926]_ ;
  assign n719 = ~\new_[975]_  | ~\new_[927]_ ;
  assign n704 = ~\new_[981]_  | ~\new_[928]_ ;
  assign n709 = ~\new_[987]_  | ~\new_[929]_ ;
  assign n684 = ~\new_[993]_  | ~\new_[930]_ ;
  assign n689 = ~\new_[998]_  | ~\new_[931]_ ;
  assign n714 = ~\new_[1002]_  | ~\new_[932]_ ;
  assign \new_[832]_  = ~\new_[2127]_  & (~\new_[940]_  | ~\new_[3857]_ );
  assign \new_[833]_  = ~\new_[2127]_  & (~\new_[941]_  | ~\new_[3858]_ );
  assign \new_[834]_  = ~\new_[2127]_  & (~\new_[942]_  | ~\new_[3763]_ );
  assign \new_[835]_  = ~\new_[2127]_  & (~\new_[943]_  | ~\new_[3859]_ );
  assign \new_[836]_  = ~\new_[2127]_  & (~\new_[944]_  | ~\new_[3764]_ );
  assign \new_[837]_  = ~\new_[2127]_  & (~\new_[945]_  | ~\new_[3860]_ );
  assign \new_[838]_  = ~\new_[2127]_  & (~\new_[946]_  | ~\new_[3861]_ );
  assign \new_[839]_  = ~\new_[2127]_  & (~\new_[947]_  | ~\new_[3864]_ );
  assign \new_[840]_  = ~\new_[2127]_  & (~\new_[948]_  | ~\new_[3865]_ );
  assign \new_[841]_  = ~\new_[2127]_  & (~\new_[949]_  | ~\new_[3765]_ );
  assign \new_[842]_  = ~\new_[2127]_  & (~\new_[950]_  | ~\new_[3866]_ );
  assign \new_[843]_  = ~\new_[2127]_  & (~\new_[951]_  | ~\new_[3766]_ );
  assign \new_[844]_  = \\i_tv80_core_F_reg[7] ;
  assign \new_[845]_  = \\i_tv80_core_SP_reg[15] ;
  assign \new_[846]_  = ~\\i_tv80_core_F_reg[3] ;
  assign \new_[847]_  = ~\\i_tv80_core_F_reg[5] ;
  assign \new_[848]_  = \\i_tv80_core_SP_reg[10] ;
  assign \new_[849]_  = \\i_tv80_core_SP_reg[13] ;
  assign \new_[850]_  = \\i_tv80_core_F_reg[4] ;
  assign \new_[851]_  = \\i_tv80_core_SP_reg[9] ;
  assign \new_[852]_  = \\i_tv80_core_SP_reg[11] ;
  assign \new_[853]_  = \\i_tv80_core_SP_reg[8] ;
  assign \new_[854]_  = ~\new_[917]_  | ~\new_[1220]_ ;
  assign n764 = ~\new_[1014]_  & ~\new_[6413]_ ;
  assign n769 = ~\new_[1013]_  | ~\new_[6393]_ ;
  assign n739 = ~\new_[1008]_  | ~\new_[6304]_ ;
  assign n754 = ~\new_[1015]_  | ~\new_[6393]_ ;
  assign n759 = ~\new_[1016]_  | ~\new_[6376]_ ;
  assign n919 = \new_[785]_  ? \new_[1180]_  : \new_[1361]_ ;
  assign n924 = \new_[786]_  ? \new_[1180]_  : \new_[1363]_ ;
  assign n929 = \new_[787]_  ? \new_[1180]_  : \new_[1364]_ ;
  assign n934 = \new_[788]_  ? \new_[1180]_  : \new_[1365]_ ;
  assign n939 = \new_[789]_  ? \new_[1180]_  : \new_[1366]_ ;
  assign n944 = \new_[790]_  ? \new_[1180]_  : \new_[1367]_ ;
  assign n974 = \new_[797]_  ? \new_[1180]_  : \new_[1368]_ ;
  assign n949 = \new_[791]_  ? \new_[1180]_  : \new_[1362]_ ;
  assign n774 = ~\new_[1026]_  & ~\new_[6424]_ ;
  assign n779 = ~\new_[1025]_  | ~\new_[6393]_ ;
  assign n784 = ~\new_[1029]_  | ~\new_[6376]_ ;
  assign n789 = ~\new_[1030]_  | ~\new_[6376]_ ;
  assign n959 = ~\new_[1009]_  | ~\new_[6393]_ ;
  assign n794 = ~\new_[1031]_  | ~\new_[6295]_ ;
  assign n964 = ~\new_[1010]_  | ~\new_[6393]_ ;
  assign n744 = ~\new_[1011]_  | ~\new_[6393]_ ;
  assign n954 = ~\new_[1012]_  | ~\new_[6393]_ ;
  assign n734 = ~\new_[1028]_  & ~\new_[6370]_ ;
  assign n814 = ~\new_[1027]_  | ~\new_[6304]_ ;
  assign n799 = ~\new_[1054]_  | ~\new_[6295]_ ;
  assign n809 = ~\new_[1056]_  | ~\new_[6295]_ ;
  assign n724 = ~\new_[1058]_  | ~\new_[6295]_ ;
  assign n804 = ~\new_[1057]_  | ~\new_[6295]_ ;
  assign n819 = ~\new_[1051]_  & ~\new_[6623]_ ;
  assign n824 = ~\new_[1050]_  | ~\new_[6376]_ ;
  assign \new_[886]_  = ~\new_[7279]_  & ~\new_[7469]_ ;
  assign \new_[887]_  = ~\new_[6739]_ ;
  assign n829 = ~\new_[962]_  | ~\new_[1036]_ ;
  assign n834 = ~\new_[968]_  | ~\new_[1037]_ ;
  assign n839 = ~\new_[976]_  | ~\new_[1038]_ ;
  assign n844 = ~\new_[959]_  | ~\new_[1039]_ ;
  assign n969 = ~\new_[986]_  | ~\new_[1041]_ ;
  assign n849 = ~\new_[992]_  | ~\new_[1043]_ ;
  assign n854 = ~\new_[960]_  | ~\new_[1045]_ ;
  assign n859 = ~\new_[972]_  | ~\new_[1047]_ ;
  assign \new_[896]_  = (~\new_[1064]_  | ~\new_[6326]_ ) & (~\new_[684]_  | ~\new_[6190]_ );
  assign n749 = ~\new_[991]_  | ~\new_[6393]_ ;
  assign \new_[898]_  = ~\new_[4007]_  | (~\new_[6805]_  & ~\new_[5495]_ );
  assign \new_[899]_  = ~\new_[4007]_  | (~\new_[6783]_  & ~\new_[5497]_ );
  assign n864 = \new_[774]_  ? \new_[1180]_  : \new_[1259]_ ;
  assign n869 = \new_[775]_  ? \new_[1180]_  : \new_[1260]_ ;
  assign \new_[902]_  = ~\new_[4007]_  | (~\new_[6788]_  & ~\new_[5496]_ );
  assign n874 = \new_[776]_  ? \new_[1105]_  : \new_[1261]_ ;
  assign \new_[904]_  = ~\new_[4007]_  | (~\new_[6794]_  & ~\new_[5493]_ );
  assign n879 = \new_[777]_  ? \new_[1105]_  : \new_[1262]_ ;
  assign n729 = \new_[737]_  ? \new_[1105]_  : \new_[1263]_ ;
  assign n884 = \new_[778]_  ? \new_[1105]_  : \new_[1264]_ ;
  assign n889 = \new_[779]_  ? \new_[1180]_  : \new_[1265]_ ;
  assign n894 = \new_[780]_  ? \new_[1180]_  : \new_[1266]_ ;
  assign n899 = ~\new_[953]_  & ~\new_[6623]_ ;
  assign n904 = ~\new_[954]_  & ~\new_[6413]_ ;
  assign n909 = ~\new_[955]_  & ~\new_[6623]_ ;
  assign n914 = ~\new_[956]_  & ~\new_[6623]_ ;
  assign \new_[914]_  = ~\new_[957]_  & ~\new_[5672]_ ;
  assign \new_[915]_  = \new_[958]_  & \new_[6055]_ ;
  assign \new_[916]_  = ~\new_[939]_ ;
  assign \new_[917]_  = ~\new_[6754]_ ;
  assign n994 = ~\new_[1102]_  | ~\new_[6393]_ ;
  assign n999 = ~\new_[1103]_  | ~\new_[6295]_ ;
  assign n989 = ~\new_[1107]_  | ~\new_[6376]_ ;
  assign \new_[921]_  = ~\new_[1101]_  | (~\new_[5444]_  & ~\new_[2127]_ );
  assign n1004 = ~\new_[1106]_  | ~\new_[6295]_ ;
  assign n979 = ~\new_[1108]_  | ~\new_[6304]_ ;
  assign n1009 = ~\new_[1109]_  | ~\new_[6376]_ ;
  assign \new_[925]_  = ~\new_[1128]_  | ~\new_[1180]_  | ~\new_[2411]_ ;
  assign \new_[926]_  = ~\new_[1129]_  | ~\new_[1105]_  | ~\new_[2417]_ ;
  assign \new_[927]_  = ~\new_[1130]_  | ~\new_[1105]_  | ~\new_[2617]_ ;
  assign \new_[928]_  = ~\new_[1131]_  | ~\new_[1105]_  | ~\new_[2245]_ ;
  assign \new_[929]_  = ~\new_[1132]_  | ~\new_[1105]_  | ~\new_[2243]_ ;
  assign \new_[930]_  = ~\new_[1133]_  | ~\new_[1180]_  | ~\new_[2508]_ ;
  assign \new_[931]_  = ~\new_[1135]_  | ~\new_[1105]_  | ~\new_[2420]_ ;
  assign \new_[932]_  = ~\new_[1134]_  | ~\new_[1105]_  | ~\new_[2500]_ ;
  assign n1014 = ~\new_[1112]_  | ~\new_[6393]_ ;
  assign n1019 = ~\new_[1060]_  | ~\new_[6393]_ ;
  assign n984 = ~\new_[1062]_  | ~\new_[6376]_ ;
  assign n1024 = ~\new_[1061]_  | ~\new_[6393]_ ;
  assign \new_[937]_  = ~\new_[1053]_ ;
  assign n1029 = ~\new_[1063]_  | ~\new_[6393]_ ;
  assign \new_[939]_  = ~\new_[3769]_  | (~\new_[1117]_  & ~\new_[7505]_ );
  assign \new_[940]_  = ~\new_[4007]_  | (~\new_[7433]_  & ~\new_[5490]_ );
  assign \new_[941]_  = ~\new_[4007]_  | (~\new_[1169]_  & ~\new_[5491]_ );
  assign \new_[942]_  = ~\new_[4007]_  | (~\new_[1170]_  & ~\new_[5487]_ );
  assign \new_[943]_  = ~\new_[4007]_  | (~\new_[1171]_  & ~\new_[5492]_ );
  assign \new_[944]_  = ~\new_[4007]_  | (~\new_[1172]_  & ~\new_[5488]_ );
  assign \new_[945]_  = ~\new_[4007]_  | (~\new_[1173]_  & ~\new_[5494]_ );
  assign \new_[946]_  = ~\new_[4007]_  | (~\new_[1174]_  & ~\new_[5510]_ );
  assign \new_[947]_  = ~\new_[4007]_  | (~\new_[1175]_  & ~\new_[5498]_ );
  assign \new_[948]_  = ~\new_[4007]_  | (~\new_[1176]_  & ~\new_[5489]_ );
  assign \new_[949]_  = ~\new_[4007]_  | (~\new_[1177]_  & ~\new_[5499]_ );
  assign \new_[950]_  = ~\new_[4007]_  | (~\new_[1178]_  & ~\new_[5502]_ );
  assign \new_[951]_  = ~\new_[4007]_  | (~\new_[1179]_  & ~\new_[5501]_ );
  assign \new_[952]_  = \\i_tv80_core_mcycle_reg[1] ;
  assign \new_[953]_  = (~\new_[1193]_  | ~\new_[6126]_ ) & (~\do[0]  | ~\new_[6239]_ );
  assign \new_[954]_  = (~\new_[1194]_  | ~\new_[6314]_ ) & (~\do[1]  | ~\new_[6322]_ );
  assign \new_[955]_  = (~\new_[1195]_  | ~\new_[6714]_ ) & (~\do[2]  | ~\new_[6225]_ );
  assign \new_[956]_  = (~\new_[1196]_  | ~\new_[6714]_ ) & (~\do[3]  | ~\new_[6225]_ );
  assign \new_[957]_  = \new_[5670]_  ? \new_[2127]_  : \new_[1197]_ ;
  assign \new_[958]_  = \new_[5562]_  ? \new_[2127]_  : \new_[1198]_ ;
  assign \new_[959]_  = ~\new_[770]_  | ~\new_[1118]_ ;
  assign \new_[960]_  = ~\new_[772]_  | ~\new_[1118]_ ;
  assign \new_[961]_  = ~\new_[533]_  | ~\new_[1119]_ ;
  assign \new_[962]_  = ~\new_[767]_  | ~\new_[1118]_ ;
  assign \new_[963]_  = ~\new_[730]_  | ~\new_[1118]_ ;
  assign \new_[964]_  = ~\new_[659]_  | ~\new_[1118]_ ;
  assign \new_[965]_  = ~\new_[650]_  | ~\new_[1118]_ ;
  assign \new_[966]_  = ~\new_[528]_  | ~\new_[1119]_ ;
  assign \new_[967]_  = ~\new_[567]_  | ~\new_[1118]_ ;
  assign \new_[968]_  = ~\new_[768]_  | ~\new_[1118]_ ;
  assign \new_[969]_  = ~\new_[731]_  | ~\new_[1118]_ ;
  assign \new_[970]_  = ~\new_[660]_  | ~\new_[1118]_ ;
  assign \new_[971]_  = ~\new_[652]_  | ~\new_[1118]_ ;
  assign \new_[972]_  = ~\new_[773]_  | ~\new_[1118]_ ;
  assign \new_[973]_  = ~\new_[529]_  | ~\new_[1119]_ ;
  assign \new_[974]_  = ~\new_[568]_  | ~\new_[1118]_ ;
  assign \new_[975]_  = ~\new_[735]_  | ~\new_[1118]_ ;
  assign \new_[976]_  = ~\new_[769]_  | ~\new_[1118]_ ;
  assign \new_[977]_  = ~\new_[661]_  | ~\new_[1119]_ ;
  assign \new_[978]_  = ~\new_[653]_  | ~\new_[1119]_ ;
  assign \new_[979]_  = ~\new_[530]_  | ~\new_[1118]_ ;
  assign \new_[980]_  = ~\new_[569]_  | ~\new_[1118]_ ;
  assign \new_[981]_  = ~\new_[732]_  | ~\new_[1118]_ ;
  assign \new_[982]_  = ~\new_[662]_  | ~\new_[1119]_ ;
  assign \new_[983]_  = ~\new_[654]_  | ~\new_[1119]_ ;
  assign \new_[984]_  = ~\new_[534]_  | ~\new_[1119]_ ;
  assign \new_[985]_  = ~\new_[570]_  | ~\new_[1118]_ ;
  assign \new_[986]_  = ~\new_[796]_  | ~\new_[1118]_ ;
  assign \new_[987]_  = ~\new_[733]_  | ~\new_[1118]_ ;
  assign \new_[988]_  = ~\new_[646]_  | ~\new_[1118]_ ;
  assign \new_[989]_  = ~\new_[535]_  | ~\new_[1118]_ ;
  assign \new_[990]_  = ~\new_[571]_  | ~\new_[1119]_ ;
  assign \new_[991]_  = (~\new_[1148]_  | ~\new_[6224]_ ) & (~\new_[6472]_  | ~\new_[6299]_ );
  assign \new_[992]_  = ~\new_[771]_  | ~\new_[1118]_ ;
  assign \new_[993]_  = ~\new_[6602]_  | ~\new_[1119]_ ;
  assign \new_[994]_  = ~\new_[665]_  | ~\new_[1118]_ ;
  assign \new_[995]_  = ~\new_[656]_  | ~\new_[1118]_ ;
  assign \new_[996]_  = ~\new_[531]_  | ~\new_[1118]_ ;
  assign \new_[997]_  = ~\new_[572]_  | ~\new_[1118]_ ;
  assign \new_[998]_  = ~\new_[686]_  | ~\new_[1119]_ ;
  assign \new_[999]_  = ~\new_[663]_  | ~\new_[1119]_ ;
  assign \new_[1000]_  = ~\new_[532]_  | ~\new_[1118]_ ;
  assign \new_[1001]_  = ~\new_[573]_  | ~\new_[1119]_ ;
  assign \new_[1002]_  = ~\new_[734]_  | ~\new_[1119]_ ;
  assign \new_[1003]_  = ~\new_[664]_  | ~\new_[1119]_ ;
  assign \new_[1004]_  = ~\new_[658]_  | ~\new_[1119]_ ;
  assign \new_[1005]_  = ~\new_[1118]_  | ~\new_[562]_ ;
  assign \new_[1006]_  = ~\new_[655]_  | ~\new_[1118]_ ;
  assign \new_[1007]_  = ~\new_[657]_  | ~\new_[1118]_ ;
  assign \new_[1008]_  = (~\new_[1203]_  | ~\new_[6326]_ ) & (~\new_[740]_  | ~\new_[6190]_ );
  assign \new_[1009]_  = (~\new_[1199]_  | ~\new_[6387]_ ) & (~\new_[793]_  | ~\new_[6334]_ );
  assign \new_[1010]_  = (~\new_[1200]_  | ~\new_[6220]_ ) & (~\new_[794]_  | ~\new_[6226]_ );
  assign \new_[1011]_  = (~\new_[1201]_  | ~\new_[6220]_ ) & (~\new_[742]_  | ~\new_[6226]_ );
  assign \new_[1012]_  = (~\new_[1202]_  | ~\new_[6326]_ ) & (~\new_[792]_  | ~\new_[6334]_ );
  assign \new_[1013]_  = (~\new_[1165]_  | ~\new_[6224]_ ) & (~\new_[755]_  | ~\new_[6226]_ );
  assign \new_[1014]_  = (~\new_[1166]_  | ~\new_[6263]_ ) & (~\do[7]  | ~\new_[6239]_ );
  assign \new_[1015]_  = (~\new_[1167]_  | ~\new_[6224]_ ) & (~\new_[6520]_  | ~\new_[6299]_ );
  assign \new_[1016]_  = (~\new_[1168]_  | ~\new_[6224]_ ) & (~\new_[753]_  | ~\new_[6334]_ );
  assign \new_[1017]_  = ~\new_[1127]_  | ~\new_[2530]_ ;
  assign \new_[1018]_  = ~\new_[1127]_  | ~\new_[7383]_ ;
  assign \new_[1019]_  = ~\new_[1127]_  | ~\new_[2710]_ ;
  assign \new_[1020]_  = ~\new_[1127]_  | ~\new_[2524]_ ;
  assign \new_[1021]_  = ~\new_[1127]_  | ~\new_[2526]_ ;
  assign \new_[1022]_  = ~\new_[1127]_  | ~\new_[7426]_ ;
  assign \new_[1023]_  = ~\new_[1127]_  | ~\new_[2624]_ ;
  assign \new_[1024]_  = ~\new_[1127]_  | ~\new_[7498]_ ;
  assign \new_[1025]_  = (~\new_[1147]_  | ~\new_[6224]_ ) & (~\new_[757]_  | ~\new_[6299]_ );
  assign \new_[1026]_  = (~\new_[1149]_  | ~\new_[6714]_ ) & (~\do[6]  | ~\new_[6225]_ );
  assign \new_[1027]_  = (~\new_[1136]_  | ~\new_[6162]_ ) & (~\new_[764]_  | ~\new_[6258]_ );
  assign \new_[1028]_  = (~\new_[1137]_  | ~\new_[6132]_ ) & (~\do[5]  | ~\new_[6438]_ );
  assign \new_[1029]_  = (~\new_[1150]_  | ~\new_[6220]_ ) & (~\new_[758]_  | ~\new_[6334]_ );
  assign \new_[1030]_  = (~\new_[1151]_  | ~\new_[6224]_ ) & (~\new_[759]_  | ~\new_[6299]_ );
  assign \new_[1031]_  = (~\new_[1152]_  | ~\new_[6220]_ ) & (~\new_[760]_  | ~\new_[6334]_ );
  assign \new_[1032]_  = \\i_tv80_core_mcycle_reg[2] ;
  assign \new_[1033]_  = ~\new_[1114]_  | ~\new_[2530]_ ;
  assign \new_[1034]_  = ~\new_[1114]_  | ~\new_[7383]_ ;
  assign \new_[1035]_  = ~\new_[1114]_  | ~\new_[2710]_ ;
  assign \new_[1036]_  = ~\new_[1139]_  | ~\new_[1180]_ ;
  assign \new_[1037]_  = ~\new_[1145]_  | ~\new_[1180]_ ;
  assign \new_[1038]_  = ~\new_[1140]_  | ~\new_[1180]_ ;
  assign \new_[1039]_  = ~\new_[1144]_  | ~\new_[1180]_ ;
  assign \new_[1040]_  = ~\new_[1114]_  | ~\new_[2524]_ ;
  assign \new_[1041]_  = ~\new_[1141]_  | ~\new_[1180]_ ;
  assign \new_[1042]_  = ~\new_[1114]_  | ~\new_[2526]_ ;
  assign \new_[1043]_  = ~\new_[1142]_  | ~\new_[1180]_ ;
  assign \new_[1044]_  = ~\new_[1114]_  | ~\new_[7426]_ ;
  assign \new_[1045]_  = ~\new_[1143]_  | ~\new_[1180]_ ;
  assign \new_[1046]_  = ~\new_[1114]_  | ~\new_[2624]_ ;
  assign \new_[1047]_  = ~\new_[1138]_  | ~\new_[1180]_ ;
  assign \new_[1048]_  = ~\new_[1114]_  | ~\new_[7498]_ ;
  assign \new_[1049]_  = ~\new_[3033]_  & (~\new_[1158]_  | ~\new_[7482]_ );
  assign \new_[1050]_  = (~\new_[1155]_  | ~\new_[6224]_ ) & (~\new_[766]_  | ~\new_[6334]_ );
  assign \new_[1051]_  = (~\new_[1156]_  | ~\new_[6714]_ ) & (~\do[4]  | ~\new_[6225]_ );
  assign \new_[1052]_  = \\i_tv80_core_mcycle_reg[0] ;
  assign \new_[1053]_  = \new_[1884]_  ? \new_[1154]_  : \new_[1833]_ ;
  assign \new_[1054]_  = (~\new_[1160]_  | ~\new_[6387]_ ) & (~\new_[761]_  | ~\new_[6334]_ );
  assign \new_[1055]_  = ~\new_[1206]_  | (~\new_[1164]_  & ~\new_[1343]_ );
  assign \new_[1056]_  = (~\new_[1161]_  | ~\new_[6387]_ ) & (~\new_[763]_  | ~\new_[6334]_ );
  assign \new_[1057]_  = (~\new_[1163]_  | ~\new_[6348]_ ) & (~\new_[762]_  | ~\new_[6226]_ );
  assign \new_[1058]_  = (~\new_[1162]_  | ~\new_[6387]_ ) & (~\new_[736]_  | ~\new_[6226]_ );
  assign \new_[1059]_  = ~\new_[1157]_  | ~\new_[1116]_ ;
  assign \new_[1060]_  = (~\new_[1218]_  | ~\new_[6348]_ ) & (~\new_[851]_  | ~\new_[6334]_ );
  assign \new_[1061]_  = (~\new_[1219]_  | ~\new_[6348]_ ) & (~\new_[852]_  | ~\new_[6334]_ );
  assign \new_[1062]_  = (~\new_[1212]_  | ~\new_[6220]_ ) & (~\new_[844]_  | ~\new_[6334]_ );
  assign \new_[1063]_  = (~\new_[1222]_  | ~\new_[6326]_ ) & (~\new_[853]_  | ~\new_[6334]_ );
  assign \new_[1064]_  = ~\new_[1274]_  | (~\new_[1224]_  & ~\new_[1547]_ );
  assign \new_[1065]_  = ~\new_[428]_  | ~\new_[1187]_ ;
  assign \new_[1066]_  = ~\new_[6491]_  | ~\new_[1187]_ ;
  assign \new_[1067]_  = ~\new_[6644]_  | ~\new_[1187]_ ;
  assign \new_[1068]_  = ~\new_[6598]_  | ~\new_[1185]_ ;
  assign \new_[1069]_  = ~\new_[575]_  | ~\new_[1192]_ ;
  assign \new_[1070]_  = ~\new_[6618]_  | ~\new_[1192]_ ;
  assign \new_[1071]_  = ~\new_[6627]_  | ~\new_[1185]_ ;
  assign \new_[1072]_  = ~\new_[576]_  | ~\new_[1192]_ ;
  assign \new_[1073]_  = ~\new_[538]_  | ~\new_[1192]_ ;
  assign \new_[1074]_  = ~\new_[6615]_  | ~\new_[1182]_ ;
  assign \new_[1075]_  = ~\new_[577]_  | ~\new_[1182]_ ;
  assign \new_[1076]_  = ~\new_[539]_  | ~\new_[1181]_ ;
  assign \new_[1077]_  = ~\new_[431]_  | ~\new_[1182]_ ;
  assign \new_[1078]_  = ~\new_[6583]_  | ~\new_[1181]_ ;
  assign \new_[1079]_  = ~\new_[6641]_  | ~\new_[1184]_ ;
  assign \new_[1080]_  = ~\new_[6556]_  | ~\new_[1188]_ ;
  assign \new_[1081]_  = ~\new_[6660]_  | ~\new_[1184]_ ;
  assign \new_[1082]_  = ~\new_[560]_  | ~\new_[1192]_ ;
  assign \new_[1083]_  = ~\new_[540]_  | ~\new_[1184]_ ;
  assign \new_[1084]_  = ~\new_[432]_  | ~\new_[1188]_ ;
  assign \new_[1085]_  = ~\new_[6639]_  | ~\new_[1192]_ ;
  assign \new_[1086]_  = ~\new_[6587]_  | ~\new_[1181]_ ;
  assign \new_[1087]_  = ~\new_[6657]_  | ~\new_[1183]_ ;
  assign \new_[1088]_  = ~\new_[6599]_  | ~\new_[1182]_ ;
  assign \new_[1089]_  = ~\new_[578]_  | ~\new_[1188]_ ;
  assign \new_[1090]_  = ~\new_[520]_  | ~\new_[1183]_ ;
  assign \new_[1091]_  = ~\new_[6612]_  | ~\new_[1182]_ ;
  assign \new_[1092]_  = ~\new_[579]_  | ~\new_[1188]_ ;
  assign \new_[1093]_  = ~\new_[6597]_  | ~\new_[1183]_ ;
  assign \new_[1094]_  = ~\new_[580]_  | ~\new_[1192]_ ;
  assign \new_[1095]_  = ~\new_[543]_  | ~\new_[1188]_ ;
  assign \new_[1096]_  = ~\new_[435]_  | ~\new_[1181]_ ;
  assign \new_[1097]_  = ~\new_[6607]_  | ~\new_[1188]_ ;
  assign \new_[1098]_  = ~\new_[6665]_  | ~\new_[1185]_ ;
  assign \new_[1099]_  = ~\new_[6673]_  | ~\new_[1181]_ ;
  assign \new_[1100]_  = ~\new_[6652]_  | ~\new_[1185]_ ;
  assign \new_[1101]_  = ~\new_[1226]_  | ~\new_[2127]_  | ~\new_[1227]_ ;
  assign \new_[1102]_  = (~\new_[1229]_  | ~\new_[6220]_ ) & (~\new_[6606]_  | ~\new_[6226]_ );
  assign \new_[1103]_  = (~\new_[1230]_  | ~\new_[6220]_ ) & (~\new_[6591]_  | ~\new_[6334]_ );
  assign \new_[1104]_  = \\i_tv80_core_TmpAddr_reg[14] ;
  assign \new_[1105]_  = ~\new_[1119]_ ;
  assign \new_[1106]_  = (~\new_[1252]_  | ~\new_[6326]_ ) & (~\new_[848]_  | ~\new_[6334]_ );
  assign \new_[1107]_  = (~\new_[1221]_  | ~\new_[6348]_ ) & (~\new_[845]_  | ~\new_[6226]_ );
  assign \new_[1108]_  = (~\new_[1208]_  | ~\new_[6326]_ ) & (~\new_[799]_  | ~\new_[6190]_ );
  assign \new_[1109]_  = (~\new_[1209]_  | ~\new_[6224]_ ) & (~\new_[849]_  | ~\new_[6334]_ );
  assign \new_[1110]_  = ~i_tv80_core_IntE_FF1_reg;
  assign \new_[1111]_  = ~i_tv80_core_IntE_FF2_reg;
  assign \new_[1112]_  = (~\new_[1211]_  | ~\new_[6220]_ ) & (~\new_[850]_  | ~\new_[6334]_ );
  assign \new_[1113]_  = ~\new_[3192]_  & (~\new_[1268]_  | ~\new_[7482]_ );
  assign \new_[1114]_  = ~\new_[1146]_ ;
  assign m1_n = i_tv80_core_m1_n_reg;
  assign \new_[1116]_  = ~\new_[1158]_ ;
  assign \new_[1117]_  = ~\new_[2523]_  & (~\new_[1269]_  | ~\new_[7482]_ );
  assign \new_[1118]_  = ~\new_[1180]_ ;
  assign \new_[1119]_  = ~\new_[1180]_ ;
  assign n1044 = ~\new_[1251]_  | ~\new_[6295]_ ;
  assign n1034 = ~\new_[5340]_  | ~\new_[1249]_ ;
  assign n1039 = ~\new_[5338]_  | ~\new_[1250]_ ;
  assign \new_[1123]_  = i_tv80_core_IntCycle_reg;
  assign \new_[1124]_  = i_tv80_core_NMICycle_reg;
  assign \new_[1125]_  = \\i_tv80_core_BusA_reg[0] ;
  assign \new_[1126]_  = \\i_tv80_core_BusA_reg[5] ;
  assign \new_[1127]_  = ~\new_[1207]_ ;
  assign \new_[1128]_  = ~\new_[1210]_  | ~\new_[7398]_ ;
  assign \new_[1129]_  = ~\new_[1210]_  | ~\new_[7383]_ ;
  assign \new_[1130]_  = ~\new_[1210]_  | ~\new_[7389]_ ;
  assign \new_[1131]_  = ~\new_[1210]_  | ~\new_[2524]_ ;
  assign \new_[1132]_  = ~\new_[1210]_  | ~\new_[2526]_ ;
  assign \new_[1133]_  = ~\new_[1210]_  | ~\new_[7426]_ ;
  assign \new_[1134]_  = ~\new_[1210]_  | ~\new_[7498]_ ;
  assign \new_[1135]_  = ~\new_[1210]_  | ~\new_[7514]_ ;
  assign \new_[1136]_  = ~\new_[1279]_  | (~\new_[1547]_  & ~\new_[1947]_ );
  assign \new_[1137]_  = ~\new_[1287]_  | (~\new_[1381]_  & ~\new_[1354]_ );
  assign \new_[1138]_  = ~\new_[2518]_  & (~\new_[1318]_  | ~\new_[7498]_ );
  assign \new_[1139]_  = ~\new_[2410]_  & (~\new_[1318]_  | ~\new_[7398]_ );
  assign \new_[1140]_  = ~\new_[2620]_  & (~\new_[1318]_  | ~\new_[7389]_ );
  assign \new_[1141]_  = ~\new_[2355]_  & (~\new_[1318]_  | ~\new_[2526]_ );
  assign \new_[1142]_  = ~\new_[2510]_  & (~\new_[1318]_  | ~\new_[7426]_ );
  assign \new_[1143]_  = ~\new_[2493]_  & (~\new_[1318]_  | ~\new_[7514]_ );
  assign \new_[1144]_  = ~\new_[2346]_  & (~\new_[1318]_  | ~\new_[2524]_ );
  assign \new_[1145]_  = ~\new_[2483]_  & (~\new_[1318]_  | ~\new_[7383]_ );
  assign \new_[1146]_  = ~\new_[3770]_  | (~\new_[1317]_  & ~\new_[7505]_ );
  assign \new_[1147]_  = ~\new_[1280]_  | (~\new_[1547]_  & ~\new_[1839]_ );
  assign \new_[1148]_  = ~\new_[1275]_  | (~\new_[1343]_  & ~\new_[1562]_ );
  assign \new_[1149]_  = ~\new_[1288]_  | (~\new_[1381]_  & ~\new_[1357]_ );
  assign \new_[1150]_  = ~\new_[1272]_  | (~\new_[1344]_  & ~\new_[1438]_ );
  assign \new_[1151]_  = ~\new_[1273]_  | (~\new_[1439]_  & ~\new_[1547]_ );
  assign \new_[1152]_  = ~\new_[1298]_  | (~\new_[1344]_  & ~\new_[1470]_ );
  assign \new_[1153]_  = ~\new_[1269]_  & ~\new_[1448]_ ;
  assign \new_[1154]_  = ~\new_[1412]_  & (~\new_[7548]_  | ~\new_[1492]_ );
  assign \new_[1155]_  = ~\new_[1278]_  | (~\new_[1547]_  & ~\new_[2042]_ );
  assign \new_[1156]_  = ~\new_[1286]_  | (~\new_[1381]_  & ~\new_[1358]_ );
  assign \new_[1157]_  = ~\new_[7476]_ ;
  assign \new_[1158]_  = \new_[1556]_  ? \new_[7547]_  : \new_[1599]_ ;
  assign n1049 = ~\new_[1270]_  & ~\new_[6323]_ ;
  assign \new_[1160]_  = ~\new_[1296]_  | (~\new_[1381]_  & ~\new_[1449]_ );
  assign \new_[1161]_  = ~\new_[1297]_  | (~\new_[1344]_  & ~\new_[1476]_ );
  assign \new_[1162]_  = ~\new_[1300]_  | (~\new_[1381]_  & ~\new_[1450]_ );
  assign \new_[1163]_  = ~\new_[1295]_  | (~\new_[1381]_  & ~\new_[1477]_ );
  assign \new_[1164]_  = \new_[3419]_  ? \new_[6243]_  : \new_[1312]_ ;
  assign \new_[1165]_  = ~\new_[1281]_  | (~\new_[1344]_  & ~\new_[1981]_ );
  assign \new_[1166]_  = ~\new_[1289]_  | (~\new_[1381]_  & ~\new_[1352]_ );
  assign \new_[1167]_  = ~\new_[1256]_  | (~\new_[1381]_  & ~\new_[1496]_ );
  assign \new_[1168]_  = ~\new_[1299]_  | (~\new_[1344]_  & ~\new_[1463]_ );
  assign \new_[1169]_  = ~\new_[7440]_  & (~\new_[1339]_  | ~\new_[4471]_ );
  assign \new_[1170]_  = ~\new_[7440]_  & (~\new_[1340]_  | ~\new_[4472]_ );
  assign \new_[1171]_  = ~\new_[7440]_  & (~\new_[1341]_  | ~\new_[4390]_ );
  assign \new_[1172]_  = ~\new_[7440]_  & (~\new_[1342]_  | ~\new_[4391]_ );
  assign \new_[1173]_  = ~\new_[7440]_  & (~\new_[1345]_  | ~\new_[4473]_ );
  assign \new_[1174]_  = ~\new_[7440]_  & (~\new_[1346]_  | ~\new_[4572]_ );
  assign \new_[1175]_  = ~\new_[7440]_  & (~\new_[1347]_  | ~\new_[4395]_ );
  assign \new_[1176]_  = ~\new_[7440]_  & (~\new_[1348]_  | ~\new_[4475]_ );
  assign \new_[1177]_  = ~\new_[7440]_  & (~\new_[1349]_  | ~\new_[4477]_ );
  assign \new_[1178]_  = ~\new_[7440]_  & (~\new_[1350]_  | ~\new_[4478]_ );
  assign \new_[1179]_  = ~\new_[7440]_  & (~\new_[1351]_  | ~\new_[4479]_ );
  assign \new_[1180]_  = ~\new_[1690]_  & (~\new_[1321]_  | ~\new_[4930]_ );
  assign \new_[1181]_  = ~\new_[7515]_ ;
  assign \new_[1182]_  = ~\new_[7515]_ ;
  assign \new_[1183]_  = ~\new_[7515]_ ;
  assign \new_[1184]_  = ~\new_[7515]_ ;
  assign \new_[1185]_  = ~\new_[7515]_ ;
  assign \new_[1186]_  = ~\new_[7515]_ ;
  assign \new_[1187]_  = ~\new_[7515]_ ;
  assign \new_[1188]_  = ~\new_[7515]_ ;
  assign \new_[1189]_  = ~\new_[7515]_ ;
  assign \new_[1190]_  = ~\new_[7515]_ ;
  assign \new_[1191]_  = ~\new_[7515]_ ;
  assign \new_[1192]_  = ~\new_[7515]_ ;
  assign \new_[1193]_  = ~\new_[1282]_  | (~\new_[1381]_  & ~\new_[1371]_ );
  assign \new_[1194]_  = ~\new_[1283]_  | (~\new_[1381]_  & ~\new_[1372]_ );
  assign \new_[1195]_  = ~\new_[1284]_  | (~\new_[1381]_  & ~\new_[1373]_ );
  assign \new_[1196]_  = ~\new_[1285]_  | (~\new_[1381]_  & ~\new_[1374]_ );
  assign \new_[1197]_  = ~\new_[1271]_  & (~\new_[1369]_  | ~\new_[597]_ );
  assign \new_[1198]_  = \new_[595]_  ^ \new_[1322]_ ;
  assign \new_[1199]_  = ~\new_[1277]_  | (~\new_[1343]_  & ~\new_[2092]_ );
  assign \new_[1200]_  = ~\new_[1290]_  | (~\new_[1344]_  & ~\new_[2452]_ );
  assign \new_[1201]_  = ~\new_[1291]_  | (~\new_[1343]_  & ~\new_[2306]_ );
  assign \new_[1202]_  = ~\new_[1276]_  | (~\new_[1344]_  & ~\new_[2149]_ );
  assign \new_[1203]_  = ~\new_[1258]_  | (~\new_[1547]_  & ~\new_[1499]_ );
  assign n1059 = ~\new_[1254]_  & ~\new_[6424]_ ;
  assign n1054 = ~\new_[6441]_  & (~\new_[3652]_  | ~\new_[1309]_ );
  assign \new_[1206]_  = ~\new_[1257]_  | ~\new_[1381]_ ;
  assign \new_[1207]_  = ~\new_[3867]_  | (~\new_[1311]_  & ~\new_[7505]_ );
  assign \new_[1208]_  = \new_[1530]_  ? \new_[1381]_  : \new_[1614]_ ;
  assign \new_[1209]_  = \new_[1568]_  ? \new_[1380]_  : \new_[1684]_ ;
  assign \new_[1210]_  = ~\new_[1267]_ ;
  assign \new_[1211]_  = \new_[1653]_  ? \new_[1380]_  : \new_[1843]_ ;
  assign \new_[1212]_  = \new_[1919]_  ? \new_[1381]_  : \new_[2081]_ ;
  assign \new_[1213]_  = ~\new_[1319]_  | ~\new_[1479]_ ;
  assign \new_[1214]_  = \new_[1319]_  & \new_[1479]_ ;
  assign \new_[1215]_  = ~\new_[1320]_  & ~\new_[1441]_ ;
  assign n1084 = \new_[1359]_  ? \new_[1690]_  : \new_[1126]_ ;
  assign n1079 = \new_[1360]_  ? \new_[6347]_  : \new_[6478]_ ;
  assign \new_[1218]_  = \new_[1731]_  ? \new_[1380]_  : \new_[1847]_ ;
  assign \new_[1219]_  = \new_[1616]_  ? \new_[1380]_  : \new_[1738]_ ;
  assign \new_[1220]_  = ~\new_[1268]_ ;
  assign \new_[1221]_  = \new_[1495]_  ? \new_[1380]_  : \new_[1571]_ ;
  assign \new_[1222]_  = \new_[1845]_  ? \new_[1380]_  : \new_[1960]_ ;
  assign \new_[1223]_  = \\i_tv80_core_PC_reg[9] ;
  assign \new_[1224]_  = ~\new_[1323]_  & (~\new_[2831]_  | ~\new_[6163]_ );
  assign \new_[1225]_  = \\i_tv80_core_PC_reg[7] ;
  assign \new_[1226]_  = ~\new_[6494]_  | ~\new_[1322]_  | ~\new_[6497]_ ;
  assign \new_[1227]_  = \new_[1322]_  | \new_[596]_ ;
  assign \new_[1228]_  = ~\\i_tv80_core_Pre_XY_F_M_reg[2] ;
  assign \new_[1229]_  = \new_[1560]_  ? \new_[1380]_  : \new_[1777]_ ;
  assign \new_[1230]_  = \new_[1561]_  ? \new_[1380]_  : \new_[1778]_ ;
  assign \new_[1231]_  = \\i_tv80_core_BusA_reg[3] ;
  assign n1069 = ~\new_[1304]_  & ~\new_[6623]_ ;
  assign \new_[1233]_  = \\i_tv80_core_PC_reg[11] ;
  assign \new_[1234]_  = \\i_tv80_core_PC_reg[12] ;
  assign \new_[1235]_  = \\i_tv80_core_PC_reg[13] ;
  assign \new_[1236]_  = \\i_tv80_core_PC_reg[1] ;
  assign \new_[1237]_  = \\i_tv80_core_PC_reg[2] ;
  assign \new_[1238]_  = \\i_tv80_core_PC_reg[3] ;
  assign \new_[1239]_  = \\i_tv80_core_PC_reg[4] ;
  assign \new_[1240]_  = \\i_tv80_core_PC_reg[5] ;
  assign \new_[1241]_  = \\i_tv80_core_PC_reg[6] ;
  assign \new_[1242]_  = \\i_tv80_core_PC_reg[8] ;
  assign n1064 = ~reset_n | (~\new_[6332]_  & ~\new_[1353]_ );
  assign \new_[1244]_  = ~\\i_tv80_core_Pre_XY_F_M_reg[0] ;
  assign \new_[1245]_  = ~\\i_tv80_core_Pre_XY_F_M_reg[1] ;
  assign \new_[1246]_  = \\i_tv80_core_BusA_reg[2] ;
  assign \new_[1247]_  = \\i_tv80_core_BusA_reg[4] ;
  assign \new_[1248]_  = \\i_tv80_core_BusA_reg[6] ;
  assign \new_[1249]_  = ~\new_[1302]_  | ~\new_[6427]_ ;
  assign \new_[1250]_  = ~\new_[1303]_  | ~\new_[6427]_ ;
  assign \new_[1251]_  = ~\new_[1301]_  & (~\new_[5672]_  | ~\new_[6442]_ );
  assign \new_[1252]_  = \new_[1466]_  ? \new_[1381]_  : \new_[1569]_ ;
  assign n1074 = ~\new_[1310]_  & ~\new_[6623]_ ;
  assign \new_[1254]_  = (~\new_[1396]_  | ~\new_[6055]_ ) & (~\new_[4186]_  | ~\new_[5614]_ );
  assign \new_[1255]_  = \\i_tv80_core_PC_reg[15] ;
  assign \new_[1256]_  = ~\new_[1380]_  | ~\new_[1564]_ ;
  assign \new_[1257]_  = ~\new_[1312]_ ;
  assign \new_[1258]_  = ~\new_[1381]_  | ~\new_[1605]_ ;
  assign \new_[1259]_  = (~\new_[1403]_  | ~\new_[7398]_ ) & (~\new_[2529]_  | ~\new_[6537]_ );
  assign \new_[1260]_  = (~\new_[1403]_  | ~\new_[7383]_ ) & (~\new_[2627]_  | ~\new_[6549]_ );
  assign \new_[1261]_  = (~\new_[1403]_  | ~\new_[7389]_ ) & (~\new_[2711]_  | ~\new_[6561]_ );
  assign \new_[1262]_  = ~\new_[2344]_  & (~\new_[1403]_  | ~\new_[2524]_ );
  assign \new_[1263]_  = ~\new_[2349]_  & (~\new_[1403]_  | ~\new_[2526]_ );
  assign \new_[1264]_  = ~\new_[2491]_  & (~\new_[1403]_  | ~\new_[7426]_ );
  assign \new_[1265]_  = ~\new_[2513]_  & (~\new_[1403]_  | ~\new_[7514]_ );
  assign \new_[1266]_  = ~\new_[2492]_  & (~\new_[1403]_  | ~\new_[7498]_ );
  assign \new_[1267]_  = ~\new_[3768]_  | (~\new_[1402]_  & ~\new_[7505]_ );
  assign \new_[1268]_  = \new_[1707]_  ? \new_[1404]_  : \new_[1755]_ ;
  assign \new_[1269]_  = \new_[1709]_  ? \new_[1405]_  : \new_[1756]_ ;
  assign \new_[1270]_  = (~\new_[1414]_  | ~\new_[6314]_ ) & (~\new_[1104]_  | ~\new_[6261]_ );
  assign \new_[1271]_  = ~\new_[6330]_  & ~\new_[1369]_ ;
  assign \new_[1272]_  = ~\new_[1550]_  | ~\new_[1547]_ ;
  assign \new_[1273]_  = ~\new_[1551]_  | ~\new_[1547]_ ;
  assign \new_[1274]_  = ~\new_[1380]_  | ~\new_[1382]_ ;
  assign \new_[1275]_  = ~\new_[1650]_  | ~\new_[1381]_ ;
  assign \new_[1276]_  = ~\new_[1380]_  | ~\new_[2378]_ ;
  assign \new_[1277]_  = ~\new_[1380]_  | ~\new_[2186]_ ;
  assign \new_[1278]_  = ~\new_[1380]_  | ~\new_[2147]_ ;
  assign \new_[1279]_  = ~\new_[1380]_  | ~\new_[2087]_ ;
  assign \new_[1280]_  = ~\new_[1380]_  | ~\new_[2012]_ ;
  assign \new_[1281]_  = ~\new_[1380]_  | ~\new_[2088]_ ;
  assign \new_[1282]_  = ~\new_[1381]_  | ~\new_[1455]_ ;
  assign \new_[1283]_  = ~\new_[1381]_  | ~\new_[1456]_ ;
  assign \new_[1284]_  = ~\new_[1381]_  | ~\new_[1457]_ ;
  assign \new_[1285]_  = ~\new_[1381]_  | ~\new_[1458]_ ;
  assign \new_[1286]_  = ~\new_[1381]_  | ~\new_[1459]_ ;
  assign \new_[1287]_  = ~\new_[1381]_  | ~\new_[1460]_ ;
  assign \new_[1288]_  = ~\new_[1381]_  | ~\new_[1461]_ ;
  assign \new_[1289]_  = ~\new_[1381]_  | ~\new_[1462]_ ;
  assign \new_[1290]_  = ~\new_[1380]_  | ~\new_[2745]_ ;
  assign \new_[1291]_  = ~\new_[1380]_  | ~\new_[2574]_ ;
  assign \new_[1292]_  = \\i_tv80_core_PC_reg[14] ;
  assign \new_[1293]_  = \\i_tv80_core_PC_reg[0] ;
  assign \new_[1294]_  = \\i_tv80_core_PC_reg[10] ;
  assign \new_[1295]_  = ~\new_[1553]_  | ~\new_[1547]_ ;
  assign \new_[1296]_  = ~\new_[1498]_  | ~\new_[1547]_ ;
  assign \new_[1297]_  = ~\new_[1557]_  | ~\new_[1547]_ ;
  assign \new_[1298]_  = ~\new_[1558]_  | ~\new_[1547]_ ;
  assign \new_[1299]_  = ~\new_[1559]_  | ~\new_[1547]_ ;
  assign \new_[1300]_  = ~\new_[1497]_  | ~\new_[1380]_ ;
  assign \new_[1301]_  = ~\new_[5672]_  & (~\new_[5449]_  | ~\new_[1434]_ );
  assign \new_[1302]_  = ~\new_[5672]_  & (~\new_[1435]_  | ~\new_[5425]_ );
  assign \new_[1303]_  = ~\new_[5672]_  & (~\new_[1436]_  | ~\new_[5427]_ );
  assign \new_[1304]_  = (~\new_[1433]_  | ~\new_[5847]_ ) & (~\new_[5614]_  | ~\new_[6523]_ );
  assign n1159 = ~\new_[1399]_  & ~\new_[6424]_ ;
  assign n1164 = ~\new_[1400]_  & ~\new_[6424]_ ;
  assign n1099 = ~\new_[1401]_  & ~\new_[6424]_ ;
  assign \new_[1308]_  = \\i_tv80_core_TmpAddr_reg[10] ;
  assign \new_[1309]_  = ~\new_[5847]_  | ~\new_[6055]_  | ~\new_[1440]_ ;
  assign \new_[1310]_  = (~\new_[1437]_  | ~\new_[5847]_ ) & (~\new_[5614]_  | ~\new_[6519]_ );
  assign \new_[1311]_  = ~\new_[2794]_  & (~\new_[1441]_  | ~\new_[7482]_ );
  assign \new_[1312]_  = ~\new_[1409]_  & (~\new_[4415]_  | ~\new_[407]_ );
  assign n1169 = \new_[1442]_  ? \new_[6258]_  : \new_[6518]_ ;
  assign n1104 = \new_[6542]_  ? \new_[6162]_  : \new_[1443]_ ;
  assign n1174 = \new_[1444]_  ? \new_[1690]_  : \new_[1247]_ ;
  assign n1179 = \new_[1445]_  ? \new_[6258]_  : \new_[1248]_ ;
  assign \new_[1317]_  = ~\new_[2807]_  & (~\new_[1448]_  | ~\new_[7482]_ );
  assign \new_[1318]_  = (~\new_[1447]_  | ~\new_[7501]_ ) & (~\new_[3937]_  | ~\new_[7505]_ );
  assign \new_[1319]_  = ~\new_[1405]_  | ~\new_[1698]_ ;
  assign \new_[1320]_  = ~\new_[1406]_  | (~\new_[7068]_  & ~\new_[1708]_ );
  assign \new_[1321]_  = \new_[1411]_  & \new_[3562]_ ;
  assign \new_[1322]_  = ~\new_[1369]_ ;
  assign \new_[1323]_  = ~\new_[1415]_  & ~\new_[5813]_ ;
  assign \new_[1324]_  = \\i_tv80_core_BusA_reg[7] ;
  assign n1109 = ~\new_[1383]_  & ~\new_[6323]_ ;
  assign n1114 = ~\new_[1384]_  & ~\new_[6403]_ ;
  assign n1119 = ~\new_[6708]_  & ~\new_[6327]_ ;
  assign n1124 = ~\new_[1385]_  & ~\new_[6424]_ ;
  assign n1129 = ~\new_[1386]_  & ~\new_[6426]_ ;
  assign n1134 = ~\new_[1387]_  & ~\new_[6323]_ ;
  assign n1139 = ~\new_[1388]_  & ~\new_[6417]_ ;
  assign n1144 = ~\new_[1389]_  & ~\new_[6623]_ ;
  assign n1149 = ~\new_[1390]_  & ~\new_[6623]_ ;
  assign n1094 = ~\new_[1391]_  & ~\new_[6424]_ ;
  assign n1154 = ~\new_[1392]_  & ~\new_[6623]_ ;
  assign n1089 = ~\new_[1393]_  & ~\new_[6424]_ ;
  assign \new_[1337]_  = ~\\i_tv80_core_TmpAddr_reg[15] ;
  assign \new_[1338]_  = \\i_tv80_core_BusA_reg[1] ;
  assign \new_[1339]_  = \new_[1417]_  | \new_[7436]_ ;
  assign \new_[1340]_  = \new_[1418]_  | \new_[7436]_ ;
  assign \new_[1341]_  = \new_[1419]_  | \new_[7436]_ ;
  assign \new_[1342]_  = \new_[1420]_  | \new_[7436]_ ;
  assign \new_[1343]_  = ~\new_[1483]_ ;
  assign \new_[1344]_  = ~\new_[1483]_ ;
  assign \new_[1345]_  = \new_[1421]_  | \new_[7436]_ ;
  assign \new_[1346]_  = \new_[1422]_  | \new_[7436]_ ;
  assign \new_[1347]_  = \new_[1423]_  | \new_[7436]_ ;
  assign \new_[1348]_  = \new_[1424]_  | \new_[7436]_ ;
  assign \new_[1349]_  = \new_[1425]_  | \new_[7436]_ ;
  assign \new_[1350]_  = \new_[1426]_  | \new_[7436]_ ;
  assign \new_[1351]_  = \new_[1427]_  | \new_[7436]_ ;
  assign \new_[1352]_  = ~\new_[1410]_  & (~\new_[2471]_  | ~\new_[6246]_ );
  assign \new_[1353]_  = (~\new_[1469]_  | ~\new_[5847]_ ) & (~\new_[3555]_  | ~\new_[5614]_ );
  assign \new_[1354]_  = \new_[1489]_  ? \new_[6246]_  : \new_[2969]_ ;
  assign \new_[1355]_  = ~\new_[1478]_  | ~\new_[1446]_ ;
  assign \new_[1356]_  = ~\new_[6842]_ ;
  assign \new_[1357]_  = \new_[1490]_  ? \new_[6246]_  : \new_[2787]_ ;
  assign \new_[1358]_  = \new_[1488]_  ? \new_[6246]_  : \new_[2977]_ ;
  assign \new_[1359]_  = ~\new_[1548]_  | ~\new_[3100]_  | ~\new_[2903]_  | ~\new_[2912]_ ;
  assign \new_[1360]_  = ~\new_[1549]_  | ~\new_[3097]_  | ~\new_[2900]_  | ~\new_[2917]_ ;
  assign \new_[1361]_  = (~\new_[1480]_  | ~\new_[7398]_ ) & (~\new_[2529]_  | ~\new_[6545]_ );
  assign \new_[1362]_  = ~\new_[2517]_  & (~\new_[1480]_  | ~\new_[7498]_ );
  assign \new_[1363]_  = (~\new_[1480]_  | ~\new_[7383]_ ) & (~\new_[2627]_  | ~\new_[6610]_ );
  assign \new_[1364]_  = (~\new_[1480]_  | ~\new_[7389]_ ) & (~\new_[2711]_  | ~\new_[6600]_ );
  assign \new_[1365]_  = ~\new_[2345]_  & (~\new_[1480]_  | ~\new_[2524]_ );
  assign \new_[1366]_  = ~\new_[2356]_  & (~\new_[1480]_  | ~\new_[2526]_ );
  assign \new_[1367]_  = ~\new_[2509]_  & (~\new_[1480]_  | ~\new_[7426]_ );
  assign \new_[1368]_  = ~\new_[2504]_  & (~\new_[1480]_  | ~\new_[7514]_ );
  assign \new_[1369]_  = \new_[1452]_  & \new_[3546]_ ;
  assign \new_[1370]_  = \new_[1451]_  & \new_[3562]_ ;
  assign \new_[1371]_  = \new_[1484]_  ? \new_[6246]_  : \new_[3840]_ ;
  assign \new_[1372]_  = \new_[1485]_  ? \new_[6246]_  : \new_[3623]_ ;
  assign \new_[1373]_  = \new_[1486]_  ? \new_[6246]_  : \new_[3419]_ ;
  assign \new_[1374]_  = \new_[1487]_  ? \new_[6246]_  : \new_[3180]_ ;
  assign n1194 = ~\new_[1428]_  & ~\new_[6424]_ ;
  assign n1199 = ~\new_[1429]_  & ~\new_[6424]_ ;
  assign n1189 = ~\new_[6623]_  & ~\new_[1430]_ ;
  assign n1184 = ~\new_[1431]_  & ~\new_[6424]_ ;
  assign \new_[1379]_  = \\i_tv80_core_TmpAddr_reg[12] ;
  assign \new_[1380]_  = ~\new_[1483]_ ;
  assign \new_[1381]_  = ~\new_[1483]_ ;
  assign \new_[1382]_  = ~\new_[1415]_ ;
  assign \new_[1383]_  = (~\new_[1518]_  | ~\new_[6099]_ ) & (~\new_[1233]_  | ~\new_[1690]_ );
  assign \new_[1384]_  = (~\new_[1519]_  | ~\new_[6714]_ ) & (~\new_[1234]_  | ~\new_[6261]_ );
  assign \new_[1385]_  = (~\new_[1520]_  | ~\new_[6099]_ ) & (~\new_[1236]_  | ~\new_[6225]_ );
  assign \new_[1386]_  = (~\new_[1521]_  | ~\new_[6132]_ ) & (~\new_[1237]_  | ~\new_[6438]_ );
  assign \new_[1387]_  = (~\new_[1522]_  | ~\new_[6714]_ ) & (~\new_[1238]_  | ~\new_[6165]_ );
  assign \new_[1388]_  = (~\new_[1523]_  | ~\new_[6129]_ ) & (~\new_[1239]_  | ~\new_[6239]_ );
  assign \new_[1389]_  = (~\new_[1524]_  | ~\new_[6132]_ ) & (~\new_[1240]_  | ~\new_[6225]_ );
  assign \new_[1390]_  = (~\new_[1525]_  | ~\new_[6129]_ ) & (~\new_[1241]_  | ~\new_[6261]_ );
  assign \new_[1391]_  = (~\new_[1526]_  | ~\new_[6129]_ ) & (~\new_[1225]_  | ~\new_[6165]_ );
  assign \new_[1392]_  = (~\new_[1527]_  | ~\new_[6314]_ ) & (~\new_[1242]_  | ~\new_[6165]_ );
  assign \new_[1393]_  = (~\new_[1528]_  | ~busak_n) & (~\new_[1223]_  | ~\new_[6438]_ );
  assign \new_[1394]_  = \\i_tv80_core_TmpAddr_reg[13] ;
  assign n1214 = ~\new_[1468]_  & ~\new_[6424]_ ;
  assign \new_[1396]_  = ~\new_[1471]_  & ~\new_[5672]_ ;
  assign n1219 = \new_[1533]_  ? \new_[1690]_  : \new_[6515]_ ;
  assign n1209 = \new_[1324]_  ? \new_[6162]_  : \new_[1534]_ ;
  assign \new_[1399]_  = (~\new_[1535]_  | ~\new_[5847]_ ) & (~\new_[6663]_  | ~\new_[5614]_ );
  assign \new_[1400]_  = (~\new_[1536]_  | ~\new_[5847]_ ) & (~\new_[6667]_  | ~\new_[5614]_ );
  assign \new_[1401]_  = (~\new_[1537]_  | ~\new_[5847]_ ) & (~\new_[6674]_  | ~\new_[5614]_ );
  assign \new_[1402]_  = ~\new_[3034]_  & (~\new_[7406]_  | ~\new_[7482]_ );
  assign \new_[1403]_  = (~\new_[1540]_  | ~\new_[7501]_ ) & (~\new_[3936]_  | ~\new_[7505]_ );
  assign \new_[1404]_  = ~\new_[1473]_  | ~\new_[1543]_ ;
  assign \new_[1405]_  = ~\new_[1474]_  | ~\new_[1820]_ ;
  assign \new_[1406]_  = ~\new_[7068]_  | ~\new_[1708]_ ;
  assign \new_[1407]_  = ~\new_[7312]_  & (~\new_[1542]_  | ~\new_[1704]_ );
  assign \new_[1408]_  = ~\new_[7069]_  | ~\new_[1697]_ ;
  assign \new_[1409]_  = ~\new_[1467]_  & ~\new_[4415]_ ;
  assign \new_[1410]_  = ~\new_[1491]_  & ~\new_[6246]_ ;
  assign \new_[1411]_  = ~\new_[6634]_  | ~\new_[1483]_  | ~\new_[6277]_ ;
  assign \new_[1412]_  = ~\new_[1482]_  | ~\new_[7327]_ ;
  assign \new_[1413]_  = i_tv80_core_BTR_r_reg;
  assign \new_[1414]_  = ~\new_[1493]_  | (~\new_[1779]_  & ~\new_[6047]_ );
  assign \new_[1415]_  = ~\new_[1494]_  & (~\new_[684]_  | ~\new_[6713]_ );
  assign n1204 = ~\new_[1465]_  & ~\new_[6424]_ ;
  assign \new_[1417]_  = ~\new_[4943]_  & (~\new_[1503]_  | ~\new_[5223]_ );
  assign \new_[1418]_  = ~\new_[4941]_  & (~\new_[1504]_  | ~\new_[5223]_ );
  assign \new_[1419]_  = ~\new_[4944]_  & (~\new_[5223]_  | ~\new_[1505]_ );
  assign \new_[1420]_  = ~\new_[4954]_  & (~\new_[5223]_  | ~\new_[1506]_ );
  assign \new_[1421]_  = ~\new_[4946]_  & (~\new_[1507]_  | ~\new_[5223]_ );
  assign \new_[1422]_  = ~\new_[4948]_  & (~\new_[1508]_  | ~\new_[5223]_ );
  assign \new_[1423]_  = ~\new_[4945]_  & (~\new_[1511]_  | ~\new_[5223]_ );
  assign \new_[1424]_  = ~\new_[4940]_  & (~\new_[1512]_  | ~\new_[5223]_ );
  assign \new_[1425]_  = ~\new_[4955]_  & (~\new_[1515]_  | ~\new_[5223]_ );
  assign \new_[1426]_  = ~\new_[4947]_  & (~\new_[1516]_  | ~\new_[5223]_ );
  assign \new_[1427]_  = ~\new_[4942]_  & (~\new_[1517]_  | ~\new_[5223]_ );
  assign \new_[1428]_  = ~\new_[1500]_  & (~\new_[1293]_  | ~\new_[6338]_ );
  assign \new_[1429]_  = (~\new_[1565]_  | ~\new_[6714]_ ) & (~\new_[1294]_  | ~\new_[1690]_ );
  assign \new_[1430]_  = (~\new_[1567]_  | ~\new_[6099]_ ) & (~\new_[1292]_  | ~\new_[6258]_ );
  assign \new_[1431]_  = ~\new_[1501]_  & (~\new_[1255]_  | ~\new_[6338]_ );
  assign n1224 = ~\new_[1529]_  & ~\new_[6402]_ ;
  assign \new_[1433]_  = ~\new_[1532]_  & ~\new_[5909]_ ;
  assign \new_[1434]_  = (~\new_[1573]_  | ~\new_[6055]_ ) & (~\new_[5654]_  | ~\new_[2127]_ );
  assign \new_[1435]_  = (~\new_[1570]_  | ~\new_[6055]_ ) & (~\new_[5625]_  | ~\new_[2127]_ );
  assign \new_[1436]_  = (~\new_[1572]_  | ~\new_[6055]_ ) & (~\new_[5622]_  | ~\new_[2127]_ );
  assign \new_[1437]_  = ~\new_[5909]_  & (~\new_[1575]_  | ~\new_[2152]_ );
  assign \new_[1438]_  = \new_[1583]_  ? \new_[6257]_  : \new_[3180]_ ;
  assign \new_[1439]_  = \new_[1584]_  ? \new_[6257]_  : \new_[2969]_ ;
  assign \new_[1440]_  = (~\new_[3817]_  & ~\new_[2211]_ ) | (~\new_[2127]_  & ~\new_[1576]_ );
  assign \new_[1441]_  = \new_[1829]_  ? \new_[6695]_  : \new_[1876]_ ;
  assign \new_[1442]_  = ~\new_[1629]_  | ~\new_[3104]_  | ~\new_[2907]_  | ~\new_[2916]_ ;
  assign \new_[1443]_  = ~\new_[1630]_  | ~\new_[3099]_  | ~\new_[2902]_  | ~\new_[2913]_ ;
  assign \new_[1444]_  = ~\new_[1631]_  | ~\new_[3103]_  | ~\new_[2906]_  | ~\new_[2911]_ ;
  assign \new_[1445]_  = ~\new_[1632]_  | ~\new_[3101]_  | ~\new_[2904]_  | ~\new_[2914]_ ;
  assign \new_[1446]_  = ~\new_[1472]_ ;
  assign \new_[1447]_  = ~\new_[3126]_  | ~\new_[1538]_ ;
  assign \new_[1448]_  = \new_[1830]_  ? \new_[7492]_  : \new_[1877]_ ;
  assign \new_[1449]_  = \new_[1555]_  ? \new_[6257]_  : \new_[3419]_ ;
  assign \new_[1450]_  = \new_[1552]_  ? \new_[6257]_  : \new_[3840]_ ;
  assign \new_[1451]_  = \new_[6245]_  | \new_[1547]_ ;
  assign \new_[1452]_  = (~\new_[1636]_  | ~\new_[1585]_ ) & (~\new_[3662]_  | ~\new_[1770]_ );
  assign \new_[1453]_  = \\i_tv80_core_TmpAddr_reg[11] ;
  assign halt_n = ~i_tv80_core_Halt_FF_reg;
  assign \new_[1455]_  = ~\new_[1484]_ ;
  assign \new_[1456]_  = ~\new_[1485]_ ;
  assign \new_[1457]_  = ~\new_[1486]_ ;
  assign \new_[1458]_  = ~\new_[1487]_ ;
  assign \new_[1459]_  = ~\new_[1488]_ ;
  assign \new_[1460]_  = ~\new_[1489]_ ;
  assign \new_[1461]_  = ~\new_[1490]_ ;
  assign \new_[1462]_  = ~\new_[1491]_ ;
  assign \new_[1463]_  = ~\new_[1546]_  & (~\new_[2471]_  | ~\new_[6257]_ );
  assign n1229 = ~\new_[1566]_  & ~\new_[6424]_ ;
  assign \new_[1465]_  = (~\new_[1609]_  | ~\new_[6129]_ ) & (~\new_[1308]_  | ~\new_[6438]_ );
  assign \new_[1466]_  = ~\new_[3354]_  | (~\new_[1611]_  & ~\new_[5813]_ );
  assign \new_[1467]_  = \new_[1603]_  ? \new_[2373]_  : \new_[5916]_ ;
  assign \new_[1468]_  = (~\new_[1613]_  | ~busak_n) & (~\new_[6580]_  | ~\new_[6258]_ );
  assign \new_[1469]_  = ~\new_[5909]_  & (~\new_[2156]_  | ~\new_[1617]_ );
  assign \new_[1470]_  = \new_[1601]_  ? \new_[6257]_  : \new_[2787]_ ;
  assign \new_[1471]_  = (~\new_[4186]_  | ~\new_[2313]_ ) & (~\new_[2674]_  | ~\new_[1618]_ );
  assign \new_[1472]_  = \new_[1634]_  & \new_[1574]_ ;
  assign \new_[1473]_  = ~\new_[1699]_  | ~\new_[7492]_ ;
  assign \new_[1474]_  = ~\new_[1577]_  | ~\new_[7493]_ ;
  assign n1234 = ~\new_[1541]_ ;
  assign \new_[1476]_  = \new_[1600]_  ? \new_[6257]_  : \new_[2977]_ ;
  assign \new_[1477]_  = \new_[1595]_  ? \new_[6257]_  : \new_[3623]_ ;
  assign \new_[1478]_  = ~\new_[1542]_ ;
  assign \new_[1479]_  = ~\new_[1544]_ ;
  assign \new_[1480]_  = (~\new_[1633]_  | ~\new_[7501]_ ) & (~\new_[3945]_  | ~\new_[7505]_ );
  assign \new_[1481]_  = ~\\i_tv80_core_Read_To_Reg_r_reg[4] ;
  assign \new_[1482]_  = ~\new_[1594]_  | ~\new_[1596]_ ;
  assign \new_[1483]_  = ~\new_[1547]_ ;
  assign \new_[1484]_  = ~\new_[1586]_  & (~\new_[1637]_  | ~\do[0] );
  assign \new_[1485]_  = ~\new_[1593]_  & (~\new_[1637]_  | ~\do[1] );
  assign \new_[1486]_  = ~\new_[1592]_  & (~\new_[1637]_  | ~\do[2] );
  assign \new_[1487]_  = ~\new_[1591]_  & (~\new_[1637]_  | ~\do[3] );
  assign \new_[1488]_  = ~\new_[1590]_  & (~\new_[1637]_  | ~\do[4] );
  assign \new_[1489]_  = ~\new_[1587]_  & (~\new_[1637]_  | ~\do[5] );
  assign \new_[1490]_  = ~\new_[1589]_  & (~\new_[1637]_  | ~\do[6] );
  assign \new_[1491]_  = ~\new_[1588]_  & (~\new_[1637]_  | ~\do[7] );
  assign \new_[1492]_  = ~\new_[1703]_  & ~\new_[1554]_ ;
  assign \new_[1493]_  = ~\new_[1563]_  | ~\new_[4864]_ ;
  assign \new_[1494]_  = ~\new_[6938]_  & ~\new_[3663]_ ;
  assign \new_[1495]_  = ~\new_[2266]_  | (~\new_[1615]_  & ~\new_[5813]_ );
  assign \new_[1496]_  = \new_[3840]_  ? \new_[6243]_  : \new_[1604]_ ;
  assign \new_[1497]_  = ~\new_[1552]_ ;
  assign \new_[1498]_  = ~\new_[1555]_ ;
  assign \new_[1499]_  = \new_[3623]_  ? \new_[6243]_  : \new_[1652]_ ;
  assign \new_[1500]_  = ~\new_[1606]_  & ~\new_[1690]_ ;
  assign \new_[1501]_  = ~\new_[1607]_  & ~\new_[6299]_ ;
  assign \new_[1502]_  = ~\new_[2271]_  | ~\new_[2192]_  | ~\new_[2290]_  | ~\new_[1655]_ ;
  assign \new_[1503]_  = ~\new_[2272]_  | ~\new_[2193]_  | ~\new_[1656]_  | ~\new_[2303]_ ;
  assign \new_[1504]_  = ~\new_[2273]_  | ~\new_[2194]_  | ~\new_[1657]_  | ~\new_[2291]_ ;
  assign \new_[1505]_  = ~\new_[2274]_  | ~\new_[2195]_  | ~\new_[1658]_  | ~\new_[2292]_ ;
  assign \new_[1506]_  = ~\new_[2275]_  | ~\new_[2196]_  | ~\new_[1659]_  | ~\new_[2293]_ ;
  assign \new_[1507]_  = ~\new_[2276]_  | ~\new_[2197]_  | ~\new_[2294]_  | ~\new_[1660]_ ;
  assign \new_[1508]_  = ~\new_[2277]_  | ~\new_[2198]_  | ~\new_[2295]_  | ~\new_[1661]_ ;
  assign \new_[1509]_  = ~\new_[2278]_  | ~\new_[2199]_  | ~\new_[1662]_  | ~\new_[2304]_ ;
  assign \new_[1510]_  = ~\new_[2279]_  | ~\new_[2200]_  | ~\new_[1663]_  | ~\new_[2296]_ ;
  assign \new_[1511]_  = ~\new_[2280]_  | ~\new_[2201]_  | ~\new_[1664]_  | ~\new_[2297]_ ;
  assign \new_[1512]_  = ~\new_[2281]_  | ~\new_[2202]_  | ~\new_[1665]_  | ~\new_[2298]_ ;
  assign \new_[1513]_  = ~\new_[2282]_  | ~\new_[2203]_  | ~\new_[1666]_  | ~\new_[2299]_ ;
  assign \new_[1514]_  = ~\new_[2283]_  | ~\new_[2204]_  | ~\new_[1667]_  | ~\new_[2300]_ ;
  assign \new_[1515]_  = ~\new_[2284]_  | ~\new_[2205]_  | ~\new_[2301]_  | ~\new_[1668]_ ;
  assign \new_[1516]_  = ~\new_[2285]_  | ~\new_[2206]_  | ~\new_[2302]_  | ~\new_[1669]_ ;
  assign \new_[1517]_  = ~\new_[2286]_  | ~\new_[2207]_  | ~\new_[1670]_  | ~\new_[2305]_ ;
  assign \new_[1518]_  = ~\new_[2239]_  | (~\new_[1671]_  & ~\new_[6712]_ );
  assign \new_[1519]_  = ~\new_[2122]_  | (~\new_[1672]_  & ~\new_[6712]_ );
  assign \new_[1520]_  = ~\new_[3110]_  | (~\new_[1673]_  & ~\new_[6712]_ );
  assign \new_[1521]_  = ~\new_[3014]_  | (~\new_[1674]_  & ~\new_[3288]_ );
  assign \new_[1522]_  = ~\new_[2817]_  | (~\new_[1675]_  & ~\new_[3288]_ );
  assign \new_[1523]_  = ~\new_[2892]_  | (~\new_[1676]_  & ~\new_[3287]_ );
  assign \new_[1524]_  = ~\new_[2428]_  | (~\new_[1677]_  & ~\new_[3287]_ );
  assign \new_[1525]_  = ~\new_[2743]_  | (~\new_[1678]_  & ~\new_[3287]_ );
  assign \new_[1526]_  = ~\new_[2632]_  | (~\new_[1679]_  & ~\new_[3234]_ );
  assign \new_[1527]_  = ~\new_[2621]_  | (~\new_[1680]_  & ~\new_[3287]_ );
  assign \new_[1528]_  = ~\new_[2240]_  | (~\new_[1681]_  & ~\new_[3287]_ );
  assign \new_[1529]_  = (~\new_[1682]_  | ~\new_[6129]_ ) & (~\new_[1379]_  | ~\new_[1690]_ );
  assign \new_[1530]_  = ~\new_[2813]_  | (~\new_[1683]_  & ~\new_[5813]_ );
  assign n1239 = ~\new_[1612]_  & ~\new_[6424]_ ;
  assign \new_[1532]_  = (~\new_[1685]_  | ~\new_[5979]_ ) & (~\new_[2313]_  | ~\new_[6523]_ );
  assign \new_[1533]_  = ~\new_[1745]_  | ~\new_[3098]_  | ~\new_[2901]_  | ~\new_[2910]_ ;
  assign \new_[1534]_  = ~\new_[1746]_  | ~\new_[3102]_  | ~\new_[2905]_  | ~\new_[2915]_ ;
  assign \new_[1535]_  = ~\new_[5909]_  & (~\new_[2153]_  | ~\new_[1686]_ );
  assign \new_[1536]_  = ~\new_[5909]_  & (~\new_[2154]_  | ~\new_[1687]_ );
  assign \new_[1537]_  = ~\new_[5909]_  & (~\new_[2155]_  | ~\new_[1688]_ );
  assign \new_[1538]_  = ~\new_[1625]_  | ~\new_[7482]_ ;
  assign n1244 = ~\new_[5270]_  | (~\new_[1695]_  & ~\new_[6441]_ );
  assign \new_[1540]_  = ~\new_[3186]_  | ~\new_[1619]_ ;
  assign \new_[1541]_  = (~\new_[1696]_  | ~\new_[6481]_ ) & (~\new_[1413]_  | ~\new_[6406]_ );
  assign \new_[1542]_  = ~\new_[1626]_  | ~\new_[7568]_ ;
  assign \new_[1543]_  = ~\new_[7524]_ ;
  assign \new_[1544]_  = ~\new_[1627]_  | ~\new_[7523]_ ;
  assign \new_[1545]_  = \\i_tv80_core_TmpAddr_reg[9] ;
  assign \new_[1546]_  = ~\new_[1602]_  & ~\new_[6257]_ ;
  assign \new_[1547]_  = \new_[1637]_  ? \new_[1623]_  : \new_[5572]_ ;
  assign \new_[1548]_  = (~\new_[2755]_  | ~\new_[1126]_ ) & (~\new_[1642]_  | ~\new_[3196]_ );
  assign \new_[1549]_  = (~\new_[2755]_  | ~\new_[6478]_ ) & (~\new_[1643]_  | ~\new_[3196]_ );
  assign \new_[1550]_  = ~\new_[1583]_ ;
  assign \new_[1551]_  = ~\new_[1584]_ ;
  assign \new_[1552]_  = (~\new_[2045]_  | ~\new_[5183]_ ) & (~\new_[1719]_  | ~\new_[4865]_ );
  assign \new_[1553]_  = ~\new_[1595]_ ;
  assign \new_[1554]_  = ~\new_[1596]_ ;
  assign \new_[1555]_  = (~\new_[2041]_  | ~\new_[5183]_ ) & (~\new_[1720]_  | ~\new_[4865]_ );
  assign \new_[1556]_  = ~\new_[1599]_ ;
  assign \new_[1557]_  = ~\new_[1600]_ ;
  assign \new_[1558]_  = ~\new_[1601]_ ;
  assign \new_[1559]_  = ~\new_[1602]_ ;
  assign \new_[1560]_  = ~\new_[1648]_  | (~\new_[6243]_  & ~\new_[3180]_ );
  assign \new_[1561]_  = ~\new_[1649]_  | (~\new_[2969]_  & ~\new_[6243]_ );
  assign \new_[1562]_  = \new_[2787]_  ? \new_[6243]_  : \new_[1718]_ ;
  assign \new_[1563]_  = \new_[4549]_  ? \new_[4042]_  : \new_[1722]_ ;
  assign \new_[1564]_  = ~\new_[1604]_ ;
  assign \new_[1565]_  = ~\new_[2267]_  | (~\new_[1726]_  & ~\new_[6712]_ );
  assign \new_[1566]_  = (~\new_[1728]_  | ~\new_[6132]_ ) & (~\new_[1394]_  | ~\new_[6225]_ );
  assign \new_[1567]_  = ~\new_[2080]_  | (~\new_[1727]_  & ~\new_[3287]_ );
  assign \new_[1568]_  = ~\new_[2884]_  | (~\new_[1730]_  & ~\new_[5813]_ );
  assign \new_[1569]_  = ~\new_[1611]_ ;
  assign \new_[1570]_  = ~\new_[2127]_  & (~\new_[1735]_  | ~\new_[5671]_ );
  assign \new_[1571]_  = ~\new_[1615]_ ;
  assign \new_[1572]_  = ~\new_[2127]_  & (~\new_[1737]_  | ~\new_[5677]_ );
  assign \new_[1573]_  = ~\new_[2127]_  & (~\new_[5691]_  | ~\new_[1736]_ );
  assign \new_[1574]_  = ~\new_[1873]_  | ~\new_[1817]_  | ~\new_[1740]_ ;
  assign \new_[1575]_  = ~\new_[1651]_  | ~\new_[2211]_ ;
  assign \new_[1576]_  = ~\new_[1694]_  | ~\new_[5979]_ ;
  assign \new_[1577]_  = ~\new_[1743]_  | ~\new_[1701]_ ;
  assign \new_[1578]_  = \\i_tv80_core_TmpAddr_reg[6] ;
  assign \new_[1579]_  = ~\\i_tv80_core_Read_To_Reg_r_reg[2] ;
  assign \new_[1580]_  = ~\\i_tv80_core_RegBusA_r_reg[0] ;
  assign \new_[1581]_  = ~\\i_tv80_core_RegBusA_r_reg[13] ;
  assign n1249 = ~\new_[1628]_ ;
  assign \new_[1583]_  = (~\new_[2043]_  | ~\new_[5183]_ ) & (~\new_[1716]_  | ~\new_[4865]_ );
  assign \new_[1584]_  = (~\new_[2044]_  | ~\new_[5183]_ ) & (~\new_[1717]_  | ~\new_[6047]_ );
  assign \new_[1585]_  = i_tv80_core_Auto_Wait_t2_reg;
  assign \new_[1586]_  = ~\new_[4574]_  & ~\new_[1637]_ ;
  assign \new_[1587]_  = ~\new_[4578]_  & ~\new_[1637]_ ;
  assign \new_[1588]_  = ~\new_[4580]_  & ~\new_[1637]_ ;
  assign \new_[1589]_  = ~\new_[4579]_  & ~\new_[1637]_ ;
  assign \new_[1590]_  = ~\new_[4577]_  & ~\new_[1637]_ ;
  assign \new_[1591]_  = ~\new_[4576]_  & ~\new_[1637]_ ;
  assign \new_[1592]_  = ~\new_[4575]_  & ~\new_[1637]_ ;
  assign \new_[1593]_  = ~\new_[4581]_  & ~\new_[1637]_ ;
  assign \new_[1594]_  = ~\new_[1640]_  | ~\new_[1836]_ ;
  assign \new_[1595]_  = (~\new_[2082]_  | ~\new_[5183]_ ) & (~\new_[1773]_  | ~\new_[4865]_ );
  assign \new_[1596]_  = ~\new_[7375]_  & ~\new_[1714]_ ;
  assign \new_[1597]_  = ~\new_[7534]_ ;
  assign \new_[1598]_  = ~\new_[1714]_  & ~\new_[1836]_ ;
  assign \new_[1599]_  = ~\new_[6686]_  | ~\new_[1715]_ ;
  assign \new_[1600]_  = (~\new_[2062]_  | ~\new_[5183]_ ) & (~\new_[1774]_  | ~\new_[6047]_ );
  assign \new_[1601]_  = (~\new_[2060]_  | ~\new_[5183]_ ) & (~\new_[1775]_  | ~\new_[6047]_ );
  assign \new_[1602]_  = (~\new_[2061]_  | ~\new_[5183]_ ) & (~\new_[1776]_  | ~\new_[6047]_ );
  assign \new_[1603]_  = ~\new_[1721]_  & (~\new_[3405]_  | ~\new_[4506]_ );
  assign \new_[1604]_  = (~\new_[1804]_  | ~\new_[4413]_ ) & (~\new_[2001]_  | ~\new_[4339]_ );
  assign \new_[1605]_  = ~\new_[1652]_ ;
  assign \new_[1606]_  = \new_[1780]_  ? \new_[6712]_  : \new_[3391]_ ;
  assign \new_[1607]_  = \new_[1781]_  ? \new_[6712]_  : \new_[2132]_ ;
  assign n1254 = ~\new_[1729]_  & ~\new_[6382]_ ;
  assign \new_[1609]_  = ~\new_[1724]_  | (~\new_[2047]_  & ~\new_[6047]_ );
  assign \new_[1610]_  = \\i_tv80_core_TmpAddr_reg[8] ;
  assign \new_[1611]_  = ~\new_[1725]_  & (~\new_[848]_  | ~\new_[3619]_ );
  assign \new_[1612]_  = (~\new_[1805]_  | ~busak_n) & (~\new_[1453]_  | ~\new_[6258]_ );
  assign \new_[1613]_  = ~\new_[1732]_  | (~\new_[2052]_  & ~\new_[4865]_ );
  assign \new_[1614]_  = ~\new_[1683]_ ;
  assign \new_[1615]_  = ~\new_[1733]_  & (~\new_[845]_  | ~\new_[3617]_ );
  assign \new_[1616]_  = ~\new_[3037]_  | (~\new_[1806]_  & ~\new_[5813]_ );
  assign \new_[1617]_  = ~\new_[5979]_  | ~\new_[1734]_  | ~\new_[3555]_ ;
  assign \new_[1618]_  = ~\new_[5991]_  & (~\new_[1870]_  | ~\new_[1813]_ );
  assign \new_[1619]_  = ~\new_[1747]_  | ~\new_[7482]_ ;
  assign \new_[1620]_  = ~\\i_tv80_core_Read_To_Reg_r_reg[0] ;
  assign \new_[1621]_  = ~\\i_tv80_core_Read_To_Reg_r_reg[1] ;
  assign \new_[1622]_  = \\i_tv80_core_ALU_Op_r_reg[1] ;
  assign \new_[1623]_  = i_tv80_core_Save_ALU_r_reg;
  assign \new_[1624]_  = \\i_tv80_core_ALU_Op_r_reg[3] ;
  assign \new_[1625]_  = \new_[1831]_  ^ \new_[1819]_ ;
  assign \new_[1626]_  = ~\new_[7345]_  | ~\new_[1824]_ ;
  assign \new_[1627]_  = ~\new_[1748]_  | ~\new_[7520]_ ;
  assign \new_[1628]_  = (~\new_[1758]_  | ~\new_[6481]_ ) & (~\new_[6649]_  | ~\new_[6406]_ );
  assign \new_[1629]_  = (~\new_[2755]_  | ~\new_[6518]_ ) & (~\new_[1765]_  | ~\new_[3196]_ );
  assign \new_[1630]_  = (~\new_[2755]_  | ~\new_[6542]_ ) & (~\new_[1762]_  | ~\new_[3196]_ );
  assign \new_[1631]_  = (~\new_[2755]_  | ~\new_[1247]_ ) & (~\new_[1763]_  | ~\new_[3196]_ );
  assign \new_[1632]_  = (~\new_[2755]_  | ~\new_[1248]_ ) & (~\new_[1764]_  | ~\new_[3196]_ );
  assign \new_[1633]_  = ~\new_[1710]_  | ~\new_[3295]_ ;
  assign \new_[1634]_  = ~\new_[7348]_  & ~\new_[7566]_ ;
  assign \new_[1635]_  = ~\new_[1772]_  & (~\new_[1834]_  | ~\new_[1771]_ );
  assign \new_[1636]_  = \new_[3903]_  | \new_[1770]_ ;
  assign \new_[1637]_  = \new_[1770]_  | \new_[6401]_ ;
  assign n1279 = \new_[1770]_  & reset_n;
  assign \new_[1639]_  = ~\new_[1703]_ ;
  assign \new_[1640]_  = ~\new_[1834]_  | ~\new_[1771]_ ;
  assign \new_[1641]_  = ~\new_[1706]_ ;
  assign \new_[1642]_  = \new_[1837]_  ? \new_[3456]_  : \new_[2067]_ ;
  assign \new_[1643]_  = \new_[6693]_  ? \new_[3456]_  : \new_[1945]_ ;
  assign n1269 = \new_[1945]_  ? \new_[6347]_  : \new_[6595]_ ;
  assign n1274 = \new_[1837]_  ? \new_[1690]_  : \new_[6558]_ ;
  assign \new_[1646]_  = \\i_tv80_core_TmpAddr_reg[7] ;
  assign \new_[1647]_  = ~\\i_tv80_core_RegBusA_r_reg[11] ;
  assign \new_[1648]_  = ~\new_[6243]_  | ~\new_[1777]_ ;
  assign \new_[1649]_  = ~\new_[6243]_  | ~\new_[1778]_ ;
  assign \new_[1650]_  = ~\new_[1718]_ ;
  assign \new_[1651]_  = \new_[3401]_  ? \new_[1980]_  : \new_[6519]_ ;
  assign \new_[1652]_  = ~\new_[2182]_  | (~\new_[1840]_  & ~\new_[4080]_ );
  assign \new_[1653]_  = \new_[3026]_  ? \new_[6243]_  : \new_[1843]_ ;
  assign n1259 = ~\new_[1786]_  & ~\new_[6426]_ ;
  assign \new_[1655]_  = ~\new_[1788]_  | ~\new_[2384]_ ;
  assign \new_[1656]_  = ~\new_[1789]_  | ~\new_[2384]_ ;
  assign \new_[1657]_  = ~\new_[1790]_  | ~\new_[2383]_ ;
  assign \new_[1658]_  = ~\new_[1791]_  | ~\new_[2383]_ ;
  assign \new_[1659]_  = ~\new_[1792]_  | ~\new_[2383]_ ;
  assign \new_[1660]_  = ~\new_[1793]_  | ~\new_[2383]_ ;
  assign \new_[1661]_  = ~\new_[1794]_  | ~\new_[2383]_ ;
  assign \new_[1662]_  = ~\new_[1795]_  | ~\new_[2383]_ ;
  assign \new_[1663]_  = ~\new_[1796]_  | ~\new_[2383]_ ;
  assign \new_[1664]_  = ~\new_[1797]_  | ~\new_[2384]_ ;
  assign \new_[1665]_  = ~\new_[1798]_  | ~\new_[2384]_ ;
  assign \new_[1666]_  = ~\new_[1799]_  | ~\new_[2383]_ ;
  assign \new_[1667]_  = ~\new_[1800]_  | ~\new_[2383]_ ;
  assign \new_[1668]_  = ~\new_[1801]_  | ~\new_[2384]_ ;
  assign \new_[1669]_  = ~\new_[1802]_  | ~\new_[2383]_ ;
  assign \new_[1670]_  = ~\new_[1803]_  | ~\new_[2384]_ ;
  assign \new_[1671]_  = \new_[1848]_  ? \new_[5724]_  : \new_[2104]_ ;
  assign \new_[1672]_  = \new_[1849]_  ? \new_[5724]_  : \new_[2105]_ ;
  assign \new_[1673]_  = \new_[1851]_  ? \new_[5724]_  : \new_[2112]_ ;
  assign \new_[1674]_  = \new_[1852]_  ? \new_[5724]_  : \new_[2113]_ ;
  assign \new_[1675]_  = \new_[1853]_  ? \new_[5724]_  : \new_[2107]_ ;
  assign \new_[1676]_  = \new_[1854]_  ? \new_[5724]_  : \new_[2108]_ ;
  assign \new_[1677]_  = \new_[1855]_  ? \new_[5724]_  : \new_[2114]_ ;
  assign \new_[1678]_  = \new_[1856]_  ? \new_[5724]_  : \new_[2115]_ ;
  assign \new_[1679]_  = \new_[1857]_  ? \new_[5724]_  : \new_[2109]_ ;
  assign \new_[1680]_  = \new_[1858]_  ? \new_[5724]_  : \new_[2110]_ ;
  assign \new_[1681]_  = \new_[1859]_  ? \new_[5724]_  : \new_[2111]_ ;
  assign \new_[1682]_  = ~\new_[1784]_  | (~\new_[2089]_  & ~\new_[4866]_ );
  assign \new_[1683]_  = ~\new_[1785]_  & (~\new_[799]_  | ~\new_[3619]_ );
  assign \new_[1684]_  = ~\new_[1730]_ ;
  assign \new_[1685]_  = ~\new_[1807]_  & ~\new_[2129]_ ;
  assign \new_[1686]_  = ~\new_[1814]_  | ~\new_[2211]_ ;
  assign \new_[1687]_  = ~\new_[1815]_  | ~\new_[2211]_ ;
  assign \new_[1688]_  = ~\new_[1816]_  | ~\new_[2211]_ ;
  assign \new_[1689]_  = \\i_tv80_core_TmpAddr_reg[5] ;
  assign \new_[1690]_  = i_tv80_core_BusAck_reg;
  assign \new_[1691]_  = ~\\i_tv80_core_RegBusA_r_reg[10] ;
  assign \new_[1692]_  = ~\\i_tv80_core_RegBusA_r_reg[12] ;
  assign \new_[1693]_  = ~\\i_tv80_core_RegBusA_r_reg[14] ;
  assign \new_[1694]_  = ~\new_[1812]_  | (~\new_[3817]_  & ~\new_[1914]_ );
  assign \new_[1695]_  = ~\new_[1818]_  & (~\new_[5382]_  | ~\new_[5588]_ );
  assign \new_[1696]_  = ~\new_[1744]_ ;
  assign \new_[1697]_  = ~\new_[7566]_  & ~\new_[7264]_ ;
  assign \new_[1698]_  = ~\new_[7495]_  & ~\new_[7519]_ ;
  assign \new_[1699]_  = ~\new_[7495]_  & ~\new_[1753]_ ;
  assign \new_[1700]_  = ~\new_[1748]_ ;
  assign \new_[1701]_  = ~\new_[1749]_ ;
  assign n1264 = ~\new_[1751]_ ;
  assign \new_[1703]_  = ~\new_[6686]_  | ~\new_[1834]_ ;
  assign \new_[1704]_  = ~\new_[7264]_ ;
  assign \new_[1705]_  = ~\new_[1754]_ ;
  assign \new_[1706]_  = \new_[7314]_  & \new_[7393]_ ;
  assign \new_[1707]_  = ~\new_[1755]_ ;
  assign \new_[1708]_  = ~\new_[1885]_  | ~\new_[7101]_ ;
  assign \new_[1709]_  = ~\new_[1756]_ ;
  assign \new_[1710]_  = (~\new_[1999]_  | ~\new_[7482]_ ) & (~\new_[6595]_  | ~\new_[5295]_ );
  assign n1304 = ~\new_[1759]_ ;
  assign n1309 = ~\new_[1760]_ ;
  assign n1299 = ~\new_[1761]_ ;
  assign \new_[1714]_  = ~\new_[7535]_ ;
  assign \new_[1715]_  = ~\new_[1771]_ ;
  assign \new_[1716]_  = ~\new_[5486]_  & (~\new_[4359]_  | ~\new_[1896]_ );
  assign \new_[1717]_  = ~\new_[5486]_  & (~\new_[4362]_  | ~\new_[1897]_ );
  assign \new_[1718]_  = ~\new_[1838]_  & (~\new_[2086]_  | ~\new_[6541]_ );
  assign \new_[1719]_  = ~\new_[5486]_  & (~\new_[4357]_  | ~\new_[1899]_ );
  assign \new_[1720]_  = ~\new_[5486]_  & (~\new_[4358]_  | ~\new_[1900]_ );
  assign \new_[1721]_  = ~\new_[4506]_  & (~\new_[3063]_  | ~\new_[1895]_ );
  assign \new_[1722]_  = ~\new_[1779]_ ;
  assign n1284 = ~\new_[1844]_  & ~\new_[6623]_ ;
  assign \new_[1724]_  = ~\new_[1846]_  | ~\new_[4864]_ ;
  assign \new_[1725]_  = ~\new_[7218]_  & ~\new_[3620]_ ;
  assign \new_[1726]_  = \new_[1907]_  ? \new_[5724]_  : \new_[2157]_ ;
  assign \new_[1727]_  = \new_[1910]_  ? \new_[5724]_  : \new_[2158]_ ;
  assign \new_[1728]_  = ~\new_[1841]_  | (~\new_[2139]_  & ~\new_[4865]_ );
  assign \new_[1729]_  = (~\new_[1905]_  | ~\new_[6129]_ ) & (~\new_[1545]_  | ~\new_[6438]_ );
  assign \new_[1730]_  = ~\new_[1842]_  & (~\new_[849]_  | ~\new_[3617]_ );
  assign \new_[1731]_  = ~\new_[3421]_  | (~\new_[1902]_  & ~\new_[5813]_ );
  assign \new_[1732]_  = ~\new_[1867]_  | ~\new_[6047]_ ;
  assign \new_[1733]_  = ~\new_[6921]_  & ~\new_[3620]_ ;
  assign \new_[1734]_  = ~\new_[2127]_  & (~\new_[3720]_  | ~\new_[1914]_ );
  assign \new_[1735]_  = ~\new_[1868]_  & (~\new_[6431]_  | ~\new_[4748]_ );
  assign \new_[1736]_  = (~\new_[1979]_  | ~\new_[5681]_ ) & (~\new_[1915]_  | ~\new_[4862]_ );
  assign \new_[1737]_  = ~\new_[1869]_  & (~\new_[6209]_  | ~\new_[4748]_ );
  assign \new_[1738]_  = ~\new_[1806]_ ;
  assign \new_[1739]_  = ~\\i_tv80_core_Read_To_Reg_r_reg[3] ;
  assign \new_[1740]_  = ~\new_[7285]_  | ~\new_[7353]_ ;
  assign \new_[1741]_  = ~\new_[1874]_  | ~\new_[7496]_ ;
  assign \new_[1742]_  = ~\new_[1872]_  | ~\new_[1827]_ ;
  assign \new_[1743]_  = ~\new_[1872]_  | ~\new_[1827]_ ;
  assign \new_[1744]_  = ~\new_[1871]_  & (~\new_[3181]_  | ~\new_[1413]_ );
  assign \new_[1745]_  = (~\new_[2755]_  | ~\new_[6515]_ ) & (~\new_[1879]_  | ~\new_[3196]_ );
  assign \new_[1746]_  = (~\new_[2755]_  | ~\new_[1324]_ ) & (~\new_[1880]_  | ~\new_[3196]_ );
  assign \new_[1747]_  = \new_[1945]_  ^ \new_[1878]_ ;
  assign \new_[1748]_  = ~\new_[1826]_  | ~\new_[7101]_ ;
  assign \new_[1749]_  = ~\new_[1828]_  | ~\new_[7374]_ ;
  assign n1289 = ~\new_[1821]_ ;
  assign \new_[1751]_  = (~\new_[1889]_  | ~reset_n) & (~\new_[6622]_  | ~\new_[6406]_ );
  assign n1294 = ~\new_[1822]_ ;
  assign \new_[1753]_  = ~\new_[7493]_ ;
  assign \new_[1754]_  = ~\new_[1932]_  | ~\new_[7075]_ ;
  assign \new_[1755]_  = ~\new_[7099]_  | ~\new_[7091]_ ;
  assign \new_[1756]_  = ~\new_[1991]_  | ~\new_[6688]_ ;
  assign \new_[1757]_  = \new_[7373]_  & \new_[1989]_ ;
  assign \new_[1758]_  = ~\new_[2035]_  | (~\new_[1940]_  & ~\new_[6347]_ );
  assign \new_[1759]_  = (~\new_[1937]_  | ~\new_[3183]_ ) & (~\new_[1623]_  | ~\new_[6406]_ );
  assign \new_[1760]_  = (~\new_[1938]_  | ~\new_[3183]_ ) & (~\new_[1624]_  | ~\new_[6406]_ );
  assign \new_[1761]_  = (~\new_[1941]_  | ~\new_[3183]_ ) & (~\new_[6429]_  | ~\new_[6406]_ );
  assign \new_[1762]_  = \new_[6690]_  ? \new_[3456]_  : \new_[6680]_ ;
  assign \new_[1763]_  = \new_[1943]_  ? \new_[3456]_  : \new_[2119]_ ;
  assign \new_[1764]_  = \new_[1944]_  ? \new_[3456]_  : \new_[7085]_ ;
  assign \new_[1765]_  = \new_[1942]_  ? \new_[3456]_  : \new_[6694]_ ;
  assign n1334 = \new_[1942]_  ? \new_[1690]_  : \new_[6643]_ ;
  assign n1319 = \new_[6690]_  ? \new_[1690]_  : \new_[6656]_ ;
  assign n1339 = \new_[1943]_  ? \new_[1690]_  : \new_[6551]_ ;
  assign n1344 = \new_[1944]_  ? \new_[1690]_  : \new_[6671]_ ;
  assign \new_[1770]_  = i_tv80_core_Auto_Wait_t1_reg;
  assign \new_[1771]_  = ~\new_[1835]_ ;
  assign \new_[1772]_  = ~\new_[1836]_ ;
  assign \new_[1773]_  = ~\new_[5486]_  & (~\new_[1948]_  | ~\new_[4361]_ );
  assign \new_[1774]_  = ~\new_[5486]_  & (~\new_[1949]_  | ~\new_[4360]_ );
  assign \new_[1775]_  = ~\new_[5486]_  & (~\new_[1950]_  | ~\new_[4363]_ );
  assign \new_[1776]_  = ~\new_[5486]_  & (~\new_[1951]_  | ~\new_[4364]_ );
  assign \new_[1777]_  = \new_[1952]_  ? \new_[4804]_  : \new_[3622]_ ;
  assign \new_[1778]_  = \new_[1953]_  ? \new_[4804]_  : \new_[4124]_ ;
  assign \new_[1779]_  = ~\new_[1898]_  & (~\new_[1104]_  | ~\new_[3619]_ );
  assign \new_[1780]_  = \new_[1957]_  ? \new_[6271]_  : \new_[2183]_ ;
  assign \new_[1781]_  = \new_[1958]_  ? \new_[6271]_  : \new_[2184]_ ;
  assign n1324 = ~\new_[1903]_  & ~\new_[6327]_ ;
  assign n1314 = ~\new_[1904]_  & ~\new_[6327]_ ;
  assign \new_[1784]_  = ~\new_[1911]_  | ~\new_[6047]_ ;
  assign \new_[1785]_  = ~\new_[1906]_  & ~\new_[3619]_ ;
  assign \new_[1786]_  = (~\new_[1961]_  | ~\new_[6129]_ ) & (~\new_[1578]_  | ~\new_[6165]_ );
  assign \new_[1787]_  = ~\\i_tv80_core_RegBusA_r_reg[15] ;
  assign \new_[1788]_  = \new_[1962]_  ? \new_[6466]_  : \new_[5833]_ ;
  assign \new_[1789]_  = \new_[1963]_  ? \new_[6466]_  : \new_[7223]_ ;
  assign \new_[1790]_  = \new_[1964]_  ? \new_[7115]_  : \new_[7339]_ ;
  assign \new_[1791]_  = \new_[1965]_  ? \new_[7115]_  : \new_[5835]_ ;
  assign \new_[1792]_  = \new_[1966]_  ? \new_[7115]_  : \new_[7188]_ ;
  assign \new_[1793]_  = \new_[1967]_  ? \new_[6466]_  : \new_[6940]_ ;
  assign \new_[1794]_  = \new_[1968]_  ? \new_[7115]_  : \new_[6926]_ ;
  assign \new_[1795]_  = \new_[1969]_  ? \new_[7115]_  : \new_[5841]_ ;
  assign \new_[1796]_  = \new_[1970]_  ? \new_[7115]_  : \new_[5837]_ ;
  assign \new_[1797]_  = \new_[1971]_  ? \new_[7115]_  : \new_[5822]_ ;
  assign \new_[1798]_  = \new_[1972]_  ? \new_[6466]_  : \new_[5832]_ ;
  assign \new_[1799]_  = \new_[1973]_  ? \new_[7115]_  : \new_[5839]_ ;
  assign \new_[1800]_  = \new_[1974]_  ? \new_[7115]_  : \new_[5834]_ ;
  assign \new_[1801]_  = \new_[1975]_  ? \new_[6466]_  : \new_[5838]_ ;
  assign \new_[1802]_  = \new_[1976]_  ? \new_[6466]_  : \new_[5836]_ ;
  assign \new_[1803]_  = \new_[1977]_  ? \new_[6466]_  : \new_[5840]_ ;
  assign \new_[1804]_  = ~\new_[1901]_  | (~\new_[2935]_  & ~\new_[3586]_ );
  assign \new_[1805]_  = ~\new_[1912]_  | (~\new_[2159]_  & ~\new_[6047]_ );
  assign \new_[1806]_  = ~\new_[1913]_  & (~\new_[852]_  | ~\new_[3617]_ );
  assign \new_[1807]_  = (~\new_[3280]_  | ~\new_[1916]_ ) & (~\new_[1980]_  | ~\new_[6523]_ );
  assign \new_[1808]_  = ~\\i_tv80_core_RegBusA_r_reg[7] ;
  assign \new_[1809]_  = ~\\i_tv80_core_RegBusA_r_reg[9] ;
  assign \new_[1810]_  = \\i_tv80_core_ALU_Op_r_reg[2] ;
  assign \new_[1811]_  = \\i_tv80_core_ALU_Op_r_reg[0] ;
  assign \new_[1812]_  = ~\new_[3534]_  | ~\new_[1914]_ ;
  assign \new_[1813]_  = ~\new_[4186]_  | ~\new_[1914]_  | ~\new_[3592]_ ;
  assign \new_[1814]_  = \new_[6442]_  ? \new_[1916]_  : \new_[6663]_ ;
  assign \new_[1815]_  = \new_[6452]_  ? \new_[1916]_  : \new_[6667]_ ;
  assign \new_[1816]_  = \new_[6504]_  ? \new_[1916]_  : \new_[6674]_ ;
  assign \new_[1817]_  = ~\new_[7353]_  | ~\new_[1875]_  | ~\new_[2032]_ ;
  assign \new_[1818]_  = ~\new_[5672]_  & (~\new_[1994]_  | ~\new_[1933]_ );
  assign \new_[1819]_  = ~\new_[1872]_ ;
  assign \new_[1820]_  = ~\new_[1874]_ ;
  assign \new_[1821]_  = (~\new_[1935]_  | ~\new_[6427]_ ) & (~\new_[6634]_  | ~\new_[6406]_ );
  assign \new_[1822]_  = (~\new_[1936]_  | ~\new_[6481]_ ) & (~\new_[6570]_  | ~\new_[6406]_ );
  assign n1329 = ~\new_[1888]_  | (~\new_[6356]_  & ~\new_[5847]_ );
  assign \new_[1824]_  = ~\new_[7102]_  & ~\new_[1927]_ ;
  assign \new_[1825]_  = ~\new_[6688]_  | ~\new_[2033]_ ;
  assign \new_[1826]_  = ~\new_[1931]_  | ~\new_[1986]_ ;
  assign \new_[1827]_  = ~\new_[1988]_  & ~\new_[1930]_ ;
  assign \new_[1828]_  = ~\new_[1928]_  | ~\new_[1989]_ ;
  assign \new_[1829]_  = ~\new_[1876]_ ;
  assign \new_[1830]_  = ~\new_[1877]_ ;
  assign \new_[1831]_  = ~\new_[7142]_  | ~\new_[1929]_ ;
  assign n1349 = ~\new_[1934]_  | (~\new_[1739]_  & ~\new_[6356]_ );
  assign \new_[1833]_  = ~\new_[1884]_ ;
  assign \new_[1834]_  = \new_[7536]_ ;
  assign \new_[1835]_  = ~\new_[6691]_  | ~\new_[3926]_ ;
  assign \new_[1836]_  = ~\new_[3854]_  | ~\new_[1943]_ ;
  assign \new_[1837]_  = ~\new_[1894]_ ;
  assign \new_[1838]_  = ~\new_[1926]_  & ~\new_[2373]_ ;
  assign \new_[1839]_  = (~\new_[2831]_  | ~\new_[6236]_ ) & (~\new_[2012]_  | ~\new_[5849]_ );
  assign \new_[1840]_  = ~\new_[1954]_  | (~\new_[4404]_  & ~\new_[4339]_ );
  assign \new_[1841]_  = ~\new_[1959]_  | ~\new_[4864]_ ;
  assign \new_[1842]_  = ~\new_[7183]_  & ~\new_[3620]_ ;
  assign \new_[1843]_  = \new_[1956]_  & \new_[2182]_ ;
  assign \new_[1844]_  = (~\new_[2015]_  | ~busak_n) & (~\new_[1610]_  | ~\new_[1690]_ );
  assign \new_[1845]_  = ~\new_[3746]_  | (~\new_[2013]_  & ~\new_[5813]_ );
  assign \new_[1846]_  = \new_[4557]_  ? \new_[4042]_  : \new_[2014]_ ;
  assign \new_[1847]_  = ~\new_[1902]_ ;
  assign \new_[1848]_  = ~\new_[2854]_  & (~\new_[2018]_  | ~\new_[4316]_ );
  assign \new_[1849]_  = ~\new_[2760]_  & (~\new_[2019]_  | ~\new_[4316]_ );
  assign \new_[1850]_  = ~\new_[2811]_  & (~\new_[2020]_  | ~\new_[4316]_ );
  assign \new_[1851]_  = ~\new_[3583]_  & (~\new_[2021]_  | ~\new_[4316]_ );
  assign \new_[1852]_  = ~\new_[3446]_  & (~\new_[2022]_  | ~\new_[4316]_ );
  assign \new_[1853]_  = ~\new_[3208]_  & (~\new_[2023]_  | ~\new_[4316]_ );
  assign \new_[1854]_  = ~\new_[3297]_  & (~\new_[2024]_  | ~\new_[4316]_ );
  assign \new_[1855]_  = ~\new_[2972]_  & (~\new_[2025]_  | ~\new_[4316]_ );
  assign \new_[1856]_  = ~\new_[3148]_  & (~\new_[2026]_  | ~\new_[4316]_ );
  assign \new_[1857]_  = ~\new_[3056]_  & (~\new_[2027]_  | ~\new_[4316]_ );
  assign \new_[1858]_  = ~\new_[3049]_  & (~\new_[2028]_  | ~\new_[4316]_ );
  assign \new_[1859]_  = ~\new_[2857]_  & (~\new_[2029]_  | ~\new_[4316]_ );
  assign \new_[1860]_  = ~\\i_tv80_core_RegBusA_r_reg[8] ;
  assign \new_[1861]_  = \\i_tv80_core_TmpAddr_reg[4] ;
  assign \new_[1862]_  = ~\\i_tv80_core_RegBusA_r_reg[1] ;
  assign \new_[1863]_  = ~\\i_tv80_core_RegBusA_r_reg[2] ;
  assign \new_[1864]_  = ~\\i_tv80_core_RegBusA_r_reg[5] ;
  assign \new_[1865]_  = ~\\i_tv80_core_RegBusA_r_reg[6] ;
  assign \new_[1866]_  = \\i_tv80_core_BusB_reg[0] ;
  assign \new_[1867]_  = \new_[4556]_  ? \new_[4042]_  : \new_[2017]_ ;
  assign \new_[1868]_  = ~\new_[3533]_  | ~\new_[1978]_ ;
  assign \new_[1869]_  = ~\new_[3536]_  | ~\new_[1978]_ ;
  assign \new_[1870]_  = ~\new_[4186]_  | ~\new_[1980]_ ;
  assign \new_[1871]_  = ~\new_[6334]_  & (~\new_[2036]_  | ~\new_[1992]_ );
  assign \new_[1872]_  = ~\new_[1917]_  | ~\new_[1987]_ ;
  assign \new_[1873]_  = ~\new_[7346]_ ;
  assign \new_[1874]_  = ~\new_[1918]_  | ~\new_[1990]_ ;
  assign \new_[1875]_  = ~\new_[1988]_  & ~\new_[1999]_ ;
  assign \new_[1876]_  = ~\new_[1990]_  | ~\new_[2031]_ ;
  assign \new_[1877]_  = ~\new_[7342]_  | ~\new_[7360]_ ;
  assign \new_[1878]_  = \new_[1987]_  & \new_[2032]_ ;
  assign \new_[1879]_  = \new_[7537]_  ? \new_[3456]_  : \new_[2065]_ ;
  assign \new_[1880]_  = \new_[2038]_  ? \new_[3456]_  : \new_[7103]_ ;
  assign n1359 = \new_[2038]_  ? \new_[1690]_  : \new_[6569]_ ;
  assign n1364 = \new_[7103]_  ? \new_[6252]_  : \new_[6596]_ ;
  assign n1369 = \new_[7537]_  ? \new_[6252]_  : \new_[6573]_ ;
  assign \new_[1884]_  = \new_[3705]_  ^ \new_[2038]_ ;
  assign \new_[1885]_  = ~\new_[1927]_ ;
  assign \new_[1886]_  = ~\new_[1932]_ ;
  assign \new_[1887]_  = ~\new_[1998]_  | ~\new_[3705]_ ;
  assign \new_[1888]_  = ~\new_[6055]_  | ~reset_n | ~\new_[1993]_  | ~\new_[5991]_ ;
  assign \new_[1889]_  = ~\new_[2035]_  | (~\new_[2127]_  & ~\new_[3303]_ );
  assign n1374 = ~\new_[6211]_  | (~\new_[2723]_  & ~\new_[2127]_ );
  assign n1379 = ~\new_[6136]_  | (~\new_[2658]_  & ~\new_[2127]_ );
  assign \new_[1892]_  = \\i_tv80_core_TmpAddr_reg[3] ;
  assign n1354 = ~\new_[1939]_ ;
  assign \new_[1894]_  = ~\new_[7525]_ ;
  assign \new_[1895]_  = ~\new_[1983]_  & ~\new_[3973]_ ;
  assign \new_[1896]_  = (~\new_[2043]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2553]_ );
  assign \new_[1897]_  = (~\new_[2044]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2552]_ );
  assign \new_[1898]_  = ~\new_[2000]_  & ~\new_[3618]_ ;
  assign \new_[1899]_  = (~\new_[2045]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2633]_ );
  assign \new_[1900]_  = (~\new_[2041]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2554]_ );
  assign \new_[1901]_  = ~\new_[2001]_  | ~\new_[3586]_ ;
  assign \new_[1902]_  = ~\new_[2009]_  & (~\new_[851]_  | ~\new_[3617]_ );
  assign \new_[1903]_  = (~\new_[2053]_  | ~busak_n) & (~\new_[1689]_  | ~\new_[6261]_ );
  assign \new_[1904]_  = (~\new_[2054]_  | ~\new_[6126]_ ) & (~\new_[1646]_  | ~\new_[6225]_ );
  assign \new_[1905]_  = ~\new_[2010]_  | (~\new_[2289]_  & ~\new_[6047]_ );
  assign \new_[1906]_  = ~\new_[2011]_  & (~\new_[5835]_  | ~\new_[7335]_ );
  assign \new_[1907]_  = ~\new_[2798]_  & (~\new_[2055]_  | ~\new_[4316]_ );
  assign \new_[1908]_  = ~\\i_tv80_core_RegBusA_r_reg[4] ;
  assign \new_[1909]_  = ~\\i_tv80_core_RegBusA_r_reg[3] ;
  assign \new_[1910]_  = (~\new_[2056]_  | ~\new_[4316]_ ) & (~\new_[2671]_  | ~\new_[4292]_ );
  assign \new_[1911]_  = \new_[4558]_  ? \new_[4042]_  : \new_[2051]_ ;
  assign \new_[1912]_  = ~\new_[2030]_  | ~\new_[6047]_ ;
  assign \new_[1913]_  = ~\new_[7333]_  & ~\new_[3620]_ ;
  assign \new_[1914]_  = ~\new_[1980]_ ;
  assign \new_[1915]_  = ~\new_[1982]_  & (~\new_[3650]_  | ~\new_[6442]_ );
  assign \new_[1916]_  = ~\new_[1982]_ ;
  assign \new_[1917]_  = ~\new_[2032]_  | ~\new_[2040]_ ;
  assign \new_[1918]_  = ~\new_[7343]_  | ~\new_[2031]_ ;
  assign \new_[1919]_  = \new_[2471]_  ? \new_[6243]_  : \new_[2081]_ ;
  assign n1394 = \new_[2065]_  ? \new_[1690]_  : \new_[6576]_ ;
  assign n1399 = \new_[6694]_  ? \new_[1690]_  : \new_[6552]_ ;
  assign n1404 = \new_[2067]_  ? \new_[6252]_  : \new_[6658]_ ;
  assign n1409 = \new_[6605]_  ? \new_[6388]_  : \new_[7085]_ ;
  assign n1384 = \new_[6560]_  ? \new_[6162]_  : \new_[6693]_ ;
  assign \new_[1925]_  = \\i_tv80_core_TmpAddr_reg[2] ;
  assign \new_[1926]_  = (~\new_[2078]_  | ~\new_[4413]_ ) & (~\new_[3473]_  | ~\new_[4339]_ );
  assign \new_[1927]_  = ~\new_[1986]_ ;
  assign \new_[1928]_  = ~\new_[7142]_ ;
  assign \new_[1929]_  = ~\new_[1988]_ ;
  assign \new_[1930]_  = ~\new_[1989]_ ;
  assign \new_[1931]_  = ~\new_[1991]_ ;
  assign \new_[1932]_  = ~\new_[3926]_  | ~\new_[7537]_ ;
  assign \new_[1933]_  = ~\new_[2037]_  | ~\new_[6055]_ ;
  assign \new_[1934]_  = ~\new_[4041]_  | ~\new_[6342]_  | ~\new_[2674]_  | ~\new_[3655]_ ;
  assign \new_[1935]_  = ~\new_[2035]_  | (~\new_[3315]_  & ~\new_[2127]_ );
  assign \new_[1936]_  = ~\new_[2035]_  | (~\new_[2127]_  & ~\new_[3361]_ );
  assign \new_[1937]_  = ~\new_[2127]_  & (~\new_[3465]_  | ~\new_[3653]_ );
  assign \new_[1938]_  = ~\new_[2127]_  & (~\new_[3329]_  | ~\new_[4201]_ );
  assign \new_[1939]_  = ~\new_[6427]_  | ~\new_[2127]_  | ~\new_[3546]_ ;
  assign \new_[1940]_  = ~\new_[1995]_ ;
  assign \new_[1941]_  = ~\new_[2127]_  & (~\new_[3211]_  | ~\new_[2864]_ );
  assign \new_[1942]_  = ~\new_[1996]_ ;
  assign \new_[1943]_  = ~\new_[1997]_ ;
  assign \new_[1944]_  = ~\new_[1998]_ ;
  assign \new_[1945]_  = ~\new_[1999]_ ;
  assign n1414 = \new_[6528]_  ? \new_[6162]_  : \new_[2076]_ ;
  assign \new_[1947]_  = (~\new_[3020]_  | ~\new_[6236]_ ) & (~\new_[2087]_  | ~\new_[5849]_ );
  assign \new_[1948]_  = (~\new_[2082]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2661]_ );
  assign \new_[1949]_  = (~\new_[2062]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2555]_ );
  assign \new_[1950]_  = (~\new_[2060]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[2551]_ );
  assign \new_[1951]_  = (~\new_[2061]_  | ~\new_[5103]_ ) & (~\new_[4626]_  | ~\new_[3285]_ );
  assign \new_[1952]_  = \new_[2079]_  ? \new_[4413]_  : \new_[3503]_ ;
  assign \new_[1953]_  = \new_[2077]_  ? \new_[4413]_  : \new_[3117]_ ;
  assign \new_[1954]_  = (~\new_[2083]_  | ~\new_[3601]_ ) & (~\new_[3556]_  | ~\new_[4339]_ );
  assign n1389 = ~\new_[2048]_  & ~\new_[6426]_ ;
  assign \new_[1956]_  = ~\new_[2046]_  | ~\new_[3353]_ ;
  assign \new_[1957]_  = ~\new_[3924]_  & (~\new_[2095]_  | ~\new_[4316]_ );
  assign \new_[1958]_  = ~\new_[2636]_  & (~\new_[2096]_  | ~\new_[4316]_ );
  assign \new_[1959]_  = \new_[4559]_  ? \new_[4042]_  : \new_[2090]_ ;
  assign \new_[1960]_  = ~\new_[2013]_ ;
  assign \new_[1961]_  = ~\new_[2050]_  | (~\new_[2379]_  & ~\new_[6047]_ );
  assign \new_[1962]_  = \new_[1293]_  ? \new_[2058]_  : \new_[2429]_ ;
  assign \new_[1963]_  = \new_[1294]_  ? \new_[2058]_  : \new_[1308]_ ;
  assign \new_[1964]_  = \new_[1233]_  ? \new_[2057]_  : \new_[1453]_ ;
  assign \new_[1965]_  = \new_[1234]_  ? \new_[2057]_  : \new_[1379]_ ;
  assign \new_[1966]_  = \new_[1235]_  ? \new_[2057]_  : \new_[1394]_ ;
  assign \new_[1967]_  = \new_[1292]_  ? \new_[2059]_  : \new_[1104]_ ;
  assign \new_[1968]_  = \new_[1255]_  ? \new_[2059]_  : \new_[6580]_ ;
  assign \new_[1969]_  = \new_[1236]_  ? \new_[2059]_  : \new_[2034]_ ;
  assign \new_[1970]_  = \new_[1237]_  ? \new_[2059]_  : \new_[1925]_ ;
  assign \new_[1971]_  = \new_[1238]_  ? \new_[2057]_  : \new_[1892]_ ;
  assign \new_[1972]_  = \new_[1239]_  ? \new_[2058]_  : \new_[1861]_ ;
  assign \new_[1973]_  = \new_[1240]_  ? \new_[2059]_  : \new_[1689]_ ;
  assign \new_[1974]_  = \new_[1241]_  ? \new_[2059]_  : \new_[1578]_ ;
  assign \new_[1975]_  = \new_[1225]_  ? \new_[2059]_  : \new_[1646]_ ;
  assign \new_[1976]_  = \new_[1242]_  ? \new_[2059]_  : \new_[1610]_ ;
  assign \new_[1977]_  = \new_[1223]_  ? \new_[2058]_  : \new_[1545]_ ;
  assign \new_[1978]_  = \new_[2059]_  | \new_[5991]_ ;
  assign \new_[1979]_  = \new_[5125]_  & \new_[2059]_ ;
  assign \new_[1980]_  = ~\new_[4996]_  | ~\new_[2059]_ ;
  assign \new_[1981]_  = (~\new_[2471]_  | ~\new_[6236]_ ) & (~\new_[2088]_  | ~\new_[5849]_ );
  assign \new_[1982]_  = ~\new_[2059]_ ;
  assign \new_[1983]_  = ~\new_[4489]_  | (~\new_[2133]_  & ~\new_[1624]_ );
  assign n1429 = \new_[6624]_  ? \new_[6388]_  : \new_[6680]_ ;
  assign n1424 = \new_[2119]_  ? \new_[6252]_  : \new_[6678]_ ;
  assign \new_[1986]_  = ~\new_[7096]_  | ~\new_[4001]_ ;
  assign \new_[1987]_  = ~\new_[7141]_ ;
  assign \new_[1988]_  = ~\new_[7140]_ ;
  assign \new_[1989]_  = ~\new_[7356]_ ;
  assign \new_[1990]_  = ~\new_[2033]_ ;
  assign \new_[1991]_  = ~\new_[7077]_  | ~\new_[7085]_ ;
  assign \new_[1992]_  = ~\new_[3402]_  | ~\new_[2063]_ ;
  assign \new_[1993]_  = ~\new_[2127]_  & ~\new_[5672]_ ;
  assign \new_[1994]_  = ~\new_[6055]_  | ~\new_[2127]_  | ~\new_[5588]_ ;
  assign \new_[1995]_  = ~\new_[2127]_  & (~\new_[3439]_  | ~\new_[3654]_ );
  assign \new_[1996]_  = ~\new_[2162]_  & ~\new_[2068]_ ;
  assign \new_[1997]_  = ~\new_[2125]_  & ~\new_[6973]_ ;
  assign \new_[1998]_  = ~\new_[7453]_  & ~\new_[2126]_ ;
  assign \new_[1999]_  = ~\new_[2040]_ ;
  assign \new_[2000]_  = (~\new_[4704]_  | ~\new_[1104]_ ) & (~\new_[2136]_  | ~\new_[5304]_ );
  assign \new_[2001]_  = \new_[2140]_  ? \new_[6713]_  : \new_[6520]_ ;
  assign \new_[2002]_  = \\i_tv80_core_BusB_reg[6] ;
  assign \new_[2003]_  = \\i_tv80_core_BusB_reg[4] ;
  assign \new_[2004]_  = \\i_tv80_core_BusB_reg[1] ;
  assign \new_[2005]_  = \\i_tv80_core_BusB_reg[3] ;
  assign \new_[2006]_  = \\i_tv80_core_BusB_reg[5] ;
  assign \new_[2007]_  = \\i_tv80_core_BusB_reg[2] ;
  assign n1419 = ~\new_[2091]_  & ~\new_[6370]_ ;
  assign \new_[2009]_  = ~\new_[2093]_  & ~\new_[3620]_ ;
  assign \new_[2010]_  = ~\new_[2097]_  | ~\new_[6047]_ ;
  assign \new_[2011]_  = ~\new_[7335]_  & ~\new_[2094]_ ;
  assign \new_[2012]_  = ~\new_[3501]_  | (~\new_[2102]_  & ~\new_[3619]_ );
  assign \new_[2013]_  = ~\new_[2084]_  & (~\new_[853]_  | ~\new_[3617]_ );
  assign \new_[2014]_  = ~\new_[2047]_ ;
  assign \new_[2015]_  = ~\new_[2085]_  | (~\new_[2441]_  & ~\new_[4866]_ );
  assign \new_[2016]_  = \\i_tv80_core_BusB_reg[7] ;
  assign \new_[2017]_  = ~\new_[2052]_ ;
  assign \new_[2018]_  = (~\new_[2104]_  | ~\new_[3318]_ ) & (~\new_[2968]_  | ~\new_[3395]_ );
  assign \new_[2019]_  = (~\new_[2105]_  | ~\new_[3318]_ ) & (~\new_[2850]_  | ~\new_[3395]_ );
  assign \new_[2020]_  = (~\new_[2106]_  | ~\new_[3318]_ ) & (~\new_[2908]_  | ~\new_[3395]_ );
  assign \new_[2021]_  = (~\new_[2112]_  | ~\new_[3318]_ ) & (~\new_[3395]_  | ~\new_[3694]_ );
  assign \new_[2022]_  = (~\new_[2113]_  | ~\new_[3318]_ ) & (~\new_[3580]_  | ~\new_[3395]_ );
  assign \new_[2023]_  = (~\new_[2107]_  | ~\new_[3318]_ ) & (~\new_[3319]_  | ~\new_[3395]_ );
  assign \new_[2024]_  = (~\new_[2108]_  | ~\new_[3318]_ ) & (~\new_[3442]_  | ~\new_[3395]_ );
  assign \new_[2025]_  = (~\new_[2114]_  | ~\new_[3318]_ ) & (~\new_[3057]_  | ~\new_[3395]_ );
  assign \new_[2026]_  = (~\new_[2115]_  | ~\new_[3318]_ ) & (~\new_[3246]_  | ~\new_[3395]_ );
  assign \new_[2027]_  = (~\new_[2109]_  | ~\new_[3318]_ ) & (~\new_[3161]_  | ~\new_[3395]_ );
  assign \new_[2028]_  = (~\new_[2110]_  | ~\new_[3318]_ ) & (~\new_[3153]_  | ~\new_[3395]_ );
  assign \new_[2029]_  = (~\new_[2111]_  | ~\new_[3318]_ ) & (~\new_[2967]_  | ~\new_[3395]_ );
  assign \new_[2030]_  = \new_[4553]_  ? \new_[4042]_  : \new_[2116]_ ;
  assign \new_[2031]_  = ~\new_[7094]_  | ~\new_[2120]_ ;
  assign \new_[2032]_  = ~\new_[2117]_  | ~\new_[4002]_ ;
  assign \new_[2033]_  = ~\new_[7094]_  & ~\new_[2120]_ ;
  assign \new_[2034]_  = \\i_tv80_core_TmpAddr_reg[1] ;
  assign \new_[2035]_  = ~\new_[3543]_  | ~\new_[2674]_ ;
  assign \new_[2036]_  = ~\new_[6711]_  | ~\new_[2127]_  | ~\new_[1413]_ ;
  assign \new_[2037]_  = ~\new_[2127]_  & (~\new_[4997]_  | ~\new_[5605]_ );
  assign \new_[2038]_  = ~\new_[2329]_  | ~\new_[2328]_  | ~\new_[2388]_  | ~\new_[2166]_ ;
  assign \new_[2039]_  = ~\new_[2237]_  | ~\new_[2165]_  | ~\new_[2130]_ ;
  assign \new_[2040]_  = ~\new_[2131]_  | ~\new_[2123]_ ;
  assign \new_[2041]_  = \new_[2174]_  ? \new_[6713]_  : \new_[761]_ ;
  assign \new_[2042]_  = (~\new_[3026]_  | ~\new_[6236]_ ) & (~\new_[2147]_  | ~\new_[5849]_ );
  assign \new_[2043]_  = \new_[2171]_  ? \new_[6713]_  : \new_[758]_ ;
  assign \new_[2044]_  = \new_[2172]_  ? \new_[6712]_  : \new_[759]_ ;
  assign \new_[2045]_  = \new_[2173]_  ? \new_[6713]_  : \new_[736]_ ;
  assign \new_[2046]_  = ~\new_[2141]_  | ~\new_[3601]_ ;
  assign \new_[2047]_  = ~\new_[2138]_  & (~\new_[1308]_  | ~\new_[6713]_ );
  assign \new_[2048]_  = (~\new_[2148]_  | ~\new_[6126]_ ) & (~\new_[1861]_  | ~\new_[1690]_ );
  assign n1434 = ~\new_[2101]_  & ~\new_[6424]_ ;
  assign \new_[2050]_  = ~\new_[2103]_  | ~\new_[4864]_ ;
  assign \new_[2051]_  = ~\new_[2089]_ ;
  assign \new_[2052]_  = ~\new_[2144]_  & (~\new_[6580]_  | ~\new_[3620]_ );
  assign \new_[2053]_  = ~\new_[2098]_  | (~\new_[2675]_  & ~\new_[4865]_ );
  assign \new_[2054]_  = ~\new_[2099]_  | (~\new_[2572]_  & ~\new_[4865]_ );
  assign \new_[2055]_  = (~\new_[2157]_  | ~\new_[3318]_ ) & (~\new_[2891]_  | ~\new_[3395]_ );
  assign \new_[2056]_  = (~\new_[2158]_  | ~\new_[3318]_ ) & (~\new_[2564]_  | ~\new_[3395]_ );
  assign \new_[2057]_  = ~\new_[2100]_ ;
  assign \new_[2058]_  = ~\new_[2100]_ ;
  assign \new_[2059]_  = ~\new_[2100]_ ;
  assign \new_[2060]_  = \new_[2259]_  ? \new_[6712]_  : \new_[760]_ ;
  assign \new_[2061]_  = \new_[2260]_  ? \new_[6712]_  : \new_[753]_ ;
  assign \new_[2062]_  = \new_[2256]_  ? \new_[6712]_  : \new_[763]_ ;
  assign \new_[2063]_  = ~\new_[2127]_  & (~\new_[4920]_  | ~\new_[4342]_ );
  assign \new_[2064]_  = ~\new_[2389]_  | ~\new_[2385]_  | ~\new_[2325]_  | ~\new_[2324]_ ;
  assign \new_[2065]_  = ~\new_[2117]_ ;
  assign \new_[2066]_  = ~\new_[2163]_  | ~\new_[2226]_ ;
  assign \new_[2067]_  = ~\new_[2120]_ ;
  assign \new_[2068]_  = ~\new_[2405]_  | ~\new_[2481]_  | ~\new_[7441]_  | ~\new_[2238]_ ;
  assign n1464 = \new_[2007]_  ? \new_[6162]_  : \new_[2247]_ ;
  assign n1449 = \new_[6548]_  ? \new_[6162]_  : \new_[2252]_ ;
  assign n1454 = \new_[2005]_  ? \new_[6162]_  : \new_[2246]_ ;
  assign n1444 = \new_[2003]_  ? \new_[6162]_  : \new_[2248]_ ;
  assign n1459 = \new_[2006]_  ? \new_[6162]_  : \new_[2249]_ ;
  assign n1439 = \new_[2002]_  ? \new_[6162]_  : \new_[2250]_ ;
  assign n1469 = \new_[2016]_  ? \new_[6388]_  : \new_[2251]_ ;
  assign \new_[2076]_  = ~\new_[2357]_  | ~\new_[2640]_  | ~\new_[2532]_  | ~\new_[2533]_ ;
  assign \new_[2077]_  = \new_[2258]_  ? \new_[6713]_  : \new_[6591]_ ;
  assign \new_[2078]_  = ~\new_[4520]_  | ~\new_[3827]_  | ~\new_[2169]_  | ~\new_[3490]_ ;
  assign \new_[2079]_  = \new_[2257]_  ? \new_[6713]_  : \new_[6606]_ ;
  assign \new_[2080]_  = ~\new_[2168]_  | ~\new_[6712]_ ;
  assign \new_[2081]_  = \new_[2208]_  ? \new_[2373]_  : \new_[4556]_ ;
  assign \new_[2082]_  = \new_[2255]_  ? \new_[6713]_  : \new_[762]_ ;
  assign \new_[2083]_  = \new_[3261]_  ? \new_[5439]_  : \new_[2178]_ ;
  assign \new_[2084]_  = ~\new_[2150]_  & ~\new_[3620]_ ;
  assign \new_[2085]_  = ~\new_[2151]_  | ~\new_[6047]_ ;
  assign \new_[2086]_  = ~\new_[2146]_  & ~\new_[4554]_ ;
  assign \new_[2087]_  = ~\new_[3358]_  | (~\new_[2189]_  & ~\new_[3620]_ );
  assign \new_[2088]_  = ~\new_[3500]_  | (~\new_[2190]_  & ~\new_[3619]_ );
  assign \new_[2089]_  = ~\new_[2177]_  & (~\new_[1379]_  | ~\new_[3619]_ );
  assign \new_[2090]_  = ~\new_[2139]_ ;
  assign \new_[2091]_  = (~\new_[2188]_  | ~busak_n) & (~\new_[1892]_  | ~\new_[6438]_ );
  assign \new_[2092]_  = (~\new_[2186]_  | ~\new_[5849]_ ) & (~\new_[3230]_  | ~\new_[6236]_ );
  assign \new_[2093]_  = ~\new_[2176]_  & (~\new_[5840]_  | ~\new_[7335]_ );
  assign \new_[2094]_  = ~\new_[2175]_  & (~\new_[6723]_  | ~\new_[799]_ );
  assign \new_[2095]_  = (~\new_[2183]_  | ~\new_[3318]_ ) & (~\new_[3395]_  | ~\new_[4064]_ );
  assign \new_[2096]_  = (~\new_[2184]_  | ~\new_[3318]_ ) & (~\new_[2763]_  | ~\new_[3395]_ );
  assign \new_[2097]_  = \new_[4554]_  ? \new_[4042]_  : \new_[2185]_ ;
  assign \new_[2098]_  = ~\new_[2209]_  | ~\new_[6047]_ ;
  assign \new_[2099]_  = ~\new_[2210]_  | ~\new_[6047]_ ;
  assign \new_[2100]_  = ~\new_[2145]_ ;
  assign \new_[2101]_  = (~\new_[2318]_  | ~busak_n) & (~\new_[1925]_  | ~\new_[6225]_ );
  assign \new_[2102]_  = ~\new_[2181]_  & (~\new_[5834]_  | ~\new_[7335]_ );
  assign \new_[2103]_  = \new_[4549]_  ? \new_[3276]_  : \new_[2317]_ ;
  assign \new_[2104]_  = ~\new_[2216]_  & (~\new_[2729]_  | ~\new_[1233]_ );
  assign \new_[2105]_  = ~\new_[2217]_  & (~\new_[2729]_  | ~\new_[1234]_ );
  assign \new_[2106]_  = ~\new_[2218]_  & (~\new_[2729]_  | ~\new_[1235]_ );
  assign \new_[2107]_  = ~\new_[2219]_  & (~\new_[2569]_  | ~\new_[1238]_ );
  assign \new_[2108]_  = ~\new_[2220]_  & (~\new_[2729]_  | ~\new_[1239]_ );
  assign \new_[2109]_  = ~\new_[2221]_  & (~\new_[2569]_  | ~\new_[1225]_ );
  assign \new_[2110]_  = ~\new_[2222]_  & (~\new_[2729]_  | ~\new_[1242]_ );
  assign \new_[2111]_  = ~\new_[2223]_  & (~\new_[2729]_  | ~\new_[1223]_ );
  assign \new_[2112]_  = ~\new_[2212]_  & (~\new_[2569]_  | ~\new_[1236]_ );
  assign \new_[2113]_  = ~\new_[2213]_  & (~\new_[2729]_  | ~\new_[1237]_ );
  assign \new_[2114]_  = ~\new_[2214]_  & (~\new_[2569]_  | ~\new_[1240]_ );
  assign \new_[2115]_  = ~\new_[2215]_  & (~\new_[2729]_  | ~\new_[1241]_ );
  assign \new_[2116]_  = ~\new_[2159]_ ;
  assign \new_[2117]_  = ~\new_[2319]_  & ~\new_[2224]_ ;
  assign \new_[2118]_  = ~\new_[2320]_  & ~\new_[2227]_ ;
  assign \new_[2119]_  = ~\new_[7362]_ ;
  assign \new_[2120]_  = ~\new_[2229]_  & ~\new_[2228]_ ;
  assign \new_[2121]_  = ~\new_[2580]_  | ~\new_[7270]_  | ~\new_[2326]_  | ~\new_[2456]_ ;
  assign \new_[2122]_  = \new_[2232]_  | \new_[6711]_ ;
  assign \new_[2123]_  = ~\new_[2234]_  & ~\new_[2233]_ ;
  assign \new_[2124]_  = ~\new_[2161]_ ;
  assign \new_[2125]_  = ~\new_[2392]_  | ~\new_[2395]_  | ~\new_[2402]_  | ~\new_[2477]_ ;
  assign \new_[2126]_  = ~\new_[2393]_  | ~\new_[2394]_  | ~\new_[2404]_  | ~\new_[2480]_ ;
  assign \new_[2127]_  = ~\new_[2674]_ ;
  assign \new_[2128]_  = ~\new_[2674]_ ;
  assign \new_[2129]_  = ~\new_[2674]_ ;
  assign \new_[2130]_  = ~\new_[2235]_  & ~\new_[7483]_ ;
  assign \new_[2131]_  = ~\new_[2164]_ ;
  assign \new_[2132]_  = ~\new_[2244]_  & (~\new_[1255]_  | ~\new_[6271]_ );
  assign \new_[2133]_  = \new_[2265]_  ? \new_[3841]_  : \new_[6659]_ ;
  assign \new_[2134]_  = \\i_tv80_core_RegAddrC_reg[1] ;
  assign \new_[2135]_  = i_tv80_core_Z16_r_reg;
  assign \new_[2136]_  = \new_[3313]_  ^ \new_[2263]_ ;
  assign \new_[2137]_  = ~\new_[6723]_  & (~\new_[3428]_  | ~\new_[2287]_ );
  assign \new_[2138]_  = ~\new_[2179]_  & ~\new_[3663]_ ;
  assign \new_[2139]_  = ~\new_[2262]_  & (~\new_[1394]_  | ~\new_[3619]_ );
  assign \new_[2140]_  = \new_[3263]_  ? \new_[5439]_  : \new_[2288]_ ;
  assign \new_[2141]_  = \new_[3265]_  ? \new_[5439]_  : \new_[2309]_ ;
  assign n1474 = ~\new_[2187]_  & ~\new_[6424]_ ;
  assign \new_[2143]_  = ~\new_[6723]_  & (~\new_[3432]_  | ~\new_[2314]_ );
  assign \new_[2144]_  = ~\new_[2191]_  & ~\new_[3618]_ ;
  assign \new_[2145]_  = ~\new_[2270]_  | ~\new_[6428]_ ;
  assign \new_[2146]_  = ~\new_[6540]_  | ~\new_[6572]_  | ~\new_[6531]_  | ~\new_[2373]_ ;
  assign \new_[2147]_  = ~\new_[3499]_  | (~\new_[2381]_  & ~\new_[3620]_ );
  assign \new_[2148]_  = ~\new_[2269]_  | (~\new_[2792]_  & ~\new_[6047]_ );
  assign \new_[2149]_  = (~\new_[3502]_  | ~\new_[6236]_ ) & (~\new_[2378]_  | ~\new_[5849]_ );
  assign \new_[2150]_  = ~\new_[2268]_  & (~\new_[5836]_  | ~\new_[7335]_ );
  assign \new_[2151]_  = \new_[4560]_  ? \new_[4042]_  : \new_[2380]_ ;
  assign \new_[2152]_  = ~\new_[2313]_  | ~\new_[6519]_ ;
  assign \new_[2153]_  = ~\new_[2313]_  | ~\new_[6663]_ ;
  assign \new_[2154]_  = ~\new_[2313]_  | ~\new_[6667]_ ;
  assign \new_[2155]_  = ~\new_[2313]_  | ~\new_[6674]_ ;
  assign \new_[2156]_  = ~\new_[2313]_  | ~\new_[3555]_ ;
  assign \new_[2157]_  = ~\new_[2315]_  & (~\new_[2569]_  | ~\new_[1294]_ );
  assign \new_[2158]_  = ~\new_[2316]_  & (~\new_[2569]_  | ~\new_[1292]_ );
  assign \new_[2159]_  = ~\new_[2312]_  & (~\new_[1453]_  | ~\new_[3620]_ );
  assign \new_[2160]_  = ~\new_[2225]_ ;
  assign \new_[2161]_  = ~\new_[2462]_  | ~\new_[2463]_  | ~\new_[2400]_  | ~\new_[2472]_ ;
  assign \new_[2162]_  = ~\new_[2396]_  | ~\new_[2464]_  | ~\new_[2473]_  | ~\new_[2397]_ ;
  assign \new_[2163]_  = ~\new_[2227]_ ;
  assign \new_[2164]_  = ~\new_[2583]_  | ~\new_[2468]_  | ~\new_[2460]_  | ~\new_[2459]_ ;
  assign \new_[2165]_  = ~\new_[2330]_  & (~\new_[7442]_  | ~\new_[6612]_ );
  assign \new_[2166]_  = (~\new_[7457]_  | ~n329) & (~\new_[7442]_  | ~n324);
  assign iorq_n = iorq_n_reg;
  assign \new_[2168]_  = \new_[2362]_  ? \new_[5724]_  : \new_[1292]_ ;
  assign \new_[2169]_  = ~\new_[2308]_  & ~\new_[3973]_ ;
  assign \new_[2170]_  = ~\new_[4423]_  | ~\new_[2264]_ ;
  assign \new_[2171]_  = \new_[3254]_  ? \new_[5439]_  : \new_[2360]_ ;
  assign \new_[2172]_  = \new_[3257]_  ? \new_[5439]_  : \new_[2361]_ ;
  assign \new_[2173]_  = \new_[3267]_  ? \new_[5439]_  : \new_[2365]_ ;
  assign \new_[2174]_  = \new_[3268]_  ? \new_[5439]_  : \new_[2366]_ ;
  assign \new_[2175]_  = ~\new_[6723]_  & (~\new_[3430]_  | ~\new_[2374]_ );
  assign \new_[2176]_  = ~\new_[2310]_  & ~\new_[7335]_ ;
  assign \new_[2177]_  = ~\new_[2307]_  & ~\new_[3618]_ ;
  assign \new_[2178]_  = ~\new_[2372]_  | ~\new_[2363]_ ;
  assign \new_[2179]_  = (~\new_[4704]_  | ~\new_[1308]_ ) & (~\new_[2444]_  | ~\new_[5304]_ );
  assign n1479 = ~\new_[2377]_  | ~\new_[4588]_ ;
  assign \new_[2181]_  = ~\new_[2382]_  & ~\new_[7335]_ ;
  assign \new_[2182]_  = ~\new_[2373]_  & ~\new_[4804]_ ;
  assign \new_[2183]_  = ~\new_[2375]_  & (~\new_[2569]_  | ~\new_[1293]_ );
  assign \new_[2184]_  = ~\new_[2376]_  & (~\new_[2569]_  | ~\new_[1255]_ );
  assign \new_[2185]_  = ~\new_[2289]_ ;
  assign \new_[2186]_  = ~\new_[3357]_  | (~\new_[2453]_  & ~\new_[3619]_ );
  assign \new_[2187]_  = (~\new_[2450]_  | ~\new_[6126]_ ) & (~\new_[2034]_  | ~\new_[6239]_ );
  assign \new_[2188]_  = ~\new_[2371]_  | (~\new_[2837]_  & ~\new_[6047]_ );
  assign \new_[2189]_  = ~\new_[2369]_  & (~\new_[5839]_  | ~\new_[7335]_ );
  assign \new_[2190]_  = ~\new_[2370]_  & (~\new_[5838]_  | ~\new_[7335]_ );
  assign \new_[2191]_  = (~\new_[4704]_  | ~\new_[6580]_ ) & (~\new_[2455]_  | ~\new_[5304]_ );
  assign \new_[2192]_  = (~\new_[2449]_  | ~\new_[4560]_ ) & (~\new_[6689]_  | ~\new_[794]_ );
  assign \new_[2193]_  = (~\new_[2449]_  | ~\new_[761]_ ) & (~\new_[6689]_  | ~\new_[848]_ );
  assign \new_[2194]_  = (~\new_[2449]_  | ~\new_[758]_ ) & (~\new_[6689]_  | ~\new_[852]_ );
  assign \new_[2195]_  = (~\new_[2449]_  | ~\new_[763]_ ) & (~\new_[6689]_  | ~\new_[799]_ );
  assign \new_[2196]_  = (~\new_[2449]_  | ~\new_[759]_ ) & (~\new_[6689]_  | ~\new_[849]_ );
  assign \new_[2197]_  = (~\new_[2449]_  | ~\new_[760]_ ) & (~\new_[6689]_  | ~\new_[684]_ );
  assign \new_[2198]_  = (~\new_[2449]_  | ~\new_[753]_ ) & (~\new_[6689]_  | ~\new_[845]_ );
  assign \new_[2199]_  = (~\new_[2449]_  | ~\new_[4554]_ ) & (~\new_[6689]_  | ~\new_[742]_ );
  assign \new_[2200]_  = (~\new_[2449]_  | ~\new_[4557]_ ) & (~\new_[6689]_  | ~\new_[792]_ );
  assign \new_[2201]_  = (~\new_[2449]_  | ~\new_[4553]_ ) & (~\new_[6689]_  | ~\new_[793]_ );
  assign \new_[2202]_  = (~\new_[2449]_  | ~\new_[4558]_ ) & (~\new_[6689]_  | ~\new_[766]_ );
  assign \new_[2203]_  = (~\new_[2449]_  | ~\new_[4559]_ ) & (~\new_[6689]_  | ~\new_[764]_ );
  assign \new_[2204]_  = (~\new_[2449]_  | ~\new_[4549]_ ) & (~\new_[6689]_  | ~\new_[757]_ );
  assign \new_[2205]_  = (~\new_[2449]_  | ~\new_[4556]_ ) & (~\new_[6689]_  | ~\new_[755]_ );
  assign \new_[2206]_  = (~\new_[2449]_  | ~\new_[736]_ ) & (~\new_[6689]_  | ~\new_[853]_ );
  assign \new_[2207]_  = (~\new_[2449]_  | ~\new_[762]_ ) & (~\new_[6689]_  | ~\new_[851]_ );
  assign \new_[2208]_  = \new_[3548]_  ? \new_[4413]_  : \new_[2525]_ ;
  assign \new_[2209]_  = ~\new_[2368]_  | (~\new_[3276]_  & ~\new_[6572]_ );
  assign \new_[2210]_  = \new_[4556]_  ? \new_[3276]_  : \new_[2451]_ ;
  assign \new_[2211]_  = ~\new_[2313]_ ;
  assign \new_[2212]_  = ~\new_[2569]_  & (~\new_[3775]_  | ~\new_[3862]_ );
  assign \new_[2213]_  = ~\new_[2569]_  & (~\new_[3776]_  | ~\new_[3863]_ );
  assign \new_[2214]_  = ~\new_[2569]_  & (~\new_[3777]_  | ~\new_[3855]_ );
  assign \new_[2215]_  = ~\new_[2569]_  & (~\new_[3778]_  | ~\new_[3856]_ );
  assign \new_[2216]_  = ~\new_[2569]_  & (~\new_[3696]_  | ~\new_[3763]_ );
  assign \new_[2217]_  = ~\new_[2569]_  & (~\new_[3697]_  | ~\new_[3859]_ );
  assign \new_[2218]_  = ~\new_[2569]_  & (~\new_[3698]_  | ~\new_[3764]_ );
  assign \new_[2219]_  = ~\new_[2569]_  & (~\new_[3699]_  | ~\new_[3864]_ );
  assign \new_[2220]_  = ~\new_[2569]_  & (~\new_[3700]_  | ~\new_[3865]_ );
  assign \new_[2221]_  = ~\new_[2569]_  & (~\new_[3701]_  | ~\new_[3765]_ );
  assign \new_[2222]_  = ~\new_[2569]_  & (~\new_[3702]_  | ~\new_[3866]_ );
  assign \new_[2223]_  = ~\new_[2569]_  & (~\new_[3703]_  | ~\new_[3766]_ );
  assign \new_[2224]_  = ~\new_[2584]_  | ~\new_[2585]_  | ~\new_[2603]_  | ~\new_[2605]_ ;
  assign \new_[2225]_  = ~\new_[2587]_  | ~\new_[2606]_  | ~\new_[2461]_  | ~\new_[2586]_ ;
  assign \new_[2226]_  = ~\new_[2320]_ ;
  assign \new_[2227]_  = ~\new_[2683]_  | ~\new_[2607]_  | ~\new_[2593]_  | ~\new_[2687]_ ;
  assign \new_[2228]_  = ~\new_[2700]_  | ~\new_[2695]_  | ~\new_[2465]_  | ~\new_[2467]_ ;
  assign \new_[2229]_  = ~\new_[2595]_  | ~\new_[2602]_  | ~\new_[2609]_  | ~\new_[2594]_ ;
  assign \new_[2230]_  = ~\new_[2458]_  & ~\new_[2386]_ ;
  assign \new_[2231]_  = ~\new_[2387]_  & ~\new_[2457]_ ;
  assign \new_[2232]_  = ~\new_[2421]_  & (~\new_[1234]_  | ~\new_[5746]_ );
  assign \new_[2233]_  = ~\new_[2398]_  | ~\new_[2604]_ ;
  assign \new_[2234]_  = ~\new_[2469]_  | ~\new_[2399]_ ;
  assign \new_[2235]_  = ~\new_[2401]_  | ~\new_[2478]_ ;
  assign \new_[2236]_  = ~\new_[2403]_  | ~\new_[2479]_ ;
  assign \new_[2237]_  = \new_[2390]_  & \new_[2391]_ ;
  assign \new_[2238]_  = ~\new_[7457]_  | ~\new_[434]_ ;
  assign \new_[2239]_  = \new_[2425]_  | \new_[6711]_ ;
  assign \new_[2240]_  = \new_[2426]_  | \new_[6711]_ ;
  assign \new_[2241]_  = ~\new_[6611]_  | ~\new_[2622]_ ;
  assign \new_[2242]_  = ~\new_[6553]_  | ~\new_[2423]_ ;
  assign \new_[2243]_  = ~\new_[2623]_  | ~\new_[6630]_ ;
  assign \new_[2244]_  = ~\new_[2424]_  & ~\new_[5746]_ ;
  assign \new_[2245]_  = ~\new_[2422]_  | ~\new_[7277]_ ;
  assign \new_[2246]_  = ~\new_[2644]_  | ~\new_[2653]_  | ~\new_[2538]_  | ~\new_[2547]_ ;
  assign \new_[2247]_  = ~\new_[2643]_  | ~\new_[2638]_  | ~\new_[2536]_  | ~\new_[2531]_ ;
  assign \new_[2248]_  = ~\new_[2645]_  | ~\new_[2652]_  | ~\new_[2539]_  | ~\new_[2540]_ ;
  assign \new_[2249]_  = ~\new_[2646]_  | ~\new_[2647]_  | ~\new_[2541]_  | ~\new_[2542]_ ;
  assign \new_[2250]_  = ~\new_[2648]_  | ~\new_[2649]_  | ~\new_[2543]_  | ~\new_[2544]_ ;
  assign \new_[2251]_  = ~\new_[2650]_  | ~\new_[2651]_  | ~\new_[2545]_  | ~\new_[2546]_ ;
  assign \new_[2252]_  = ~\new_[2641]_  | ~\new_[2642]_  | ~\new_[2535]_  | ~\new_[2537]_ ;
  assign n1484 = ~\new_[6441]_  & (~\new_[6023]_  | ~\new_[2549]_ );
  assign \new_[2254]_  = \\i_tv80_core_RegAddrB_r_reg[2] ;
  assign \new_[2255]_  = \new_[3260]_  ? \new_[5439]_  : \new_[2432]_ ;
  assign \new_[2256]_  = \new_[3269]_  ? \new_[5439]_  : \new_[2433]_ ;
  assign \new_[2257]_  = \new_[3262]_  ? \new_[5439]_  : \new_[2436]_ ;
  assign \new_[2258]_  = \new_[3251]_  ? \new_[5439]_  : \new_[2437]_ ;
  assign \new_[2259]_  = \new_[3270]_  ? \new_[5439]_  : \new_[2434]_ ;
  assign \new_[2260]_  = \new_[3271]_  ? \new_[5439]_  : \new_[2435]_ ;
  assign \new_[2261]_  = ~\new_[6723]_  & (~\new_[3431]_  | ~\new_[2440]_ );
  assign \new_[2262]_  = ~\new_[2367]_  & ~\new_[3618]_ ;
  assign \new_[2263]_  = ~\new_[2563]_  | ~\new_[3527]_  | ~\new_[3095]_ ;
  assign \new_[2264]_  = ~\new_[3434]_  | ~\new_[2471]_ ;
  assign \new_[2265]_  = ~\new_[2931]_  & (~\new_[2630]_  | ~\new_[5687]_ );
  assign \new_[2266]_  = ~\new_[2471]_  | ~\new_[6163]_ ;
  assign \new_[2267]_  = ~\new_[2442]_  | ~\new_[6712]_ ;
  assign \new_[2268]_  = ~\new_[2443]_  & ~\new_[7335]_ ;
  assign \new_[2269]_  = ~\new_[2445]_  | ~\new_[6047]_ ;
  assign \new_[2270]_  = ~\new_[6889]_  | ~\new_[2568]_  | ~\new_[4279]_ ;
  assign \new_[2271]_  = ~\new_[6820]_  | ~\new_[5833]_ ;
  assign \new_[2272]_  = ~\new_[6820]_  | ~\new_[7223]_ ;
  assign \new_[2273]_  = ~\new_[6820]_  | ~\new_[7339]_ ;
  assign \new_[2274]_  = ~\new_[6820]_  | ~\new_[5835]_ ;
  assign \new_[2275]_  = ~\new_[6820]_  | ~\new_[7188]_ ;
  assign \new_[2276]_  = ~\new_[6820]_  | ~\new_[6940]_ ;
  assign \new_[2277]_  = ~\new_[6820]_  | ~\new_[6926]_ ;
  assign \new_[2278]_  = ~\new_[6820]_  | ~\new_[5841]_ ;
  assign \new_[2279]_  = ~\new_[6820]_  | ~\new_[5837]_ ;
  assign \new_[2280]_  = ~\new_[6820]_  | ~\new_[5822]_ ;
  assign \new_[2281]_  = ~\new_[6820]_  | ~\new_[5832]_ ;
  assign \new_[2282]_  = ~\new_[6820]_  | ~\new_[5839]_ ;
  assign \new_[2283]_  = ~\new_[6820]_  | ~\new_[5834]_ ;
  assign \new_[2284]_  = ~\new_[6820]_  | ~\new_[5838]_ ;
  assign \new_[2285]_  = ~\new_[6820]_  | ~\new_[5836]_ ;
  assign \new_[2286]_  = ~\new_[6820]_  | ~\new_[5840]_ ;
  assign \new_[2287]_  = ~\new_[2444]_  | ~\new_[3509]_ ;
  assign \new_[2288]_  = ~\new_[2364]_ ;
  assign \new_[2289]_  = ~\new_[2439]_  & (~\new_[1545]_  | ~\new_[6713]_ );
  assign \new_[2290]_  = (~\new_[2570]_  | ~\new_[4660]_ ) & (~\new_[6724]_  | ~\new_[1293]_ );
  assign \new_[2291]_  = (~\new_[2570]_  | ~\new_[4774]_ ) & (~\new_[6724]_  | ~\new_[1233]_ );
  assign \new_[2292]_  = (~\new_[2570]_  | ~\new_[4775]_ ) & (~\new_[6724]_  | ~\new_[1234]_ );
  assign \new_[2293]_  = (~\new_[2570]_  | ~\new_[4649]_ ) & (~\new_[6724]_  | ~\new_[1235]_ );
  assign \new_[2294]_  = (~\new_[2570]_  | ~\new_[4768]_ ) & (~\new_[6724]_  | ~\new_[1292]_ );
  assign \new_[2295]_  = (~\new_[2570]_  | ~\new_[4771]_ ) & (~\new_[6724]_  | ~\new_[1255]_ );
  assign \new_[2296]_  = (~\new_[2570]_  | ~\new_[4789]_ ) & (~\new_[6724]_  | ~\new_[1237]_ );
  assign \new_[2297]_  = (~\new_[2570]_  | ~\new_[4780]_ ) & (~\new_[6724]_  | ~\new_[1238]_ );
  assign \new_[2298]_  = (~\new_[2570]_  | ~\new_[4658]_ ) & (~\new_[6724]_  | ~\new_[1239]_ );
  assign \new_[2299]_  = (~\new_[2570]_  | ~\new_[4659]_ ) & (~\new_[6724]_  | ~\new_[1240]_ );
  assign \new_[2300]_  = (~\new_[2570]_  | ~\new_[4776]_ ) & (~\new_[6724]_  | ~\new_[1241]_ );
  assign \new_[2301]_  = (~\new_[2570]_  | ~\new_[4879]_ ) & (~\new_[6724]_  | ~\new_[1225]_ );
  assign \new_[2302]_  = (~\new_[2570]_  | ~\new_[4778]_ ) & (~\new_[6724]_  | ~\new_[1242]_ );
  assign \new_[2303]_  = (~\new_[2570]_  | ~\new_[4826]_ ) & (~\new_[6724]_  | ~\new_[1294]_ );
  assign \new_[2304]_  = (~\new_[2570]_  | ~\new_[4792]_ ) & (~\new_[6724]_  | ~\new_[1236]_ );
  assign \new_[2305]_  = (~\new_[2570]_  | ~\new_[4791]_ ) & (~\new_[6724]_  | ~\new_[1223]_ );
  assign \new_[2306]_  = (~\new_[2574]_  | ~\new_[5849]_ ) & (~\new_[3672]_  | ~\new_[6236]_ );
  assign \new_[2307]_  = (~\new_[4704]_  | ~\new_[1379]_ ) & (~\new_[2577]_  | ~\new_[5304]_ );
  assign \new_[2308]_  = ~\new_[4491]_  | (~\new_[2631]_  & ~\new_[1624]_ );
  assign \new_[2309]_  = \new_[4148]_  ? \new_[2569]_  : \new_[850]_ ;
  assign \new_[2310]_  = ~\new_[2438]_  & (~\new_[6723]_  | ~\new_[851]_ );
  assign \new_[2311]_  = ~\new_[6723]_  & (~\new_[3429]_  | ~\new_[2579]_ );
  assign \new_[2312]_  = ~\new_[2454]_  & ~\new_[3618]_ ;
  assign \new_[2313]_  = ~\new_[2674]_  | ~\new_[5979]_ ;
  assign \new_[2314]_  = ~\new_[2455]_  | ~\new_[3509]_ ;
  assign \new_[2315]_  = ~\new_[2569]_  & (~\new_[3757]_  | ~\new_[3858]_ );
  assign \new_[2316]_  = ~\new_[2569]_  & (~\new_[3758]_  | ~\new_[3860]_ );
  assign \new_[2317]_  = ~\new_[2379]_ ;
  assign \new_[2318]_  = ~\new_[2446]_  | (~\new_[2888]_  & ~\new_[4866]_ );
  assign \new_[2319]_  = ~\new_[2703]_  | ~\new_[2696]_  | ~\new_[2697]_  | ~\new_[2682]_ ;
  assign \new_[2320]_  = ~\new_[2698]_  | ~\new_[2588]_  | ~\new_[2589]_  | ~\new_[2684]_ ;
  assign \new_[2321]_  = ~\new_[2699]_  | ~\new_[2685]_  | ~\new_[2590]_  | ~\new_[2591]_ ;
  assign \new_[2322]_  = ~\new_[2686]_  | ~\new_[2688]_  | ~\new_[2592]_  | ~\new_[2608]_ ;
  assign \new_[2323]_  = ~\new_[2522]_  & (~\new_[1235]_  | ~\new_[5746]_ );
  assign \new_[2324]_  = ~\new_[2476]_  & (~\new_[2753]_  | ~\new_[580]_ );
  assign \new_[2325]_  = ~\new_[2470]_  & (~\new_[7443]_  | ~\new_[578]_ );
  assign \new_[2326]_  = ~\new_[2475]_  & (~\new_[2756]_  | ~\new_[6602]_ );
  assign \new_[2327]_  = ~\new_[2474]_  | ~\new_[2466]_ ;
  assign \new_[2328]_  = (~\new_[2709]_  | ~n319) & (~\new_[2628]_  | ~n334);
  assign \new_[2329]_  = (~\new_[2712]_  | ~n314) & (~\new_[2713]_  | ~n309);
  assign \new_[2330]_  = ~\new_[511]_  & ~\new_[6684]_ ;
  assign \new_[2331]_  = \new_[539]_  | \new_[2524]_ ;
  assign \new_[2332]_  = \new_[431]_  | \new_[2524]_ ;
  assign \new_[2333]_  = \new_[6583]_  | \new_[2524]_ ;
  assign \new_[2334]_  = \new_[6641]_  | \new_[2524]_ ;
  assign \new_[2335]_  = \new_[6556]_  | \new_[2524]_ ;
  assign \new_[2336]_  = \new_[6660]_  | \new_[2524]_ ;
  assign \new_[2337]_  = \new_[2524]_  | \new_[654]_ ;
  assign \new_[2338]_  = \new_[540]_  | \new_[2526]_ ;
  assign \new_[2339]_  = \new_[432]_  | \new_[2526]_ ;
  assign \new_[2340]_  = \new_[6639]_  | \new_[2526]_ ;
  assign \new_[2341]_  = \new_[6587]_  | \new_[2526]_ ;
  assign \new_[2342]_  = \new_[6657]_  | \new_[2526]_ ;
  assign \new_[2343]_  = \new_[6599]_  | \new_[2526]_ ;
  assign \new_[2344]_  = ~\new_[2524]_  & ~\new_[777]_ ;
  assign \new_[2345]_  = ~\new_[2524]_  & ~\new_[788]_ ;
  assign \new_[2346]_  = ~\new_[2524]_  & ~\new_[770]_ ;
  assign \new_[2347]_  = \new_[2524]_  | \new_[534]_ ;
  assign \new_[2348]_  = \new_[2524]_  | \new_[570]_ ;
  assign \new_[2349]_  = ~\new_[2526]_  & ~\new_[737]_ ;
  assign \new_[2350]_  = \new_[2526]_  | \new_[535]_ ;
  assign \new_[2351]_  = \new_[2526]_  | \new_[571]_ ;
  assign \new_[2352]_  = \new_[2526]_  | \new_[646]_ ;
  assign \new_[2353]_  = \new_[2526]_  | \new_[655]_ ;
  assign \new_[2354]_  = \new_[2524]_  | \new_[662]_ ;
  assign \new_[2355]_  = ~\new_[2526]_  & ~\new_[796]_ ;
  assign \new_[2356]_  = ~\new_[2526]_  & ~\new_[789]_ ;
  assign \new_[2357]_  = ~\new_[2534]_  & (~\new_[2815]_  | ~\new_[1293]_ );
  assign n1489 = ~\new_[2719]_  | ~\new_[5182]_  | ~\new_[3558]_  | ~reset_n;
  assign mreq_n = mreq_n_reg;
  assign \new_[2360]_  = ~\new_[2557]_  | (~\new_[2730]_  & ~\new_[4844]_ );
  assign \new_[2361]_  = ~\new_[2558]_  | (~\new_[2729]_  & ~\new_[4847]_ );
  assign \new_[2362]_  = \new_[2671]_  ? \new_[3925]_  : \new_[1292]_ ;
  assign \new_[2363]_  = ~\new_[4965]_  | ~\new_[2562]_  | ~\new_[4966]_ ;
  assign \new_[2364]_  = ~\new_[2561]_  & (~\new_[2729]_  | ~\new_[6520]_ );
  assign \new_[2365]_  = ~\new_[2559]_  | (~\new_[2730]_  & ~\new_[4623]_ );
  assign \new_[2366]_  = ~\new_[2560]_  | (~\new_[2730]_  & ~\new_[4620]_ );
  assign \new_[2367]_  = (~\new_[4704]_  | ~\new_[1394]_ ) & (~\new_[2676]_  | ~\new_[5304]_ );
  assign \new_[2368]_  = ~\new_[2573]_  | ~\new_[3276]_ ;
  assign \new_[2369]_  = ~\new_[2575]_  & ~\new_[7335]_ ;
  assign \new_[2370]_  = ~\new_[2576]_  & ~\new_[7335]_ ;
  assign \new_[2371]_  = ~\new_[2578]_  | ~\new_[4864]_ ;
  assign \new_[2372]_  = ~\new_[2729]_  | ~\new_[740]_ ;
  assign \new_[2373]_  = ~\new_[4281]_  & ~\new_[2729]_ ;
  assign \new_[2374]_  = ~\new_[2577]_  | ~\new_[3509]_ ;
  assign \new_[2375]_  = ~\new_[2569]_  & (~\new_[3851]_  | ~\new_[3857]_ );
  assign \new_[2376]_  = ~\new_[2569]_  & (~\new_[3852]_  | ~\new_[3861]_ );
  assign \new_[2377]_  = ~\new_[2571]_  & (~\new_[2134]_  | ~\new_[6252]_ );
  assign \new_[2378]_  = ~\new_[3498]_  | (~\new_[2680]_  & ~\new_[3620]_ );
  assign \new_[2379]_  = ~\new_[2567]_  & (~\new_[1578]_  | ~\new_[6712]_ );
  assign \new_[2380]_  = ~\new_[2441]_ ;
  assign \new_[2381]_  = ~\new_[2566]_  & (~\new_[5832]_  | ~\new_[7335]_ );
  assign \new_[2382]_  = ~\new_[2565]_  & (~\new_[6723]_  | ~\new_[757]_ );
  assign \new_[2383]_  = ~\new_[2447]_ ;
  assign \new_[2384]_  = ~\new_[2447]_ ;
  assign \new_[2385]_  = ~\new_[2581]_  & (~\new_[7485]_  | ~\new_[574]_ );
  assign \new_[2386]_  = ~\new_[2600]_  | ~\new_[2599]_ ;
  assign \new_[2387]_  = ~\new_[2601]_  | ~\new_[2611]_ ;
  assign \new_[2388]_  = (~\new_[2706]_  | ~n304) & (~\new_[7489]_  | ~n299);
  assign \new_[2389]_  = ~\new_[2582]_  & (~\new_[7275]_  | ~\new_[576]_ );
  assign \new_[2390]_  = ~\new_[2713]_  | ~\new_[6615]_ ;
  assign \new_[2391]_  = ~\new_[2712]_  | ~\new_[6583]_ ;
  assign \new_[2392]_  = ~\new_[2713]_  | ~\new_[6645]_ ;
  assign \new_[2393]_  = ~\new_[2713]_  | ~\new_[6564]_ ;
  assign \new_[2394]_  = ~\new_[2712]_  | ~\new_[6660]_ ;
  assign \new_[2395]_  = ~\new_[2712]_  | ~\new_[6641]_ ;
  assign \new_[2396]_  = ~\new_[2713]_  | ~\new_[430]_ ;
  assign \new_[2397]_  = ~\new_[2712]_  | ~\new_[431]_ ;
  assign \new_[2398]_  = ~\new_[2753]_  | ~\new_[791]_ ;
  assign \new_[2399]_  = ~\new_[7459]_  | ~\new_[797]_ ;
  assign \new_[2400]_  = ~\new_[6976]_  | ~\new_[542]_ ;
  assign \new_[2401]_  = ~\new_[2628]_  | ~\new_[6607]_ ;
  assign \new_[2402]_  = ~\new_[2628]_  | ~\new_[6665]_ ;
  assign \new_[2403]_  = ~\new_[2628]_  | ~\new_[6673]_ ;
  assign \new_[2404]_  = ~\new_[2628]_  | ~\new_[6652]_ ;
  assign \new_[2405]_  = ~\new_[2628]_  | ~\new_[435]_ ;
  assign \new_[2406]_  = \new_[6644]_  | \new_[7398]_ ;
  assign \new_[2407]_  = \new_[428]_  | \new_[7398]_ ;
  assign \new_[2408]_  = \new_[6491]_  | \new_[7398]_ ;
  assign \new_[2409]_  = ~\new_[6638]_  | ~\new_[2627]_ ;
  assign \new_[2410]_  = ~\new_[7398]_  & ~\new_[767]_ ;
  assign \new_[2411]_  = \new_[7398]_  | \new_[730]_ ;
  assign \new_[2412]_  = \new_[7398]_  | \new_[659]_ ;
  assign \new_[2413]_  = \new_[6598]_  | \new_[7398]_ ;
  assign \new_[2414]_  = \new_[7398]_  | \new_[650]_ ;
  assign \new_[2415]_  = \new_[7398]_  | \new_[528]_ ;
  assign \new_[2416]_  = \new_[7398]_  | \new_[567]_ ;
  assign \new_[2417]_  = ~\new_[6846]_  | ~\new_[6609]_ ;
  assign \new_[2418]_  = ~\new_[6555]_  | ~\new_[6853]_ ;
  assign \new_[2419]_  = ~\new_[511]_  | ~\new_[6853]_ ;
  assign \new_[2420]_  = ~\new_[7419]_  | ~\new_[6563]_ ;
  assign \new_[2421]_  = ~\new_[2629]_  & ~\new_[5746]_ ;
  assign \new_[2422]_  = ~\new_[2524]_ ;
  assign \new_[2423]_  = ~\new_[2526]_ ;
  assign \new_[2424]_  = ~\new_[2635]_  & (~\new_[3925]_  | ~\new_[1255]_ );
  assign \new_[2425]_  = ~\new_[2634]_  & (~\new_[1233]_  | ~\new_[5746]_ );
  assign \new_[2426]_  = ~\new_[2637]_  & (~\new_[1223]_  | ~\new_[5746]_ );
  assign n1494 = \new_[2717]_  ? \new_[1690]_  : \new_[2254]_ ;
  assign \new_[2428]_  = \new_[2656]_  | \new_[6711]_ ;
  assign \new_[2429]_  = \\i_tv80_core_TmpAddr_reg[0] ;
  assign \new_[2430]_  = \\i_tv80_core_RegAddrB_r_reg[0] ;
  assign \new_[2431]_  = \\i_tv80_core_RegAddrB_r_reg[1] ;
  assign \new_[2432]_  = ~\new_[2667]_  | (~\new_[2730]_  & ~\new_[4624]_ );
  assign \new_[2433]_  = ~\new_[2668]_  | (~\new_[2730]_  & ~\new_[4621]_ );
  assign \new_[2434]_  = ~\new_[2669]_  | (~\new_[2730]_  & ~\new_[4622]_ );
  assign \new_[2435]_  = ~\new_[2670]_  | (~\new_[2729]_  & ~\new_[4618]_ );
  assign \new_[2436]_  = \new_[4078]_  ? \new_[2729]_  : \new_[6606]_ ;
  assign \new_[2437]_  = \new_[4079]_  ? \new_[2729]_  : \new_[6591]_ ;
  assign \new_[2438]_  = ~\new_[6723]_  & (~\new_[3425]_  | ~\new_[2735]_ );
  assign \new_[2439]_  = ~\new_[3663]_  & (~\new_[2737]_  | ~\new_[4680]_ );
  assign \new_[2440]_  = ~\new_[2676]_  | ~\new_[3509]_ ;
  assign \new_[2441]_  = ~\new_[2673]_  & (~\new_[1610]_  | ~\new_[6713]_ );
  assign \new_[2442]_  = \new_[2740]_  ? \new_[5724]_  : \new_[1294]_ ;
  assign \new_[2443]_  = ~\new_[2672]_  & (~\new_[6723]_  | ~\new_[853]_ );
  assign \new_[2444]_  = \new_[3387]_  ^ \new_[2731]_ ;
  assign \new_[2445]_  = \new_[4558]_  ? \new_[3276]_  : \new_[2738]_ ;
  assign \new_[2446]_  = ~\new_[2681]_  | ~\new_[6047]_ ;
  assign \new_[2447]_  = \new_[2568]_ ;
  assign \new_[2448]_  = \new_[2679]_  & \new_[2955]_ ;
  assign \new_[2449]_  = \new_[6821]_  & \new_[2679]_ ;
  assign \new_[2450]_  = ~\new_[2678]_  | (~\new_[3000]_  & ~\new_[4866]_ );
  assign \new_[2451]_  = ~\new_[2572]_ ;
  assign \new_[2452]_  = (~\new_[3919]_  | ~\new_[6236]_ ) & (~\new_[2745]_  | ~\new_[5849]_ );
  assign \new_[2453]_  = ~\new_[2677]_  & (~\new_[5822]_  | ~\new_[7335]_ );
  assign \new_[2454]_  = (~\new_[4704]_  | ~\new_[1453]_ ) & (~\new_[2746]_  | ~\new_[5304]_ );
  assign \new_[2455]_  = \new_[3314]_  ^ \new_[2744]_ ;
  assign \new_[2456]_  = ~\new_[2704]_  & (~\new_[2752]_  | ~\new_[734]_ );
  assign \new_[2457]_  = ~\new_[2702]_  | ~\new_[2694]_ ;
  assign \new_[2458]_  = ~\new_[2692]_  | ~\new_[2693]_ ;
  assign \new_[2459]_  = ~\new_[2712]_  | ~\new_[788]_ ;
  assign \new_[2460]_  = ~\new_[2707]_  | ~\new_[786]_ ;
  assign \new_[2461]_  = ~\new_[2707]_  | ~\new_[6547]_ ;
  assign \new_[2462]_  = ~\new_[2713]_  | ~\new_[538]_ ;
  assign \new_[2463]_  = ~\new_[2712]_  | ~\new_[539]_ ;
  assign \new_[2464]_  = ~\new_[2706]_  | ~\new_[429]_ ;
  assign \new_[2465]_  = ~\new_[7275]_  | ~\new_[653]_ ;
  assign \new_[2466]_  = ~\new_[2706]_  | ~\new_[6566]_ ;
  assign \new_[2467]_  = ~\new_[7272]_  | ~\new_[654]_ ;
  assign \new_[2468]_  = ~\new_[2713]_  | ~\new_[787]_ ;
  assign \new_[2469]_  = ~\new_[7443]_  | ~\new_[790]_ ;
  assign \new_[2470]_  = ~\new_[7458]_  & ~\new_[6555]_ ;
  assign \new_[2471]_  = \new_[2016]_  ? \new_[4760]_  : \new_[2775]_ ;
  assign \new_[2472]_  = ~\new_[7443]_  | ~\new_[520]_ ;
  assign \new_[2473]_  = ~\new_[7489]_  | ~\new_[428]_ ;
  assign \new_[2474]_  = ~\new_[7489]_  | ~\new_[6644]_ ;
  assign \new_[2475]_  = ~\new_[6563]_  & ~\new_[6682]_ ;
  assign \new_[2476]_  = ~\new_[2708]_  & ~\new_[6553]_ ;
  assign \new_[2477]_  = ~\new_[2709]_  | ~\new_[6587]_ ;
  assign \new_[2478]_  = ~\new_[2709]_  | ~\new_[6639]_ ;
  assign \new_[2479]_  = ~\new_[2709]_  | ~\new_[6657]_ ;
  assign \new_[2480]_  = ~\new_[2709]_  | ~\new_[6599]_ ;
  assign \new_[2481]_  = ~\new_[2709]_  | ~\new_[432]_ ;
  assign \new_[2482]_  = \new_[6627]_  | \new_[7383]_ ;
  assign \new_[2483]_  = ~\new_[7383]_  & ~\new_[768]_ ;
  assign \new_[2484]_  = \new_[7383]_  | \new_[660]_ ;
  assign \new_[2485]_  = \new_[7383]_  | \new_[652]_ ;
  assign \new_[2486]_  = \new_[7383]_  | \new_[529]_ ;
  assign \new_[2487]_  = \new_[7383]_  | \new_[568]_ ;
  assign \new_[2488]_  = \new_[6618]_  | \new_[7383]_ ;
  assign \new_[2489]_  = \new_[7514]_  | \new_[657]_ ;
  assign \new_[2490]_  = \new_[664]_  | \new_[7498]_ ;
  assign \new_[2491]_  = ~\new_[7426]_  & ~\new_[778]_ ;
  assign \new_[2492]_  = ~\new_[780]_  & ~\new_[7498]_ ;
  assign \new_[2493]_  = ~\new_[7514]_  & ~\new_[772]_ ;
  assign \new_[2494]_  = \new_[578]_  | \new_[7426]_ ;
  assign \new_[2495]_  = \new_[520]_  | \new_[7426]_ ;
  assign \new_[2496]_  = \new_[6612]_  | \new_[7426]_ ;
  assign \new_[2497]_  = \new_[580]_  | \new_[7498]_ ;
  assign \new_[2498]_  = \new_[543]_  | \new_[7498]_ ;
  assign \new_[2499]_  = \new_[7426]_  | \new_[656]_ ;
  assign \new_[2500]_  = \new_[734]_  | \new_[7498]_ ;
  assign \new_[2501]_  = \new_[435]_  | \new_[7498]_ ;
  assign \new_[2502]_  = \new_[6607]_  | \new_[7498]_ ;
  assign \new_[2503]_  = \new_[6665]_  | \new_[7498]_ ;
  assign \new_[2504]_  = ~\new_[7514]_  & ~\new_[797]_ ;
  assign \new_[2505]_  = \new_[658]_  | \new_[7498]_ ;
  assign \new_[2506]_  = \new_[6673]_  | \new_[7498]_ ;
  assign \new_[2507]_  = \new_[6652]_  | \new_[7498]_ ;
  assign \new_[2508]_  = \new_[7426]_  | \new_[6602]_ ;
  assign \new_[2509]_  = ~\new_[7426]_  & ~\new_[790]_ ;
  assign \new_[2510]_  = ~\new_[7426]_  & ~\new_[771]_ ;
  assign \new_[2511]_  = \new_[7426]_  | \new_[531]_ ;
  assign \new_[2512]_  = \new_[7426]_  | \new_[572]_ ;
  assign \new_[2513]_  = ~\new_[7514]_  & ~\new_[779]_ ;
  assign \new_[2514]_  = \new_[7514]_  | \new_[532]_ ;
  assign \new_[2515]_  = \new_[7426]_  | \new_[665]_ ;
  assign \new_[2516]_  = \new_[7514]_  | \new_[573]_ ;
  assign \new_[2517]_  = ~\new_[791]_  & ~\new_[7498]_ ;
  assign \new_[2518]_  = ~\new_[773]_  & ~\new_[7498]_ ;
  assign \new_[2519]_  = \new_[533]_  | \new_[7498]_ ;
  assign \new_[2520]_  = \new_[7498]_  | \new_[562]_ ;
  assign \new_[2521]_  = \new_[7514]_  | \new_[663]_ ;
  assign \new_[2522]_  = ~\new_[2715]_  & ~\new_[5746]_ ;
  assign \new_[2523]_  = \new_[4529]_  | \new_[2720]_ ;
  assign \new_[2524]_  = ~\new_[2622]_ ;
  assign \new_[2525]_  = ~\new_[2830]_  | ~\new_[4312]_  | ~\new_[4525]_  | ~\new_[4056]_ ;
  assign \new_[2526]_  = ~\new_[2623]_ ;
  assign \new_[2529]_  = ~\new_[7398]_ ;
  assign \new_[2530]_  = \new_[7398]_ ;
  assign \new_[2531]_  = (~\new_[2861]_  | ~\new_[2957]_ ) & (~\new_[2766]_  | ~\new_[792]_ );
  assign \new_[2532]_  = (~\new_[2765]_  | ~\new_[6520]_ ) & (~\new_[2818]_  | ~\new_[853]_ );
  assign \new_[2533]_  = (~\new_[2861]_  | ~\new_[2959]_ ) & (~\new_[2766]_  | ~\new_[794]_ );
  assign \new_[2534]_  = ~\new_[2639]_ ;
  assign \new_[2535]_  = (~\new_[2765]_  | ~\new_[740]_ ) & (~\new_[2818]_  | ~\new_[851]_ );
  assign \new_[2536]_  = (~\new_[2765]_  | ~\new_[6521]_ ) & (~\new_[2818]_  | ~\new_[848]_ );
  assign \new_[2537]_  = (~\new_[2861]_  | ~\new_[2956]_ ) & (~\new_[2766]_  | ~\new_[742]_ );
  assign \new_[2538]_  = (~\new_[2765]_  | ~\new_[6606]_ ) & (~\new_[2818]_  | ~\new_[852]_ );
  assign \new_[2539]_  = (~\new_[2765]_  | ~\new_[850]_ ) & (~\new_[2818]_  | ~\new_[799]_ );
  assign \new_[2540]_  = (~\new_[2861]_  | ~\new_[2963]_ ) & (~\new_[2766]_  | ~\new_[766]_ );
  assign \new_[2541]_  = (~\new_[2861]_  | ~\new_[2960]_ ) & (~\new_[2766]_  | ~\new_[764]_ );
  assign \new_[2542]_  = (~\new_[2765]_  | ~\new_[6591]_ ) & (~\new_[2818]_  | ~\new_[849]_ );
  assign \new_[2543]_  = (~\new_[2765]_  | ~\new_[6472]_ ) & (~\new_[2818]_  | ~\new_[684]_ );
  assign \new_[2544]_  = (~\new_[2861]_  | ~\new_[2961]_ ) & (~\new_[2766]_  | ~\new_[757]_ );
  assign \new_[2545]_  = (~\new_[2765]_  | ~\new_[844]_ ) & (~\new_[2818]_  | ~\new_[845]_ );
  assign \new_[2546]_  = (~\new_[2861]_  | ~\new_[2962]_ ) & (~\new_[2766]_  | ~\new_[755]_ );
  assign \new_[2547]_  = (~\new_[2861]_  | ~\new_[2958]_ ) & (~\new_[2766]_  | ~\new_[793]_ );
  assign n1499 = ~\new_[6363]_  | ~\new_[2718]_  | ~\new_[3417]_ ;
  assign \new_[2549]_  = ~\new_[4373]_  | ~\new_[4564]_  | ~\new_[2774]_  | ~\new_[2777]_ ;
  assign \new_[2550]_  = \\i_tv80_core_RegAddrC_reg[0] ;
  assign \new_[2551]_  = \\i_tv80_core_R_reg[6] ;
  assign \new_[2552]_  = \\i_tv80_core_R_reg[5] ;
  assign \new_[2553]_  = \\i_tv80_core_R_reg[3] ;
  assign \new_[2554]_  = \\i_tv80_core_R_reg[2] ;
  assign \new_[2555]_  = \\i_tv80_core_R_reg[4] ;
  assign \new_[2556]_  = \\i_tv80_core_IR_reg[2] ;
  assign \new_[2557]_  = ~\new_[2728]_  | ~\new_[758]_ ;
  assign \new_[2558]_  = ~\new_[2728]_  | ~\new_[759]_ ;
  assign \new_[2559]_  = ~\new_[2730]_  | ~\new_[736]_ ;
  assign \new_[2560]_  = ~\new_[2730]_  | ~\new_[761]_ ;
  assign \new_[2561]_  = ~\new_[2729]_  & (~\new_[4612]_  | ~\new_[4966]_ );
  assign \new_[2562]_  = ~\new_[2729]_  & (~\new_[5221]_  | ~\new_[6625]_ );
  assign \new_[2563]_  = ~\new_[3528]_  | ~\new_[3526]_  | ~\new_[2731]_  | ~\new_[3444]_ ;
  assign \new_[2564]_  = ~\new_[2671]_ ;
  assign \new_[2565]_  = ~\new_[6723]_  & (~\new_[3370]_  | ~\new_[2797]_ );
  assign \new_[2566]_  = ~\new_[2741]_  & ~\new_[7335]_ ;
  assign \new_[2567]_  = ~\new_[2739]_  & ~\new_[3618]_ ;
  assign \new_[2568]_  = ~\new_[2734]_  | ~\new_[2944]_ ;
  assign \new_[2569]_  = ~\new_[2674]_ ;
  assign \new_[2570]_  = \new_[2734]_  & \new_[2886]_ ;
  assign \new_[2571]_  = ~\new_[1690]_  & (~\new_[7539]_  | ~\new_[5197]_ );
  assign \new_[2572]_  = ~\new_[2736]_  & (~\new_[1646]_  | ~\new_[6713]_ );
  assign \new_[2573]_  = ~\new_[2675]_ ;
  assign \new_[2574]_  = ~\new_[3355]_  | (~\new_[2800]_  & ~\new_[3619]_ );
  assign \new_[2575]_  = ~\new_[2732]_  & (~\new_[6723]_  | ~\new_[764]_ );
  assign \new_[2576]_  = ~\new_[2733]_  & (~\new_[6723]_  | ~\new_[755]_ );
  assign \new_[2577]_  = \new_[3209]_  ^ \new_[2795]_ ;
  assign \new_[2578]_  = \new_[4553]_  ? \new_[3276]_  : \new_[2799]_ ;
  assign \new_[2579]_  = ~\new_[2746]_  | ~\new_[3509]_ ;
  assign \new_[2580]_  = ~\new_[2742]_  & (~\new_[7486]_  | ~\new_[730]_ );
  assign \new_[2581]_  = ~\new_[6638]_  & ~\new_[2747]_ ;
  assign \new_[2582]_  = ~\new_[2750]_  & ~\new_[6611]_ ;
  assign \new_[2583]_  = ~\new_[7485]_  | ~\new_[785]_ ;
  assign \new_[2584]_  = ~\new_[7444]_  | ~\new_[778]_ ;
  assign \new_[2585]_  = ~\new_[6977]_  | ~\new_[779]_ ;
  assign \new_[2586]_  = ~\new_[7485]_  | ~\new_[536]_ ;
  assign \new_[2587]_  = ~\new_[2753]_  | ~\new_[543]_ ;
  assign \new_[2588]_  = ~\new_[6977]_  | ~\new_[772]_ ;
  assign \new_[2589]_  = ~\new_[2756]_  | ~\new_[771]_ ;
  assign \new_[2590]_  = ~\new_[7444]_  | ~\new_[665]_ ;
  assign \new_[2591]_  = ~\new_[6977]_  | ~\new_[663]_ ;
  assign \new_[2592]_  = ~\new_[2752]_  | ~\new_[664]_ ;
  assign \new_[2593]_  = ~\new_[2754]_  | ~\new_[773]_ ;
  assign \new_[2594]_  = ~\new_[2753]_  | ~\new_[658]_ ;
  assign \new_[2595]_  = ~\new_[656]_  | ~\new_[2756]_ ;
  assign \new_[2596]_  = ~\new_[2754]_  | ~\new_[533]_ ;
  assign \new_[2597]_  = ~\new_[7444]_  | ~\new_[531]_ ;
  assign \new_[2598]_  = ~\new_[6683]_  | ~\new_[532]_ ;
  assign \new_[2599]_  = ~\new_[7459]_  | ~\new_[573]_ ;
  assign \new_[2600]_  = ~\new_[2756]_  | ~\new_[572]_ ;
  assign \new_[2601]_  = ~\new_[2752]_  | ~\new_[6546]_ ;
  assign \new_[2602]_  = ~\new_[7459]_  | ~\new_[657]_ ;
  assign \new_[2603]_  = ~\new_[2752]_  | ~\new_[780]_ ;
  assign \new_[2604]_  = ~\new_[2749]_  | ~\new_[789]_ ;
  assign \new_[2605]_  = ~\new_[2748]_  | ~\new_[737]_ ;
  assign \new_[2606]_  = ~\new_[2749]_  | ~\new_[540]_ ;
  assign \new_[2607]_  = ~\new_[2748]_  | ~\new_[796]_ ;
  assign \new_[2608]_  = ~\new_[2748]_  | ~\new_[646]_ ;
  assign \new_[2609]_  = ~\new_[2749]_  | ~\new_[655]_ ;
  assign \new_[2610]_  = ~\new_[2748]_  | ~\new_[535]_ ;
  assign \new_[2611]_  = ~\new_[2748]_  | ~\new_[571]_ ;
  assign \new_[2612]_  = \new_[576]_  | \new_[7389]_ ;
  assign \new_[2613]_  = \new_[538]_  | \new_[7389]_ ;
  assign \new_[2614]_  = \new_[7389]_  | \new_[653]_ ;
  assign \new_[2615]_  = \new_[6615]_  | \new_[7389]_ ;
  assign \new_[2616]_  = \new_[7389]_  | \new_[661]_ ;
  assign \new_[2617]_  = \new_[7389]_  | \new_[735]_ ;
  assign \new_[2618]_  = \new_[7389]_  | \new_[530]_ ;
  assign \new_[2619]_  = \new_[7389]_  | \new_[569]_ ;
  assign \new_[2620]_  = ~\new_[7389]_  & ~\new_[769]_ ;
  assign \new_[2621]_  = \new_[2757]_  | \new_[6711]_ ;
  assign \new_[2622]_  = \new_[2849]_  | \new_[2846]_ ;
  assign \new_[2623]_  = ~\new_[2849]_  | ~\new_[2758]_ ;
  assign \new_[2624]_  = \new_[7514]_ ;
  assign \new_[2625]_  = ~\new_[7498]_ ;
  assign \new_[2626]_  = ~\new_[7498]_ ;
  assign \new_[2627]_  = ~\new_[7383]_ ;
  assign \new_[2628]_  = ~\new_[2714]_ ;
  assign \new_[2629]_  = ~\new_[2759]_  & (~\new_[3925]_  | ~\new_[1234]_ );
  assign \new_[2630]_  = ~\new_[2771]_  | (~\new_[2873]_  & ~\new_[3155]_ );
  assign \new_[2631]_  = ~\new_[2772]_  & (~\new_[3841]_  | ~\new_[6472]_ );
  assign \new_[2632]_  = \new_[2761]_  | \new_[6711]_ ;
  assign \new_[2633]_  = \\i_tv80_core_R_reg[0] ;
  assign \new_[2634]_  = ~\new_[2762]_  & ~\new_[5746]_ ;
  assign \new_[2635]_  = ~\new_[3925]_  & ~\new_[2763]_ ;
  assign \new_[2636]_  = ~\new_[2763]_  & ~\new_[4316]_ ;
  assign \new_[2637]_  = ~\new_[2764]_  & ~\new_[5724]_ ;
  assign \new_[2638]_  = (~\new_[2851]_  | ~\new_[1294]_ ) & (~\new_[2815]_  | ~\new_[1237]_ );
  assign \new_[2639]_  = (~\new_[3112]_  | ~\new_[2821]_ ) & (~\new_[2851]_  | ~\new_[1242]_ );
  assign \new_[2640]_  = (~\new_[2852]_  | ~\new_[4560]_ ) & (~\new_[2816]_  | ~\new_[736]_ );
  assign \new_[2641]_  = (~\new_[2851]_  | ~\new_[1223]_ ) & (~\new_[2815]_  | ~\new_[1236]_ );
  assign \new_[2642]_  = (~\new_[2852]_  | ~\new_[4554]_ ) & (~\new_[2816]_  | ~\new_[762]_ );
  assign \new_[2643]_  = (~\new_[2852]_  | ~\new_[4557]_ ) & (~\new_[2816]_  | ~\new_[761]_ );
  assign \new_[2644]_  = (~\new_[2851]_  | ~\new_[1233]_ ) & (~\new_[2815]_  | ~\new_[1238]_ );
  assign \new_[2645]_  = (~\new_[2851]_  | ~\new_[1234]_ ) & (~\new_[2815]_  | ~\new_[1239]_ );
  assign \new_[2646]_  = (~\new_[2851]_  | ~\new_[1235]_ ) & (~\new_[2815]_  | ~\new_[1240]_ );
  assign \new_[2647]_  = (~\new_[2852]_  | ~\new_[4559]_ ) & (~\new_[2816]_  | ~\new_[759]_ );
  assign \new_[2648]_  = (~\new_[2852]_  | ~\new_[4549]_ ) & (~\new_[2816]_  | ~\new_[760]_ );
  assign \new_[2649]_  = (~\new_[2851]_  | ~\new_[1292]_ ) & (~\new_[2815]_  | ~\new_[1241]_ );
  assign \new_[2650]_  = (~\new_[2852]_  | ~\new_[4556]_ ) & (~\new_[2816]_  | ~\new_[753]_ );
  assign \new_[2651]_  = (~\new_[2851]_  | ~\new_[1255]_ ) & (~\new_[2815]_  | ~\new_[1225]_ );
  assign \new_[2652]_  = (~\new_[2852]_  | ~\new_[4558]_ ) & (~\new_[2816]_  | ~\new_[763]_ );
  assign \new_[2653]_  = (~\new_[2852]_  | ~\new_[4553]_ ) & (~\new_[2816]_  | ~\new_[758]_ );
  assign n1509 = ~\new_[2773]_  | ~\new_[2768]_ ;
  assign n1514 = ~\new_[2922]_  | ~\new_[2768]_ ;
  assign \new_[2656]_  = ~\new_[2767]_  & (~\new_[1240]_  | ~\new_[5746]_ );
  assign n1504 = ~\new_[2770]_  & ~\new_[6426]_ ;
  assign \new_[2658]_  = ~\new_[2777]_  | ~\new_[3183]_ ;
  assign rd_n = rd_n_reg;
  assign \new_[2660]_  = \\i_tv80_core_ISet_reg[0] ;
  assign \new_[2661]_  = \\i_tv80_core_R_reg[1] ;
  assign \new_[2662]_  = \\i_tv80_core_IR_reg[0] ;
  assign \new_[2663]_  = \\i_tv80_core_IR_reg[1] ;
  assign \new_[2664]_  = \\i_tv80_core_IR_reg[5] ;
  assign \new_[2665]_  = \\i_tv80_core_IR_reg[6] ;
  assign \new_[2666]_  = \\i_tv80_core_IR_reg[7] ;
  assign \new_[2667]_  = ~\new_[2790]_  | ~\new_[762]_ ;
  assign \new_[2668]_  = ~\new_[2790]_  | ~\new_[763]_ ;
  assign \new_[2669]_  = ~\new_[2790]_  | ~\new_[760]_ ;
  assign \new_[2670]_  = ~\new_[2790]_  | ~\new_[753]_ ;
  assign \new_[2671]_  = \new_[3721]_  ^ \new_[2833]_ ;
  assign \new_[2672]_  = ~\new_[6723]_  & (~\new_[3426]_  | ~\new_[2836]_ );
  assign \new_[2673]_  = ~\new_[2793]_  & ~\new_[3617]_ ;
  assign \new_[2674]_  = ~\new_[2729]_ ;
  assign \new_[2675]_  = (~\new_[2838]_  | ~\new_[6711]_ ) & (~\new_[1689]_  | ~\new_[6712]_ );
  assign \new_[2676]_  = \new_[3253]_  ^ \new_[2834]_ ;
  assign \new_[2677]_  = ~\new_[2801]_  & ~\new_[7335]_ ;
  assign \new_[2678]_  = ~\new_[2802]_  | ~\new_[6047]_ ;
  assign \new_[2679]_  = \new_[2992]_  & \new_[7539]_ ;
  assign \new_[2680]_  = ~\new_[2796]_  & (~\new_[5837]_  | ~\new_[7335]_ );
  assign \new_[2681]_  = \new_[4557]_  ? \new_[3276]_  : \new_[2843]_ ;
  assign \new_[2682]_  = ~\new_[7272]_  | ~\new_[777]_ ;
  assign \new_[2683]_  = ~\new_[7275]_  | ~\new_[769]_ ;
  assign \new_[2684]_  = ~\new_[768]_  | ~\new_[2804]_ ;
  assign \new_[2685]_  = ~\new_[2804]_  | ~\new_[660]_ ;
  assign \new_[2686]_  = ~\new_[7275]_  | ~\new_[661]_ ;
  assign \new_[2687]_  = ~\new_[7272]_  | ~\new_[770]_ ;
  assign \new_[2688]_  = ~\new_[7272]_  | ~\new_[662]_ ;
  assign \new_[2689]_  = ~\new_[529]_  | ~\new_[2803]_ ;
  assign \new_[2690]_  = ~\new_[7272]_  | ~\new_[534]_ ;
  assign \new_[2691]_  = ~\new_[7275]_  | ~\new_[530]_ ;
  assign \new_[2692]_  = ~\new_[7275]_  | ~\new_[569]_ ;
  assign \new_[2693]_  = ~\new_[7272]_  | ~\new_[570]_ ;
  assign \new_[2694]_  = ~\new_[2803]_  | ~\new_[568]_ ;
  assign \new_[2695]_  = ~\new_[2803]_  | ~\new_[652]_ ;
  assign \new_[2696]_  = ~\new_[7275]_  | ~\new_[776]_ ;
  assign \new_[2697]_  = ~\new_[2804]_  | ~\new_[775]_ ;
  assign \new_[2698]_  = ~\new_[7486]_  | ~\new_[767]_ ;
  assign \new_[2699]_  = ~\new_[7486]_  | ~\new_[659]_ ;
  assign \new_[2700]_  = ~\new_[7486]_  | ~\new_[650]_ ;
  assign \new_[2701]_  = ~\new_[7486]_  | ~\new_[528]_ ;
  assign \new_[2702]_  = ~\new_[7486]_  | ~\new_[567]_ ;
  assign \new_[2703]_  = ~\new_[7486]_  | ~\new_[774]_ ;
  assign \new_[2704]_  = ~\new_[2805]_  & ~\new_[6630]_ ;
  assign n1519 = ~\new_[2812]_  | ~\new_[4588]_ ;
  assign \new_[2706]_  = ~\new_[2747]_ ;
  assign \new_[2707]_  = ~\new_[2747]_ ;
  assign \new_[2708]_  = ~\new_[2748]_ ;
  assign \new_[2709]_  = \new_[2749]_ ;
  assign \new_[2710]_  = \new_[7389]_ ;
  assign \new_[2711]_  = ~\new_[7389]_ ;
  assign \new_[2712]_  = ~\new_[2750]_ ;
  assign \new_[2713]_  = ~\new_[2751]_ ;
  assign \new_[2714]_  = ~\new_[2753]_ ;
  assign \new_[2715]_  = ~\new_[2810]_  & (~\new_[3925]_  | ~\new_[1235]_ );
  assign \new_[2716]_  = \\i_tv80_core_ISet_reg[1] ;
  assign \new_[2717]_  = \new_[3029]_  ? \new_[2860]_  : \new_[2780]_ ;
  assign \new_[2718]_  = ~\new_[2820]_  & (~\new_[3825]_  | ~\new_[3061]_ );
  assign \new_[2719]_  = ~\new_[2819]_  & (~\new_[3903]_  | ~\new_[3061]_ );
  assign \new_[2720]_  = \new_[3434]_  & \new_[2831]_ ;
  assign n1524 = ~\new_[2822]_  & ~\new_[6329]_ ;
  assign n1529 = ~\new_[2824]_  & ~\new_[6623]_ ;
  assign \new_[2723]_  = ~\new_[2823]_  | ~\new_[3183]_ ;
  assign n1534 = ~\new_[2825]_  & ~\new_[6424]_ ;
  assign n1539 = ~\new_[2827]_  & ~\new_[6327]_ ;
  assign n1544 = ~\new_[2828]_  & ~\new_[6417]_ ;
  assign \new_[2727]_  = \\i_tv80_core_IR_reg[4] ;
  assign \new_[2728]_  = \new_[6706]_  | \new_[5221]_ ;
  assign \new_[2729]_  = ~\new_[2789]_ ;
  assign \new_[2730]_  = ~\new_[2791]_ ;
  assign \new_[2731]_  = ~\new_[3379]_  | (~\new_[2887]_  & ~\new_[3519]_ );
  assign \new_[2732]_  = ~\new_[6723]_  & (~\new_[3371]_  | ~\new_[2881]_ );
  assign \new_[2733]_  = ~\new_[6723]_  & (~\new_[3369]_  | ~\new_[2882]_ );
  assign \new_[2734]_  = ~\new_[7540]_  & ~\new_[6725]_ ;
  assign \new_[2735]_  = ~\new_[2840]_  | ~\new_[3509]_ ;
  assign \new_[2736]_  = ~\new_[2839]_  & ~\new_[3617]_ ;
  assign \new_[2737]_  = ~\new_[2840]_  | ~\new_[5304]_ ;
  assign \new_[2738]_  = ~\new_[2792]_ ;
  assign \new_[2739]_  = (~\new_[4704]_  | ~\new_[1578]_ ) & (~\new_[2890]_  | ~\new_[5304]_ );
  assign \new_[2740]_  = ~\new_[3803]_  | (~\new_[3925]_  & ~\new_[2891]_ );
  assign \new_[2741]_  = ~\new_[2835]_  & (~\new_[6723]_  | ~\new_[766]_ );
  assign \new_[2742]_  = ~\new_[2841]_  & ~\new_[6609]_ ;
  assign \new_[2743]_  = \new_[2844]_  | \new_[6711]_ ;
  assign \new_[2744]_  = ~\new_[3054]_  & (~\new_[3249]_  | ~\new_[2895]_ );
  assign \new_[2745]_  = ~\new_[3359]_  | (~\new_[2896]_  & ~\new_[3620]_ );
  assign \new_[2746]_  = \new_[3389]_  ^ \new_[2895]_ ;
  assign \new_[2747]_  = ~\new_[2803]_ ;
  assign \new_[2748]_  = ~\new_[2805]_ ;
  assign \new_[2749]_  = ~\new_[2805]_ ;
  assign \new_[2750]_  = ~\new_[7272]_ ;
  assign \new_[2751]_  = ~\new_[7275]_ ;
  assign \new_[2752]_  = ~\new_[2806]_ ;
  assign \new_[2753]_  = ~\new_[2806]_ ;
  assign \new_[2754]_  = ~\new_[2806]_ ;
  assign \new_[2755]_  = ~\new_[3105]_  & ~\new_[2848]_ ;
  assign \new_[2756]_  = ~\new_[7445]_ ;
  assign \new_[2757]_  = ~\new_[2847]_  & (~\new_[1242]_  | ~\new_[5746]_ );
  assign \new_[2758]_  = ~\new_[2951]_  & ~\new_[2954]_ ;
  assign \new_[2759]_  = ~\new_[3925]_  & ~\new_[2850]_ ;
  assign \new_[2760]_  = ~\new_[2850]_  & ~\new_[4316]_ ;
  assign \new_[2761]_  = ~\new_[2855]_  & (~\new_[1225]_  | ~\new_[5746]_ );
  assign \new_[2762]_  = ~\new_[2853]_  & (~\new_[3925]_  | ~\new_[1233]_ );
  assign \new_[2763]_  = \new_[3807]_  ^ \new_[2921]_ ;
  assign \new_[2764]_  = ~\new_[2856]_  & (~\new_[3925]_  | ~\new_[1223]_ );
  assign \new_[2765]_  = ~\new_[3112]_  & ~\new_[2859]_ ;
  assign \new_[2766]_  = \new_[3112]_  & \new_[2858]_ ;
  assign \new_[2767]_  = ~\new_[2862]_  & ~\new_[5724]_ ;
  assign \new_[2768]_  = \new_[2860]_  | \new_[6258]_ ;
  assign n1559 = ~\new_[2974]_  | ~\new_[3558]_  | ~\new_[3836]_  | ~reset_n;
  assign \new_[2770]_  = (~\new_[2924]_  | ~\new_[6099]_ ) & (~\new_[2429]_  | ~\new_[1690]_ );
  assign \new_[2771]_  = ~\new_[2873]_  | ~\new_[3155]_ ;
  assign \new_[2772]_  = ~\new_[2867]_  & ~\new_[3841]_ ;
  assign \new_[2773]_  = (~\new_[3027]_  | ~\new_[6348]_ ) & (~\new_[2430]_  | ~\new_[6299]_ );
  assign \new_[2774]_  = ~\new_[2823]_ ;
  assign \new_[2775]_  = \new_[4556]_  ? \new_[1623]_  : \new_[2933]_ ;
  assign n1554 = ~\new_[2866]_  & ~\new_[6417]_ ;
  assign \new_[2777]_  = ~\new_[3069]_  | ~\new_[2865]_ ;
  assign n1564 = ~\new_[2869]_  & ~\new_[6441]_ ;
  assign \new_[2779]_  = \\i_tv80_core_IR_reg[3] ;
  assign \new_[2780]_  = i_tv80_core_Alternate_reg;
  assign n1574 = ~\new_[2874]_  & ~\new_[6424]_ ;
  assign n1579 = ~\new_[2875]_  & ~\new_[6623]_ ;
  assign n1549 = ~\new_[2876]_  & ~\new_[6424]_ ;
  assign n1584 = ~\new_[2877]_  & ~\new_[6424]_ ;
  assign n1589 = ~\new_[2878]_  & ~\new_[6424]_ ;
  assign n1594 = ~\new_[2879]_  & ~\new_[6424]_ ;
  assign \new_[2787]_  = ~\new_[2831]_ ;
  assign n1569 = ~\new_[2868]_  & ~\new_[6323]_ ;
  assign \new_[2789]_  = ~\new_[7194]_ ;
  assign \new_[2790]_  = \new_[6706]_ ;
  assign \new_[2791]_  = ~\new_[7194]_ ;
  assign \new_[2792]_  = (~\new_[2945]_  | ~\new_[3616]_ ) & (~\new_[1861]_  | ~\new_[6712]_ );
  assign \new_[2793]_  = (~\new_[4704]_  | ~\new_[1610]_ ) & (~\new_[2946]_  | ~\new_[5304]_ );
  assign \new_[2794]_  = ~\new_[4426]_  | ~\new_[2883]_ ;
  assign \new_[2795]_  = ~\new_[3143]_  | ~\new_[3378]_  | ~\new_[2949]_ ;
  assign \new_[2796]_  = ~\new_[2889]_  & ~\new_[7335]_ ;
  assign \new_[2797]_  = ~\new_[2890]_  | ~\new_[3509]_ ;
  assign \new_[2798]_  = ~\new_[2891]_  & ~\new_[4316]_ ;
  assign \new_[2799]_  = ~\new_[2837]_ ;
  assign \new_[2800]_  = ~\new_[2885]_  & (~\new_[5841]_  | ~\new_[7335]_ );
  assign \new_[2801]_  = ~\new_[2880]_  & (~\new_[6723]_  | ~\new_[793]_ );
  assign \new_[2802]_  = \new_[4554]_  ? \new_[3276]_  : \new_[2950]_ ;
  assign \new_[2803]_  = ~\new_[2841]_ ;
  assign \new_[2804]_  = ~\new_[2841]_ ;
  assign \new_[2805]_  = ~\new_[2898]_  | ~\new_[2947]_ ;
  assign \new_[2806]_  = ~\new_[2893]_  | ~\new_[2899]_ ;
  assign \new_[2807]_  = ~\new_[4424]_  | ~\new_[2897]_ ;
  assign \new_[2808]_  = ~\new_[2846]_ ;
  assign \new_[2809]_  = ~\new_[2951]_  | ~\new_[2909]_ ;
  assign \new_[2810]_  = ~\new_[3925]_  & ~\new_[2908]_ ;
  assign \new_[2811]_  = ~\new_[2908]_  & ~\new_[4316]_ ;
  assign \new_[2812]_  = (~\new_[4921]_  | ~\new_[2955]_ ) & (~\new_[2550]_  | ~\new_[6190]_ );
  assign \new_[2813]_  = ~\new_[3026]_  | ~\new_[6163]_ ;
  assign \new_[2814]_  = ~\new_[2849]_ ;
  assign \new_[2815]_  = \new_[2920]_  & \new_[3112]_ ;
  assign \new_[2816]_  = ~\new_[2919]_  & ~\new_[3112]_ ;
  assign \new_[2817]_  = \new_[2923]_  | \new_[6711]_ ;
  assign \new_[2818]_  = ~\new_[3112]_  & ~\new_[2918]_ ;
  assign \new_[2819]_  = ~\new_[4371]_  & (~\new_[3062]_  | ~\new_[2975]_ );
  assign \new_[2820]_  = ~\new_[4371]_  & (~\new_[3060]_  | ~\new_[2975]_ );
  assign \new_[2821]_  = ~\new_[2859]_ ;
  assign \new_[2822]_  = (~\new_[2979]_  | ~\new_[6099]_ ) & (~\new_[2551]_  | ~\new_[1690]_ );
  assign \new_[2823]_  = ~\new_[3068]_  | ~\new_[2927]_ ;
  assign \new_[2824]_  = (~\new_[2981]_  | ~\new_[6099]_ ) & (~\new_[2552]_  | ~\new_[6165]_ );
  assign \new_[2825]_  = (~\new_[2980]_  | ~busak_n) & (~\new_[2553]_  | ~\new_[6258]_ );
  assign \new_[2826]_  = i_tv80_core_XY_Ind_reg;
  assign \new_[2827]_  = (~\new_[2984]_  | ~busak_n) & (~\new_[2554]_  | ~\new_[6258]_ );
  assign \new_[2828]_  = (~\new_[2985]_  | ~busak_n) & (~\new_[2555]_  | ~\new_[1690]_ );
  assign n1599 = ~\new_[2932]_  & ~\new_[6424]_ ;
  assign \new_[2830]_  = ~\new_[2934]_  & (~\new_[4682]_  | ~\new_[844]_ );
  assign \new_[2831]_  = \new_[2002]_  ? \new_[4760]_  : \new_[2943]_ ;
  assign wr_n = wr_n_reg;
  assign \new_[2833]_  = ~\new_[2993]_  | ~\new_[3948]_  | ~\new_[3397]_ ;
  assign \new_[2834]_  = ~\new_[3042]_  | ~\new_[3250]_  | ~\new_[2998]_ ;
  assign \new_[2835]_  = ~\new_[6723]_  & (~\new_[3367]_  | ~\new_[2995]_ );
  assign \new_[2836]_  = ~\new_[2946]_  | ~\new_[3509]_ ;
  assign \new_[2837]_  = (~\new_[3001]_  | ~\new_[3616]_ ) & (~\new_[1892]_  | ~\new_[6713]_ );
  assign \new_[2838]_  = \new_[4508]_  ? \new_[5304]_  : \new_[3004]_ ;
  assign \new_[2839]_  = (~\new_[4704]_  | ~\new_[1646]_ ) & (~\new_[3005]_  | ~\new_[5304]_ );
  assign \new_[2840]_  = \new_[3382]_  ^ \new_[2997]_ ;
  assign \new_[2841]_  = ~\new_[3015]_  | ~\new_[7447]_  | ~\new_[2952]_ ;
  assign \new_[2842]_  = ~\new_[2886]_ ;
  assign \new_[2843]_  = ~\new_[2888]_ ;
  assign \new_[2844]_  = ~\new_[2948]_  & (~\new_[1241]_  | ~\new_[5746]_ );
  assign \new_[2845]_  = ~\new_[3009]_  | ~\new_[2954]_ ;
  assign \new_[2846]_  = ~\new_[2951]_  | ~\new_[2954]_ ;
  assign \new_[2847]_  = ~\new_[2953]_  & ~\new_[5724]_ ;
  assign \new_[2848]_  = ~\new_[3157]_  | ~\new_[3052]_  | ~\new_[3152]_  | ~\new_[3051]_ ;
  assign \new_[2849]_  = \new_[2899]_ ;
  assign \new_[2850]_  = \new_[3717]_  ^ \new_[3018]_ ;
  assign \new_[2851]_  = ~\new_[2965]_  & ~\new_[3112]_ ;
  assign \new_[2852]_  = \new_[2964]_  & \new_[3112]_ ;
  assign \new_[2853]_  = ~\new_[3925]_  & ~\new_[2968]_ ;
  assign \new_[2854]_  = ~\new_[2968]_  & ~\new_[4316]_ ;
  assign \new_[2855]_  = ~\new_[2966]_  & ~\new_[5724]_ ;
  assign \new_[2856]_  = ~\new_[3925]_  & ~\new_[2967]_ ;
  assign \new_[2857]_  = ~\new_[2967]_  & ~\new_[4316]_ ;
  assign \new_[2858]_  = ~\new_[2918]_ ;
  assign \new_[2859]_  = \new_[3064]_  | \new_[2970]_ ;
  assign \new_[2860]_  = ~\new_[6428]_  | ~\new_[3064]_  | ~\new_[3160]_ ;
  assign \new_[2861]_  = ~\new_[3383]_  & (~\new_[3027]_  | ~\new_[3160]_ );
  assign \new_[2862]_  = ~\new_[2971]_  & (~\new_[3925]_  | ~\new_[1240]_ );
  assign \new_[2863]_  = \\i_tv80_core_mcycles_reg[0] ;
  assign \new_[2864]_  = ~\new_[3282]_  & (~\new_[3031]_  | ~\new_[6193]_ );
  assign \new_[2865]_  = (~\new_[3470]_  | ~\new_[6272]_ ) & (~\new_[3030]_  | ~\new_[6193]_ );
  assign \new_[2866]_  = ~\new_[2982]_  & (~\new_[2633]_  | ~\new_[6338]_ );
  assign \new_[2867]_  = ~\new_[3039]_  | ~\new_[3610]_  | ~\new_[3996]_  | ~\new_[6410]_ ;
  assign \new_[2868]_  = ~\new_[2983]_  & (~\new_[2661]_  | ~\new_[6338]_ );
  assign \new_[2869]_  = (~\new_[3032]_  | ~\new_[6388]_ ) & (~\new_[2660]_  | ~\new_[6252]_ );
  assign n1609 = ~\new_[2986]_  & ~\new_[6424]_ ;
  assign n1604 = ~\new_[2987]_  & ~\new_[6424]_ ;
  assign n1614 = ~\new_[2936]_  & ~\new_[6403]_ ;
  assign \new_[2873]_  = \new_[3554]_  ? \new_[2991]_  : \new_[3497]_ ;
  assign \new_[2874]_  = ~\new_[2937]_  & (~\new_[6113]_  | ~\new_[1690]_ );
  assign \new_[2875]_  = ~\new_[2938]_  & (~\new_[6227]_  | ~\new_[1690]_ );
  assign \new_[2876]_  = ~\new_[2939]_  & (~\new_[7549]_  | ~\new_[6338]_ );
  assign \new_[2877]_  = ~\new_[2940]_  & (~\new_[6128]_  | ~\new_[6338]_ );
  assign \new_[2878]_  = ~\new_[2941]_  & (~\new_[6152]_  | ~\new_[1690]_ );
  assign \new_[2879]_  = ~\new_[2942]_  & (~\new_[6120]_  | ~\new_[1690]_ );
  assign \new_[2880]_  = ~\new_[6723]_  & (~\new_[3368]_  | ~\new_[3043]_ );
  assign \new_[2881]_  = ~\new_[3004]_  | ~\new_[3509]_ ;
  assign \new_[2882]_  = ~\new_[3005]_  | ~\new_[3509]_ ;
  assign \new_[2883]_  = ~\new_[3434]_  | ~\new_[3020]_ ;
  assign \new_[2884]_  = ~\new_[3020]_  | ~\new_[6163]_ ;
  assign \new_[2885]_  = ~\new_[3003]_  & ~\new_[7335]_ ;
  assign \new_[2886]_  = ~\new_[2944]_ ;
  assign \new_[2887]_  = ~\new_[3437]_  & (~\new_[3045]_  | ~\new_[3518]_ );
  assign \new_[2888]_  = ~\new_[2996]_  & (~\new_[1925]_  | ~\new_[6712]_ );
  assign \new_[2889]_  = ~\new_[2994]_  & (~\new_[6723]_  | ~\new_[792]_ );
  assign \new_[2890]_  = \new_[3513]_  ^ \new_[3045]_ ;
  assign \new_[2891]_  = \new_[3798]_  ^ \new_[3046]_ ;
  assign \new_[2892]_  = \new_[3010]_  | \new_[6711]_ ;
  assign \new_[2893]_  = ~\new_[7448]_  & ~\new_[3017]_ ;
  assign \new_[2894]_  = ~\new_[3044]_  & ~\new_[3016]_ ;
  assign \new_[2895]_  = ~\new_[3380]_  | ~\new_[3006]_  | ~\new_[3299]_ ;
  assign \new_[2896]_  = ~\new_[3007]_  & (~\new_[5833]_  | ~\new_[7335]_ );
  assign \new_[2897]_  = ~\new_[3434]_  | ~\new_[3026]_ ;
  assign \new_[2898]_  = ~\new_[7446]_ ;
  assign \new_[2899]_  = ~\new_[2952]_ ;
  assign \new_[2900]_  = (~\new_[3106]_  | ~\new_[4560]_ ) & (~\new_[3198]_  | ~\new_[794]_ );
  assign \new_[2901]_  = (~\new_[3106]_  | ~\new_[4554]_ ) & (~\new_[3198]_  | ~\new_[742]_ );
  assign \new_[2902]_  = (~\new_[3106]_  | ~\new_[4553]_ ) & (~\new_[3198]_  | ~\new_[793]_ );
  assign \new_[2903]_  = (~\new_[3106]_  | ~\new_[4559]_ ) & (~\new_[3198]_  | ~\new_[764]_ );
  assign \new_[2904]_  = (~\new_[3106]_  | ~\new_[4549]_ ) & (~\new_[3198]_  | ~\new_[757]_ );
  assign \new_[2905]_  = (~\new_[3106]_  | ~\new_[4556]_ ) & (~\new_[3198]_  | ~\new_[755]_ );
  assign \new_[2906]_  = (~\new_[3106]_  | ~\new_[4558]_ ) & (~\new_[3198]_  | ~\new_[766]_ );
  assign \new_[2907]_  = (~\new_[3106]_  | ~\new_[4557]_ ) & (~\new_[3198]_  | ~\new_[792]_ );
  assign \new_[2908]_  = \new_[3718]_  ^ \new_[3053]_ ;
  assign \new_[2909]_  = ~\new_[2954]_ ;
  assign \new_[2910]_  = ~\new_[3019]_  | ~\new_[762]_ ;
  assign \new_[2911]_  = ~\new_[3019]_  | ~\new_[763]_ ;
  assign \new_[2912]_  = ~\new_[3019]_  | ~\new_[759]_ ;
  assign \new_[2913]_  = ~\new_[3019]_  | ~\new_[758]_ ;
  assign \new_[2914]_  = ~\new_[3019]_  | ~\new_[760]_ ;
  assign \new_[2915]_  = ~\new_[3019]_  | ~\new_[753]_ ;
  assign \new_[2916]_  = ~\new_[3019]_  | ~\new_[761]_ ;
  assign \new_[2917]_  = ~\new_[3019]_  | ~\new_[736]_ ;
  assign \new_[2918]_  = ~\new_[3064]_  | ~\new_[3021]_ ;
  assign \new_[2919]_  = ~\new_[2964]_ ;
  assign \new_[2920]_  = ~\new_[2965]_ ;
  assign \new_[2921]_  = ~\new_[3022]_  | ~\new_[3453]_ ;
  assign \new_[2922]_  = (~\new_[3160]_  | ~\new_[6326]_ ) & (~\new_[2431]_  | ~\new_[6299]_ );
  assign \new_[2923]_  = ~\new_[3023]_  & (~\new_[1238]_  | ~\new_[5746]_ );
  assign \new_[2924]_  = ~\new_[3025]_  | (~\new_[3399]_  & ~\new_[6047]_ );
  assign n1619 = ~\new_[3028]_  & ~\new_[6329]_ ;
  assign \new_[2926]_  = \\i_tv80_core_mcycles_reg[2] ;
  assign \new_[2927]_  = ~\new_[3468]_  & (~\new_[3066]_  | ~\new_[6193]_ );
  assign \new_[2928]_  = \\i_tv80_core_RegAddrA_r_reg[1] ;
  assign \new_[2929]_  = \\i_tv80_core_mcycles_reg[1] ;
  assign \new_[2930]_  = \\i_tv80_core_RegAddrA_r_reg[2] ;
  assign \new_[2931]_  = ~\new_[5687]_  & (~\new_[5667]_  | ~\new_[3038]_ );
  assign \new_[2932]_  = (~\new_[3074]_  | ~\new_[6263]_ ) & (~\new_[6193]_  | ~\new_[6165]_ );
  assign \new_[2933]_  = ~\new_[4755]_  | ~\new_[3914]_  | ~\new_[2989]_  | ~\new_[4525]_ ;
  assign \new_[2934]_  = ~\new_[2990]_  & ~\new_[1624]_ ;
  assign \new_[2935]_  = ~\new_[2988]_  & (~\new_[4492]_  | ~\new_[6520]_ );
  assign \new_[2936]_  = (~\new_[3076]_  | ~\new_[6714]_ ) & (~\new_[2780]_  | ~\new_[1690]_ );
  assign \new_[2937]_  = ~\new_[6225]_  & (~\new_[3223]_  | ~\new_[3077]_ );
  assign \new_[2938]_  = ~\new_[6225]_  & (~\new_[3224]_  | ~\new_[3078]_ );
  assign \new_[2939]_  = ~\new_[6225]_  & (~\new_[3229]_  | ~\new_[3079]_ );
  assign \new_[2940]_  = ~\new_[6258]_  & (~\new_[3222]_  | ~\new_[3080]_ );
  assign \new_[2941]_  = ~\new_[1690]_  & (~\new_[3227]_  | ~\new_[3081]_ );
  assign \new_[2942]_  = ~\new_[6299]_  & (~\new_[3228]_  | ~\new_[3082]_ );
  assign \new_[2943]_  = \new_[4549]_  ? \new_[1623]_  : \new_[3083]_ ;
  assign \new_[2944]_  = ~\new_[2992]_ ;
  assign \new_[2945]_  = \new_[4509]_  ? \new_[5304]_  : \new_[3092]_ ;
  assign \new_[2946]_  = \new_[3386]_  ^ \new_[3089]_ ;
  assign \new_[2947]_  = ~\new_[3044]_  & ~\new_[7451]_ ;
  assign \new_[2948]_  = ~\new_[3047]_  & ~\new_[5724]_ ;
  assign \new_[2949]_  = ~\new_[2999]_ ;
  assign \new_[2950]_  = ~\new_[3000]_ ;
  assign \new_[2951]_  = ~\new_[3009]_ ;
  assign \new_[2952]_  = ~\new_[7544]_ ;
  assign \new_[2953]_  = ~\new_[3048]_  & (~\new_[3925]_  | ~\new_[1242]_ );
  assign \new_[2954]_  = ~\new_[7450]_ ;
  assign \new_[2955]_  = ~\new_[6821]_ ;
  assign \new_[2956]_  = \new_[3936]_  ? \new_[3112]_  : \new_[3932]_ ;
  assign \new_[2957]_  = \new_[3937]_  ? \new_[3112]_  : \new_[3938]_ ;
  assign \new_[2958]_  = \new_[3939]_  ? \new_[3112]_  : \new_[3940]_ ;
  assign \new_[2959]_  = \new_[3945]_  ? \new_[3112]_  : \new_[3935]_ ;
  assign \new_[2960]_  = \new_[4013]_  ? \new_[3112]_  : \new_[3942]_ ;
  assign \new_[2961]_  = \new_[3943]_  ? \new_[3112]_  : \new_[3944]_ ;
  assign \new_[2962]_  = \new_[3933]_  ? \new_[3112]_  : \new_[6747]_ ;
  assign \new_[2963]_  = \new_[3941]_  ? \new_[3112]_  : \new_[3934]_ ;
  assign \new_[2964]_  = ~\new_[3064]_  & ~\new_[3111]_ ;
  assign \new_[2965]_  = ~\new_[3160]_  | ~\new_[3064]_  | ~\new_[3383]_ ;
  assign \new_[2966]_  = ~\new_[3055]_  & (~\new_[3925]_  | ~\new_[1225]_ );
  assign \new_[2967]_  = \new_[3794]_  ^ \new_[3114]_ ;
  assign \new_[2968]_  = \new_[3802]_  ^ \new_[3113]_ ;
  assign \new_[2969]_  = ~\new_[3020]_ ;
  assign \new_[2970]_  = ~\new_[3021]_ ;
  assign \new_[2971]_  = ~\new_[3925]_  & ~\new_[3057]_ ;
  assign \new_[2972]_  = ~\new_[3057]_  & ~\new_[4316]_ ;
  assign n1629 = ~\new_[3059]_  & ~\new_[6623]_ ;
  assign \new_[2974]_  = ~\new_[3058]_  | ~\new_[7209]_ ;
  assign \new_[2975]_  = ~\new_[3058]_  | ~\new_[3165]_ ;
  assign \new_[2976]_  = \\i_tv80_core_RegAddrA_r_reg[0] ;
  assign \new_[2977]_  = ~\new_[3026]_ ;
  assign n1624 = ~\new_[6363]_  | ~\new_[7209]_  | ~\new_[3119]_ ;
  assign \new_[2979]_  = ~\new_[3065]_  | (~\new_[3542]_  & ~\new_[5247]_ );
  assign \new_[2980]_  = ~\new_[3067]_  | (~\new_[3331]_  & ~\new_[5247]_ );
  assign \new_[2981]_  = ~\new_[3040]_  | (~\new_[3467]_  & ~\new_[5247]_ );
  assign \new_[2982]_  = ~\new_[3070]_  & ~\new_[6299]_ ;
  assign \new_[2983]_  = ~\new_[3073]_  & ~\new_[6299]_ ;
  assign \new_[2984]_  = ~\new_[3071]_  | (~\new_[3352]_  & ~\new_[5247]_ );
  assign \new_[2985]_  = ~\new_[3072]_  | (~\new_[3472]_  & ~\new_[5247]_ );
  assign \new_[2986]_  = ~\new_[3035]_  & (~\new_[5772]_  | ~\new_[6258]_ );
  assign \new_[2987]_  = ~\new_[3036]_  & (~\new_[6084]_  | ~\new_[6258]_ );
  assign \new_[2988]_  = ~\new_[3745]_  | (~\new_[3142]_  & ~\new_[1624]_ );
  assign \new_[2989]_  = (~\new_[6873]_  | ~\new_[6589]_ ) & (~\new_[4831]_  | ~\new_[6040]_ );
  assign \new_[2990]_  = (~\new_[6873]_  | ~\new_[6655]_ ) & (~\new_[3841]_  | ~\new_[844]_ );
  assign \new_[2991]_  = \new_[5133]_  ? \new_[6874]_  : \new_[5014]_ ;
  assign \new_[2992]_  = ~\new_[3084]_  & ~\new_[6825]_ ;
  assign \new_[2993]_  = ~\new_[3885]_  | ~\new_[3884]_  | ~\new_[3090]_  | ~\new_[3877]_ ;
  assign \new_[2994]_  = ~\new_[6723]_  & (~\new_[3424]_  | ~\new_[3146]_ );
  assign \new_[2995]_  = ~\new_[3092]_  | ~\new_[3509]_ ;
  assign \new_[2996]_  = ~\new_[3091]_  & ~\new_[3618]_ ;
  assign \new_[2997]_  = ~\new_[3292]_  & (~\new_[3144]_  | ~\new_[3377]_ );
  assign \new_[2998]_  = ~\new_[3041]_ ;
  assign \new_[2999]_  = ~\new_[3385]_  & (~\new_[3145]_  | ~\new_[3379]_ );
  assign \new_[3000]_  = ~\new_[3086]_  & (~\new_[2034]_  | ~\new_[6712]_ );
  assign \new_[3001]_  = \new_[4414]_  ? \new_[5304]_  : \new_[3151]_ ;
  assign \new_[3002]_  = \\i_tv80_core_XY_State_reg[0] ;
  assign \new_[3003]_  = ~\new_[3085]_  & (~\new_[6723]_  | ~\new_[742]_ );
  assign \new_[3004]_  = \new_[3567]_  ^ \new_[3144]_ ;
  assign \new_[3005]_  = \new_[3512]_  ^ \new_[3150]_ ;
  assign \new_[3006]_  = ~\new_[3515]_  | ~\new_[3094]_  | ~\new_[3388]_ ;
  assign \new_[3007]_  = ~\new_[3096]_  & ~\new_[7335]_ ;
  assign \new_[3008]_  = ~\new_[7448]_ ;
  assign \new_[3009]_  = ~\new_[3044]_ ;
  assign \new_[3010]_  = ~\new_[3093]_  & (~\new_[1239]_  | ~\new_[5746]_ );
  assign n1649 = \new_[2930]_  ? \new_[6326]_  : \new_[3154]_ ;
  assign n1644 = ~\new_[3107]_  & ~\new_[6623]_ ;
  assign n1639 = ~\new_[3108]_  | ~\new_[3303]_ ;
  assign \new_[3014]_  = \new_[3109]_  | \new_[6711]_ ;
  assign \new_[3015]_  = ~\new_[7451]_ ;
  assign \new_[3016]_  = ~\new_[7451]_ ;
  assign \new_[3017]_  = ~\new_[7451]_ ;
  assign \new_[3018]_  = ~\new_[3381]_  | ~\new_[3715]_  | ~\new_[3162]_ ;
  assign \new_[3019]_  = ~\new_[3052]_ ;
  assign \new_[3020]_  = \new_[2006]_  ? \new_[4760]_  : \new_[3167]_ ;
  assign \new_[3021]_  = \new_[3383]_  & \new_[3203]_ ;
  assign \new_[3022]_  = ~\new_[3760]_  | ~\new_[3113]_  | ~\new_[3793]_ ;
  assign \new_[3023]_  = ~\new_[3115]_  & ~\new_[5724]_ ;
  assign n1634 = ~\new_[6297]_  | (~\new_[3163]_  & ~\new_[6412]_ );
  assign \new_[3025]_  = ~\new_[3118]_  | ~\new_[4864]_ ;
  assign \new_[3026]_  = \new_[2003]_  ? \new_[4760]_  : \new_[3171]_ ;
  assign \new_[3027]_  = ~\new_[3064]_ ;
  assign \new_[3028]_  = (~\new_[3168]_  | ~\new_[6132]_ ) & (~\new_[2826]_  | ~\new_[6225]_ );
  assign \new_[3029]_  = \\i_tv80_core_XY_State_reg[1] ;
  assign \new_[3030]_  = ~\new_[3121]_  | ~\new_[3551]_ ;
  assign \new_[3031]_  = ~\new_[4738]_  | ~\new_[5636]_  | ~\new_[3120]_  | ~\new_[4596]_ ;
  assign \new_[3032]_  = ~\new_[3233]_  | ~\new_[3348]_  | ~\new_[3185]_  | ~\new_[3122]_ ;
  assign \new_[3033]_  = ~\new_[3123]_  | (~\new_[1647]_  & ~\new_[5184]_ );
  assign \new_[3034]_  = ~\new_[3123]_  | (~\new_[1909]_  & ~\new_[5184]_ );
  assign \new_[3035]_  = ~\new_[6258]_  & (~\new_[3225]_  | ~\new_[3178]_ );
  assign \new_[3036]_  = ~\new_[6258]_  & (~\new_[3226]_  | ~\new_[3179]_ );
  assign \new_[3037]_  = ~\new_[3230]_  | ~\new_[6163]_ ;
  assign \new_[3038]_  = (~\new_[3187]_  | ~\new_[5783]_ ) & (~\new_[5959]_  | ~\new_[6521]_ );
  assign \new_[3039]_  = ~\new_[3400]_  & ~\new_[6873]_ ;
  assign \new_[3040]_  = ~\new_[3169]_  | ~\new_[6047]_ ;
  assign \new_[3041]_  = ~\new_[3390]_  & (~\new_[3188]_  | ~\new_[3380]_ );
  assign \new_[3042]_  = ~\new_[3388]_  | ~\new_[3377]_  | ~\new_[3144]_  | ~\new_[3312]_ ;
  assign \new_[3043]_  = ~\new_[3151]_  | ~\new_[3509]_ ;
  assign \new_[3044]_  = \new_[7449]_ ;
  assign \new_[3045]_  = ~\new_[3149]_  | ~\new_[3436]_ ;
  assign \new_[3046]_  = ~\new_[3090]_ ;
  assign \new_[3047]_  = ~\new_[3147]_  & (~\new_[3925]_  | ~\new_[1241]_ );
  assign \new_[3048]_  = ~\new_[3925]_  & ~\new_[3153]_ ;
  assign \new_[3049]_  = ~\new_[3153]_  & ~\new_[4316]_ ;
  assign n1654 = ~\new_[3210]_  | ~\new_[3158]_ ;
  assign \new_[3051]_  = ~\new_[3106]_ ;
  assign \new_[3052]_  = ~\new_[3456]_  | ~\new_[3156]_ ;
  assign \new_[3053]_  = ~\new_[3205]_  | ~\new_[3594]_  | ~\new_[3255]_ ;
  assign \new_[3054]_  = ~\new_[3159]_  | (~\new_[3250]_  & ~\new_[3384]_ );
  assign \new_[3055]_  = ~\new_[3925]_  & ~\new_[3161]_ ;
  assign \new_[3056]_  = ~\new_[3161]_  & ~\new_[4316]_ ;
  assign \new_[3057]_  = \new_[3796]_  ^ \new_[3316]_ ;
  assign \new_[3058]_  = ~\new_[5844]_  | ~\new_[3810]_  | ~\new_[3212]_ ;
  assign \new_[3059]_  = ~\new_[3164]_  & (~\new_[2863]_  | ~\new_[6338]_ );
  assign \new_[3060]_  = ~\new_[3825]_  | ~\new_[3165]_ ;
  assign \new_[3061]_  = ~\new_[4371]_  & ~\new_[3165]_ ;
  assign \new_[3062]_  = ~\new_[3903]_  | ~\new_[3165]_ ;
  assign \new_[3063]_  = ~\new_[3521]_  & (~\new_[3215]_  | ~\new_[5459]_ );
  assign \new_[3064]_  = ~\new_[3166]_  & (~\new_[5676]_  | ~\new_[6227]_ );
  assign \new_[3065]_  = ~\new_[3125]_  | ~\new_[6047]_ ;
  assign \new_[3066]_  = ~\new_[3274]_  | ~\new_[5193]_  | ~\new_[4527]_  | ~\new_[3608]_ ;
  assign \new_[3067]_  = ~\new_[3170]_  | ~\new_[6047]_ ;
  assign \new_[3068]_  = ~\new_[5969]_  | (~\new_[3175]_  & ~\new_[4032]_ );
  assign \new_[3069]_  = ~\new_[5969]_  | (~\new_[3174]_  & ~\new_[4070]_ );
  assign \new_[3070]_  = (~\new_[3218]_  | ~\new_[6047]_ ) & (~\new_[3485]_  | ~\new_[5183]_ );
  assign \new_[3071]_  = ~\new_[3172]_  | ~\new_[6047]_ ;
  assign \new_[3072]_  = ~\new_[3173]_  | ~\new_[6047]_ ;
  assign \new_[3073]_  = (~\new_[3176]_  | ~\new_[6047]_ ) & (~\new_[3496]_  | ~\new_[5183]_ );
  assign \new_[3074]_  = ~\new_[3232]_  | ~\new_[3349]_  | ~\new_[3184]_  | ~\new_[3177]_ ;
  assign n1664 = ~\new_[3214]_  & ~\new_[6417]_ ;
  assign \new_[3076]_  = ~\new_[3182]_  | (~\new_[3981]_  & ~\new_[3360]_ );
  assign \new_[3077]_  = (~\new_[5176]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[6113]_ );
  assign \new_[3078]_  = (~\new_[5177]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[6227]_ );
  assign \new_[3079]_  = (~\new_[5174]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[7549]_ );
  assign \new_[3080]_  = (~\new_[5053]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[6128]_ );
  assign \new_[3081]_  = (~\new_[5175]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[6152]_ );
  assign \new_[3082]_  = (~\new_[5178]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[6120]_ );
  assign \new_[3083]_  = ~\new_[5368]_  | ~\new_[3320]_  | ~\new_[3669]_  | ~\new_[4693]_ ;
  assign \new_[3084]_  = ~\new_[5052]_  & (~\new_[3238]_  | ~\new_[6041]_ );
  assign \new_[3085]_  = ~\new_[6723]_  & (~\new_[3372]_  | ~\new_[3243]_ );
  assign \new_[3086]_  = ~\new_[3190]_  & ~\new_[3618]_ ;
  assign \new_[3087]_  = ~\new_[4282]_  & (~\new_[3240]_  | ~\new_[5641]_ );
  assign \new_[3088]_  = ~\new_[6364]_  & ~\new_[3189]_ ;
  assign \new_[3089]_  = ~\new_[3239]_  & (~\new_[3242]_  | ~\new_[3376]_ );
  assign \new_[3090]_  = ~\new_[3713]_  | (~\new_[3244]_  & ~\new_[3873]_ );
  assign \new_[3091]_  = (~\new_[4704]_  | ~\new_[1925]_ ) & (~\new_[3245]_  | ~\new_[5304]_ );
  assign \new_[3092]_  = \new_[3511]_  ^ \new_[3242]_ ;
  assign \new_[3093]_  = ~\new_[3194]_  & ~\new_[5724]_ ;
  assign \new_[3094]_  = ~\new_[3150]_ ;
  assign \new_[3095]_  = ~\new_[3528]_  | (~\new_[3247]_  & ~\new_[3393]_ );
  assign \new_[3096]_  = ~\new_[3191]_  & (~\new_[6723]_  | ~\new_[794]_ );
  assign \new_[3097]_  = ~\new_[3197]_  | ~\new_[853]_ ;
  assign \new_[3098]_  = ~\new_[3197]_  | ~\new_[851]_ ;
  assign \new_[3099]_  = ~\new_[3197]_  | ~\new_[852]_ ;
  assign \new_[3100]_  = ~\new_[3197]_  | ~\new_[849]_ ;
  assign \new_[3101]_  = ~\new_[3197]_  | ~\new_[684]_ ;
  assign \new_[3102]_  = ~\new_[3197]_  | ~\new_[845]_ ;
  assign \new_[3103]_  = ~\new_[3197]_  | ~\new_[799]_ ;
  assign \new_[3104]_  = ~\new_[3197]_  | ~\new_[848]_ ;
  assign \new_[3105]_  = \new_[3197]_  | \new_[3196]_ ;
  assign \new_[3106]_  = ~\new_[3456]_  & ~\new_[3195]_ ;
  assign \new_[3107]_  = ~\new_[3201]_  & (~\new_[2929]_  | ~\new_[6338]_ );
  assign \new_[3108]_  = ~\new_[3200]_  & (~\new_[2928]_  | ~\new_[6252]_ );
  assign \new_[3109]_  = ~\new_[3199]_  & (~\new_[1237]_  | ~\new_[5746]_ );
  assign \new_[3110]_  = \new_[3204]_  | \new_[6711]_ ;
  assign \new_[3111]_  = \new_[3383]_  | \new_[3203]_ ;
  assign \new_[3112]_  = ~\new_[3202]_  & (~\new_[5676]_  | ~\new_[6113]_ );
  assign \new_[3113]_  = ~\new_[3206]_  | ~\new_[3588]_ ;
  assign \new_[3114]_  = ~\new_[3589]_  | (~\new_[3256]_  & ~\new_[3643]_ );
  assign \new_[3115]_  = ~\new_[3207]_  & (~\new_[3925]_  | ~\new_[1238]_ );
  assign n1659 = ~\new_[3213]_  & ~\new_[6441]_ ;
  assign \new_[3117]_  = ~\new_[3327]_  | ~\new_[4406]_  | ~\new_[4583]_  | ~\new_[3992]_ ;
  assign \new_[3118]_  = \new_[4560]_  ? \new_[3276]_  : \new_[3325]_ ;
  assign \new_[3119]_  = ~\new_[3165]_ ;
  assign \new_[3120]_  = ~\new_[3658]_  & ~\new_[3217]_ ;
  assign \new_[3121]_  = ~\new_[3216]_  & (~\new_[5607]_  | ~\new_[5772]_ );
  assign \new_[3122]_  = ~\new_[6711]_  | ~\new_[5962]_  | ~\new_[4095]_ ;
  assign \new_[3123]_  = ~\new_[3434]_  | ~\new_[3230]_ ;
  assign \new_[3124]_  = ~\new_[5266]_  | ~\new_[6712]_ ;
  assign \new_[3125]_  = ~\new_[3272]_  & ~\new_[5486]_ ;
  assign \new_[3126]_  = ~\new_[3231]_  & (~\new_[6552]_  | ~\new_[5295]_ );
  assign \new_[3127]_  = ~\new_[5317]_  | ~\new_[6712]_ ;
  assign \new_[3128]_  = ~\new_[5290]_  | ~\new_[6712]_ ;
  assign \new_[3129]_  = ~\new_[5254]_  | ~\new_[6712]_ ;
  assign \new_[3130]_  = ~\new_[5321]_  | ~\new_[6712]_ ;
  assign \new_[3131]_  = ~\new_[5324]_  | ~\new_[6712]_ ;
  assign \new_[3132]_  = ~\new_[5323]_  | ~\new_[6712]_ ;
  assign \new_[3133]_  = ~\new_[5325]_  | ~\new_[6712]_ ;
  assign \new_[3134]_  = ~\new_[5329]_  | ~\new_[6712]_ ;
  assign \new_[3135]_  = ~\new_[5251]_  | ~\new_[6712]_ ;
  assign \new_[3136]_  = ~\new_[5322]_  | ~\new_[6712]_ ;
  assign \new_[3137]_  = ~\new_[5316]_  | ~\new_[6712]_ ;
  assign \new_[3138]_  = ~\new_[5328]_  | ~\new_[6712]_ ;
  assign \new_[3139]_  = ~\new_[5319]_  | ~\new_[6712]_ ;
  assign \new_[3140]_  = ~\new_[5320]_  | ~\new_[6712]_ ;
  assign \new_[3141]_  = ~\new_[5252]_  | ~\new_[6712]_ ;
  assign \new_[3142]_  = ~\new_[3236]_  & (~\new_[7289]_  | ~\new_[6952]_ );
  assign \new_[3143]_  = ~\new_[3444]_  | ~\new_[3376]_  | ~\new_[3242]_  | ~\new_[3569]_ ;
  assign \new_[3144]_  = ~\new_[3301]_  | ~\new_[3507]_  | ~\new_[3300]_ ;
  assign \new_[3145]_  = ~\new_[3239]_  | ~\new_[3569]_ ;
  assign \new_[3146]_  = ~\new_[3245]_  | ~\new_[3509]_ ;
  assign \new_[3147]_  = ~\new_[3925]_  & ~\new_[3246]_ ;
  assign \new_[3148]_  = ~\new_[3246]_  & ~\new_[4316]_ ;
  assign \new_[3149]_  = ~\new_[3242]_  | ~\new_[3517]_ ;
  assign \new_[3150]_  = ~\new_[3291]_  & (~\new_[3298]_  | ~\new_[3375]_ );
  assign \new_[3151]_  = \new_[3514]_  ^ \new_[3298]_ ;
  assign \new_[3152]_  = ~\new_[3307]_  | ~\new_[3761]_  | ~\new_[4041]_ ;
  assign \new_[3153]_  = \new_[3874]_  ^ \new_[3302]_ ;
  assign \new_[3154]_  = \new_[3029]_  ? \new_[3308]_  : \new_[2780]_ ;
  assign \new_[3155]_  = \new_[3412]_  ^ \new_[3323]_ ;
  assign \new_[3156]_  = ~\new_[3195]_ ;
  assign \new_[3157]_  = ~\new_[3198]_ ;
  assign \new_[3158]_  = ~\new_[3200]_ ;
  assign \new_[3159]_  = ~\new_[3252]_  | (~\new_[5591]_  & ~\new_[3450]_ );
  assign \new_[3160]_  = ~\new_[3203]_ ;
  assign \new_[3161]_  = \new_[3805]_  ^ \new_[3317]_ ;
  assign \new_[3162]_  = ~\new_[3258]_  | ~\new_[3877]_ ;
  assign \new_[3163]_  = ~\new_[4276]_  & (~\new_[3278]_  | ~\new_[6348]_ );
  assign \new_[3164]_  = ~\new_[6252]_  & (~\new_[3324]_  | ~\new_[4861]_ );
  assign \new_[3165]_  = \new_[3221]_  | \new_[6365]_ ;
  assign \new_[3166]_  = ~\new_[5676]_  & (~\new_[3326]_  | ~\new_[5706]_ );
  assign \new_[3167]_  = \new_[4559]_  ? \new_[1623]_  : \new_[3328]_ ;
  assign \new_[3168]_  = \new_[3538]_  ? \new_[6711]_  : \new_[4880]_ ;
  assign \new_[3169]_  = ~\new_[3273]_  & ~\new_[5486]_ ;
  assign \new_[3170]_  = ~\new_[3275]_  & ~\new_[5486]_ ;
  assign \new_[3171]_  = \new_[4558]_  ? \new_[1623]_  : \new_[3277]_ ;
  assign \new_[3172]_  = ~\new_[3220]_  & ~\new_[5486]_ ;
  assign \new_[3173]_  = ~\new_[3219]_  & ~\new_[5486]_ ;
  assign \new_[3174]_  = ~\new_[4366]_  | ~\new_[3905]_  | ~\new_[4266]_  | ~\new_[3351]_ ;
  assign \new_[3175]_  = ~\new_[4528]_  | ~\new_[3418]_  | ~\new_[4332]_  | ~\new_[3830]_ ;
  assign \new_[3176]_  = ~\new_[3283]_  & ~\new_[5486]_ ;
  assign \new_[3177]_  = ~\new_[5962]_  | ~\new_[6193]_  | ~\new_[4273]_  | ~\new_[6711]_ ;
  assign \new_[3178]_  = (~\new_[5054]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[5772]_ );
  assign \new_[3179]_  = (~\new_[5051]_  | ~\new_[6712]_ ) & (~\new_[5724]_  | ~\new_[6084]_ );
  assign \new_[3180]_  = ~\new_[3230]_ ;
  assign \new_[3181]_  = ~\new_[6711]_  & ~\new_[6438]_ ;
  assign \new_[3182]_  = ~\new_[6712]_  | ~\new_[2780]_ ;
  assign \new_[3183]_  = \new_[6342]_  & \new_[6711]_ ;
  assign \new_[3184]_  = ~\new_[6193]_  | ~\new_[6711]_  | ~\new_[5641]_ ;
  assign \new_[3185]_  = ~\new_[2660]_  | ~\new_[6711]_  | ~\new_[5641]_ ;
  assign \new_[3186]_  = ~\new_[3289]_  & (~\new_[6576]_  | ~\new_[5295]_ );
  assign \new_[3187]_  = \new_[7295]_  ^ \new_[7289]_ ;
  assign \new_[3188]_  = ~\new_[3292]_  | ~\new_[3388]_ ;
  assign \new_[3189]_  = ~\new_[4059]_  | ~\new_[3293]_ ;
  assign \new_[3190]_  = (~\new_[4704]_  | ~\new_[2034]_ ) & (~\new_[3366]_  | ~\new_[5304]_ );
  assign \new_[3191]_  = ~\new_[6723]_  & (~\new_[3427]_  | ~\new_[3374]_ );
  assign \new_[3192]_  = ~\new_[3295]_  | (~\new_[1860]_  & ~\new_[5184]_ );
  assign \new_[3193]_  = ~\new_[3294]_  | ~\new_[3363]_ ;
  assign \new_[3194]_  = ~\new_[3296]_  & (~\new_[3925]_  | ~\new_[1239]_ );
  assign \new_[3195]_  = \new_[4041]_  | \new_[3309]_ ;
  assign \new_[3196]_  = \new_[4082]_  & \new_[3309]_ ;
  assign \new_[3197]_  = \new_[3306]_  & \new_[3456]_ ;
  assign \new_[3198]_  = \new_[3307]_  & \new_[3469]_ ;
  assign \new_[3199]_  = ~\new_[3310]_  & ~\new_[5724]_ ;
  assign \new_[3200]_  = ~\new_[3308]_  & ~\new_[6347]_ ;
  assign \new_[3201]_  = ~\new_[6225]_  & (~\new_[3392]_  | ~\new_[4380]_ );
  assign \new_[3202]_  = ~\new_[5676]_  & (~\new_[3396]_  | ~\new_[5780]_ );
  assign \new_[3203]_  = (~\new_[3394]_  | ~\new_[6216]_ ) & (~\new_[5676]_  | ~\new_[7549]_ );
  assign \new_[3204]_  = ~\new_[3311]_  & (~\new_[1236]_  | ~\new_[5746]_ );
  assign \new_[3205]_  = ~\new_[3876]_  | ~\new_[3710]_  | ~\new_[3316]_  | ~\new_[3793]_ ;
  assign \new_[3206]_  = ~\new_[3880]_  | ~\new_[3317]_  | ~\new_[3876]_ ;
  assign \new_[3207]_  = ~\new_[3925]_  & ~\new_[3319]_ ;
  assign \new_[3208]_  = ~\new_[3319]_  & ~\new_[4316]_ ;
  assign \new_[3209]_  = ~\new_[3393]_  & ~\new_[3449]_ ;
  assign \new_[3210]_  = ~\new_[3290]_  & (~\new_[2976]_  | ~\new_[6252]_ );
  assign \new_[3211]_  = ~\new_[3322]_  | ~\new_[5969]_ ;
  assign \new_[3212]_  = ~\new_[3284]_  & (~\new_[6730]_  | ~\new_[5188]_ );
  assign \new_[3213]_  = (~\new_[3404]_  | ~\new_[6388]_ ) & (~\new_[3002]_  | ~\new_[6347]_ );
  assign \new_[3214]_  = (~\new_[3403]_  | ~\new_[6129]_ ) & (~\new_[3029]_  | ~\new_[6165]_ );
  assign \new_[3215]_  = \new_[3667]_  ^ \new_[3350]_ ;
  assign \new_[3216]_  = ~\new_[4269]_  | ~\new_[3414]_  | ~\new_[4402]_  | ~\new_[4084]_ ;
  assign \new_[3217]_  = ~\new_[4510]_  | ~\new_[3413]_  | ~\new_[3494]_  | ~\new_[6016]_ ;
  assign \new_[3218]_  = ~\new_[3279]_  & ~\new_[5486]_ ;
  assign \new_[3219]_  = (~\new_[763]_  | ~\new_[4538]_ ) & (~\new_[3415]_  | ~\new_[4428]_ );
  assign \new_[3220]_  = (~\new_[761]_  | ~\new_[4538]_ ) & (~\new_[3416]_  | ~\new_[4428]_ );
  assign \new_[3221]_  = ~\new_[3284]_ ;
  assign \new_[3222]_  = ~\new_[4285]_  | ~\new_[3356]_ ;
  assign \new_[3223]_  = ~\new_[4630]_  | ~\new_[3356]_ ;
  assign \new_[3224]_  = ~\new_[5149]_  | ~\new_[3356]_ ;
  assign \new_[3225]_  = ~\new_[4286]_  | ~\new_[3356]_ ;
  assign \new_[3226]_  = ~\new_[4568]_  | ~\new_[3356]_ ;
  assign \new_[3227]_  = ~\new_[5326]_  | ~\new_[3356]_ ;
  assign \new_[3228]_  = ~\new_[5327]_  | ~\new_[3356]_ ;
  assign \new_[3229]_  = ~\new_[4750]_  | ~\new_[3356]_ ;
  assign \new_[3230]_  = \new_[2005]_  ? \new_[4760]_  : \new_[3420]_ ;
  assign \new_[3231]_  = ~\new_[3286]_ ;
  assign \new_[3232]_  = ~\new_[6193]_  | ~\new_[6712]_  | ~\new_[5724]_ ;
  assign \new_[3233]_  = ~\new_[2660]_  | ~\new_[6712]_  | ~\new_[5724]_ ;
  assign \new_[3234]_  = ~\new_[6711]_ ;
  assign \new_[3235]_  = ~\new_[3289]_ ;
  assign \new_[3236]_  = ~\new_[7289]_  & ~\new_[5842]_ ;
  assign \new_[3237]_  = ~\new_[4282]_  & (~\new_[3422]_  | ~\new_[5641]_ );
  assign \new_[3238]_  = ~\new_[4319]_  | ~\new_[3423]_  | ~\new_[4212]_ ;
  assign \new_[3239]_  = ~\new_[3506]_  | (~\new_[3436]_  & ~\new_[3568]_ );
  assign \new_[3240]_  = ~\new_[4033]_  | ~\new_[3364]_ ;
  assign \new_[3241]_  = ~\new_[7265]_ ;
  assign \new_[3242]_  = ~\new_[3365]_  | ~\new_[3505]_ ;
  assign \new_[3243]_  = ~\new_[3366]_  | ~\new_[3509]_ ;
  assign \new_[3244]_  = ~\new_[3780]_  & (~\new_[3441]_  | ~\new_[3872]_ );
  assign \new_[3245]_  = \new_[3504]_  ^ \new_[3443]_ ;
  assign \new_[3246]_  = \new_[3804]_  ^ \new_[3441]_ ;
  assign \new_[3247]_  = ~\new_[3378]_  & ~\new_[3449]_ ;
  assign \new_[3248]_  = ~\new_[3373]_  | ~\new_[3849]_ ;
  assign \new_[3249]_  = ~\new_[3390]_  & ~\new_[3384]_ ;
  assign \new_[3250]_  = ~\new_[3393]_  & (~\new_[3526]_  | ~\new_[3573]_ );
  assign \new_[3251]_  = \\i_tv80_core_Fp_reg[5] ;
  assign \new_[3252]_  = (~\new_[3636]_  | ~\new_[3527]_ ) & (~\new_[3451]_  | ~\new_[3452]_ );
  assign \new_[3253]_  = \new_[3527]_  & \new_[3528]_ ;
  assign \new_[3254]_  = \\i_tv80_core_Ap_reg[3] ;
  assign \new_[3255]_  = ~\new_[3793]_  | (~\new_[3455]_  & ~\new_[3784]_ );
  assign \new_[3256]_  = ~\new_[3316]_ ;
  assign \new_[3257]_  = \\i_tv80_core_Ap_reg[5] ;
  assign \new_[3258]_  = ~\new_[3713]_  | (~\new_[3458]_  & ~\new_[3873]_ );
  assign \new_[3259]_  = \\i_tv80_core_Fp_reg[7] ;
  assign \new_[3260]_  = \\i_tv80_core_Ap_reg[1] ;
  assign \new_[3261]_  = \\i_tv80_core_Fp_reg[1] ;
  assign \new_[3262]_  = \\i_tv80_core_Fp_reg[3] ;
  assign \new_[3263]_  = \\i_tv80_core_Fp_reg[0] ;
  assign \new_[3264]_  = \\i_tv80_core_Fp_reg[2] ;
  assign \new_[3265]_  = \\i_tv80_core_Fp_reg[4] ;
  assign \new_[3266]_  = \\i_tv80_core_Fp_reg[6] ;
  assign \new_[3267]_  = \\i_tv80_core_Ap_reg[0] ;
  assign \new_[3268]_  = \\i_tv80_core_Ap_reg[2] ;
  assign \new_[3269]_  = \\i_tv80_core_Ap_reg[4] ;
  assign \new_[3270]_  = \\i_tv80_core_Ap_reg[6] ;
  assign \new_[3271]_  = \\i_tv80_core_Ap_reg[7] ;
  assign \new_[3272]_  = (~\new_[760]_  | ~\new_[4538]_ ) & (~\new_[3466]_  | ~\new_[4428]_ );
  assign \new_[3273]_  = (~\new_[759]_  | ~\new_[4538]_ ) & (~\new_[3408]_  | ~\new_[4428]_ );
  assign \new_[3274]_  = ~\new_[3406]_  & (~\new_[6961]_  | ~\new_[6128]_ );
  assign \new_[3275]_  = (~\new_[758]_  | ~\new_[4538]_ ) & (~\new_[3410]_  | ~\new_[4428]_ );
  assign \new_[3276]_  = ~\new_[3330]_  & (~\new_[4354]_  | ~\new_[6193]_ );
  assign \new_[3277]_  = ~\new_[4637]_  | ~\new_[3553]_  | ~\new_[4642]_  | ~\new_[4355]_ ;
  assign \new_[3278]_  = ~\new_[3540]_  | ~\new_[3899]_  | ~\new_[3886]_ ;
  assign \new_[3279]_  = (~\new_[736]_  | ~\new_[4538]_ ) & (~\new_[3485]_  | ~\new_[4428]_ );
  assign \new_[3280]_  = ~\new_[5125]_  & (~\new_[3537]_  | ~\new_[3592]_ );
  assign \new_[3281]_  = \\i_tv80_core_IStatus_reg[1] ;
  assign \new_[3282]_  = ~\new_[5995]_  & (~\new_[3495]_  | ~\new_[3737]_ );
  assign \new_[3283]_  = (~\new_[762]_  | ~\new_[4538]_ ) & (~\new_[3496]_  | ~\new_[4428]_ );
  assign \new_[3284]_  = ~\new_[4368]_  | ~\new_[3463]_ ;
  assign \new_[3285]_  = \\i_tv80_core_R_reg[7] ;
  assign \new_[3286]_  = ~\new_[3434]_  | ~\new_[3502]_ ;
  assign \new_[3287]_  = ~\new_[6711]_ ;
  assign \new_[3288]_  = ~\new_[6711]_ ;
  assign \new_[3289]_  = \new_[3434]_  & \new_[3672]_ ;
  assign \new_[3290]_  = ~\new_[3361]_ ;
  assign \new_[3291]_  = ~\new_[3508]_  | (~\new_[3507]_  & ~\new_[3520]_ );
  assign \new_[3292]_  = ~\new_[3440]_  | (~\new_[3508]_  & ~\new_[3565]_ );
  assign \new_[3293]_  = ~\new_[6313]_  | (~\new_[7018]_  & ~\new_[6998]_ );
  assign \new_[3294]_  = ~\new_[3433]_  | ~\new_[4910]_ ;
  assign \new_[3295]_  = ~\new_[3434]_  | ~\new_[3919]_ ;
  assign \new_[3296]_  = ~\new_[3925]_  & ~\new_[3442]_ ;
  assign \new_[3297]_  = ~\new_[3442]_  & ~\new_[4316]_ ;
  assign \new_[3298]_  = ~\new_[3435]_  | ~\new_[3438]_ ;
  assign \new_[3299]_  = \new_[3440]_  | \new_[3447]_ ;
  assign \new_[3300]_  = \new_[3438]_  | \new_[3566]_ ;
  assign \new_[3301]_  = ~\new_[3678]_  | ~\new_[3627]_  | ~\new_[3516]_ ;
  assign \new_[3302]_  = ~\new_[3458]_  | (~\new_[3634]_  & ~\new_[3593]_ );
  assign \new_[3303]_  = ~\new_[3448]_  | ~\new_[6314]_ ;
  assign \new_[3304]_  = ~\new_[6697]_ ;
  assign \new_[3305]_  = ~\new_[6697]_ ;
  assign \new_[3306]_  = ~\new_[3448]_  & ~\new_[3561]_ ;
  assign \new_[3307]_  = ~\new_[3456]_  & ~\new_[3448]_ ;
  assign \new_[3308]_  = ~\new_[6428]_  | ~\new_[3448]_  | ~\new_[3704]_ ;
  assign \new_[3309]_  = ~\new_[3448]_  | ~\new_[3761]_ ;
  assign \new_[3310]_  = ~\new_[3445]_  & (~\new_[3925]_  | ~\new_[1237]_ );
  assign \new_[3311]_  = ~\new_[3454]_  & ~\new_[5746]_ ;
  assign \new_[3312]_  = ~\new_[3390]_ ;
  assign \new_[3313]_  = \new_[3451]_  & \new_[3529]_ ;
  assign \new_[3314]_  = \new_[5146]_  ^ \new_[3636]_ ;
  assign \new_[3315]_  = ~\new_[3456]_  | ~\new_[6326]_ ;
  assign \new_[3316]_  = ~\new_[3457]_  | ~\new_[3714]_ ;
  assign \new_[3317]_  = ~\new_[3587]_  | (~\new_[3531]_  & ~\new_[3709]_ );
  assign \new_[3318]_  = ~\new_[3395]_ ;
  assign \new_[3319]_  = \new_[3879]_  ^ \new_[3531]_ ;
  assign \new_[3320]_  = ~\new_[5344]_  & (~\new_[3541]_  | ~\new_[6589]_ );
  assign \new_[3321]_  = \\i_tv80_core_IStatus_reg[0] ;
  assign \new_[3322]_  = ~\new_[4679]_  | ~\new_[4417]_  | ~\new_[3462]_  | ~\new_[4653]_ ;
  assign \new_[3323]_  = \new_[4769]_  ^ \new_[3541]_ ;
  assign \new_[3324]_  = (~\new_[3539]_  | ~\new_[5969]_ ) & (~\new_[4103]_  | ~\new_[6193]_ );
  assign \new_[3325]_  = ~\new_[3399]_ ;
  assign \new_[3326]_  = ~\new_[3464]_  & (~\new_[3897]_  | ~\new_[6193]_ );
  assign \new_[3327]_  = ~\new_[3411]_  | ~\new_[6589]_ ;
  assign \new_[3328]_  = ~\new_[4633]_  | ~\new_[3838]_  | ~\new_[3409]_  | ~\new_[4583]_ ;
  assign \new_[3329]_  = \new_[3407]_  & \new_[4116]_ ;
  assign \new_[3330]_  = ~\new_[6031]_  & (~\new_[3547]_  | ~\new_[4334]_ );
  assign \new_[3331]_  = ~\new_[3410]_ ;
  assign n1729 = ~\new_[3483]_  | ~\new_[6363]_ ;
  assign n1704 = ~\new_[3491]_  | ~reset_n;
  assign n1694 = ~\new_[3476]_  | ~reset_n;
  assign n1709 = ~\new_[3477]_  | ~reset_n;
  assign n1699 = ~\new_[3478]_  | ~reset_n;
  assign n1714 = ~\new_[3479]_  | ~reset_n;
  assign n1669 = ~\new_[3480]_  | ~reset_n;
  assign n1719 = ~\new_[3481]_  | ~reset_n;
  assign n1684 = ~\new_[3482]_  | ~\new_[6304]_ ;
  assign n1724 = ~\new_[3486]_  | ~\new_[6363]_ ;
  assign n1689 = ~\new_[3488]_  | ~\new_[6363]_ ;
  assign n1674 = ~\new_[3474]_  | ~\new_[6363]_ ;
  assign n1734 = ~\new_[3487]_  | ~\new_[6363]_ ;
  assign n1679 = ~\new_[3475]_  | ~\new_[6363]_ ;
  assign n1739 = ~\new_[3484]_  | ~\new_[6363]_ ;
  assign n1744 = ~\new_[3489]_  | ~reset_n;
  assign \new_[3348]_  = ~\new_[4194]_  | ~\new_[3471]_  | ~\new_[4427]_ ;
  assign \new_[3349]_  = ~\new_[4194]_  | ~\new_[3471]_  | ~\new_[4737]_ ;
  assign \new_[3350]_  = \new_[3993]_  ^ \new_[3552]_ ;
  assign \new_[3351]_  = ~\new_[3493]_  & (~\new_[5644]_  | ~\new_[5772]_ );
  assign \new_[3352]_  = ~\new_[3416]_ ;
  assign \new_[3353]_  = (~\new_[3559]_  | ~\new_[4413]_ ) & (~\new_[3613]_  | ~\new_[4339]_ );
  assign \new_[3354]_  = ~\new_[3502]_  | ~\new_[6163]_ ;
  assign \new_[3355]_  = ~\new_[742]_  | ~\new_[3620]_ ;
  assign \new_[3356]_  = ~\new_[6713]_  & ~\new_[5724]_ ;
  assign \new_[3357]_  = ~\new_[793]_  | ~\new_[3620]_ ;
  assign \new_[3358]_  = ~\new_[764]_  | ~\new_[6713]_ ;
  assign \new_[3359]_  = ~\new_[794]_  | ~\new_[6713]_ ;
  assign \new_[3360]_  = ~\new_[6711]_ ;
  assign \new_[3361]_  = ~\new_[3761]_  | ~\new_[6314]_ ;
  assign \new_[3362]_  = ~\new_[7266]_ ;
  assign \new_[3363]_  = ~\new_[6698]_  | ~\new_[6994]_ ;
  assign \new_[3364]_  = (~\new_[7255]_  | ~\new_[5969]_ ) & (~\new_[4139]_  | ~\new_[6471]_ );
  assign \new_[3365]_  = ~\new_[3678]_  | ~\new_[3504]_  | ~\new_[3677]_ ;
  assign \new_[3366]_  = \new_[5253]_  ^ \new_[3570]_ ;
  assign \new_[3367]_  = ~\new_[3563]_  | ~\new_[766]_ ;
  assign \new_[3368]_  = ~\new_[3563]_  | ~\new_[793]_ ;
  assign \new_[3369]_  = ~\new_[3563]_  | ~\new_[755]_ ;
  assign \new_[3370]_  = ~\new_[3563]_  | ~\new_[757]_ ;
  assign \new_[3371]_  = ~\new_[3563]_  | ~\new_[764]_ ;
  assign \new_[3372]_  = ~\new_[3563]_  | ~\new_[742]_ ;
  assign \new_[3373]_  = ~\new_[7267]_ ;
  assign \new_[3374]_  = ~\new_[5139]_  | ~\new_[3509]_ ;
  assign \new_[3375]_  = ~\new_[3566]_  & ~\new_[3520]_ ;
  assign \new_[3376]_  = \new_[3517]_  & \new_[3518]_ ;
  assign \new_[3377]_  = ~\new_[3520]_  & ~\new_[3565]_ ;
  assign \new_[3378]_  = ~\new_[3573]_  & (~\new_[3578]_  | ~\new_[3576]_ );
  assign \new_[3379]_  = ~\new_[3572]_  & (~\new_[3575]_  | ~\new_[3688]_ );
  assign \new_[3380]_  = ~\new_[3576]_  & (~\new_[3577]_  | ~\new_[3572]_ );
  assign \new_[3381]_  = ~\new_[3642]_  | ~\new_[3510]_  | ~\new_[3877]_ ;
  assign \new_[3382]_  = ~\new_[3688]_  | ~\new_[3522]_ ;
  assign \new_[3383]_  = ~\new_[5676]_  & (~\new_[3730]_  | ~\new_[3581]_ );
  assign \new_[3384]_  = ~\new_[3528]_  | ~\new_[3529]_ ;
  assign \new_[3385]_  = ~\new_[3444]_ ;
  assign \new_[3386]_  = ~\new_[3523]_  | ~\new_[3675]_ ;
  assign \new_[3387]_  = ~\new_[3576]_  & ~\new_[3524]_ ;
  assign \new_[3388]_  = ~\new_[3447]_ ;
  assign \new_[3389]_  = ~\new_[3525]_  & ~\new_[3573]_ ;
  assign \new_[3390]_  = ~\new_[3578]_  | ~\new_[3526]_ ;
  assign \new_[3391]_  = ~\new_[3530]_  & (~\new_[1293]_  | ~\new_[6271]_ );
  assign \new_[3392]_  = (~\new_[4657]_  | ~\new_[6039]_ ) & (~\new_[3584]_  | ~\new_[5969]_ );
  assign \new_[3393]_  = ~\new_[5256]_  & ~\new_[3636]_ ;
  assign \new_[3394]_  = ~\new_[5962]_  & (~\new_[3711]_  | ~\new_[3544]_ );
  assign \new_[3395]_  = ~\new_[5160]_  | ~\new_[3640]_  | ~\new_[5641]_  | ~\new_[4932]_ ;
  assign \new_[3396]_  = (~\new_[3564]_  | ~\new_[5969]_ ) & (~\new_[4045]_  | ~\new_[6193]_ );
  assign \new_[3397]_  = ~\new_[3532]_  | ~\new_[3885]_ ;
  assign rfsh_n = i_tv80_core_rfsh_n_reg;
  assign \new_[3399]_  = ~\new_[3535]_  & (~\new_[2429]_  | ~\new_[6712]_ );
  assign \new_[3400]_  = \new_[3541]_  | \new_[3605]_ ;
  assign \new_[3401]_  = \new_[6519]_  ? \new_[3720]_  : \new_[4096]_ ;
  assign \new_[3402]_  = ~\new_[3619]_  & ~\new_[3808]_ ;
  assign \new_[3403]_  = \new_[3029]_  ? \new_[3661]_  : \new_[3731]_ ;
  assign \new_[3404]_  = \new_[3002]_  ? \new_[3661]_  : \new_[3823]_ ;
  assign \new_[3405]_  = \new_[3545]_  ? \new_[5183]_  : \new_[3734]_ ;
  assign \new_[3406]_  = ~\new_[4706]_  | ~\new_[3607]_  | ~\new_[4149]_  | ~\new_[4619]_ ;
  assign \new_[3407]_  = (~\new_[3602]_  | ~\new_[6272]_ ) & (~\new_[5082]_  | ~\new_[4867]_ );
  assign \new_[3408]_  = ~\new_[3467]_ ;
  assign \new_[3409]_  = ~\new_[4544]_  & (~\new_[3605]_  | ~\new_[6589]_ );
  assign \new_[3410]_  = \new_[6105]_  ? \new_[3744]_  : \new_[2553]_ ;
  assign \new_[3411]_  = \new_[2006]_  ? \new_[5708]_  : \new_[3605]_ ;
  assign \new_[3412]_  = \new_[4121]_  ^ \new_[3605]_ ;
  assign \new_[3413]_  = ~\new_[3549]_  & (~\new_[5087]_  | ~\new_[6084]_ );
  assign \new_[3414]_  = ~\new_[3550]_  & (~\new_[4962]_  | ~\new_[5772]_ );
  assign \new_[3415]_  = ~\new_[3472]_ ;
  assign \new_[3416]_  = \new_[6285]_  ? \new_[3744]_  : \new_[2554]_ ;
  assign \new_[3417]_  = ~\new_[4371]_  | ~\new_[6264]_  | ~\new_[5471]_ ;
  assign \new_[3418]_  = ~\new_[3557]_  & (~\new_[5300]_  | ~\new_[6128]_ );
  assign \new_[3419]_  = ~\new_[3502]_ ;
  assign \new_[3420]_  = \new_[4553]_  ? \new_[1623]_  : \new_[3622]_ ;
  assign \new_[3421]_  = ~\new_[3672]_  | ~\new_[6163]_ ;
  assign \new_[3422]_  = ~\new_[3625]_  | ~\new_[4033]_  | ~\new_[3759]_ ;
  assign \new_[3423]_  = ~\new_[6313]_  | (~\new_[7148]_  & ~\new_[4379]_ );
  assign \new_[3424]_  = ~\new_[3563]_  | ~\new_[792]_ ;
  assign \new_[3425]_  = ~\new_[3563]_  | ~\new_[851]_ ;
  assign \new_[3426]_  = ~\new_[3563]_  | ~\new_[853]_ ;
  assign \new_[3427]_  = ~\new_[3563]_  | ~\new_[794]_ ;
  assign \new_[3428]_  = ~\new_[3563]_  | ~\new_[848]_ ;
  assign \new_[3429]_  = ~\new_[3563]_  | ~\new_[852]_ ;
  assign \new_[3430]_  = ~\new_[3563]_  | ~\new_[799]_ ;
  assign \new_[3431]_  = ~\new_[3563]_  | ~\new_[849]_ ;
  assign \new_[3432]_  = ~\new_[3563]_  | ~\new_[845]_ ;
  assign \new_[3433]_  = ~\new_[6698]_ ;
  assign \new_[3434]_  = ~\new_[3571]_  & ~\new_[5295]_ ;
  assign \new_[3435]_  = ~\new_[3678]_  | ~\new_[5253]_  | ~\new_[3749]_ ;
  assign \new_[3436]_  = ~\new_[3683]_  & (~\new_[3682]_  | ~\new_[3630]_ );
  assign \new_[3437]_  = ~\new_[3506]_ ;
  assign \new_[3438]_  = ~\new_[3679]_  & (~\new_[3678]_  | ~\new_[3750]_ );
  assign \new_[3439]_  = (~\new_[3641]_  | ~\new_[5969]_ ) & (~\new_[3657]_  | ~\new_[6193]_ );
  assign \new_[3440]_  = ~\new_[3575]_  & (~\new_[3686]_  | ~\new_[3675]_ );
  assign \new_[3441]_  = ~\new_[3712]_  | (~\new_[3634]_  & ~\new_[3871]_ );
  assign \new_[3442]_  = \new_[3869]_  ^ \new_[3634]_ ;
  assign \new_[3443]_  = ~\new_[3679]_  & ~\new_[3574]_ ;
  assign \new_[3444]_  = \new_[3578]_  & \new_[3577]_ ;
  assign \new_[3445]_  = ~\new_[3925]_  & ~\new_[3580]_ ;
  assign \new_[3446]_  = ~\new_[3580]_  & ~\new_[4316]_ ;
  assign \new_[3447]_  = ~\new_[3577]_  | ~\new_[3688]_ ;
  assign \new_[3448]_  = ~\new_[3579]_  | ~\new_[5472]_ ;
  assign \new_[3449]_  = ~\new_[3526]_ ;
  assign \new_[3450]_  = ~\new_[3527]_ ;
  assign \new_[3451]_  = ~\new_[5591]_  | ~\new_[3585]_ ;
  assign \new_[3452]_  = ~\new_[3529]_ ;
  assign \new_[3453]_  = (~\new_[3646]_  | ~\new_[3760]_ ) & (~\new_[3692]_  | ~\new_[3693]_ );
  assign \new_[3454]_  = ~\new_[3582]_  & (~\new_[3925]_  | ~\new_[1236]_ );
  assign \new_[3455]_  = ~\new_[3589]_  & ~\new_[3801]_ ;
  assign \new_[3456]_  = ~\new_[3590]_  | ~\new_[5780]_ ;
  assign \new_[3457]_  = (~\new_[3708]_  | ~\new_[3999]_ ) & (~\new_[3645]_  | ~\new_[3868]_ );
  assign \new_[3458]_  = ~\new_[3780]_  & (~\new_[3644]_  | ~\new_[3872]_ );
  assign n1754 = ~\new_[3595]_  & ~\new_[6424]_ ;
  assign n1759 = ~\new_[3596]_  & ~\new_[6623]_ ;
  assign n1749 = ~\new_[3597]_  & ~\new_[6623]_ ;
  assign \new_[3462]_  = ~\new_[3591]_  & (~\new_[5055]_  | ~\new_[6084]_ );
  assign \new_[3463]_  = (~\new_[3648]_  | ~\new_[5969]_ ) & (~\new_[4071]_  | ~\new_[6193]_ );
  assign \new_[3464]_  = ~\new_[3599]_  & ~\new_[6031]_ ;
  assign \new_[3465]_  = \new_[3598]_  & \new_[3654]_ ;
  assign \new_[3466]_  = ~\new_[3542]_ ;
  assign \new_[3467]_  = (~\new_[5918]_  | ~\new_[3661]_ ) & (~\new_[2552]_  | ~\new_[3744]_ );
  assign \new_[3468]_  = ~\new_[3604]_  & ~\new_[5995]_ ;
  assign \new_[3469]_  = ~\new_[3561]_ ;
  assign \new_[3470]_  = ~\new_[4343]_  | ~\new_[4964]_  | ~\new_[3609]_  | ~\new_[3828]_ ;
  assign \new_[3471]_  = ~\new_[4270]_  & ~\new_[3744]_ ;
  assign \new_[3472]_  = (~\new_[6092]_  | ~\new_[3661]_ ) & (~\new_[2555]_  | ~\new_[3744]_ );
  assign \new_[3473]_  = \new_[6472]_  ? \new_[6711]_  : \new_[5075]_ ;
  assign \new_[3474]_  = (~\new_[5070]_  | ~\new_[3660]_ ) & (~\new_[3254]_  | ~\new_[3735]_ );
  assign \new_[3475]_  = (~\new_[5072]_  | ~\new_[3660]_ ) & (~\new_[3257]_  | ~\new_[3735]_ );
  assign \new_[3476]_  = (~\new_[5060]_  | ~\new_[3660]_ ) & (~\new_[3261]_  | ~\new_[3735]_ );
  assign \new_[3477]_  = (~\new_[5074]_  | ~\new_[3660]_ ) & (~\new_[3264]_  | ~\new_[3735]_ );
  assign \new_[3478]_  = (~\new_[5063]_  | ~\new_[3660]_ ) & (~\new_[3262]_  | ~\new_[3735]_ );
  assign \new_[3479]_  = (~\new_[5067]_  | ~\new_[3660]_ ) & (~\new_[3265]_  | ~\new_[3735]_ );
  assign \new_[3480]_  = (~\new_[5064]_  | ~\new_[3660]_ ) & (~\new_[3251]_  | ~\new_[3735]_ );
  assign \new_[3481]_  = (~\new_[5065]_  | ~\new_[3660]_ ) & (~\new_[3266]_  | ~\new_[3735]_ );
  assign \new_[3482]_  = (~\new_[5066]_  | ~\new_[3660]_ ) & (~\new_[3735]_  | ~\new_[3259]_ );
  assign \new_[3483]_  = (~\new_[5069]_  | ~\new_[3660]_ ) & (~\new_[3268]_  | ~\new_[3735]_ );
  assign \new_[3484]_  = (~\new_[5073]_  | ~\new_[3660]_ ) & (~\new_[3270]_  | ~\new_[3735]_ );
  assign \new_[3485]_  = \new_[2633]_  ? \new_[6713]_  : \new_[5535]_ ;
  assign \new_[3486]_  = (~\new_[5061]_  | ~\new_[3660]_ ) & (~\new_[3267]_  | ~\new_[3735]_ );
  assign \new_[3487]_  = (~\new_[5071]_  | ~\new_[3660]_ ) & (~\new_[3269]_  | ~\new_[3735]_ );
  assign \new_[3488]_  = (~\new_[5068]_  | ~\new_[3660]_ ) & (~\new_[3260]_  | ~\new_[3735]_ );
  assign \new_[3489]_  = (~\new_[5059]_  | ~\new_[3660]_ ) & (~\new_[3271]_  | ~\new_[3735]_ );
  assign \new_[3490]_  = ~\new_[5365]_  | ~\new_[5467]_  | ~\new_[3611]_  | ~\new_[5135]_ ;
  assign \new_[3491]_  = (~\new_[5062]_  | ~\new_[3660]_ ) & (~\new_[3263]_  | ~\new_[3735]_ );
  assign n1764 = ~\new_[6363]_  | (~\new_[5505]_  & ~\new_[3666]_ );
  assign \new_[3493]_  = ~\new_[3668]_  | ~\new_[4531]_  | ~\new_[3990]_ ;
  assign \new_[3494]_  = ~\new_[3614]_  & (~\new_[7315]_  | ~\new_[6084]_ );
  assign \new_[3495]_  = ~\new_[3612]_  & (~\new_[5525]_  | ~\new_[3665]_ );
  assign \new_[3496]_  = \new_[2661]_  ? \new_[6713]_  : \new_[5652]_ ;
  assign \new_[3497]_  = ~\new_[3554]_ ;
  assign \new_[3498]_  = ~\new_[792]_  | ~\new_[3663]_ ;
  assign \new_[3499]_  = ~\new_[766]_  | ~\new_[3663]_ ;
  assign \new_[3500]_  = ~\new_[755]_  | ~\new_[3663]_ ;
  assign \new_[3501]_  = ~\new_[757]_  | ~\new_[3663]_ ;
  assign \new_[3502]_  = \new_[2007]_  ? \new_[4760]_  : \new_[3671]_ ;
  assign \new_[3503]_  = ~\new_[3743]_  | ~\new_[4405]_  | ~\new_[4573]_  | ~\new_[5245]_ ;
  assign \new_[3504]_  = \new_[3627]_  | \new_[3750]_ ;
  assign \new_[3505]_  = ~\new_[3674]_  & (~\new_[3677]_  | ~\new_[3679]_ );
  assign \new_[3506]_  = ~\new_[3686]_  & (~\new_[3684]_  | ~\new_[3687]_ );
  assign \new_[3507]_  = ~\new_[3682]_  & (~\new_[3674]_  | ~\new_[3680]_ );
  assign \new_[3508]_  = ~\new_[3687]_  & (~\new_[3685]_  | ~\new_[3683]_ );
  assign \new_[3509]_  = ~\new_[3563]_ ;
  assign \new_[3510]_  = ~\new_[3634]_  & ~\new_[3873]_ ;
  assign \new_[3511]_  = ~\new_[3682]_  & ~\new_[3629]_ ;
  assign \new_[3512]_  = ~\new_[3632]_  | ~\new_[3684]_ ;
  assign \new_[3513]_  = ~\new_[3687]_  & ~\new_[3631]_ ;
  assign \new_[3514]_  = ~\new_[3674]_  & ~\new_[3628]_ ;
  assign \new_[3515]_  = ~\new_[3565]_ ;
  assign \new_[3516]_  = ~\new_[3566]_ ;
  assign \new_[3517]_  = ~\new_[3629]_  & ~\new_[3681]_ ;
  assign \new_[3518]_  = ~\new_[3568]_ ;
  assign \new_[3519]_  = ~\new_[3569]_ ;
  assign \new_[3520]_  = ~\new_[3630]_  | ~\new_[3685]_ ;
  assign \new_[3521]_  = ~\new_[3633]_  | (~\new_[5220]_  & ~\new_[5318]_ );
  assign \new_[3522]_  = ~\new_[3572]_ ;
  assign \new_[3523]_  = ~\new_[3575]_ ;
  assign \new_[3524]_  = ~\new_[3577]_ ;
  assign \new_[3525]_  = ~\new_[3578]_ ;
  assign \new_[3526]_  = ~\new_[5256]_  | ~\new_[3636]_ ;
  assign \new_[3527]_  = \new_[5258]_  | \new_[3636]_ ;
  assign \new_[3528]_  = ~\new_[5258]_  | ~\new_[3636]_ ;
  assign \new_[3529]_  = \new_[5591]_  | \new_[3635]_ ;
  assign \new_[3530]_  = ~\new_[3637]_  & ~\new_[5746]_ ;
  assign \new_[3531]_  = ~\new_[3645]_  & (~\new_[3799]_  | ~\new_[4133]_ );
  assign \new_[3532]_  = ~\new_[3961]_  | (~\new_[3715]_  & ~\new_[3960]_ );
  assign \new_[3533]_  = ~\new_[5964]_  | ~\new_[5979]_  | ~\new_[3650]_  | ~\new_[4996]_ ;
  assign \new_[3534]_  = ~\new_[3817]_  & (~\new_[3820]_  | ~\new_[3720]_ );
  assign \new_[3535]_  = ~\new_[4444]_  & ~\new_[3618]_ ;
  assign \new_[3536]_  = ~\new_[6302]_  | ~\new_[6216]_  | ~\new_[3650]_  | ~\new_[4862]_ ;
  assign \new_[3537]_  = ~\new_[3650]_  | ~\new_[6523]_ ;
  assign \new_[3538]_  = ~\new_[3649]_  & (~\new_[6670]_  | ~\new_[5724]_ );
  assign \new_[3539]_  = ~\new_[3895]_  | ~\new_[3809]_  | ~\new_[3811]_  | ~\new_[3722]_ ;
  assign \new_[3540]_  = ~\new_[3647]_  | ~\new_[5969]_ ;
  assign \new_[3541]_  = ~\new_[3733]_  | ~\new_[5858]_  | ~\new_[3656]_  | ~\new_[5732]_ ;
  assign \new_[3542]_  = ~\new_[3651]_  & (~\new_[2551]_  | ~\new_[3744]_ );
  assign \new_[3543]_  = ~\new_[3655]_  & ~\new_[6438]_ ;
  assign \new_[3544]_  = ~\new_[3707]_  | ~\new_[5969]_ ;
  assign \new_[3545]_  = \new_[6675]_  ? \new_[5103]_  : \new_[3734]_ ;
  assign \new_[3546]_  = ~\new_[3903]_  | ~\new_[3662]_ ;
  assign \new_[3547]_  = (~\new_[3736]_  | ~\new_[5894]_ ) & (~\new_[4926]_  | ~\new_[5116]_ );
  assign \new_[3548]_  = \new_[5076]_  ? \new_[6713]_  : \new_[844]_ ;
  assign \new_[3549]_  = ~\new_[5127]_  | (~\new_[5872]_  & ~\new_[3739]_ );
  assign \new_[3550]_  = ~\new_[4751]_  | (~\new_[5872]_  & ~\new_[3738]_ );
  assign \new_[3551]_  = ~\new_[3659]_  & (~\new_[5799]_  | ~\new_[5772]_ );
  assign \new_[3552]_  = \new_[3915]_  ^ \new_[3742]_ ;
  assign \new_[3553]_  = ~\new_[4543]_  & (~\new_[3740]_  | ~\new_[6589]_ );
  assign \new_[3554]_  = \new_[4439]_  ^ \new_[3740]_ ;
  assign \new_[3555]_  = \new_[3666]_  | m1_n;
  assign \new_[3556]_  = ~\new_[6711]_  & ~\new_[6625]_ ;
  assign \new_[3557]_  = ~\new_[4117]_  | ~\new_[3670]_ ;
  assign \new_[3558]_  = \new_[7209]_  | \new_[5844]_ ;
  assign \new_[3559]_  = ~\new_[3839]_  | ~\new_[6011]_  | ~\new_[4441]_  | ~\new_[4490]_ ;
  assign \new_[3560]_  = ~\new_[3752]_  | ~\new_[3673]_ ;
  assign \new_[3561]_  = ~\new_[3704]_  | ~\new_[4041]_ ;
  assign \new_[3562]_  = ~\new_[3690]_  | (~\new_[3748]_  & ~\new_[3751]_ );
  assign \new_[3563]_  = \new_[3922]_  | \new_[3690]_ ;
  assign \new_[3564]_  = \new_[4314]_  | \new_[3706]_ ;
  assign \new_[3565]_  = ~\new_[3684]_  | ~\new_[3675]_ ;
  assign \new_[3566]_  = ~\new_[3677]_  | ~\new_[3680]_ ;
  assign \new_[3567]_  = ~\new_[3681]_  & ~\new_[3683]_ ;
  assign \new_[3568]_  = ~\new_[3684]_  | ~\new_[3685]_ ;
  assign \new_[3569]_  = \new_[3675]_  & \new_[3688]_ ;
  assign \new_[3570]_  = ~\new_[3676]_  & ~\new_[3750]_ ;
  assign \new_[3571]_  = ~\new_[3689]_  | (~\new_[3986]_  & ~\new_[3922]_ );
  assign \new_[3572]_  = ~\new_[5485]_  & ~\new_[3691]_ ;
  assign \new_[3573]_  = ~\new_[5593]_  & ~\new_[3691]_ ;
  assign \new_[3574]_  = ~\new_[3678]_ ;
  assign \new_[3575]_  = ~\new_[5484]_  & ~\new_[3691]_ ;
  assign \new_[3576]_  = ~\new_[5477]_  & ~\new_[3691]_ ;
  assign \new_[3577]_  = ~\new_[5477]_  | ~\new_[3691]_ ;
  assign \new_[3578]_  = ~\new_[5593]_  | ~\new_[3691]_ ;
  assign \new_[3579]_  = (~\new_[4336]_  | ~\new_[6193]_ ) & (~\new_[3756]_  | ~\new_[5969]_ );
  assign \new_[3580]_  = \new_[3806]_  ^ \new_[3881]_ ;
  assign \new_[3581]_  = ~\new_[3695]_  & (~\new_[5216]_  | ~\new_[4547]_ );
  assign \new_[3582]_  = ~\new_[3925]_  & ~\new_[3694]_ ;
  assign \new_[3583]_  = ~\new_[3694]_  & ~\new_[4316]_ ;
  assign \new_[3584]_  = ~\new_[3814]_  | ~\new_[3970]_  | ~\new_[3724]_  | ~\new_[3762]_ ;
  assign \new_[3585]_  = ~\new_[3636]_ ;
  assign \new_[3586]_  = i_tv80_core_PreserveC_r_reg;
  assign \new_[3587]_  = ~\new_[3781]_  & (~\new_[3782]_  | ~\new_[3875]_ );
  assign \new_[3588]_  = ~\new_[3784]_  & (~\new_[3783]_  | ~\new_[3876]_ );
  assign \new_[3589]_  = ~\new_[3783]_  & (~\new_[3781]_  | ~\new_[3880]_ );
  assign \new_[3590]_  = (~\new_[3773]_  | ~\new_[5969]_ ) & (~\new_[4481]_  | ~\new_[6193]_ );
  assign \new_[3591]_  = ~\new_[3831]_  | ~\new_[4260]_  | ~\new_[4584]_  | ~\new_[4051]_ ;
  assign \new_[3592]_  = ~\new_[3816]_  | ~\new_[3720]_ ;
  assign \new_[3593]_  = ~\new_[3642]_ ;
  assign \new_[3594]_  = ~\new_[3646]_ ;
  assign \new_[3595]_  = ~\new_[3719]_  & (~\new_[3285]_  | ~\new_[6338]_ );
  assign \new_[3596]_  = (~\new_[3726]_  | ~busak_n) & (~\new_[3321]_  | ~\new_[6258]_ );
  assign \new_[3597]_  = (~\new_[3727]_  | ~busak_n) & (~\new_[3281]_  | ~\new_[6258]_ );
  assign \new_[3598]_  = ~\new_[4207]_  & (~\new_[3728]_  | ~\new_[5969]_ );
  assign \new_[3599]_  = ~\new_[3723]_  & (~\new_[5575]_  | ~\new_[6227]_ );
  assign \new_[3600]_  = \\i_tv80_core_I_reg[5] ;
  assign \new_[3601]_  = ~\new_[4413]_  & ~\new_[6713]_ ;
  assign \new_[3602]_  = ~\new_[4964]_  | ~\new_[3732]_  | ~\new_[4052]_ ;
  assign \new_[3603]_  = \\i_tv80_core_I_reg[2] ;
  assign \new_[3604]_  = (~\new_[5206]_  | ~\new_[4288]_ ) & (~\new_[5157]_  | ~\new_[3835]_ );
  assign \new_[3605]_  = ~\new_[3910]_  | ~\new_[5738]_  | ~\new_[3832]_  | ~\new_[5828]_ ;
  assign \new_[3606]_  = \\i_tv80_core_I_reg[4] ;
  assign \new_[3607]_  = (~\new_[5994]_  | ~\new_[6128]_ ) & (~\new_[5782]_  | ~\new_[3835]_ );
  assign \new_[3608]_  = (~\new_[5895]_  | ~\new_[3835]_ ) & (~\new_[5799]_  | ~\new_[6128]_ );
  assign \new_[3609]_  = (~\new_[5526]_  | ~\new_[3834]_ ) & (~\new_[5656]_  | ~\new_[4115]_ );
  assign \new_[3610]_  = ~\new_[4555]_  & ~\new_[3740]_ ;
  assign \new_[3611]_  = ~\new_[3741]_  & ~\new_[4055]_ ;
  assign \new_[3612]_  = ~\new_[5402]_  & ~\new_[3739]_ ;
  assign \new_[3613]_  = \new_[6712]_  & \new_[850]_ ;
  assign \new_[3614]_  = ~\new_[5602]_  & ~\new_[3739]_ ;
  assign \new_[3615]_  = \\i_tv80_core_I_reg[7] ;
  assign \new_[3616]_  = ~\new_[3663]_ ;
  assign \new_[3617]_  = ~\new_[3664]_ ;
  assign \new_[3618]_  = ~\new_[3664]_ ;
  assign \new_[3619]_  = ~\new_[3664]_ ;
  assign \new_[3620]_  = ~\new_[3664]_ ;
  assign \new_[3621]_  = \\i_tv80_core_I_reg[6] ;
  assign \new_[3622]_  = ~\new_[4756]_  | ~\new_[3916]_  | ~\new_[4573]_  | ~\new_[4443]_ ;
  assign \new_[3623]_  = ~\new_[3672]_ ;
  assign \new_[3624]_  = ~\new_[4585]_  | ~\new_[4610]_  | ~\new_[3747]_  | ~\new_[4309]_ ;
  assign \new_[3625]_  = ~\new_[6313]_  | (~\new_[3850]_  & ~\new_[3920]_ );
  assign \new_[3626]_  = \\i_tv80_core_I_reg[0] ;
  assign \new_[3627]_  = \new_[5253]_  & \new_[3749]_ ;
  assign \new_[3628]_  = ~\new_[3677]_ ;
  assign \new_[3629]_  = ~\new_[3680]_ ;
  assign \new_[3630]_  = ~\new_[3681]_ ;
  assign \new_[3631]_  = ~\new_[3685]_ ;
  assign \new_[3632]_  = ~\new_[3686]_ ;
  assign \new_[3633]_  = ~\new_[3755]_  | ~\new_[6040]_ ;
  assign \new_[3634]_  = ~\new_[3779]_  & (~\new_[3881]_  | ~\new_[3870]_ );
  assign \new_[3635]_  = ~\new_[3691]_ ;
  assign \new_[3636]_  = \new_[3691]_ ;
  assign \new_[3637]_  = ~\new_[3795]_  & (~\new_[3925]_  | ~\new_[1293]_ );
  assign \new_[3638]_  = \\i_tv80_core_I_reg[1] ;
  assign \new_[3639]_  = \\i_tv80_core_I_reg[3] ;
  assign \new_[3640]_  = ~\new_[3772]_  | ~\new_[5969]_ ;
  assign \new_[3641]_  = ~\new_[5903]_  | ~\new_[3774]_  | ~\new_[5373]_ ;
  assign \new_[3642]_  = \new_[3797]_  & \new_[3872]_ ;
  assign \new_[3643]_  = ~\new_[3710]_ ;
  assign \new_[3644]_  = ~\new_[3712]_ ;
  assign \new_[3645]_  = ~\new_[3800]_  | ~\new_[4017]_ ;
  assign \new_[3646]_  = ~\new_[3961]_  | (~\new_[3960]_  & ~\new_[3883]_ );
  assign \new_[3647]_  = ~\new_[3818]_  | ~\new_[3725]_ ;
  assign \new_[3648]_  = ~\new_[5217]_  | ~\new_[5078]_  | ~\new_[3812]_  | ~\new_[6937]_ ;
  assign \new_[3649]_  = ~\new_[5724]_  & (~\new_[3822]_  | ~\new_[2826]_ );
  assign \new_[3650]_  = ~\new_[3720]_ ;
  assign \new_[3651]_  = ~\new_[5913]_  & ~\new_[3744]_ ;
  assign \new_[3652]_  = ~\new_[3729]_  | ~\new_[5614]_ ;
  assign \new_[3653]_  = ~\new_[6193]_  | (~\new_[3901]_  & ~\new_[3904]_ );
  assign \new_[3654]_  = ~\new_[3824]_  | ~\new_[6272]_ ;
  assign \new_[3655]_  = ~\new_[3826]_  & (~\new_[5351]_  | ~\new_[5123]_ );
  assign \new_[3656]_  = (~\new_[3906]_  | ~\new_[6952]_ ) & (~\new_[6324]_  | ~\new_[5959]_ );
  assign \new_[3657]_  = \new_[4600]_  | \new_[3829]_ ;
  assign \new_[3658]_  = ~\new_[3833]_  | ~\new_[5201]_ ;
  assign \new_[3659]_  = \new_[5895]_  & \new_[3834]_ ;
  assign \new_[3660]_  = ~\new_[3735]_ ;
  assign \new_[3661]_  = ~\new_[3744]_ ;
  assign \new_[3662]_  = ~\new_[3908]_  & (~\new_[4371]_  | ~\new_[6519]_ );
  assign \new_[3663]_  = \new_[6713]_ ;
  assign \new_[3664]_  = ~\new_[6713]_ ;
  assign \new_[3665]_  = \new_[7209]_  & \new_[6084]_ ;
  assign \new_[3666]_  = ~\new_[7209]_  & ~\new_[5746]_ ;
  assign \new_[3667]_  = \new_[5135]_  ^ \new_[3911]_ ;
  assign \new_[3668]_  = ~\new_[5772]_  | ~\new_[7209]_  | ~\new_[5447]_ ;
  assign \new_[3669]_  = ~\new_[3837]_  & (~\new_[4663]_  | ~\new_[6040]_ );
  assign \new_[3670]_  = ~\new_[6128]_  | ~\new_[7209]_  | ~\new_[5447]_ ;
  assign \new_[3671]_  = \new_[4557]_  ? \new_[1623]_  : \new_[3912]_ ;
  assign \new_[3672]_  = \new_[6548]_  ? \new_[4760]_  : \new_[3918]_ ;
  assign \new_[3673]_  = ~\new_[6313]_  | (~\new_[4455]_  & ~\new_[7037]_ );
  assign \new_[3674]_  = ~\new_[5586]_  & ~\new_[3844]_ ;
  assign \new_[3675]_  = ~\new_[5484]_  | ~\new_[3848]_ ;
  assign \new_[3676]_  = ~\new_[3749]_ ;
  assign \new_[3677]_  = ~\new_[5586]_  | ~\new_[3844]_ ;
  assign \new_[3678]_  = ~\new_[5478]_  | ~\new_[3845]_ ;
  assign \new_[3679]_  = ~\new_[5478]_  & ~\new_[3845]_ ;
  assign \new_[3680]_  = ~\new_[5481]_  | ~\new_[3846]_ ;
  assign \new_[3681]_  = \new_[5482]_  & \new_[3847]_ ;
  assign \new_[3682]_  = ~\new_[5481]_  & ~\new_[3846]_ ;
  assign \new_[3683]_  = ~\new_[5482]_  & ~\new_[3847]_ ;
  assign \new_[3684]_  = ~\new_[5563]_  | ~\new_[3848]_ ;
  assign \new_[3685]_  = ~\new_[5483]_  | ~\new_[3843]_ ;
  assign \new_[3686]_  = ~\new_[5563]_  & ~\new_[3848]_ ;
  assign \new_[3687]_  = ~\new_[5483]_  & ~\new_[3843]_ ;
  assign \new_[3688]_  = ~\new_[5485]_  | ~\new_[3848]_ ;
  assign \new_[3689]_  = ~\new_[3751]_ ;
  assign \new_[3690]_  = ~\new_[6994]_  | ~\new_[3849]_ ;
  assign \new_[3691]_  = ~\new_[3753]_ ;
  assign \new_[3692]_  = (~\new_[3967]_  | ~\new_[3948]_ ) & (~\new_[3963]_  | ~\new_[6629]_ );
  assign \new_[3693]_  = (~\new_[3967]_  | ~\new_[3963]_ ) & (~\new_[3948]_  | ~\new_[6629]_ );
  assign \new_[3694]_  = \new_[4133]_  ^ \new_[3930]_ ;
  assign \new_[3695]_  = ~\new_[6031]_  & (~\new_[3928]_  | ~\new_[6800]_ );
  assign \new_[3696]_  = ~\new_[4007]_  | (~\new_[4300]_  & ~\new_[5487]_ );
  assign \new_[3697]_  = ~\new_[4007]_  | (~\new_[4214]_  & ~\new_[5492]_ );
  assign \new_[3698]_  = ~\new_[4007]_  | (~\new_[4211]_  & ~\new_[5488]_ );
  assign \new_[3699]_  = ~\new_[4007]_  | (~\new_[4215]_  & ~\new_[5498]_ );
  assign \new_[3700]_  = ~\new_[4007]_  | (~\new_[4302]_  & ~\new_[5489]_ );
  assign \new_[3701]_  = ~\new_[4007]_  | (~\new_[4303]_  & ~\new_[5499]_ );
  assign \new_[3702]_  = ~\new_[4007]_  | (~\new_[4304]_  & ~\new_[5502]_ );
  assign \new_[3703]_  = ~\new_[4007]_  | (~\new_[4305]_  & ~\new_[5501]_ );
  assign \new_[3704]_  = ~\new_[3761]_ ;
  assign \new_[3705]_  = ~\new_[3854]_ ;
  assign \new_[3706]_  = ~\new_[4012]_  | ~\new_[5233]_  | ~\new_[4987]_  | ~\new_[4973]_ ;
  assign \new_[3707]_  = ~\new_[3977]_  | ~\new_[6800]_  | ~\new_[4010]_  | ~\new_[4809]_ ;
  assign \new_[3708]_  = \new_[3868]_  & \new_[3951]_ ;
  assign \new_[3709]_  = ~\new_[3868]_  | ~\new_[3875]_ ;
  assign \new_[3710]_  = \new_[3875]_  & \new_[3880]_ ;
  assign \new_[3711]_  = ~\new_[5378]_  & (~\new_[3964]_  | ~\new_[6193]_ );
  assign \new_[3712]_  = ~\new_[3950]_  & (~\new_[4021]_  | ~\new_[3952]_ );
  assign \new_[3713]_  = ~\new_[3958]_  & (~\new_[4027]_  | ~\new_[3956]_ );
  assign \new_[3714]_  = ~\new_[3782]_ ;
  assign \new_[3715]_  = ~\new_[3878]_  & ~\new_[3949]_ ;
  assign n1769 = ~\new_[3813]_  & ~\new_[6623]_ ;
  assign \new_[3717]_  = ~\new_[3961]_  | ~\new_[3884]_ ;
  assign \new_[3718]_  = ~\new_[3948]_  | ~\new_[3885]_ ;
  assign \new_[3719]_  = ~\new_[3815]_  & ~\new_[1690]_ ;
  assign \new_[3720]_  = ~\new_[5653]_  | ~\new_[3882]_  | ~\new_[4507]_ ;
  assign \new_[3721]_  = ~\new_[3963]_  & (~\new_[4075]_  | ~\new_[1292]_ );
  assign \new_[3722]_  = ~\new_[3821]_  & (~\new_[3997]_  | ~\new_[3971]_ );
  assign \new_[3723]_  = ~\new_[5233]_  | ~\new_[4973]_  | ~\new_[3896]_  | ~\new_[3902]_ ;
  assign \new_[3724]_  = ~\new_[3819]_  & ~\new_[3971]_ ;
  assign \new_[3725]_  = ~\new_[6104]_  | ~\new_[6812]_  | ~\new_[5887]_  | ~\new_[3968]_ ;
  assign \new_[3726]_  = \new_[3321]_  ? \new_[3969]_  : \new_[4098]_ ;
  assign \new_[3727]_  = \new_[3281]_  ? \new_[3969]_  : \new_[4101]_ ;
  assign \new_[3728]_  = ~\new_[4907]_  | ~\new_[5297]_  | ~\new_[7159]_  | ~\new_[3978]_ ;
  assign \new_[3729]_  = ~\new_[3817]_ ;
  assign \new_[3730]_  = ~\new_[6193]_  | (~\new_[4411]_  & ~\new_[3982]_ );
  assign \new_[3731]_  = ~\new_[3900]_  | (~\new_[4043]_  & ~\new_[4048]_ );
  assign \new_[3732]_  = ~\new_[3824]_ ;
  assign \new_[3733]_  = ~\new_[3906]_  | ~\new_[6953]_ ;
  assign \new_[3734]_  = \new_[5020]_  ? \new_[6713]_  : \new_[6521]_ ;
  assign \new_[3735]_  = ~\new_[3664]_  | ~\new_[6714]_ ;
  assign \new_[3736]_  = ~\new_[3909]_  | ~\new_[5983]_ ;
  assign \new_[3737]_  = ~\new_[3907]_  & (~\new_[5536]_  | ~\new_[4308]_ );
  assign \new_[3738]_  = ~\new_[3834]_ ;
  assign \new_[3739]_  = ~\new_[4371]_  & ~\new_[6084]_ ;
  assign \new_[3740]_  = ~\new_[4054]_  | ~\new_[5856]_  | ~\new_[3991]_  | ~\new_[5797]_ ;
  assign \new_[3741]_  = ~\new_[3989]_  | ~\new_[4120]_  | ~\new_[5243]_ ;
  assign \new_[3742]_  = \new_[5365]_  ^ \new_[3989]_ ;
  assign \new_[3743]_  = ~\new_[3917]_  | ~\new_[6589]_ ;
  assign \new_[3744]_  = \new_[3664]_  | \new_[6271]_ ;
  assign \new_[3745]_  = (~\new_[3994]_  | ~\new_[5459]_ ) & (~\new_[4608]_  | ~\new_[6040]_ );
  assign \new_[3746]_  = ~\new_[3919]_  | ~\new_[6163]_ ;
  assign \new_[3747]_  = ~\new_[3921]_  & (~\new_[5301]_  | ~\new_[5455]_ );
  assign \new_[3748]_  = ~\new_[4370]_  & ~\new_[3922]_ ;
  assign \new_[3749]_  = ~\new_[5480]_  | ~\new_[3923]_ ;
  assign \new_[3750]_  = ~\new_[5480]_  & ~\new_[3923]_ ;
  assign \new_[3751]_  = ~\new_[7304]_ ;
  assign \new_[3752]_  = ~\new_[4393]_  & (~\new_[7224]_  | ~\new_[6471]_ );
  assign \new_[3753]_  = ~\new_[3848]_ ;
  assign \new_[3754]_  = ~\new_[3849]_ ;
  assign \new_[3755]_  = (~\new_[4005]_  & ~\new_[5969]_ ) | (~\new_[6659]_  & ~\new_[6031]_ );
  assign \new_[3756]_  = ~\new_[4061]_  | ~\new_[5189]_  | ~\new_[5690]_  | ~\new_[5292]_ ;
  assign \new_[3757]_  = ~\new_[4132]_  | (~\new_[4298]_  & ~\new_[5491]_ );
  assign \new_[3758]_  = ~\new_[4132]_  | (~\new_[4296]_  & ~\new_[5494]_ );
  assign \new_[3759]_  = ~\new_[6193]_  | (~\new_[4006]_  & ~\new_[4310]_ );
  assign \new_[3760]_  = ~\new_[3962]_  & ~\new_[3963]_ ;
  assign \new_[3761]_  = ~\new_[3929]_  | ~\new_[5706]_ ;
  assign \new_[3762]_  = (~\new_[4009]_  | ~\new_[3968]_ ) & (~\new_[5310]_  | ~\new_[4036]_ );
  assign \new_[3763]_  = ~\new_[4062]_  | ~\new_[4553]_ ;
  assign \new_[3764]_  = ~\new_[4062]_  | ~\new_[4559]_ ;
  assign \new_[3765]_  = ~\new_[4062]_  | ~\new_[1646]_ ;
  assign \new_[3766]_  = ~\new_[4062]_  | ~\new_[4554]_ ;
  assign \new_[3767]_  = ~\new_[3935]_  | ~\new_[7466]_ ;
  assign \new_[3768]_  = ~\new_[3939]_  | ~\new_[6745]_ ;
  assign \new_[3769]_  = ~\new_[3943]_  | ~\new_[6745]_ ;
  assign \new_[3770]_  = ~\new_[3941]_  | ~\new_[6745]_ ;
  assign \new_[3771]_  = ~\new_[3940]_  | ~\new_[7466]_ ;
  assign \new_[3772]_  = ~\new_[5233]_  | ~\new_[3947]_  | ~\new_[4369]_ ;
  assign \new_[3773]_  = ~\new_[5430]_  | ~\new_[3931]_  | ~\new_[5690]_ ;
  assign \new_[3774]_  = ~\new_[3946]_  & ~\new_[3980]_ ;
  assign \new_[3775]_  = ~\new_[4007]_  | (~\new_[4145]_  & ~\new_[5495]_ );
  assign \new_[3776]_  = ~\new_[4007]_  | (~\new_[4146]_  & ~\new_[5497]_ );
  assign \new_[3777]_  = ~\new_[4007]_  | (~\new_[4147]_  & ~\new_[5496]_ );
  assign \new_[3778]_  = ~\new_[4007]_  | (~\new_[4144]_  & ~\new_[5493]_ );
  assign \new_[3779]_  = ~\new_[4067]_  | (~\new_[4066]_  & ~\new_[4017]_ );
  assign \new_[3780]_  = ~\new_[4014]_  | (~\new_[4022]_  & ~\new_[4024]_ );
  assign \new_[3781]_  = ~\new_[4024]_  | (~\new_[4023]_  & ~\new_[4015]_ );
  assign \new_[3782]_  = ~\new_[3953]_  | (~\new_[4067]_  & ~\new_[4019]_ );
  assign \new_[3783]_  = ~\new_[3957]_  | (~\new_[4014]_  & ~\new_[4026]_ );
  assign \new_[3784]_  = ~\new_[4029]_  | (~\new_[4030]_  & ~\new_[4028]_ );
  assign n1799 = ~\new_[3887]_  & ~\new_[6403]_ ;
  assign n1804 = ~\new_[3888]_  & ~\new_[6382]_ ;
  assign n1779 = ~\new_[3889]_  & ~\new_[6413]_ ;
  assign n1809 = ~\new_[3890]_  & ~\new_[6424]_ ;
  assign n1784 = ~\new_[3891]_  & ~\new_[6424]_ ;
  assign n1774 = ~\new_[3892]_  & ~\new_[6402]_ ;
  assign n1794 = ~\new_[3893]_  & ~\new_[6402]_ ;
  assign n1789 = ~\new_[3894]_  & ~\new_[6424]_ ;
  assign \new_[3793]_  = ~\new_[4031]_  & ~\new_[3960]_ ;
  assign \new_[3794]_  = ~\new_[3956]_  | ~\new_[4028]_ ;
  assign \new_[3795]_  = ~\new_[3925]_  & ~\new_[4064]_ ;
  assign \new_[3796]_  = ~\new_[3952]_  | ~\new_[4015]_ ;
  assign \new_[3797]_  = ~\new_[3871]_ ;
  assign \new_[3798]_  = ~\new_[3959]_  & ~\new_[4030]_ ;
  assign \new_[3799]_  = \new_[4134]_  & \new_[3951]_ ;
  assign \new_[3800]_  = ~\new_[3951]_  | ~\new_[4135]_ ;
  assign \new_[3801]_  = ~\new_[3876]_ ;
  assign \new_[3802]_  = \new_[4031]_  | \new_[3949]_ ;
  assign \new_[3803]_  = ~\new_[3925]_  | ~\new_[1294]_ ;
  assign \new_[3804]_  = ~\new_[4024]_  | ~\new_[3955]_ ;
  assign \new_[3805]_  = ~\new_[4014]_  | ~\new_[3954]_ ;
  assign \new_[3806]_  = ~\new_[4017]_  | ~\new_[3951]_ ;
  assign \new_[3807]_  = \new_[1255]_  ^ \new_[3967]_ ;
  assign \new_[3808]_  = ~\new_[3882]_ ;
  assign \new_[3809]_  = ~\new_[4036]_  & (~\new_[4340]_  | ~\new_[3968]_ );
  assign \new_[3810]_  = ~\new_[4331]_  & (~\new_[3975]_  | ~\new_[6193]_ );
  assign \new_[3811]_  = (~\new_[4008]_  | ~\new_[3972]_ ) & (~\new_[3995]_  | ~\new_[4038]_ );
  assign \new_[3812]_  = ~\new_[3898]_  & (~\new_[5865]_  | ~\new_[6284]_ );
  assign \new_[3813]_  = ~\new_[3965]_  & (~\new_[3586]_  | ~\new_[6338]_ );
  assign \new_[3814]_  = (~\new_[4035]_  | ~\new_[6519]_ ) & (~\new_[4037]_  | ~\new_[5148]_ );
  assign \new_[3815]_  = (~\new_[4039]_  | ~\new_[6047]_ ) & (~\new_[5183]_  | ~\new_[3285]_ );
  assign \new_[3816]_  = ~\new_[3974]_  & ~\new_[4096]_ ;
  assign \new_[3817]_  = ~\new_[3976]_  | ~\new_[4418]_ ;
  assign \new_[3818]_  = ~\new_[4487]_  | ~\new_[3968]_ ;
  assign \new_[3819]_  = \new_[4038]_  | \new_[3972]_ ;
  assign \new_[3820]_  = ~\new_[3974]_  | ~\new_[4044]_ ;
  assign \new_[3821]_  = ~\new_[3970]_  & (~\new_[6520]_  | ~\new_[5116]_ );
  assign \new_[3822]_  = ~\new_[4047]_  | (~\new_[4048]_  & ~\new_[4270]_ );
  assign \new_[3823]_  = (~\new_[4271]_  & ~\new_[4193]_  & ~\new_[6128]_ ) | (~\new_[4048]_  & ~\new_[4270]_  & ~\new_[6669]_ );
  assign \new_[3824]_  = ~\new_[4111]_  | ~\new_[4825]_  | ~\new_[4114]_  | ~\new_[4746]_ ;
  assign \new_[3825]_  = ~\new_[3903]_ ;
  assign \new_[3826]_  = ~\new_[6031]_  & (~\new_[4050]_  | ~\new_[4650]_ );
  assign \new_[3827]_  = \new_[4004]_  | \new_[5925]_ ;
  assign \new_[3828]_  = \new_[3983]_  & \new_[4114]_ ;
  assign \new_[3829]_  = \new_[3984]_  | \new_[3982]_ ;
  assign \new_[3830]_  = ~\new_[3985]_  & (~\new_[5203]_  | ~\new_[6128]_ );
  assign \new_[3831]_  = ~\new_[4185]_  & (~\new_[4046]_  | ~\new_[6084]_ );
  assign \new_[3832]_  = (~\new_[4053]_  | ~\new_[6952]_ ) & (~\new_[6476]_  | ~\new_[5959]_ );
  assign \new_[3833]_  = ~\new_[3988]_  & (~\new_[5429]_  | ~\new_[6084]_ );
  assign \new_[3834]_  = \new_[7209]_  & \new_[5772]_ ;
  assign \new_[3835]_  = \new_[7209]_  & \new_[6128]_ ;
  assign \new_[3836]_  = ~\new_[3908]_ ;
  assign \new_[3837]_  = ~\new_[3989]_  & ~\new_[5877]_ ;
  assign \new_[3838]_  = \new_[4545]_  & \new_[3992]_ ;
  assign \new_[3839]_  = ~\new_[3913]_ ;
  assign \new_[3840]_  = ~\new_[3919]_ ;
  assign \new_[3841]_  = i_tv80_core_Arith16_r_reg;
  assign \new_[3842]_  = ~\new_[3922]_ ;
  assign \new_[3843]_  = ~\new_[7545]_  & (~\new_[4549]_  | ~\new_[6215]_ );
  assign \new_[3844]_  = ~\new_[7545]_  & (~\new_[4553]_  | ~\new_[6384]_ );
  assign \new_[3845]_  = ~\new_[7545]_  & (~\new_[4557]_  | ~\new_[6384]_ );
  assign \new_[3846]_  = ~\new_[7545]_  & (~\new_[4558]_  | ~\new_[6215]_ );
  assign \new_[3847]_  = ~\new_[7545]_  & (~\new_[4559]_  | ~\new_[6215]_ );
  assign \new_[3848]_  = ~\new_[7545]_  & (~\new_[4556]_  | ~\new_[6215]_ );
  assign \new_[3849]_  = ~\new_[7302]_ ;
  assign \new_[3850]_  = ~\new_[4685]_  | ~\new_[7262]_  | ~\new_[4000]_  | ~\new_[4514]_ ;
  assign \new_[3851]_  = ~\new_[4007]_  | (~\new_[4299]_  & ~\new_[5490]_ );
  assign \new_[3852]_  = ~\new_[4007]_  | (~\new_[4301]_  & ~\new_[5510]_ );
  assign \new_[3853]_  = ~\new_[3926]_ ;
  assign \new_[3854]_  = ~\new_[4001]_ ;
  assign \new_[3855]_  = ~\new_[4062]_  | ~\new_[1689]_ ;
  assign \new_[3856]_  = ~\new_[4062]_  | ~\new_[1578]_ ;
  assign \new_[3857]_  = ~\new_[4062]_  | ~\new_[2429]_ ;
  assign \new_[3858]_  = ~\new_[4062]_  | ~\new_[4557]_ ;
  assign \new_[3859]_  = ~\new_[4062]_  | ~\new_[4558]_ ;
  assign \new_[3860]_  = ~\new_[4062]_  | ~\new_[4549]_ ;
  assign \new_[3861]_  = ~\new_[4062]_  | ~\new_[4556]_ ;
  assign \new_[3862]_  = ~\new_[4062]_  | ~\new_[2034]_ ;
  assign \new_[3863]_  = ~\new_[4062]_  | ~\new_[1925]_ ;
  assign \new_[3864]_  = ~\new_[4062]_  | ~\new_[1892]_ ;
  assign \new_[3865]_  = ~\new_[4062]_  | ~\new_[1861]_ ;
  assign \new_[3866]_  = ~\new_[4062]_  | ~\new_[4560]_ ;
  assign \new_[3867]_  = ~\new_[4013]_  | ~\new_[6745]_ ;
  assign \new_[3868]_  = ~\new_[4066]_  & ~\new_[4019]_ ;
  assign \new_[3869]_  = ~\new_[4021]_  & ~\new_[4019]_ ;
  assign \new_[3870]_  = ~\new_[4066]_  & ~\new_[4016]_ ;
  assign \new_[3871]_  = \new_[4019]_  | \new_[4020]_ ;
  assign \new_[3872]_  = ~\new_[4022]_  & ~\new_[4023]_ ;
  assign \new_[3873]_  = \new_[4026]_  | \new_[4025]_ ;
  assign \new_[3874]_  = \new_[4027]_  | \new_[4026]_ ;
  assign \new_[3875]_  = ~\new_[4020]_  & ~\new_[4023]_ ;
  assign \new_[3876]_  = ~\new_[4030]_  & ~\new_[4025]_ ;
  assign \new_[3877]_  = ~\new_[4031]_  & ~\new_[4030]_ ;
  assign \new_[3878]_  = ~\new_[4031]_  & ~\new_[4029]_ ;
  assign \new_[3879]_  = ~\new_[4018]_  & ~\new_[4066]_ ;
  assign \new_[3880]_  = ~\new_[4022]_  & ~\new_[4026]_ ;
  assign \new_[3881]_  = \new_[3999]_  | \new_[4135]_ ;
  assign \new_[3882]_  = ~i_tv80_core_No_BTR_reg;
  assign \new_[3883]_  = ~\new_[3949]_ ;
  assign \new_[3884]_  = ~\new_[3960]_ ;
  assign \new_[3885]_  = ~\new_[3962]_ ;
  assign \new_[3886]_  = ~\new_[5969]_  | ~\new_[6378]_  | ~\new_[4035]_ ;
  assign \new_[3887]_  = (~\new_[4085]_  | ~\new_[6126]_ ) & (~\new_[3626]_  | ~\new_[6225]_ );
  assign \new_[3888]_  = (~\new_[4086]_  | ~\new_[6714]_ ) & (~\new_[3638]_  | ~\new_[6165]_ );
  assign \new_[3889]_  = (~\new_[4087]_  | ~\new_[6714]_ ) & (~\new_[3603]_  | ~\new_[1690]_ );
  assign \new_[3890]_  = (~\new_[4088]_  | ~\new_[6714]_ ) & (~\new_[3639]_  | ~\new_[6225]_ );
  assign \new_[3891]_  = (~\new_[4089]_  | ~\new_[6099]_ ) & (~\new_[3606]_  | ~\new_[1690]_ );
  assign \new_[3892]_  = (~\new_[4090]_  | ~\new_[6099]_ ) & (~\new_[3600]_  | ~\new_[6165]_ );
  assign \new_[3893]_  = (~\new_[4091]_  | ~\new_[6314]_ ) & (~\new_[3621]_  | ~\new_[6239]_ );
  assign \new_[3894]_  = (~\new_[4092]_  | ~\new_[6314]_ ) & (~\new_[3615]_  | ~\new_[6239]_ );
  assign \new_[3895]_  = ~\new_[4035]_  & ~\new_[4037]_ ;
  assign \new_[3896]_  = ~\new_[4040]_  & (~\new_[5770]_  | ~\new_[5727]_ );
  assign \new_[3897]_  = ~\new_[5207]_  | ~\new_[4819]_  | ~\new_[4496]_  | ~\new_[4108]_ ;
  assign \new_[3898]_  = ~\new_[4337]_  | ~\new_[4855]_  | ~\new_[4422]_  | ~\new_[4102]_ ;
  assign \new_[3899]_  = ~\new_[5969]_  | ~\new_[4037]_  | ~\new_[5259]_ ;
  assign \new_[3900]_  = ~\new_[6128]_  | ~\new_[4194]_  | ~\new_[4270]_ ;
  assign \new_[3901]_  = ~\new_[4112]_  | ~\new_[6016]_  | ~\new_[4936]_ ;
  assign \new_[3902]_  = ~\new_[4049]_  & (~\new_[5353]_  | ~\new_[5958]_ );
  assign \new_[3903]_  = (~\new_[4106]_  | ~\new_[6193]_ ) & (~\new_[4539]_  | ~\new_[5969]_ );
  assign \new_[3904]_  = ~\new_[5193]_  | ~\new_[4849]_  | ~\new_[4109]_ ;
  assign \new_[3905]_  = ~\new_[4278]_  & (~\new_[4115]_  | ~\new_[7121]_ );
  assign \new_[3906]_  = \new_[5025]_  ^ \new_[4118]_ ;
  assign \new_[3907]_  = ~\new_[4057]_  & ~\new_[5255]_ ;
  assign \new_[3908]_  = \new_[4371]_  & \new_[6523]_ ;
  assign \new_[3909]_  = ~\new_[4371]_  | ~\new_[6378]_ ;
  assign \new_[3910]_  = ~\new_[4053]_  | ~\new_[6953]_ ;
  assign \new_[3911]_  = \new_[5243]_  ^ \new_[4120]_ ;
  assign \new_[3912]_  = ~\new_[4860]_  | ~\new_[4208]_  | ~\new_[4643]_  | ~\new_[4419]_ ;
  assign \new_[3913]_  = ~\new_[1624]_  & (~\new_[4123]_  | ~\new_[5821]_ );
  assign \new_[3914]_  = \new_[4779]_  & \new_[4056]_ ;
  assign \new_[3915]_  = \new_[6478]_  ^ \new_[4122]_ ;
  assign \new_[3916]_  = ~\new_[4635]_  & (~\new_[4121]_  | ~\new_[6589]_ );
  assign \new_[3917]_  = \new_[2005]_  ? \new_[5708]_  : \new_[4121]_ ;
  assign \new_[3918]_  = \new_[4554]_  ? \new_[1623]_  : \new_[4124]_ ;
  assign \new_[3919]_  = \new_[6528]_  ? \new_[4760]_  : \new_[4125]_ ;
  assign \new_[3920]_  = ~\new_[7120]_  | ~\new_[5704]_  | ~\new_[4143]_  | ~\new_[4127]_ ;
  assign \new_[3921]_  = ~\new_[4816]_  | ~\new_[4689]_  | ~\new_[4128]_ ;
  assign \new_[3922]_  = ~\new_[6702]_ ;
  assign \new_[3923]_  = ~\new_[7546]_  & (~\new_[4554]_  | ~\new_[6384]_ );
  assign \new_[3924]_  = ~\new_[4064]_  & ~\new_[4316]_ ;
  assign \new_[3925]_  = ~\new_[7173]_  | ~\new_[4997]_  | ~\new_[6100]_  | ~\new_[4132]_ ;
  assign \new_[3926]_  = ~\new_[4001]_ ;
  assign \new_[3927]_  = ~\new_[7094]_ ;
  assign \new_[3928]_  = ~\new_[4063]_  & ~\new_[5500]_ ;
  assign \new_[3929]_  = (~\new_[4140]_  | ~\new_[5969]_ ) & (~\new_[4403]_  | ~\new_[6193]_ );
  assign \new_[3930]_  = ~\new_[4134]_  | ~\new_[4065]_ ;
  assign \new_[3931]_  = ~\new_[4034]_  & (~\new_[5017]_  | ~\new_[5910]_ );
  assign \new_[3932]_  = ~\new_[4154]_  | ~\new_[4184]_  | ~\new_[4257]_  | ~\new_[4235]_ ;
  assign \new_[3933]_  = ~\new_[4176]_  | ~\new_[4177]_  | ~\new_[4246]_  | ~\new_[4255]_ ;
  assign \new_[3934]_  = ~\new_[4166]_  | ~\new_[4167]_  | ~\new_[4258]_  | ~\new_[4241]_ ;
  assign \new_[3935]_  = ~\new_[4180]_  | ~\new_[4234]_  | ~\new_[4233]_  | ~\new_[4159]_ ;
  assign \new_[3936]_  = ~\new_[4182]_  | ~\new_[4161]_  | ~\new_[4228]_  | ~\new_[4227]_ ;
  assign \new_[3937]_  = ~\new_[4155]_  | ~\new_[4157]_  | ~\new_[4256]_  | ~\new_[4236]_ ;
  assign \new_[3938]_  = ~\new_[4153]_  | ~\new_[4162]_  | ~\new_[4229]_  | ~\new_[4237]_ ;
  assign \new_[3939]_  = ~\new_[4253]_  | ~\new_[4181]_  | ~\new_[4156]_  | ~\new_[4239]_ ;
  assign \new_[3940]_  = ~\new_[4250]_  | ~\new_[4164]_  | ~\new_[4163]_  | ~\new_[4230]_ ;
  assign \new_[3941]_  = ~\new_[4160]_  | ~\new_[4165]_  | ~\new_[4252]_  | ~\new_[4240]_ ;
  assign \new_[3942]_  = ~\new_[4170]_  | ~\new_[4171]_  | ~\new_[4243]_  | ~\new_[4232]_ ;
  assign \new_[3943]_  = ~\new_[4173]_  | ~\new_[4244]_  | ~\new_[4172]_  | ~\new_[4231]_ ;
  assign \new_[3944]_  = ~\new_[4175]_  | ~\new_[4254]_  | ~\new_[4174]_  | ~\new_[4245]_ ;
  assign \new_[3945]_  = ~\new_[4183]_  | ~\new_[4158]_  | ~\new_[4251]_  | ~\new_[4249]_ ;
  assign \new_[3946]_  = ~\new_[4150]_  | ~\new_[5741]_  | ~\new_[7159]_  | ~\new_[6932]_ ;
  assign \new_[3947]_  = ~\new_[4069]_  & (~\new_[4850]_  | ~\new_[5116]_ );
  assign \new_[3948]_  = ~\new_[4075]_  | ~\new_[1235]_ ;
  assign \new_[3949]_  = \new_[4075]_  & \new_[1233]_ ;
  assign \new_[3950]_  = ~\new_[4015]_ ;
  assign \new_[3951]_  = ~\new_[4016]_ ;
  assign \new_[3952]_  = ~\new_[4020]_ ;
  assign \new_[3953]_  = ~\new_[4021]_ ;
  assign \new_[3954]_  = ~\new_[4022]_ ;
  assign \new_[3955]_  = ~\new_[4023]_ ;
  assign \new_[3956]_  = ~\new_[4025]_ ;
  assign \new_[3957]_  = ~\new_[4027]_ ;
  assign \new_[3958]_  = ~\new_[4028]_ ;
  assign \new_[3959]_  = ~\new_[4029]_ ;
  assign \new_[3960]_  = ~\new_[4075]_  & ~\new_[1234]_ ;
  assign \new_[3961]_  = ~\new_[4075]_  | ~\new_[1234]_ ;
  assign \new_[3962]_  = ~\new_[4075]_  & ~\new_[1235]_ ;
  assign \new_[3963]_  = ~\new_[4075]_  & ~\new_[1292]_ ;
  assign \new_[3964]_  = ~\new_[4503]_  | ~\new_[4856]_  | ~\new_[4496]_  | ~\new_[4107]_ ;
  assign \new_[3965]_  = ~\new_[4083]_  & ~\new_[1690]_ ;
  assign n1819 = ~\new_[6441]_  & (~\new_[4345]_  | ~\new_[4191]_ );
  assign \new_[3967]_  = ~\new_[4075]_ ;
  assign \new_[3968]_  = ~\new_[4705]_  & ~\new_[4099]_ ;
  assign \new_[3969]_  = ~\new_[4098]_  | ~\new_[4101]_ ;
  assign \new_[3970]_  = ~\new_[4705]_  | ~\new_[4094]_ ;
  assign \new_[3971]_  = ~\new_[4705]_  & ~\new_[4097]_ ;
  assign \new_[3972]_  = ~\new_[4705]_  & ~\new_[4093]_ ;
  assign \new_[3973]_  = ~\new_[4100]_  & ~\new_[4636]_ ;
  assign \new_[3974]_  = ~\new_[5432]_  | ~\new_[4271]_  | ~\new_[6035]_  | ~\new_[6635]_ ;
  assign \new_[3975]_  = ~\new_[4829]_  | ~\new_[5420]_  | ~\new_[5415]_  | ~\new_[4198]_ ;
  assign \new_[3976]_  = ~\new_[6020]_  | (~\new_[4195]_  & ~\new_[6365]_ );
  assign \new_[3977]_  = (~\new_[4197]_  | ~\new_[5865]_ ) & (~\new_[4283]_  | ~\new_[5514]_ );
  assign \new_[3978]_  = \new_[4104]_  & \new_[5700]_ ;
  assign n1814 = ~\new_[4105]_  | (~\new_[6655]_  & ~\new_[6356]_ );
  assign \new_[3980]_  = ~\new_[5366]_  | ~\new_[4104]_  | ~\new_[5189]_ ;
  assign \new_[3981]_  = \new_[2780]_  ^ \new_[4200]_ ;
  assign \new_[3982]_  = ~\new_[4112]_  | ~\new_[4109]_ ;
  assign \new_[3983]_  = ~\new_[4081]_  & (~\new_[5330]_  | ~\new_[5772]_ );
  assign \new_[3984]_  = ~\new_[4110]_  | ~\new_[4974]_ ;
  assign \new_[3985]_  = \new_[4841]_  | \new_[4113]_ ;
  assign \new_[3986]_  = \new_[4371]_  | \new_[6365]_ ;
  assign \new_[3987]_  = ~\new_[5025]_  | ~\new_[4118]_ ;
  assign \new_[3988]_  = ~\new_[5669]_  & (~\new_[4204]_  | ~\new_[5356]_ );
  assign \new_[3989]_  = ~\new_[4119]_  & (~\new_[5237]_  | ~\new_[740]_ );
  assign \new_[3990]_  = ~\new_[4115]_  | ~\new_[5924]_ ;
  assign \new_[3991]_  = (~\new_[4206]_  | ~\new_[6953]_ ) & (~\new_[6509]_  | ~\new_[5959]_ );
  assign \new_[3992]_  = \new_[4120]_  | \new_[5877]_ ;
  assign \new_[3993]_  = \new_[5467]_  ^ \new_[4205]_ ;
  assign \new_[3994]_  = ~\new_[4122]_  | ~\new_[6584]_ ;
  assign \new_[3995]_  = ~\new_[6584]_  | ~\new_[5116]_ ;
  assign \new_[3996]_  = ~\new_[4121]_  & ~\new_[4439]_ ;
  assign \new_[3997]_  = ~\new_[6472]_  | ~\new_[5116]_ ;
  assign \new_[3998]_  = ~\new_[6994]_ ;
  assign \new_[3999]_  = \new_[4133]_  & \new_[4134]_ ;
  assign \new_[4000]_  = ~\new_[4130]_  & ~\new_[5154]_ ;
  assign \new_[4001]_  = ~\new_[7357]_ ;
  assign \new_[4002]_  = ~\new_[7357]_ ;
  assign \new_[4003]_  = ~\new_[4131]_  & ~\new_[5032]_ ;
  assign \new_[4004]_  = (~\new_[4213]_  | ~\new_[4668]_ ) & (~\new_[6472]_  | ~\new_[5969]_ );
  assign \new_[4005]_  = \new_[4219]_  ^ \new_[4217]_ ;
  assign \new_[4006]_  = ~\new_[4933]_  | ~\new_[4138]_  | ~\new_[5721]_ ;
  assign \new_[4007]_  = ~\new_[4062]_ ;
  assign \new_[4008]_  = ~\new_[6513]_  | ~\new_[5116]_ ;
  assign \new_[4009]_  = ~\new_[4265]_  | ~\new_[4852]_  | ~\new_[4532]_  | ~\new_[4521]_ ;
  assign \new_[4010]_  = ~\new_[4141]_  & ~\new_[4603]_ ;
  assign \new_[4011]_  = ~\new_[4607]_  | ~\new_[4611]_  | ~\new_[4142]_  | ~\new_[4224]_ ;
  assign \new_[4012]_  = ~\new_[4136]_  & (~\new_[6070]_  | ~\new_[7208]_ );
  assign \new_[4013]_  = ~\new_[4238]_  | ~\new_[4242]_  | ~\new_[4168]_  | ~\new_[4169]_ ;
  assign \new_[4014]_  = ~\new_[4075]_  | ~\new_[1225]_ ;
  assign \new_[4015]_  = ~\new_[4074]_  | ~\new_[1240]_ ;
  assign \new_[4016]_  = ~\new_[4073]_  & ~\new_[1237]_ ;
  assign \new_[4017]_  = ~\new_[4073]_  | ~\new_[1237]_ ;
  assign \new_[4018]_  = ~\new_[4067]_ ;
  assign \new_[4019]_  = ~\new_[4072]_  & ~\new_[1239]_ ;
  assign \new_[4020]_  = ~\new_[4074]_  & ~\new_[1240]_ ;
  assign \new_[4021]_  = \new_[4072]_  & \new_[1239]_ ;
  assign \new_[4022]_  = ~\new_[4075]_  & ~\new_[1225]_ ;
  assign \new_[4023]_  = ~\new_[4076]_  & ~\new_[1241]_ ;
  assign \new_[4024]_  = ~\new_[4076]_  | ~\new_[1241]_ ;
  assign \new_[4025]_  = ~\new_[4075]_  & ~\new_[1223]_ ;
  assign \new_[4026]_  = ~\new_[4075]_  & ~\new_[1242]_ ;
  assign \new_[4027]_  = \new_[4075]_  & \new_[1242]_ ;
  assign \new_[4028]_  = ~\new_[4075]_  | ~\new_[1223]_ ;
  assign \new_[4029]_  = ~\new_[4075]_  | ~\new_[1294]_ ;
  assign \new_[4030]_  = ~\new_[4075]_  & ~\new_[1294]_ ;
  assign \new_[4031]_  = ~\new_[4075]_  & ~\new_[1233]_ ;
  assign \new_[4032]_  = ~\new_[4196]_  | ~\new_[4386]_  | ~\new_[4412]_ ;
  assign \new_[4033]_  = ~\new_[4077]_  | ~\new_[6272]_ ;
  assign \new_[4034]_  = ~\new_[5173]_  | ~\new_[4329]_  | ~\new_[5194]_  | ~\new_[5335]_ ;
  assign \new_[4035]_  = ~\new_[4705]_  & ~\new_[4188]_ ;
  assign \new_[4036]_  = \new_[4705]_  & \new_[4189]_ ;
  assign \new_[4037]_  = \new_[4705]_  & \new_[4187]_ ;
  assign \new_[4038]_  = \new_[4705]_  & \new_[4190]_ ;
  assign \new_[4039]_  = ~\new_[4192]_  & ~\new_[5486]_ ;
  assign \new_[4040]_  = ~\new_[5213]_  | ~\new_[4979]_  | ~\new_[4203]_  | ~\new_[4526]_ ;
  assign \new_[4041]_  = ~\new_[4082]_ ;
  assign \new_[4042]_  = (~\new_[4272]_  | ~\new_[5969]_ ) & (~\new_[5522]_  | ~\new_[4867]_ );
  assign \new_[4043]_  = ~\new_[4193]_  | ~\new_[3029]_ ;
  assign \new_[4044]_  = ~\new_[4096]_ ;
  assign \new_[4045]_  = ~\new_[4892]_  | ~\new_[4767]_  | ~\new_[4199]_  | ~\new_[6016]_ ;
  assign \new_[4046]_  = ~\new_[4202]_  | ~\new_[7155]_ ;
  assign \new_[4047]_  = ~\new_[4194]_  | ~\new_[4270]_ ;
  assign \new_[4048]_  = ~\new_[4194]_  | (~\new_[4427]_  & ~\new_[4833]_ );
  assign \new_[4049]_  = ~\new_[5097]_  | ~\new_[5373]_  | ~\new_[5366]_  | ~\new_[4267]_ ;
  assign \new_[4050]_  = (~\new_[5542]_  | ~\new_[5116]_ ) & (~\new_[5771]_  | ~\new_[6359]_ );
  assign \new_[4051]_  = (~\new_[4989]_  | ~\new_[5443]_ ) & (~\new_[4308]_  | ~\new_[7121]_ );
  assign \new_[4052]_  = ~\new_[4081]_ ;
  assign \new_[4053]_  = \new_[5506]_  ^ \new_[4291]_ ;
  assign \new_[4054]_  = ~\new_[4206]_  | ~\new_[6952]_ ;
  assign \new_[4055]_  = \new_[5346]_  | \new_[4205]_ ;
  assign \new_[4056]_  = ~\new_[4205]_  | ~\new_[5459]_ ;
  assign \new_[4057]_  = ~\new_[6084]_  | ~\new_[5688]_ ;
  assign \new_[4058]_  = ~\new_[6935]_  & (~\new_[4295]_  | ~\new_[5144]_ );
  assign \new_[4059]_  = ~\new_[6471]_  | (~\new_[4307]_  & ~\new_[4672]_ );
  assign \new_[4060]_  = ~\new_[4592]_  | ~\new_[4670]_  | ~\new_[4216]_  | ~\new_[4911]_ ;
  assign \new_[4061]_  = ~\new_[4210]_  & (~\new_[4761]_  | ~\new_[5910]_ );
  assign \new_[4062]_  = ~\new_[4132]_ ;
  assign \new_[4063]_  = ~\new_[4961]_  | ~\new_[4786]_  | ~\new_[4907]_  | ~\new_[4267]_ ;
  assign \new_[4064]_  = \new_[1293]_  ^ \new_[4225]_ ;
  assign \new_[4065]_  = ~\new_[4135]_ ;
  assign \new_[4066]_  = ~\new_[4151]_  & ~\new_[1238]_ ;
  assign \new_[4067]_  = ~\new_[4151]_  | ~\new_[1238]_ ;
  assign \new_[4068]_  = ~\new_[4178]_  | ~\new_[4179]_ ;
  assign \new_[4069]_  = ~\new_[4152]_  | ~\new_[4548]_ ;
  assign \new_[4070]_  = ~\new_[4275]_  | ~\new_[4259]_  | ~\new_[4341]_ ;
  assign \new_[4071]_  = ~\new_[4694]_  | ~\new_[5620]_  | ~\new_[4284]_  | ~\new_[5850]_ ;
  assign \new_[4072]_  = ~\new_[4263]_  | ~\new_[4320]_ ;
  assign \new_[4073]_  = ~\new_[4262]_  | ~\new_[4320]_ ;
  assign \new_[4074]_  = ~\new_[4320]_  | (~\new_[4589]_  & ~\new_[6572]_ );
  assign \new_[4075]_  = ~\new_[4261]_  | ~\new_[4320]_ ;
  assign \new_[4076]_  = ~\new_[4264]_  | ~\new_[4320]_ ;
  assign \new_[4077]_  = ~\new_[4429]_  | ~\new_[4522]_  | ~\new_[5167]_  | ~\new_[4524]_ ;
  assign \new_[4078]_  = \new_[758]_  ? \new_[4966]_  : \new_[4313]_ ;
  assign \new_[4079]_  = \new_[759]_  ? \new_[4966]_  : \new_[4338]_ ;
  assign \new_[4080]_  = ~\new_[5111]_  & ~\new_[4339]_ ;
  assign \new_[4081]_  = \new_[5617]_  & \new_[5116]_ ;
  assign \new_[4082]_  = (~\new_[4367]_  | ~\new_[5969]_ ) & (~\new_[4805]_  | ~\new_[6193]_ );
  assign \new_[4083]_  = (~\new_[4807]_  | ~\new_[5969]_ ) & (~\new_[5574]_  | ~\new_[6193]_ );
  assign \new_[4084]_  = ~\new_[4268]_  & (~\new_[6961]_  | ~\new_[5772]_ );
  assign \new_[4085]_  = \new_[3626]_  ? \new_[5247]_  : \new_[4347]_ ;
  assign \new_[4086]_  = \new_[3638]_  ? \new_[5247]_  : \new_[4346]_ ;
  assign \new_[4087]_  = \new_[3603]_  ? \new_[5247]_  : \new_[4348]_ ;
  assign \new_[4088]_  = \new_[3639]_  ? \new_[5247]_  : \new_[4352]_ ;
  assign \new_[4089]_  = \new_[3606]_  ? \new_[5247]_  : \new_[4349]_ ;
  assign \new_[4090]_  = \new_[3600]_  ? \new_[5247]_  : \new_[4350]_ ;
  assign \new_[4091]_  = \new_[3621]_  ? \new_[5247]_  : \new_[4351]_ ;
  assign \new_[4092]_  = \new_[3615]_  ? \new_[5247]_  : \new_[4353]_ ;
  assign \new_[4093]_  = ~\new_[4187]_ ;
  assign \new_[4094]_  = ~\new_[4188]_ ;
  assign \new_[4095]_  = ~\new_[4273]_  | ~\new_[6640]_ ;
  assign \new_[4096]_  = \new_[5124]_  & \new_[4271]_ ;
  assign \new_[4097]_  = ~\new_[4189]_ ;
  assign \new_[4098]_  = ~\new_[4274]_  | ~\new_[5995]_ ;
  assign \new_[4099]_  = ~\new_[4190]_ ;
  assign \new_[4100]_  = \new_[5010]_  | \new_[4451]_  | \new_[6011]_  | \new_[5568]_ ;
  assign \new_[4101]_  = ~\new_[4277]_  | ~\new_[5995]_ ;
  assign \new_[4102]_  = ~\new_[4280]_  & (~\new_[5518]_  | ~\new_[6405]_ );
  assign \new_[4103]_  = ~\new_[6080]_  | ~\new_[7162]_  | ~\new_[4287]_  | ~\new_[6034]_ ;
  assign \new_[4104]_  = \new_[4267]_  & \new_[5335]_ ;
  assign \new_[4105]_  = ~\new_[5969]_  | ~\new_[6342]_  | ~\new_[5560]_ ;
  assign \new_[4106]_  = ~\new_[5850]_  | ~\new_[4442]_  | ~\new_[4435]_  | ~\new_[4856]_ ;
  assign \new_[4107]_  = (~\new_[5695]_  | ~\new_[5209]_ ) & (~\new_[4371]_  | ~\new_[5362]_ );
  assign \new_[4108]_  = (~\new_[5695]_  | ~\new_[5147]_ ) & (~\new_[4371]_  | ~\new_[5609]_ );
  assign \new_[4109]_  = ~\new_[5782]_  | ~\new_[4371]_ ;
  assign \new_[4110]_  = ~\new_[5438]_  | ~\new_[5116]_ ;
  assign \new_[4111]_  = ~\new_[5656]_  | ~\new_[5116]_ ;
  assign \new_[4112]_  = ~\new_[5895]_  | ~\new_[4371]_ ;
  assign \new_[4113]_  = \new_[4288]_  & \new_[7121]_ ;
  assign \new_[4114]_  = ~\new_[5786]_  | ~\new_[5116]_ ;
  assign \new_[4115]_  = ~\new_[5884]_  & ~\new_[5116]_ ;
  assign \new_[4116]_  = ~\new_[4207]_ ;
  assign \new_[4117]_  = ~\new_[4288]_  | ~\new_[5924]_ ;
  assign \new_[4118]_  = ~\new_[5506]_  & ~\new_[4291]_ ;
  assign \new_[4119]_  = ~\new_[4289]_  & ~\new_[740]_ ;
  assign \new_[4120]_  = \new_[4374]_  ? \new_[740]_  : \new_[5355]_ ;
  assign \new_[4121]_  = ~\new_[4375]_  | ~\new_[4376]_  | ~\new_[5737]_ ;
  assign \new_[4122]_  = (~\new_[4377]_  | ~\new_[6625]_ ) & (~\new_[4875]_  | ~\new_[740]_ );
  assign \new_[4123]_  = ~\new_[4290]_  & (~\new_[4438]_  | ~\new_[6952]_ );
  assign \new_[4124]_  = ~\new_[5453]_  | ~\new_[4440]_  | ~\new_[4687]_  | ~\new_[4566]_ ;
  assign \new_[4125]_  = \new_[4560]_  ? \new_[1623]_  : \new_[4321]_ ;
  assign \new_[4126]_  = \\i_tv80_core_RegAddrC_reg[2] ;
  assign \new_[4127]_  = ~\new_[4293]_  & ~\new_[4708]_ ;
  assign \new_[4128]_  = (~\new_[4378]_  | ~\new_[5894]_ ) & (~\new_[5399]_  | ~\new_[5937]_ );
  assign \new_[4129]_  = ~\new_[4294]_  & ~\new_[4781]_ ;
  assign \new_[4130]_  = ~\new_[5080]_  | ~\new_[5299]_  | ~\new_[4297]_  | ~\new_[4928]_ ;
  assign \new_[4131]_  = ~\new_[4935]_  | ~\new_[4450]_  | ~\new_[4913]_  | ~\new_[5386]_ ;
  assign \new_[4132]_  = ~\new_[4634]_  & (~\new_[4311]_  | ~\new_[5969]_ );
  assign \new_[4133]_  = ~\new_[4225]_  & ~\new_[6631]_ ;
  assign \new_[4134]_  = ~\new_[4226]_  | ~\new_[6592]_ ;
  assign \new_[4135]_  = ~\new_[4226]_  & ~\new_[6592]_ ;
  assign \new_[4136]_  = ~\new_[4315]_  | ~\new_[5194]_  | ~\new_[5282]_ ;
  assign \new_[4137]_  = ~\new_[4247]_  | ~\new_[4248]_ ;
  assign \new_[4138]_  = ~\new_[4220]_  & ~\new_[4519]_ ;
  assign \new_[4139]_  = \new_[4505]_  | \new_[4518]_  | \new_[7232]_  | \new_[4333]_ ;
  assign \new_[4140]_  = ~\new_[5690]_  | ~\new_[5395]_  | ~\new_[4222]_  | ~\new_[4823]_ ;
  assign \new_[4141]_  = ~\new_[4673]_  | ~\new_[4416]_  | ~\new_[4835]_  | ~\new_[4786]_ ;
  assign \new_[4142]_  = ~\new_[4410]_  & ~\new_[4221]_ ;
  assign \new_[4143]_  = ~\new_[4223]_  & ~\new_[4323]_ ;
  assign \new_[4144]_  = ~\new_[7440]_  & (~\new_[4328]_  | ~\new_[6799]_ );
  assign \new_[4145]_  = ~\new_[7440]_  & (~\new_[4326]_  | ~\new_[6809]_ );
  assign \new_[4146]_  = ~\new_[7440]_  & (~\new_[4322]_  | ~\new_[6787]_ );
  assign \new_[4147]_  = ~\new_[7440]_  & (~\new_[4327]_  | ~\new_[6793]_ );
  assign \new_[4148]_  = \new_[4330]_  & \new_[4966]_ ;
  assign \new_[4149]_  = ~\new_[4582]_  & ~\new_[4318]_ ;
  assign \new_[4150]_  = ~\new_[4480]_  & (~\new_[5710]_  | ~\new_[5116]_ );
  assign \new_[4151]_  = ~\new_[4317]_  | ~\new_[4320]_ ;
  assign \new_[4152]_  = ~\new_[4325]_  & (~\new_[5296]_  | ~\new_[6284]_ );
  assign \new_[4153]_  = (~\new_[433]_  | ~\new_[4409]_ ) & (~\new_[432]_  | ~\new_[4499]_ );
  assign \new_[4154]_  = (~\new_[520]_  | ~\new_[4409]_ ) & (~\new_[540]_  | ~\new_[4499]_ );
  assign \new_[4155]_  = (~\new_[771]_  | ~\new_[4409]_ ) & (~\new_[796]_  | ~\new_[4499]_ );
  assign \new_[4156]_  = (~\new_[686]_  | ~\new_[4494]_ ) & (~\new_[734]_  | ~\new_[4408]_ );
  assign \new_[4157]_  = (~\new_[772]_  | ~\new_[4494]_ ) & (~\new_[773]_  | ~\new_[4408]_ );
  assign \new_[4158]_  = (~\new_[797]_  | ~\new_[4494]_ ) & (~\new_[791]_  | ~\new_[4408]_ );
  assign \new_[4159]_  = (~\new_[578]_  | ~\new_[4409]_ ) & (~\new_[560]_  | ~\new_[4499]_ );
  assign \new_[4160]_  = (~\new_[663]_  | ~\new_[4494]_ ) & (~\new_[664]_  | ~\new_[4408]_ );
  assign \new_[4161]_  = (~\new_[779]_  | ~\new_[4494]_ ) & (~\new_[780]_  | ~\new_[4408]_ );
  assign \new_[4162]_  = (~\new_[434]_  | ~\new_[4494]_ ) & (~\new_[435]_  | ~\new_[4408]_ );
  assign \new_[4163]_  = (~\new_[6612]_  | ~\new_[4409]_ ) & (~\new_[6639]_  | ~\new_[4499]_ );
  assign \new_[4164]_  = (~\new_[6597]_  | ~\new_[4494]_ ) & (~\new_[6607]_  | ~\new_[4408]_ );
  assign \new_[4165]_  = (~\new_[665]_  | ~\new_[4409]_ ) & (~\new_[646]_  | ~\new_[4499]_ );
  assign \new_[4166]_  = (~\new_[6496]_  | ~\new_[4409]_ ) & (~\new_[6587]_  | ~\new_[4499]_ );
  assign \new_[4167]_  = (~\new_[6512]_  | ~\new_[4494]_ ) & (~\new_[6665]_  | ~\new_[4408]_ );
  assign \new_[4168]_  = (~\new_[657]_  | ~\new_[4494]_ ) & (~\new_[658]_  | ~\new_[4408]_ );
  assign \new_[4169]_  = (~\new_[656]_  | ~\new_[4409]_ ) & (~\new_[655]_  | ~\new_[4499]_ );
  assign \new_[4170]_  = (~\new_[6672]_  | ~\new_[4409]_ ) & (~\new_[6657]_  | ~\new_[4499]_ );
  assign \new_[4171]_  = (~\new_[7513]_  | ~\new_[4494]_ ) & (~\new_[6673]_  | ~\new_[4408]_ );
  assign \new_[4172]_  = (~\new_[531]_  | ~\new_[4409]_ ) & (~\new_[535]_  | ~\new_[4499]_ );
  assign \new_[4173]_  = (~\new_[532]_  | ~\new_[4494]_ ) & (~\new_[533]_  | ~\new_[4408]_ );
  assign \new_[4174]_  = (~\new_[6482]_  | ~\new_[4494]_ ) & (~\new_[6652]_  | ~\new_[4408]_ );
  assign \new_[4175]_  = (~\new_[6559]_  | ~\new_[4409]_ ) & (~\new_[6599]_  | ~\new_[4499]_ );
  assign \new_[4176]_  = (~\new_[4499]_  | ~\new_[571]_ ) & (~\new_[4409]_  | ~\new_[572]_ );
  assign \new_[4177]_  = (~\new_[4408]_  | ~\new_[562]_ ) & (~\new_[4494]_  | ~\new_[573]_ );
  assign \new_[4178]_  = (~n319 | ~\new_[4499]_ ) & (~n324 | ~\new_[4409]_ );
  assign \new_[4179]_  = (~n329 | ~\new_[4494]_ ) & (~n334 | ~\new_[4408]_ );
  assign \new_[4180]_  = (~\new_[579]_  | ~\new_[4494]_ ) & (~\new_[580]_  | ~\new_[4408]_ );
  assign \new_[4181]_  = (~\new_[6602]_  | ~\new_[4409]_ ) & (~\new_[733]_  | ~\new_[4499]_ );
  assign \new_[4182]_  = (~\new_[778]_  | ~\new_[4409]_ ) & (~\new_[737]_  | ~\new_[4499]_ );
  assign \new_[4183]_  = (~\new_[790]_  | ~\new_[4409]_ ) & (~\new_[789]_  | ~\new_[4499]_ );
  assign \new_[4184]_  = (~\new_[542]_  | ~\new_[4494]_ ) & (~\new_[543]_  | ~\new_[4408]_ );
  assign \new_[4185]_  = ~\new_[4267]_ ;
  assign \new_[4186]_  = ~\new_[4938]_  & ~\new_[4344]_ ;
  assign \new_[4187]_  = ~\new_[4839]_  & ~\new_[4356]_ ;
  assign \new_[4188]_  = ~\new_[4839]_  | ~\new_[4356]_ ;
  assign \new_[4189]_  = \new_[4939]_  & \new_[4356]_ ;
  assign \new_[4190]_  = ~\new_[4939]_  & ~\new_[4356]_ ;
  assign \new_[4191]_  = (~\new_[4436]_  | ~\new_[4598]_ ) & (~\new_[5168]_  | ~\new_[4639]_ );
  assign \new_[4192]_  = (~\new_[4538]_  | ~\new_[753]_ ) & (~\new_[4428]_  | ~\new_[3285]_ );
  assign \new_[4193]_  = ~\new_[4270]_ ;
  assign \new_[4194]_  = ~\new_[4271]_ ;
  assign \new_[4195]_  = ~\new_[4430]_  | (~\new_[4431]_  & ~\new_[6635]_ );
  assign \new_[4196]_  = ~\new_[4365]_  & (~\new_[5777]_  | ~\new_[6128]_ );
  assign \new_[4197]_  = ~\new_[5348]_  | (~\new_[7209]_  & ~\new_[5578]_ );
  assign \new_[4198]_  = (~\new_[7015]_  | ~\new_[6359]_ ) & (~\new_[6961]_  | ~\new_[5116]_ );
  assign \new_[4199]_  = ~\new_[5015]_  & (~\new_[7208]_  | ~\new_[5463]_ );
  assign \new_[4200]_  = ~\new_[5772]_  | ~\new_[6113]_  | ~\new_[4858]_  | ~\new_[5969]_ ;
  assign \new_[4201]_  = ~\new_[5712]_  | ~\new_[5969]_ ;
  assign \new_[4202]_  = ~\new_[5924]_  | ~\new_[5688]_ ;
  assign \new_[4203]_  = ~\new_[6227]_  | ~\new_[5514]_  | ~\new_[7208]_ ;
  assign \new_[4204]_  = ~\new_[4308]_ ;
  assign \new_[4205]_  = \new_[4437]_  ? \new_[740]_  : \new_[5006]_ ;
  assign \new_[4206]_  = \new_[5905]_  ^ \new_[4438]_ ;
  assign \new_[4207]_  = ~\new_[5903]_  & ~\new_[6031]_ ;
  assign \new_[4208]_  = ~\new_[4754]_  & (~\new_[4439]_  | ~\new_[6589]_ );
  assign \new_[4209]_  = \new_[4453]_  | \new_[7349]_  | \new_[5531]_  | \new_[5661]_ ;
  assign \new_[4210]_  = ~\new_[5335]_  | ~\new_[5179]_  | ~\new_[4384]_ ;
  assign \new_[4211]_  = ~\new_[7440]_  & (~\new_[4459]_  | ~\new_[4391]_ );
  assign \new_[4212]_  = ~\new_[6471]_  | (~\new_[4467]_  & ~\new_[4446]_ );
  assign \new_[4213]_  = ~\new_[4381]_  & ~\new_[4906]_ ;
  assign \new_[4214]_  = ~\new_[7440]_  & (~\new_[4458]_  | ~\new_[4390]_ );
  assign \new_[4215]_  = ~\new_[7440]_  & (~\new_[4462]_  | ~\new_[4395]_ );
  assign \new_[4216]_  = ~\new_[4382]_  & (~\new_[5214]_  | ~\new_[5455]_ );
  assign \new_[4217]_  = \new_[4387]_  ^ \new_[4587]_ ;
  assign n1824 = \new_[4126]_  ? \new_[6326]_  : \new_[4485]_ ;
  assign \new_[4219]_  = \new_[4488]_  ^ \new_[4586]_ ;
  assign \new_[4220]_  = ~\new_[5872]_  | ~\new_[5507]_  | ~\new_[4398]_  | ~\new_[4822]_ ;
  assign \new_[4221]_  = ~\new_[4523]_  | ~\new_[4392]_  | ~\new_[4827]_ ;
  assign \new_[4222]_  = ~\new_[4484]_  & ~\new_[4389]_ ;
  assign \new_[4223]_  = ~\new_[5988]_  | ~\new_[7263]_  | ~\new_[4502]_ ;
  assign \new_[4224]_  = ~\new_[4516]_  & ~\new_[4396]_ ;
  assign \new_[4225]_  = ~\new_[4388]_  & (~\new_[4666]_  | ~\new_[4560]_ );
  assign \new_[4226]_  = ~\new_[4394]_  & (~\new_[4500]_  | ~\new_[4554]_ );
  assign \new_[4227]_  = (~\new_[776]_  | ~\new_[4498]_ ) & (~\new_[777]_  | ~\new_[4495]_ );
  assign \new_[4228]_  = (~\new_[774]_  | ~\new_[4493]_ ) & (~\new_[775]_  | ~\new_[4497]_ );
  assign \new_[4229]_  = (~\new_[428]_  | ~\new_[4493]_ ) & (~\new_[429]_  | ~\new_[4497]_ );
  assign \new_[4230]_  = (~\new_[6491]_  | ~\new_[4493]_ ) & (~\new_[6618]_  | ~\new_[4497]_ );
  assign \new_[4231]_  = (~\new_[530]_  | ~\new_[4498]_ ) & (~\new_[534]_  | ~\new_[4495]_ );
  assign \new_[4232]_  = (~\new_[6642]_  | ~\new_[4498]_ ) & (~\new_[6556]_  | ~\new_[4495]_ );
  assign \new_[4233]_  = (~\new_[574]_  | ~\new_[4493]_ ) & (~\new_[575]_  | ~\new_[4497]_ );
  assign \new_[4234]_  = (~\new_[576]_  | ~\new_[4498]_ ) & (~\new_[577]_  | ~\new_[4495]_ );
  assign \new_[4235]_  = (~\new_[538]_  | ~\new_[4498]_ ) & (~\new_[539]_  | ~\new_[4495]_ );
  assign \new_[4236]_  = (~\new_[769]_  | ~\new_[4498]_ ) & (~\new_[770]_  | ~\new_[4495]_ );
  assign \new_[4237]_  = (~\new_[430]_  | ~\new_[4498]_ ) & (~\new_[431]_  | ~\new_[4495]_ );
  assign \new_[4238]_  = (~\new_[650]_  | ~\new_[4493]_ ) & (~\new_[652]_  | ~\new_[4497]_ );
  assign \new_[4239]_  = (~\new_[730]_  | ~\new_[4493]_ ) & (~\new_[731]_  | ~\new_[4497]_ );
  assign \new_[4240]_  = (~\new_[661]_  | ~\new_[4498]_ ) & (~\new_[662]_  | ~\new_[4495]_ );
  assign \new_[4241]_  = (~\new_[6645]_  | ~\new_[4498]_ ) & (~\new_[6641]_  | ~\new_[4495]_ );
  assign \new_[4242]_  = (~\new_[653]_  | ~\new_[4498]_ ) & (~\new_[654]_  | ~\new_[4495]_ );
  assign \new_[4243]_  = (~\new_[6644]_  | ~\new_[4493]_ ) & (~\new_[6566]_  | ~\new_[4497]_ );
  assign \new_[4244]_  = (~\new_[528]_  | ~\new_[4493]_ ) & (~\new_[529]_  | ~\new_[4497]_ );
  assign \new_[4245]_  = (~\new_[6598]_  | ~\new_[4493]_ ) & (~\new_[6590]_  | ~\new_[4497]_ );
  assign \new_[4246]_  = (~\new_[4497]_  | ~\new_[568]_ ) & (~\new_[4493]_  | ~\new_[567]_ );
  assign \new_[4247]_  = (~n314 | ~\new_[4495]_ ) & (~n309 | ~\new_[4498]_ );
  assign \new_[4248]_  = (~n304 | ~\new_[4497]_ ) & (~n299 | ~\new_[4493]_ );
  assign \new_[4249]_  = (~\new_[787]_  | ~\new_[4498]_ ) & (~\new_[788]_  | ~\new_[4495]_ );
  assign \new_[4250]_  = (~\new_[6615]_  | ~\new_[4498]_ ) & (~\new_[6583]_  | ~\new_[4495]_ );
  assign \new_[4251]_  = (~\new_[785]_  | ~\new_[4493]_ ) & (~\new_[786]_  | ~\new_[4497]_ );
  assign \new_[4252]_  = (~\new_[659]_  | ~\new_[4493]_ ) & (~\new_[660]_  | ~\new_[4497]_ );
  assign \new_[4253]_  = (~\new_[735]_  | ~\new_[4498]_ ) & (~\new_[732]_  | ~\new_[4495]_ );
  assign \new_[4254]_  = (~\new_[6564]_  | ~\new_[4498]_ ) & (~\new_[6660]_  | ~\new_[4495]_ );
  assign \new_[4255]_  = (~\new_[4495]_  | ~\new_[570]_ ) & (~\new_[4498]_  | ~\new_[569]_ );
  assign \new_[4256]_  = (~\new_[767]_  | ~\new_[4493]_ ) & (~\new_[768]_  | ~\new_[4497]_ );
  assign \new_[4257]_  = (~\new_[536]_  | ~\new_[4493]_ ) & (~\new_[537]_  | ~\new_[4497]_ );
  assign \new_[4258]_  = (~\new_[6633]_  | ~\new_[4493]_ ) & (~\new_[6627]_  | ~\new_[4497]_ );
  assign \new_[4259]_  = (~\new_[5416]_  | ~\new_[5772]_ ) & (~\new_[4897]_  | ~\new_[5772]_ );
  assign \new_[4260]_  = ~\new_[4407]_  & (~\new_[4606]_  | ~\new_[6084]_ );
  assign \new_[4261]_  = ~\new_[4500]_  | ~\new_[4556]_ ;
  assign \new_[4262]_  = ~\new_[4500]_  | ~\new_[4557]_ ;
  assign \new_[4263]_  = ~\new_[4500]_  | ~\new_[4558]_ ;
  assign \new_[4264]_  = ~\new_[4500]_  | ~\new_[4549]_ ;
  assign \new_[4265]_  = ~\new_[4324]_ ;
  assign \new_[4266]_  = (~\new_[4605]_  | ~\new_[5772]_ ) & (~\new_[4912]_  | ~\new_[5772]_ );
  assign \new_[4267]_  = ~\new_[7200]_  | ~\new_[5447]_ ;
  assign \new_[4268]_  = ~\new_[5636]_  | ~\new_[4420]_  | ~\new_[5448]_ ;
  assign \new_[4269]_  = ~\new_[4421]_  & (~\new_[4918]_  | ~\new_[5772]_ );
  assign \new_[4270]_  = \new_[4427]_  & \new_[4737]_ ;
  assign \new_[4271]_  = ~\new_[4427]_  & ~\new_[4737]_ ;
  assign \new_[4272]_  = ~\new_[4899]_  | ~\new_[4432]_  | ~\new_[4987]_ ;
  assign \new_[4273]_  = ~\new_[4427]_  | ~\new_[4833]_ ;
  assign \new_[4274]_  = ~\new_[5969]_  & (~\new_[4628]_  | ~\new_[6193]_ );
  assign \new_[4275]_  = ~\new_[5293]_  & (~\new_[5647]_  | ~\new_[5772]_ );
  assign \new_[4276]_  = ~\new_[4434]_  & ~\new_[4645]_ ;
  assign \new_[4277]_  = ~\new_[5969]_  & (~\new_[5339]_  | ~\new_[6193]_ );
  assign \new_[4278]_  = ~\new_[5947]_  & (~\new_[4985]_  | ~\new_[5356]_ );
  assign \new_[4279]_  = ~\new_[5876]_  | ~\new_[6171]_  | ~\new_[7208]_  | ~\new_[5996]_ ;
  assign \new_[4280]_  = ~\new_[4546]_  | ~\new_[4433]_ ;
  assign \new_[4281]_  = \new_[4435]_  | \new_[6495]_ ;
  assign \new_[4282]_  = ~\new_[7200]_  & ~\new_[5962]_ ;
  assign \new_[4283]_  = ~\new_[7209]_  & ~\new_[7550]_ ;
  assign \new_[4284]_  = \new_[5663]_  & \new_[4442]_ ;
  assign \new_[4285]_  = \new_[6128]_  ? \new_[5680]_  : \di[5] ;
  assign \new_[4286]_  = \new_[5772]_  ? \new_[5680]_  : \di[3] ;
  assign \new_[4287]_  = ~\new_[4372]_ ;
  assign \new_[4288]_  = ~\new_[6143]_  & ~\new_[5116]_ ;
  assign \new_[4289]_  = (~\new_[5702]_  | ~\new_[4551]_ ) & (~\new_[4770]_  | ~\new_[5454]_ );
  assign \new_[4290]_  = ~\new_[4438]_  & ~\new_[5842]_ ;
  assign \new_[4291]_  = ~\new_[5905]_  | ~\new_[4438]_ ;
  assign \new_[4292]_  = ~\new_[4316]_ ;
  assign \new_[4293]_  = ~\new_[4562]_  | ~\new_[6013]_  | ~\new_[5047]_ ;
  assign \new_[4294]_  = ~\new_[5410]_  | ~\new_[5414]_  | ~\new_[4567]_  | ~\new_[5898]_ ;
  assign \new_[4295]_  = ~\new_[5517]_  & ~\new_[4445]_ ;
  assign \new_[4296]_  = ~\new_[7440]_  & (~\new_[4460]_  | ~\new_[4473]_ );
  assign \new_[4297]_  = ~\new_[4452]_  & ~\new_[5447]_ ;
  assign \new_[4298]_  = ~\new_[7440]_  & (~\new_[4454]_  | ~\new_[4471]_ );
  assign \new_[4299]_  = ~\new_[7440]_  & (~\new_[4456]_  | ~\new_[7439]_ );
  assign \new_[4300]_  = ~\new_[7440]_  & (~\new_[4457]_  | ~\new_[4472]_ );
  assign \new_[4301]_  = ~\new_[7440]_  & (~\new_[4461]_  | ~\new_[4572]_ );
  assign \new_[4302]_  = ~\new_[7440]_  & (~\new_[4463]_  | ~\new_[4475]_ );
  assign \new_[4303]_  = ~\new_[7440]_  & (~\new_[4464]_  | ~\new_[4477]_ );
  assign \new_[4304]_  = ~\new_[7440]_  & (~\new_[4465]_  | ~\new_[4478]_ );
  assign \new_[4305]_  = ~\new_[7440]_  & (~\new_[4466]_  | ~\new_[4479]_ );
  assign \new_[4306]_  = ~\new_[5264]_  & ~\new_[4449]_ ;
  assign \new_[4307]_  = ~\new_[4571]_  | ~\new_[5280]_  | ~\new_[5694]_  | ~\new_[5441]_ ;
  assign \new_[4308]_  = ~\new_[6400]_  | ~\new_[5688]_ ;
  assign \new_[4309]_  = ~\new_[4385]_  & (~\new_[5426]_  | ~\new_[5455]_ );
  assign \new_[4310]_  = ~\new_[7233]_  | ~\new_[7236]_  | ~\new_[4476]_  | ~\new_[5170]_ ;
  assign \new_[4311]_  = ~\new_[4483]_  | (~\new_[5411]_  & ~\new_[5356]_ );
  assign \new_[4312]_  = ~\new_[4486]_  | ~\new_[6040]_ ;
  assign \new_[4313]_  = \new_[758]_  ? \new_[4965]_  : \new_[4616]_ ;
  assign \new_[4314]_  = ~\new_[4718]_  | ~\new_[4899]_  | ~\new_[6915]_  | ~\new_[4979]_ ;
  assign \new_[4315]_  = ~\new_[4504]_  & (~\new_[5379]_  | ~\new_[7208]_ );
  assign \new_[4316]_  = \new_[4388]_ ;
  assign \new_[4317]_  = ~\new_[4500]_  | ~\new_[4553]_ ;
  assign \new_[4318]_  = ~\new_[4741]_  | ~\new_[5636]_  | ~\new_[5201]_  | ~\new_[4846]_ ;
  assign \new_[4319]_  = ~\new_[4393]_ ;
  assign \new_[4320]_  = ~\new_[4394]_ ;
  assign \new_[4321]_  = ~\new_[4874]_  | ~\new_[4749]_  | ~\new_[4777]_  | ~\new_[4691]_ ;
  assign \new_[4322]_  = ~\new_[4397]_ ;
  assign \new_[4323]_  = ~\new_[4709]_  | ~\new_[4710]_  | ~\new_[4811]_  | ~\new_[4968]_ ;
  assign \new_[4324]_  = ~\new_[6113]_  & (~\new_[4604]_  | ~\new_[6034]_ );
  assign \new_[4325]_  = ~\new_[4824]_  | ~\new_[5700]_  | ~\new_[4513]_  | ~\new_[5580]_ ;
  assign \new_[4326]_  = ~\new_[4399]_ ;
  assign \new_[4327]_  = ~\new_[4400]_ ;
  assign \new_[4328]_  = ~\new_[4401]_ ;
  assign \new_[4329]_  = ~\new_[4501]_  & (~\new_[5608]_  | ~\new_[5772]_ );
  assign \new_[4330]_  = ~\new_[4534]_  | (~\new_[4965]_  & ~\new_[6584]_ );
  assign \new_[4331]_  = ~\new_[6031]_  & (~\new_[4914]_  | ~\new_[5693]_ );
  assign \new_[4332]_  = (~\new_[4605]_  | ~\new_[6128]_ ) & (~\new_[4912]_  | ~\new_[6128]_ );
  assign \new_[4333]_  = ~\new_[4684]_  | ~\new_[5507]_  | ~\new_[4688]_  | ~\new_[5026]_ ;
  assign \new_[4334]_  = ~\new_[4915]_  | ~\new_[5116]_ ;
  assign \new_[4335]_  = ~\new_[4746]_  | ~\new_[4964]_  | ~\new_[4922]_  | ~\new_[4825]_ ;
  assign \new_[4336]_  = ~\new_[5058]_  | ~\new_[4515]_  | ~\new_[5389]_ ;
  assign \new_[4337]_  = ~\new_[4512]_  & (~\new_[6070]_  | ~\new_[6284]_ );
  assign \new_[4338]_  = \new_[759]_  ? \new_[4965]_  : \new_[4617]_ ;
  assign \new_[4339]_  = ~\new_[4413]_ ;
  assign \new_[4340]_  = ~\new_[4851]_  | ~\new_[4537]_  | ~\new_[5218]_ ;
  assign \new_[4341]_  = ~\new_[5055]_  | ~\new_[5772]_ ;
  assign \new_[4342]_  = ~\new_[4415]_ ;
  assign \new_[4343]_  = \new_[4535]_  & \new_[4746]_ ;
  assign \new_[4344]_  = ~\new_[4418]_ ;
  assign \new_[4345]_  = \new_[4541]_  | \new_[4920]_ ;
  assign \new_[4346]_  = \new_[762]_  ? \new_[4627]_  : \new_[3638]_ ;
  assign \new_[4347]_  = \new_[736]_  ? \new_[4627]_  : \new_[3626]_ ;
  assign \new_[4348]_  = \new_[761]_  ? \new_[4627]_  : \new_[3603]_ ;
  assign \new_[4349]_  = \new_[763]_  ? \new_[4627]_  : \new_[3606]_ ;
  assign \new_[4350]_  = \new_[759]_  ? \new_[4627]_  : \new_[3600]_ ;
  assign \new_[4351]_  = \new_[760]_  ? \new_[4627]_  : \new_[3621]_ ;
  assign \new_[4352]_  = \new_[758]_  ? \new_[4627]_  : \new_[3639]_ ;
  assign \new_[4353]_  = \new_[753]_  ? \new_[4627]_  : \new_[3615]_ ;
  assign \new_[4354]_  = \new_[5284]_  & \new_[5116]_ ;
  assign \new_[4355]_  = ~\new_[4542]_  & (~\new_[5092]_  | ~\new_[1247]_ );
  assign \new_[4356]_  = (~\new_[6461]_  & ~\new_[6034]_  & ~\new_[6113]_ ) | (~\new_[6113]_  & ~\new_[4762]_  & ~\new_[6461]_ );
  assign \new_[4357]_  = ~\new_[4536]_  | ~\new_[3626]_ ;
  assign \new_[4358]_  = ~\new_[4536]_  | ~\new_[3603]_ ;
  assign \new_[4359]_  = ~\new_[4536]_  | ~\new_[3639]_ ;
  assign \new_[4360]_  = ~\new_[4536]_  | ~\new_[3606]_ ;
  assign \new_[4361]_  = ~\new_[4536]_  | ~\new_[3638]_ ;
  assign \new_[4362]_  = ~\new_[4536]_  | ~\new_[3600]_ ;
  assign \new_[4363]_  = ~\new_[4536]_  | ~\new_[3621]_ ;
  assign \new_[4364]_  = ~\new_[4536]_  | ~\new_[3615]_ ;
  assign \new_[4365]_  = ~\new_[4540]_  | ~\new_[5292]_ ;
  assign \new_[4366]_  = ~\new_[5203]_  | ~\new_[5772]_ ;
  assign \new_[4367]_  = ~\new_[4972]_  | ~\new_[4561]_ ;
  assign \new_[4368]_  = ~\new_[6272]_  | ~\new_[5283]_  | ~\new_[5595]_ ;
  assign \new_[4369]_  = (~\new_[5558]_  | ~\new_[5116]_ ) & (~\new_[5992]_  | ~\new_[5894]_ );
  assign \new_[4370]_  = ~\new_[4857]_  | ~\new_[6156]_ ;
  assign \new_[4371]_  = ~\new_[7209]_ ;
  assign \new_[4372]_  = ~\new_[6358]_  | ~\new_[6415]_  | ~\new_[5004]_  | ~\new_[4640]_ ;
  assign \new_[4373]_  = ~\new_[5356]_  & ~\new_[2660]_ ;
  assign \new_[4374]_  = \new_[4550]_  & \new_[4551]_ ;
  assign \new_[4375]_  = (~\new_[6300]_  | ~\new_[6037]_ ) & (~\new_[4641]_  | ~\new_[6952]_ );
  assign \new_[4376]_  = (~\new_[4641]_  | ~\new_[6953]_ ) & (~\new_[6306]_  | ~\new_[5959]_ );
  assign \new_[4377]_  = ~\new_[4552]_  | (~\new_[4770]_  & ~\new_[5818]_ );
  assign \new_[4378]_  = ~\new_[4648]_  | (~\new_[4646]_  & ~\new_[6519]_ );
  assign \new_[4379]_  = ~\new_[5476]_  | ~\new_[4565]_  | ~\new_[5528]_ ;
  assign \new_[4380]_  = (~\new_[4638]_  | ~\new_[5823]_ ) & (~\new_[5123]_  | ~\new_[4873]_ );
  assign \new_[4381]_  = \new_[4665]_  | \new_[4902]_  | \new_[4470]_  | \new_[4831]_ ;
  assign \new_[4382]_  = ~\new_[4664]_  | ~\new_[5721]_  | ~\new_[4474]_  | ~\new_[4818]_ ;
  assign \new_[4383]_  = ~\new_[4980]_  | ~\new_[4468]_ ;
  assign \new_[4384]_  = ~\new_[4654]_  & ~\new_[4602]_ ;
  assign \new_[4385]_  = ~\new_[4931]_  | (~\new_[4669]_  & ~\new_[6133]_ );
  assign \new_[4386]_  = (~\new_[4897]_  | ~\new_[6128]_ ) & (~\new_[5055]_  | ~\new_[6128]_ );
  assign \new_[4387]_  = \new_[4663]_  ^ \new_[4906]_ ;
  assign \new_[4388]_  = ~\new_[4469]_ ;
  assign \new_[4389]_  = ~\new_[4978]_  | ~\new_[4594]_  | ~\new_[4975]_ ;
  assign \new_[4390]_  = ~\new_[7174]_  | ~\new_[1379]_ ;
  assign \new_[4391]_  = ~\new_[7174]_  | ~\new_[1394]_ ;
  assign \new_[4392]_  = ~\new_[4593]_  & (~\new_[5646]_  | ~\new_[7208]_ );
  assign \new_[4393]_  = ~\new_[4597]_  & ~\new_[6411]_ ;
  assign \new_[4394]_  = \new_[1413]_  & \new_[4589]_ ;
  assign \new_[4395]_  = ~\new_[7174]_  | ~\new_[1892]_ ;
  assign \new_[4396]_  = ~\new_[4830]_  | ~\new_[4973]_  | ~\new_[4609]_  | ~\new_[4695]_ ;
  assign \new_[4397]_  = ~\new_[7174]_  & (~\new_[4724]_  | ~\new_[7171]_ );
  assign \new_[4398]_  = ~\new_[4595]_  & (~\new_[5895]_  | ~\new_[5044]_ );
  assign \new_[4399]_  = ~\new_[7174]_  & (~\new_[4731]_  | ~\new_[7171]_ );
  assign \new_[4400]_  = ~\new_[7174]_  & (~\new_[4732]_  | ~\new_[7171]_ );
  assign \new_[4401]_  = ~\new_[7174]_  & (~\new_[4733]_  | ~\new_[7171]_ );
  assign \new_[4402]_  = ~\new_[5085]_  & (~\new_[4810]_  | ~\new_[5772]_ );
  assign \new_[4403]_  = ~\new_[4936]_  | ~\new_[5193]_  | ~\new_[4601]_  | ~\new_[6016]_ ;
  assign \new_[4404]_  = (~\new_[4682]_  | ~\new_[740]_ ) & (~\new_[6953]_  | ~\new_[6589]_ );
  assign \new_[4405]_  = ~\new_[5336]_  & (~\new_[4682]_  | ~\new_[6606]_ );
  assign \new_[4406]_  = ~\new_[5333]_  & (~\new_[4682]_  | ~\new_[6591]_ );
  assign \new_[4407]_  = ~\new_[5373]_  | ~\new_[5090]_  | ~\new_[4686]_ ;
  assign \new_[4408]_  = ~\new_[4909]_  & ~\new_[4599]_ ;
  assign \new_[4409]_  = \new_[4808]_  & \new_[4675]_ ;
  assign \new_[4410]_  = ~\new_[5883]_  | ~\new_[4683]_  | ~\new_[4712]_ ;
  assign \new_[4411]_  = ~\new_[4690]_  | (~\new_[5686]_  & ~\new_[4670]_ );
  assign \new_[4412]_  = (~\new_[4711]_  | ~\new_[6128]_ ) & (~\new_[5515]_  | ~\new_[6128]_ );
  assign \new_[4413]_  = ~\new_[4506]_ ;
  assign \new_[4414]_  = \new_[4743]_  ? \new_[6271]_  : \new_[1892]_ ;
  assign \new_[4415]_  = \new_[5168]_  | \new_[4598]_ ;
  assign \new_[4416]_  = ~\new_[4615]_  & ~\new_[5093]_ ;
  assign \new_[4417]_  = ~\new_[5294]_  & (~\new_[4747]_  | ~\new_[6084]_ );
  assign \new_[4418]_  = ~\new_[6047]_  | ~\new_[5969]_  | ~\new_[5112]_  | ~\new_[6104]_ ;
  assign \new_[4419]_  = ~\new_[4631]_  & (~\new_[5092]_  | ~\new_[6278]_ );
  assign \new_[4420]_  = (~\new_[5697]_  | ~\new_[5772]_ ) & (~\new_[5566]_  | ~\new_[4744]_ );
  assign \new_[4421]_  = ~\new_[5896]_  & ~\new_[4625]_ ;
  assign \new_[4422]_  = ~\new_[5514]_  | ~\new_[5116]_ ;
  assign \new_[4423]_  = ~\new_[6596]_  | ~\new_[5295]_ ;
  assign \new_[4424]_  = ~\new_[6678]_  | ~\new_[5295]_ ;
  assign \new_[4426]_  = ~\new_[6658]_  | ~\new_[5295]_ ;
  assign \new_[4427]_  = ~\new_[4629]_  | ~\new_[4994]_ ;
  assign \new_[4428]_  = ~\new_[5103]_  | ~\new_[4627]_ ;
  assign \new_[4429]_  = ~\new_[4533]_ ;
  assign \new_[4430]_  = ~\new_[1111]_  | ~\new_[4634]_ ;
  assign \new_[4431]_  = \new_[5360]_  | \new_[4634]_ ;
  assign \new_[4432]_  = ~\new_[5595]_  | (~\new_[5954]_  & ~\new_[6064]_ );
  assign \new_[4433]_  = ~\new_[5116]_  | (~\new_[7070]_  & ~\new_[6060]_ );
  assign \new_[4434]_  = (~\new_[4740]_  | ~\new_[6465]_ ) & (~\new_[7125]_  | ~\new_[6434]_ );
  assign \new_[4435]_  = ~\new_[6032]_  | ~\new_[5116]_ ;
  assign \new_[4436]_  = \new_[4639]_  | \new_[6472]_ ;
  assign \new_[4437]_  = \new_[5613]_  ? \new_[4770]_  : \new_[5011]_ ;
  assign \new_[4438]_  = \new_[5137]_  ? \new_[4655]_  : \new_[5019]_ ;
  assign \new_[4439]_  = ~\new_[4876]_  | ~\new_[5750]_  | ~\new_[4773]_  | ~\new_[5899]_ ;
  assign \new_[4440]_  = ~\new_[5332]_  & (~\new_[4769]_  | ~\new_[6589]_ );
  assign \new_[4441]_  = \new_[4644]_  | \new_[5877]_ ;
  assign \new_[4442]_  = ~\new_[5116]_  | ~\new_[6137]_ ;
  assign \new_[4443]_  = \new_[4632]_  & \new_[5245]_ ;
  assign \new_[4444]_  = (~\new_[4704]_  | ~\new_[2429]_ ) & (~\new_[5139]_  | ~\new_[5304]_ );
  assign \new_[4445]_  = ~\new_[5375]_  | ~\new_[6937]_  | ~\new_[6936]_ ;
  assign \new_[4446]_  = ~\new_[4814]_  | ~\new_[5814]_  | ~\new_[5037]_  | ~\new_[5851]_ ;
  assign \new_[4447]_  = ~\new_[4821]_  | ~\new_[7120]_  | ~\new_[4692]_  | ~\new_[4782]_ ;
  assign \new_[4448]_  = ~\new_[5648]_  | ~\new_[5140]_  | ~\new_[4786]_  | ~\new_[7564]_ ;
  assign \new_[4449]_  = ~\new_[5554]_  | ~\new_[4569]_  | ~\new_[5664]_ ;
  assign \new_[4450]_  = ~\new_[4570]_  & ~\new_[5196]_ ;
  assign \new_[4451]_  = ~\new_[6000]_  | ~\new_[5000]_  | ~\new_[4766]_  | ~\new_[4764]_ ;
  assign \new_[4452]_  = ~\new_[5715]_  | ~\new_[5843]_  | ~\new_[4790]_  | ~\new_[6003]_ ;
  assign \new_[4453]_  = ~\new_[5791]_  | ~\new_[5790]_  | ~\new_[4787]_ ;
  assign \new_[4454]_  = \new_[4728]_  | \new_[7436]_ ;
  assign \new_[4455]_  = ~\new_[5553]_  | ~\new_[5545]_  | ~\new_[7149]_  | ~\new_[4793]_ ;
  assign \new_[4456]_  = \new_[4719]_  | \new_[7436]_ ;
  assign \new_[4457]_  = \new_[4717]_  | \new_[7436]_ ;
  assign \new_[4458]_  = \new_[4723]_  | \new_[7436]_ ;
  assign \new_[4459]_  = \new_[4729]_  | \new_[7436]_ ;
  assign \new_[4460]_  = \new_[4730]_  | \new_[7436]_ ;
  assign \new_[4461]_  = \new_[4716]_  | \new_[7436]_ ;
  assign \new_[4462]_  = \new_[4720]_  | \new_[7436]_ ;
  assign \new_[4463]_  = \new_[4715]_  | \new_[7436]_ ;
  assign \new_[4464]_  = \new_[4727]_  | \new_[7436]_ ;
  assign \new_[4465]_  = \new_[4734]_  | \new_[7436]_ ;
  assign \new_[4466]_  = \new_[4735]_  | \new_[7436]_ ;
  assign \new_[4467]_  = ~\new_[5639]_  | ~\new_[5548]_  | ~\new_[4652]_  | ~\new_[5698]_ ;
  assign \new_[4468]_  = ~\new_[5050]_  & (~\new_[4803]_  | ~\new_[6064]_ );
  assign \new_[4469]_  = \new_[1413]_  | \new_[4666]_ ;
  assign \new_[4470]_  = \new_[5039]_  | \new_[4663]_ ;
  assign \new_[4471]_  = ~\new_[7174]_  | ~\new_[1308]_ ;
  assign \new_[4472]_  = ~\new_[7174]_  | ~\new_[1453]_ ;
  assign \new_[4473]_  = ~\new_[7174]_  | ~\new_[1104]_ ;
  assign \new_[4474]_  = ~\new_[4661]_  & ~\new_[5759]_ ;
  assign \new_[4475]_  = ~\new_[7174]_  | ~\new_[1861]_ ;
  assign \new_[4476]_  = \new_[4671]_  & \new_[5694]_ ;
  assign \new_[4477]_  = ~\new_[7174]_  | ~\new_[1646]_ ;
  assign \new_[4478]_  = ~\new_[7174]_  | ~\new_[1610]_ ;
  assign \new_[4479]_  = ~\new_[7174]_  | ~\new_[1545]_ ;
  assign \new_[4480]_  = ~\new_[5788]_  | ~\new_[5700]_  | ~\new_[4667]_  | ~\new_[5104]_ ;
  assign \new_[4481]_  = ~\new_[5056]_  | ~\new_[5302]_  | ~\new_[4677]_  | ~\new_[4843]_ ;
  assign \new_[4482]_  = \new_[4662]_  | \new_[5267]_ ;
  assign \new_[4483]_  = ~\new_[4739]_  & (~\new_[6919]_  | ~\new_[6002]_ );
  assign \new_[4484]_  = ~\new_[4908]_  | ~\new_[5898]_  | ~\new_[5700]_  | ~\new_[5335]_ ;
  assign \new_[4485]_  = \new_[2780]_  ? \new_[4813]_  : \new_[3029]_ ;
  assign \new_[4486]_  = \new_[844]_  ? \new_[6031]_  : \new_[4831]_ ;
  assign \new_[4487]_  = ~\new_[4753]_  | (~\new_[4988]_  & ~\new_[5692]_ );
  assign \new_[4488]_  = \new_[5039]_  ^ \new_[4831]_ ;
  assign \new_[4489]_  = ~\new_[4682]_  | ~\new_[6521]_ ;
  assign \new_[4490]_  = ~\new_[4682]_  | ~\new_[850]_ ;
  assign \new_[4491]_  = ~\new_[4682]_  | ~\new_[6472]_ ;
  assign \new_[4492]_  = \new_[4927]_  | \new_[4682]_ ;
  assign \new_[4493]_  = \new_[4909]_  & \new_[4678]_ ;
  assign \new_[4494]_  = ~\new_[4909]_  & ~\new_[4674]_ ;
  assign \new_[4495]_  = \new_[4909]_  & \new_[4676]_ ;
  assign \new_[4496]_  = \new_[4677]_  & \new_[6016]_ ;
  assign \new_[4497]_  = \new_[4909]_  & \new_[4675]_ ;
  assign \new_[4498]_  = ~\new_[4808]_  & ~\new_[4674]_ ;
  assign \new_[4499]_  = \new_[4808]_  & \new_[4678]_ ;
  assign \new_[4500]_  = ~\new_[4589]_ ;
  assign \new_[4501]_  = ~\new_[5311]_  | ~\new_[5700]_  | ~\new_[4742]_  | ~\new_[5749]_ ;
  assign \new_[4502]_  = ~\new_[4681]_  & (~\new_[5307]_  | ~\new_[6050]_ );
  assign \new_[4503]_  = ~\new_[4752]_  & (~\new_[5782]_  | ~\new_[5116]_ );
  assign \new_[4504]_  = (~\new_[4832]_  & ~\new_[5988]_ ) | (~\new_[4977]_  & ~\new_[5666]_ );
  assign \new_[4505]_  = ~\new_[4933]_  | ~\new_[5077]_  | ~\new_[5101]_  | ~\new_[5195]_ ;
  assign \new_[4506]_  = (~\new_[4828]_  | ~\new_[1623]_ ) & (~\new_[5611]_  | ~\new_[6351]_ );
  assign \new_[4507]_  = ~\new_[6357]_  | ~\new_[6452]_  | ~\new_[4722]_  | ~\new_[407]_ ;
  assign \new_[4508]_  = \new_[4838]_  ? \new_[6271]_  : \new_[1689]_ ;
  assign \new_[4509]_  = \new_[4837]_  ? \new_[6271]_  : \new_[1861]_ ;
  assign \new_[4510]_  = (~\new_[4870]_  | ~\new_[6084]_ ) & (~\new_[5607]_  | ~\new_[6084]_ );
  assign \new_[4511]_  = ~\new_[4722]_  | ~\new_[1623]_ ;
  assign \new_[4512]_  = ~\new_[5308]_  | (~\new_[5524]_  & ~\new_[5356]_ );
  assign \new_[4513]_  = ~\new_[4721]_  & ~\new_[4956]_ ;
  assign \new_[4514]_  = \new_[4714]_  & \new_[7023]_ ;
  assign \new_[4515]_  = ~\new_[4600]_ ;
  assign \new_[4516]_  = ~\new_[4979]_  | ~\new_[7059]_  | ~\new_[4853]_ ;
  assign \new_[4517]_  = \new_[4714]_  & \new_[7045]_ ;
  assign \new_[4518]_  = ~\new_[4959]_  | ~\new_[4963]_  | ~\new_[5086]_  | ~\new_[4848]_ ;
  assign \new_[4519]_  = ~\new_[4963]_  | ~\new_[5079]_  | ~\new_[4848]_  | ~\new_[4959]_ ;
  assign \new_[4520]_  = ~\new_[6161]_  | ~\new_[6310]_  | ~\new_[4713]_  | ~\new_[6340]_ ;
  assign \new_[4521]_  = ~\new_[4736]_  & (~\new_[5584]_  | ~\new_[6167]_ );
  assign \new_[4522]_  = (~\new_[5617]_  | ~\new_[5928]_ ) & (~\new_[5713]_  | ~\new_[4857]_ );
  assign \new_[4523]_  = (~\new_[5805]_  | ~\new_[5083]_ ) & (~\new_[5399]_  | ~\new_[6050]_ );
  assign \new_[4524]_  = (~\new_[5864]_  | ~\new_[5928]_ ) & (~\new_[7209]_  | ~\new_[5845]_ );
  assign \new_[4525]_  = ~\new_[4656]_  & (~\new_[5092]_  | ~\new_[1324]_ );
  assign \new_[4526]_  = ~\new_[4707]_  & (~\new_[5147]_  | ~\new_[5862]_ );
  assign \new_[4527]_  = ~\new_[5417]_  | ~\new_[6128]_ ;
  assign \new_[4528]_  = ~\new_[5644]_  | ~\new_[6128]_ ;
  assign \new_[4529]_  = ~\new_[1865]_  & ~\new_[5184]_ ;
  assign \new_[4530]_  = ~\new_[1693]_  & ~\new_[5184]_ ;
  assign \new_[4531]_  = ~\new_[5300]_  | ~\new_[5772]_ ;
  assign \new_[4532]_  = ~\new_[4745]_  & (~\new_[4995]_  | ~\new_[6113]_ );
  assign \new_[4533]_  = ~\new_[7208]_  & (~\new_[5792]_  | ~\new_[5768]_ );
  assign \new_[4534]_  = ~\new_[4965]_  | (~\new_[5018]_  & ~\new_[850]_ );
  assign \new_[4535]_  = ~\new_[5577]_  | ~\new_[5772]_ ;
  assign \new_[4536]_  = ~\new_[5103]_  & ~\new_[4759]_ ;
  assign \new_[4537]_  = ~\new_[5242]_  & (~\new_[4869]_  | ~\new_[7550]_ );
  assign \new_[4538]_  = \new_[5103]_  & \new_[4759]_ ;
  assign \new_[4539]_  = ~\new_[4650]_  | ~\new_[4855]_ ;
  assign \new_[4540]_  = \new_[4758]_  & \new_[5903]_ ;
  assign \new_[4541]_  = ~\new_[6472]_  & ~\new_[6400]_ ;
  assign \new_[4542]_  = ~\new_[6011]_  & ~\new_[4766]_ ;
  assign \new_[4543]_  = ~\new_[4765]_  & ~\new_[5458]_ ;
  assign \new_[4544]_  = ~\new_[6011]_  & ~\new_[4764]_ ;
  assign \new_[4545]_  = \new_[4763]_  | \new_[5458]_ ;
  assign \new_[4546]_  = ~\new_[5958]_  | ~\new_[5595]_ ;
  assign \new_[4547]_  = ~\new_[6031]_  & ~\new_[5688]_ ;
  assign \new_[4548]_  = (~\new_[5771]_  | ~\new_[6284]_ ) & (~\new_[5958]_  | ~\new_[5116]_ );
  assign \new_[4549]_  = \\di_reg_reg[6] ;
  assign \new_[4550]_  = \new_[5610]_  | \new_[4770]_ ;
  assign \new_[4551]_  = ~\new_[5610]_  | ~\new_[4770]_ ;
  assign \new_[4552]_  = ~\new_[4770]_  | ~\new_[4772]_ ;
  assign \new_[4553]_  = \\di_reg_reg[3] ;
  assign \new_[4554]_  = \\di_reg_reg[1] ;
  assign \new_[4555]_  = \new_[4769]_  | \new_[5133]_ ;
  assign \new_[4556]_  = \\di_reg_reg[7] ;
  assign \new_[4557]_  = \\di_reg_reg[2] ;
  assign \new_[4558]_  = \\di_reg_reg[4] ;
  assign \new_[4559]_  = \\di_reg_reg[5] ;
  assign \new_[4560]_  = \\di_reg_reg[0] ;
  assign \new_[4561]_  = ~\new_[5116]_  | ~\new_[5910]_  | ~\new_[6325]_ ;
  assign \new_[4562]_  = (~\new_[4783]_  | ~\new_[5894]_ ) & (~\new_[5307]_  | ~\new_[5937]_ );
  assign \new_[4563]_  = ~\new_[4651]_  & ~\new_[5854]_ ;
  assign \new_[4564]_  = ~\new_[4645]_ ;
  assign \new_[4565]_  = ~\new_[4647]_  & ~\new_[5262]_ ;
  assign \new_[4566]_  = ~\new_[5249]_  & (~\new_[4906]_  | ~\new_[6040]_ );
  assign \new_[4567]_  = \new_[4788]_  & \new_[5658]_ ;
  assign \new_[4568]_  = \new_[6084]_  ? \new_[5680]_  : \di[4] ;
  assign \new_[4569]_  = ~\new_[4785]_  & ~\new_[5596]_ ;
  assign \new_[4570]_  = ~\new_[5413]_  | ~\new_[5299]_  | ~\new_[5306]_  | ~\new_[4894]_ ;
  assign \new_[4571]_  = ~\new_[4802]_  & ~\new_[5159]_ ;
  assign \new_[4572]_  = ~\new_[7174]_  | ~\new_[6580]_ ;
  assign \new_[4573]_  = ~\new_[4998]_  & (~\new_[4900]_  | ~\new_[6040]_ );
  assign \new_[4574]_  = ~\new_[4794]_  & (~\new_[5088]_  | ~\new_[2003]_ );
  assign \new_[4575]_  = ~\new_[4801]_  & (~\new_[5088]_  | ~\new_[2002]_ );
  assign \new_[4576]_  = ~\new_[4800]_  & (~\new_[5088]_  | ~\new_[2016]_ );
  assign \new_[4577]_  = ~\new_[4795]_  & (~\new_[5088]_  | ~\new_[6478]_ );
  assign \new_[4578]_  = ~\new_[4784]_  & (~\new_[5088]_  | ~\new_[6515]_ );
  assign \new_[4579]_  = ~\new_[4796]_  & (~\new_[5088]_  | ~\new_[6518]_ );
  assign \new_[4580]_  = ~\new_[4797]_  & (~\new_[5088]_  | ~\new_[6542]_ );
  assign \new_[4581]_  = ~\new_[4799]_  & (~\new_[5088]_  | ~\new_[2006]_ );
  assign \new_[4582]_  = ~\new_[5246]_  | ~\new_[4820]_  | ~\new_[4905]_ ;
  assign \new_[4583]_  = (~\new_[4904]_  | ~\new_[6040]_ ) & (~\new_[5092]_  | ~\new_[1126]_ );
  assign \new_[4584]_  = (~\new_[4912]_  | ~\new_[6084]_ ) & (~\new_[5203]_  | ~\new_[6084]_ );
  assign \new_[4585]_  = (~\new_[4903]_  | ~\new_[5455]_ ) & (~\new_[7208]_  | ~\new_[5635]_ );
  assign \new_[4586]_  = \new_[4902]_  ^ \new_[4901]_ ;
  assign \new_[4587]_  = \new_[4904]_  ^ \new_[4900]_ ;
  assign \new_[4588]_  = ~\new_[4813]_  | ~\new_[6348]_ ;
  assign \new_[4589]_  = ~\new_[4666]_ ;
  assign \new_[4590]_  = ~\new_[4812]_  | ~\new_[4968]_ ;
  assign \new_[4591]_  = ~\new_[5042]_  & (~\new_[5805]_  | ~\new_[4982]_ );
  assign \new_[4592]_  = ~\new_[4817]_  & (~\new_[5455]_  | ~\new_[6032]_ );
  assign \new_[4593]_  = ~\new_[4815]_  | (~\new_[5893]_  & ~\new_[5598]_ );
  assign \new_[4594]_  = ~\new_[4840]_  & (~\new_[5172]_  | ~\new_[6084]_ );
  assign \new_[4595]_  = ~\new_[5195]_  | ~\new_[5077]_  | ~\new_[5869]_  | ~\new_[5101]_ ;
  assign \new_[4596]_  = (~\new_[4919]_  | ~\new_[6084]_ ) & (~\new_[5645]_  | ~\new_[6084]_ );
  assign \new_[4597]_  = ~\new_[4806]_  & (~\new_[5656]_  | ~\new_[5456]_ );
  assign \new_[4598]_  = \new_[5697]_  & \new_[4867]_ ;
  assign \new_[4599]_  = ~\new_[4676]_ ;
  assign \new_[4600]_  = ~\new_[4937]_  | ~\new_[4849]_ ;
  assign \new_[4601]_  = \new_[4834]_  & \new_[5637]_ ;
  assign \new_[4602]_  = ~\new_[4836]_  | ~\new_[5788]_ ;
  assign \new_[4603]_  = ~\new_[4979]_  | ~\new_[5213]_  | ~\new_[7175]_ ;
  assign \new_[4604]_  = ~\new_[5242]_  & (~\new_[4884]_  | ~\new_[6227]_ );
  assign \new_[4605]_  = ~\new_[4990]_  | ~\new_[5286]_  | ~\new_[7163]_ ;
  assign \new_[4606]_  = ~\new_[4990]_  | ~\new_[5286]_  | ~\new_[5848]_ ;
  assign \new_[4607]_  = (~\new_[5455]_  | ~\new_[6002]_ ) & (~\new_[5760]_  | ~\new_[7121]_ );
  assign \new_[4608]_  = ~\new_[5699]_  | ~\new_[5108]_  | ~\new_[5345]_  | ~\new_[5870]_ ;
  assign \new_[4609]_  = (~\new_[4371]_  | ~\new_[6995]_ ) & (~\new_[5399]_  | ~\new_[5601]_ );
  assign \new_[4610]_  = (~\new_[5455]_  | ~\new_[5752]_ ) & (~\new_[5399]_  | ~\new_[5570]_ );
  assign \new_[4611]_  = (~\new_[5751]_  | ~\new_[5455]_ ) & (~\new_[5760]_  | ~\new_[5862]_ );
  assign \new_[4612]_  = \new_[6520]_  ^ \new_[4965]_ ;
  assign \new_[4613]_  = ~\new_[6551]_  | ~\new_[5295]_ ;
  assign \new_[4614]_  = ~\new_[6558]_  | ~\new_[5295]_ ;
  assign \new_[4615]_  = ~\new_[5013]_  | ~\new_[4854]_ ;
  assign \new_[4616]_  = ~\new_[4725]_ ;
  assign \new_[4617]_  = ~\new_[4726]_ ;
  assign \new_[4618]_  = \new_[753]_  ^ \new_[5221]_ ;
  assign \new_[4619]_  = ~\new_[4842]_  & (~\new_[5860]_  | ~\new_[6128]_ );
  assign \new_[4620]_  = \new_[761]_  ^ \new_[5221]_ ;
  assign \new_[4621]_  = \new_[763]_  ^ \new_[5221]_ ;
  assign \new_[4622]_  = \new_[760]_  ^ \new_[5221]_ ;
  assign \new_[4623]_  = \new_[736]_  ^ \new_[5221]_ ;
  assign \new_[4624]_  = \new_[762]_  ^ \new_[5221]_ ;
  assign \new_[4625]_  = ~\new_[4744]_ ;
  assign \new_[4626]_  = ~\new_[5103]_  & ~\new_[4859]_ ;
  assign \new_[4627]_  = ~\new_[5103]_  | ~\new_[4859]_ ;
  assign \new_[4628]_  = ~\new_[5119]_  | ~\new_[5115]_  | ~\new_[5684]_  | ~\new_[5107]_ ;
  assign \new_[4629]_  = ~\new_[5571]_  | ~\new_[5118]_  | ~\new_[5969]_  | ~\new_[6113]_ ;
  assign \new_[4630]_  = \new_[6113]_  ? \new_[5680]_  : \di[0] ;
  assign \new_[4631]_  = ~\new_[6011]_  & ~\new_[4868]_ ;
  assign \new_[4632]_  = \new_[4863]_  | \new_[5458]_ ;
  assign \new_[4633]_  = ~\new_[5779]_  | ~\new_[4878]_  | ~\new_[2006]_ ;
  assign \new_[4634]_  = \new_[5994]_  & \new_[4867]_ ;
  assign \new_[4635]_  = ~\new_[6011]_  & ~\new_[4871]_ ;
  assign \new_[4636]_  = ~\new_[4868]_  | ~\new_[4871]_ ;
  assign \new_[4637]_  = ~\new_[5779]_  | ~\new_[4872]_  | ~\new_[2003]_ ;
  assign \new_[4638]_  = \new_[6917]_  & \new_[6193]_ ;
  assign \new_[4639]_  = ~\new_[6521]_  | ~\new_[6084]_ ;
  assign \new_[4640]_  = (~\new_[6084]_  | ~\new_[7549]_ ) & (~\new_[6143]_  | ~\new_[6120]_ );
  assign \new_[4641]_  = \new_[5244]_  ^ \new_[5016]_ ;
  assign \new_[4642]_  = ~\new_[5009]_  & (~\new_[4902]_  | ~\new_[6040]_ );
  assign \new_[4643]_  = ~\new_[4877]_  & (~\new_[4901]_  | ~\new_[6040]_ );
  assign \new_[4644]_  = (~\new_[5024]_  | ~\new_[6625]_ ) & (~\new_[4881]_  | ~\new_[740]_ );
  assign \new_[4645]_  = ~\new_[6193]_  | ~\new_[6314]_ ;
  assign \new_[4646]_  = ~\new_[5248]_  & (~\new_[4882]_  | ~\new_[6523]_ );
  assign \new_[4647]_  = ~\new_[5942]_  | ~\new_[5981]_  | ~\new_[4898]_  | ~\new_[5725]_ ;
  assign \new_[4648]_  = ~\new_[4882]_  | ~\new_[6519]_ ;
  assign \new_[4649]_  = ~\new_[4888]_  | (~\new_[5152]_  & ~\new_[5474]_ );
  assign \new_[4650]_  = ~\new_[5809]_  | ~\new_[5595]_ ;
  assign \new_[4651]_  = ~\new_[5736]_  | ~\new_[5764]_  | ~\new_[5145]_  | ~\new_[5843]_ ;
  assign \new_[4652]_  = ~\new_[5169]_  & ~\new_[4896]_ ;
  assign \new_[4653]_  = ~\new_[4897]_  | ~\new_[6084]_ ;
  assign \new_[4654]_  = ~\new_[5700]_  | ~\new_[5153]_  | ~\new_[5040]_ ;
  assign \new_[4655]_  = ~\new_[5016]_  | ~\new_[5244]_ ;
  assign \new_[4656]_  = ~\new_[6011]_  & ~\new_[5000]_ ;
  assign \new_[4657]_  = ~\new_[6113]_  & ~\new_[5995]_ ;
  assign \new_[4658]_  = ~\new_[4883]_  | (~\new_[5152]_  & ~\new_[6170]_ );
  assign \new_[4659]_  = ~\new_[4891]_  | (~\new_[5152]_  & ~\new_[6086]_ );
  assign \new_[4660]_  = ~\new_[4885]_  | (~\new_[5152]_  & ~\new_[2429]_ );
  assign \new_[4661]_  = ~\new_[4916]_  | (~\new_[5418]_  & ~\new_[5428]_ );
  assign \new_[4662]_  = ~\new_[6731]_  & (~\new_[5156]_  | ~\new_[5049]_ );
  assign \new_[4663]_  = ~\new_[5204]_  | ~\new_[6138]_  | ~\new_[5761]_  | ~\new_[5337]_ ;
  assign \new_[4664]_  = ~\new_[4917]_  & (~\new_[5576]_  | ~\new_[7017]_ );
  assign \new_[4665]_  = \new_[4904]_  | \new_[5969]_ ;
  assign \new_[4666]_  = ~\new_[4914]_  & ~\new_[6935]_ ;
  assign \new_[4667]_  = ~\new_[5043]_  & ~\new_[4956]_ ;
  assign \new_[4668]_  = ~\new_[4901]_  & ~\new_[4900]_ ;
  assign \new_[4669]_  = ~\new_[4371]_  & (~\new_[5393]_  | ~\new_[5595]_ );
  assign \new_[4670]_  = ~\new_[5455]_  | ~\new_[6137]_ ;
  assign \new_[4671]_  = ~\new_[7561]_  | (~\new_[5044]_  & ~\new_[5595]_ );
  assign \new_[4672]_  = ~\new_[5669]_  | ~\new_[5170]_  | ~\new_[5793]_  | ~\new_[5660]_ ;
  assign \new_[4673]_  = \new_[5926]_  & \new_[4973]_ ;
  assign \new_[4674]_  = ~\new_[4924]_  | ~\new_[5001]_ ;
  assign \new_[4675]_  = ~\new_[4924]_  & ~\new_[5001]_ ;
  assign \new_[4676]_  = ~\new_[5045]_  & ~\new_[5001]_ ;
  assign \new_[4677]_  = \new_[5389]_  & \new_[4937]_ ;
  assign \new_[4678]_  = \new_[5045]_  & \new_[5001]_ ;
  assign \new_[4679]_  = ~\new_[5431]_  | ~\new_[6084]_ ;
  assign \new_[4680]_  = \new_[4929]_  | \new_[4957]_ ;
  assign \new_[4681]_  = ~\new_[5769]_  & (~\new_[5083]_  | ~\new_[6233]_ );
  assign \new_[4682]_  = ~\new_[4927]_  & ~\new_[5550]_ ;
  assign \new_[4683]_  = ~\new_[5875]_  & (~\new_[5668]_  | ~\new_[5331]_ );
  assign \new_[4684]_  = ~\new_[5298]_  | ~\new_[5782]_  | ~\new_[7209]_ ;
  assign \new_[4685]_  = ~\new_[4986]_  & (~\new_[5534]_  | ~\new_[5928]_ );
  assign \new_[4686]_  = ~\new_[5003]_  | ~\new_[6084]_ ;
  assign \new_[4687]_  = ~\new_[5377]_  & (~\new_[5092]_  | ~\new_[6110]_ );
  assign \new_[4688]_  = \new_[4934]_  & \new_[5079]_ ;
  assign \new_[4689]_  = ~\new_[4371]_  | (~\new_[5401]_  & ~\new_[5631]_ );
  assign \new_[4690]_  = (~\new_[5094]_  | ~\new_[5239]_ ) & (~\new_[5385]_  | ~\new_[6325]_ );
  assign \new_[4691]_  = ~\new_[4923]_  & (~\new_[6478]_  | ~\new_[5459]_ );
  assign \new_[4692]_  = ~\new_[4925]_  & (~\new_[5598]_  | ~\new_[5631]_ );
  assign \new_[4693]_  = ~\new_[5852]_  & (~\new_[5092]_  | ~\new_[1248]_ );
  assign \new_[4694]_  = (~\new_[5082]_  | ~\new_[6359]_ ) & (~\new_[7315]_  | ~\new_[6405]_ );
  assign \new_[4695]_  = (~\new_[5608]_  | ~\new_[5331]_ ) & (~\new_[5760]_  | ~\new_[5924]_ );
  assign n1839 = ~\new_[6424]_  & (~\new_[5099]_  | ~\new_[5589]_ );
  assign n1834 = ~\new_[6424]_  & (~\new_[5128]_  | ~\new_[5423]_ );
  assign n1859 = ~\new_[6424]_  & (~\new_[5110]_  | ~\new_[5422]_ );
  assign n1854 = ~\new_[6424]_  & (~\new_[5131]_  | ~\new_[5424]_ );
  assign n1829 = ~\new_[6424]_  & (~\new_[5100]_  | ~\new_[5539]_ );
  assign n1844 = ~\new_[6424]_  & (~\new_[5121]_  | ~\new_[5540]_ );
  assign n1849 = ~\new_[6424]_  & (~\new_[5105]_  | ~\new_[5537]_ );
  assign n1864 = ~\new_[6424]_  & (~\new_[5102]_  | ~\new_[5585]_ );
  assign \new_[4704]_  = ~\new_[4957]_  & ~\new_[5304]_ ;
  assign \new_[4705]_  = ~\new_[4983]_  & ~\new_[6113]_ ;
  assign \new_[4706]_  = ~\new_[5087]_  | ~\new_[6128]_ ;
  assign \new_[4707]_  = ~\new_[5880]_  | ~\new_[5462]_  | ~\new_[5098]_ ;
  assign \new_[4708]_  = ~\new_[4821]_ ;
  assign \new_[4709]_  = ~\new_[5084]_  & ~\new_[4976]_ ;
  assign \new_[4710]_  = ~\new_[4970]_  & ~\new_[4951]_ ;
  assign \new_[4711]_  = ~\new_[4971]_  | ~\new_[5874]_ ;
  assign \new_[4712]_  = ~\new_[5547]_  | ~\new_[7208]_ ;
  assign \new_[4713]_  = ~\new_[5220]_  & ~\new_[5935]_ ;
  assign \new_[4714]_  = ~\new_[5638]_  & (~\new_[5751]_  | ~\new_[7209]_ );
  assign \new_[4715]_  = ~\new_[4940]_  & (~\new_[5223]_  | ~\new_[1239]_ );
  assign \new_[4716]_  = ~\new_[4948]_  & (~\new_[5223]_  | ~\new_[1255]_ );
  assign \new_[4717]_  = ~\new_[4941]_  & (~\new_[5223]_  | ~\new_[1233]_ );
  assign \new_[4718]_  = \new_[4960]_  & \new_[5213]_ ;
  assign \new_[4719]_  = ~\new_[4950]_  & (~\new_[5223]_  | ~\new_[1293]_ );
  assign \new_[4720]_  = ~\new_[4945]_  & (~\new_[5223]_  | ~\new_[1238]_ );
  assign \new_[4721]_  = \new_[4993]_  | \new_[5186]_ ;
  assign \new_[4722]_  = ~\new_[4828]_ ;
  assign \new_[4723]_  = ~\new_[4944]_  & (~\new_[5223]_  | ~\new_[1234]_ );
  assign \new_[4724]_  = ~\new_[4952]_  & (~\new_[5223]_  | ~\new_[1237]_ );
  assign \new_[4725]_  = ~\new_[4967]_  & (~\new_[5221]_  | ~\new_[6606]_ );
  assign \new_[4726]_  = ~\new_[4981]_  & (~\new_[5221]_  | ~\new_[6591]_ );
  assign \new_[4727]_  = ~\new_[4955]_  & (~\new_[5223]_  | ~\new_[1225]_ );
  assign \new_[4728]_  = ~\new_[4943]_  & (~\new_[5223]_  | ~\new_[1294]_ );
  assign \new_[4729]_  = ~\new_[4954]_  & (~\new_[5223]_  | ~\new_[1235]_ );
  assign \new_[4730]_  = ~\new_[4946]_  & (~\new_[5223]_  | ~\new_[1292]_ );
  assign \new_[4731]_  = ~\new_[4949]_  & (~\new_[5223]_  | ~\new_[1236]_ );
  assign \new_[4732]_  = ~\new_[4953]_  & (~\new_[5223]_  | ~\new_[1240]_ );
  assign \new_[4733]_  = ~\new_[4984]_  & (~\new_[5223]_  | ~\new_[1241]_ );
  assign \new_[4734]_  = ~\new_[4947]_  & (~\new_[5223]_  | ~\new_[1242]_ );
  assign \new_[4735]_  = ~\new_[4942]_  & (~\new_[5223]_  | ~\new_[1223]_ );
  assign \new_[4736]_  = (~\new_[5106]_  & ~\new_[6461]_ ) | (~\new_[5776]_  & ~\new_[5772]_ );
  assign \new_[4737]_  = ~\new_[4833]_ ;
  assign \new_[4738]_  = ~\new_[5609]_  & (~\new_[5697]_  | ~\new_[6084]_ );
  assign \new_[4739]_  = ~\new_[5205]_  | (~\new_[6013]_  & ~\new_[5356]_ );
  assign \new_[4740]_  = \new_[5005]_  & \new_[5823]_ ;
  assign \new_[4741]_  = (~\new_[5697]_  | ~\new_[6128]_ ) & (~\new_[5566]_  | ~\new_[5091]_ );
  assign \new_[4742]_  = ~\new_[4958]_  & (~\new_[5751]_  | ~\new_[6009]_ );
  assign \new_[4743]_  = \new_[5772]_  ? \new_[7172]_  : \new_[1892]_ ;
  assign \new_[4744]_  = ~\new_[4985]_  | ~\new_[5443]_ ;
  assign \new_[4745]_  = (~\new_[5675]_  & ~\new_[7549]_ ) | (~\new_[5775]_  & ~\new_[5772]_ );
  assign \new_[4746]_  = ~\new_[4371]_  | ~\new_[5845]_ ;
  assign \new_[4747]_  = ~\new_[5640]_  | ~\new_[5955]_  | ~\new_[5874]_ ;
  assign \new_[4748]_  = ~\new_[4996]_  & ~\new_[5991]_ ;
  assign \new_[4749]_  = ~\new_[4992]_  & (~\new_[5579]_  | ~\new_[5350]_ );
  assign \new_[4750]_  = \new_[7549]_  ? \new_[5680]_  : \di[2] ;
  assign \new_[4751]_  = ~\new_[5759]_  | ~\new_[5772]_ ;
  assign \new_[4752]_  = ~\new_[5163]_  | (~\new_[5669]_  & ~\new_[5095]_ );
  assign \new_[4753]_  = ~\new_[5597]_  | ~\new_[5008]_ ;
  assign \new_[4754]_  = ~\new_[5458]_  & (~\new_[5119]_  | ~\new_[6654]_ );
  assign \new_[4755]_  = ~\new_[2016]_  | ~\new_[5779]_  | ~\new_[5115]_ ;
  assign \new_[4756]_  = ~\new_[5779]_  | ~\new_[5012]_  | ~\new_[2005]_ ;
  assign \new_[4757]_  = ~\new_[4976]_  & ~\new_[4970]_ ;
  assign \new_[4758]_  = \new_[5948]_  | \new_[6143]_ ;
  assign \new_[4759]_  = ~\new_[4859]_ ;
  assign \new_[4760]_  = ~\new_[5773]_  | ~\new_[5969]_  | ~\new_[5823]_  | ~\new_[7170]_ ;
  assign \new_[4761]_  = ~\new_[5348]_  | (~\new_[5578]_  & ~\new_[5356]_ );
  assign \new_[4762]_  = ~\new_[5002]_  & (~\new_[6812]_  | ~\new_[5972]_ );
  assign \new_[4763]_  = ~\new_[4991]_  & ~\new_[2006]_ ;
  assign \new_[4764]_  = ~\new_[4991]_  | ~\new_[2006]_ ;
  assign \new_[4765]_  = ~\new_[5007]_  & ~\new_[2003]_ ;
  assign \new_[4766]_  = ~\new_[5007]_  | ~\new_[2003]_ ;
  assign \new_[4767]_  = ~\new_[7315]_  | (~\new_[5117]_  & ~\new_[6124]_ );
  assign \new_[4768]_  = ~\new_[4889]_  | (~\new_[5152]_  & ~\new_[5785]_ );
  assign \new_[4769]_  = ~\new_[5130]_  | ~\new_[5129]_  | ~\new_[5747]_ ;
  assign \new_[4770]_  = ~\new_[6584]_  | ~\new_[5818]_  | ~\new_[5126]_ ;
  assign \new_[4771]_  = ~\new_[4890]_  | (~\new_[5152]_  & ~\new_[5594]_ );
  assign \new_[4772]_  = \new_[5818]_  ^ \new_[5126]_ ;
  assign \new_[4773]_  = (~\new_[5132]_  | ~\new_[6953]_ ) & (~\new_[6339]_  | ~\new_[5959]_ );
  assign \new_[4774]_  = ~\new_[4886]_  | (~\new_[5152]_  & ~\new_[5604]_ );
  assign \new_[4775]_  = ~\new_[4887]_  | (~\new_[5152]_  & ~\new_[5600]_ );
  assign \new_[4776]_  = ~\new_[4893]_  | (~\new_[5152]_  & ~\new_[6131]_ );
  assign \new_[4777]_  = (~\new_[5133]_  | ~\new_[6589]_ ) & (~\new_[5039]_  | ~\new_[6040]_ );
  assign \new_[4778]_  = ~\new_[4895]_  | (~\new_[5152]_  & ~\new_[5806]_ );
  assign \new_[4779]_  = \new_[4999]_  | \new_[5458]_ ;
  assign \new_[4780]_  = \new_[6287]_  ? \new_[5152]_  : \new_[1892]_ ;
  assign \new_[4781]_  = \new_[5022]_  | \new_[5516]_ ;
  assign \new_[4782]_  = ~\new_[5894]_  | (~\new_[5191]_  & ~\new_[5230]_ );
  assign \new_[4783]_  = \new_[5023]_  | \new_[5191]_ ;
  assign \new_[4784]_  = ~\new_[5088]_  & (~\new_[5275]_  | ~\new_[5161]_ );
  assign \new_[4785]_  = ~\new_[5915]_  | ~\new_[5634]_  | ~\new_[5041]_  | ~\new_[7023]_ ;
  assign \new_[4786]_  = ~\new_[6913]_ ;
  assign \new_[4787]_  = ~\new_[5021]_  | ~\new_[6116]_ ;
  assign \new_[4788]_  = ~\new_[5029]_  | ~\new_[6064]_ ;
  assign \new_[4789]_  = \new_[6290]_  ? \new_[5152]_  : \new_[1925]_ ;
  assign \new_[4790]_  = ~\new_[5030]_  & (~\new_[5307]_  | ~\new_[5601]_ );
  assign \new_[4791]_  = \new_[5940]_  ? \new_[5152]_  : \new_[4554]_ ;
  assign \new_[4792]_  = \new_[6449]_  ? \new_[5152]_  : \new_[2034]_ ;
  assign \new_[4793]_  = ~\new_[5181]_  & ~\new_[5038]_ ;
  assign \new_[4794]_  = ~\new_[5088]_  & (~\new_[5269]_  | ~\new_[5158]_ );
  assign \new_[4795]_  = ~\new_[5088]_  & (~\new_[5274]_  | ~\new_[5164]_ );
  assign \new_[4796]_  = ~\new_[5088]_  & (~\new_[5276]_  | ~\new_[5222]_ );
  assign \new_[4797]_  = ~\new_[5088]_  & (~\new_[5277]_  | ~\new_[5224]_ );
  assign \new_[4798]_  = ~\new_[5035]_  & ~\new_[5994]_ ;
  assign \new_[4799]_  = ~\new_[5088]_  & (~\new_[5271]_  | ~\new_[5166]_ );
  assign \new_[4800]_  = ~\new_[5088]_  & (~\new_[5273]_  | ~\new_[5165]_ );
  assign \new_[4801]_  = ~\new_[5088]_  & (~\new_[5272]_  | ~\new_[5136]_ );
  assign \new_[4802]_  = ~\new_[5651]_  | ~\new_[5034]_  | ~\new_[5354]_ ;
  assign \new_[4803]_  = ~\new_[5399]_  | (~\new_[5226]_  & ~\new_[5393]_ );
  assign \new_[4804]_  = ~\new_[5048]_  & ~\new_[6401]_ ;
  assign \new_[4805]_  = ~\new_[5302]_  | ~\new_[6016]_  | ~\new_[5202]_ ;
  assign \new_[4806]_  = ~\new_[5046]_  | ~\new_[5268]_ ;
  assign \new_[4807]_  = ~\new_[4907]_ ;
  assign \new_[4808]_  = ~\new_[4909]_ ;
  assign \new_[4809]_  = ~\new_[5081]_  & (~\new_[5575]_  | ~\new_[7549]_ );
  assign \new_[4810]_  = ~\new_[5851]_  | ~\new_[5890]_  | ~\new_[5441]_ ;
  assign \new_[4811]_  = ~\new_[5089]_  & (~\new_[5307]_  | ~\new_[5570]_ );
  assign \new_[4812]_  = ~\new_[5089]_  & (~\new_[5187]_  | ~\new_[5570]_ );
  assign \new_[4813]_  = ~\new_[5641]_  | (~\new_[5197]_  & ~\new_[7115]_ );
  assign \new_[4814]_  = ~\new_[5057]_  & (~\new_[7015]_  | ~\new_[6085]_ );
  assign \new_[4815]_  = ~\new_[5447]_  | (~\new_[7017]_  & ~\new_[5399]_ );
  assign \new_[4816]_  = (~\new_[7349]_  | ~\new_[5455]_ ) & (~\new_[5399]_  | ~\new_[5984]_ );
  assign \new_[4817]_  = (~\new_[5660]_  & ~\new_[5187]_ ) | (~\new_[5669]_  & ~\new_[5928]_ );
  assign \new_[4818]_  = (~\new_[5257]_  | ~\new_[5895]_ ) & (~\new_[5399]_  | ~\new_[6961]_ );
  assign \new_[4819]_  = (~\new_[5566]_  | ~\new_[5147]_ ) & (~\new_[5385]_  | ~\new_[5831]_ );
  assign \new_[4820]_  = ~\new_[5530]_  | ~\new_[6128]_ ;
  assign \new_[4821]_  = ~\new_[5401]_  | ~\new_[7209]_ ;
  assign \new_[4822]_  = \new_[5086]_  & \new_[5026]_ ;
  assign \new_[4823]_  = ~\new_[5910]_  | (~\new_[5210]_  & ~\new_[5239]_ );
  assign \new_[4824]_  = \new_[5312]_  & \new_[5104]_ ;
  assign \new_[4825]_  = ~\new_[5526]_  | ~\new_[5455]_ ;
  assign \new_[4826]_  = \new_[5907]_  ? \new_[5152]_  : \new_[4557]_ ;
  assign \new_[4827]_  = ~\new_[5421]_  | ~\new_[5455]_ ;
  assign \new_[4828]_  = ~\new_[5969]_  | ~\new_[5760]_  | ~\new_[5447]_ ;
  assign \new_[4829]_  = ~\new_[5096]_  & (~\new_[5697]_  | ~\new_[5802]_ );
  assign \new_[4830]_  = ~\new_[5529]_  | ~\new_[5331]_ ;
  assign \new_[4831]_  = ~\new_[5359]_  | ~\new_[5870]_  | ~\new_[5857]_  | ~\new_[5665]_ ;
  assign \new_[4832]_  = ~\new_[5927]_  & (~\new_[7017]_  | ~\new_[6325]_ );
  assign \new_[4833]_  = ~\new_[6267]_  | ~\new_[6113]_  | ~\new_[5341]_  | ~\new_[5969]_ ;
  assign \new_[4834]_  = (~\new_[5757]_  | ~\new_[7378]_ ) & (~\new_[5438]_  | ~\new_[5231]_ );
  assign \new_[4835]_  = (~\new_[5228]_  | ~\new_[6075]_ ) & (~\new_[5209]_  | ~\new_[5862]_ );
  assign \new_[4836]_  = (~\new_[5751]_  | ~\new_[6128]_ ) & (~\new_[5209]_  | ~\new_[5767]_ );
  assign \new_[4837]_  = \new_[6084]_  ? \new_[7172]_  : \new_[1861]_ ;
  assign \new_[4838]_  = \new_[6128]_  ? \new_[7172]_  : \new_[1689]_ ;
  assign \new_[4839]_  = ~\new_[4939]_ ;
  assign \new_[4840]_  = ~\new_[7163]_  & ~\new_[5114]_ ;
  assign \new_[4841]_  = \new_[5091]_  & \new_[5862]_ ;
  assign \new_[4842]_  = \new_[5695]_  & \new_[5091]_ ;
  assign \new_[4843]_  = ~\new_[5094]_  | ~\new_[5116]_ ;
  assign \new_[4844]_  = ~\new_[4967]_ ;
  assign \new_[4845]_  = ~\new_[4951]_ ;
  assign \new_[4846]_  = ~\new_[5429]_  | ~\new_[6128]_ ;
  assign \new_[4847]_  = ~\new_[4981]_ ;
  assign \new_[4848]_  = ~\new_[5607]_  | ~\new_[7209]_ ;
  assign \new_[4849]_  = ~\new_[5096]_  & ~\new_[5549]_ ;
  assign \new_[4850]_  = ~\new_[5640]_  | ~\new_[5826]_  | ~\new_[5863]_  | ~\new_[5901]_ ;
  assign \new_[4851]_  = (~\new_[5683]_  | ~\new_[5229]_ ) & (~\new_[5208]_  | ~\new_[6113]_ );
  assign \new_[4852]_  = ~\new_[5582]_  & (~\new_[5225]_  | ~\new_[6227]_ );
  assign \new_[4853]_  = ~\new_[5331]_  | (~\new_[5767]_  & ~\new_[5933]_ );
  assign \new_[4854]_  = (~\new_[5228]_  | ~\new_[6995]_ ) & (~\new_[5802]_  | ~\new_[7116]_ );
  assign \new_[4855]_  = \new_[6986]_  | \new_[5356]_ ;
  assign \new_[4856]_  = ~\new_[5895]_  | ~\new_[5116]_ ;
  assign \new_[4857]_  = ~\new_[7208]_ ;
  assign \new_[4858]_  = ~\new_[5109]_  & ~\new_[6461]_ ;
  assign \new_[4859]_  = ~\new_[5772]_  | ~\new_[5227]_  | ~\new_[5800]_ ;
  assign \new_[4860]_  = ~\new_[5779]_  | ~\new_[5119]_  | ~\new_[2007]_ ;
  assign \new_[4861]_  = ~\new_[5122]_  | ~\new_[6272]_ ;
  assign \new_[4862]_  = ~\new_[5125]_  & ~\new_[5991]_ ;
  assign \new_[4863]_  = ~\new_[5134]_  & ~\new_[2005]_ ;
  assign \new_[4864]_  = ~\new_[6264]_ ;
  assign \new_[4865]_  = ~\new_[6264]_ ;
  assign \new_[4866]_  = ~\new_[6264]_ ;
  assign \new_[4867]_  = ~\new_[5356]_  & ~\new_[6495]_ ;
  assign \new_[4868]_  = \new_[5119]_  | \new_[6654]_ ;
  assign \new_[4869]_  = \new_[6989]_  | \new_[6120]_  | \new_[6967]_  | \new_[5232]_ ;
  assign \new_[4870]_  = ~\new_[5673]_  | ~\new_[5418]_  | ~\new_[5235]_ ;
  assign \new_[4871]_  = ~\new_[5134]_  | ~\new_[2005]_ ;
  assign \new_[4872]_  = ~\new_[5007]_ ;
  assign \new_[4873]_  = ~\new_[4988]_ ;
  assign \new_[4874]_  = \new_[5113]_  | \new_[6011]_ ;
  assign \new_[4875]_  = ~\new_[5696]_  & (~\new_[5241]_  | ~\new_[5659]_ );
  assign \new_[4876]_  = ~\new_[5132]_  | ~\new_[6952]_ ;
  assign \new_[4877]_  = ~\new_[5135]_  & ~\new_[5877]_ ;
  assign \new_[4878]_  = ~\new_[4991]_ ;
  assign \new_[4879]_  = \new_[5912]_  ? \new_[5152]_  : \new_[1646]_ ;
  assign \new_[4880]_  = ~\new_[6670]_  | ~\new_[5641]_ ;
  assign \new_[4881]_  = ~\new_[5142]_  | ~\new_[5376]_ ;
  assign \new_[4882]_  = ~\new_[5928]_  | ~\new_[6107]_  | ~\new_[5261]_ ;
  assign \new_[4883]_  = ~\new_[5152]_  | ~\new_[1861]_ ;
  assign \new_[4884]_  = (~\new_[5394]_  & ~\new_[7550]_ ) | (~\new_[6128]_  & ~\new_[6080]_ );
  assign \new_[4885]_  = ~\new_[5152]_  | ~\new_[2429]_ ;
  assign \new_[4886]_  = ~\new_[5152]_  | ~\new_[4553]_ ;
  assign \new_[4887]_  = ~\new_[5152]_  | ~\new_[4558]_ ;
  assign \new_[4888]_  = ~\new_[5152]_  | ~\new_[4559]_ ;
  assign \new_[4889]_  = ~\new_[5152]_  | ~\new_[4549]_ ;
  assign \new_[4890]_  = ~\new_[5152]_  | ~\new_[4556]_ ;
  assign \new_[4891]_  = ~\new_[5152]_  | ~\new_[1689]_ ;
  assign \new_[4892]_  = \new_[5219]_  | \new_[5669]_ ;
  assign \new_[4893]_  = ~\new_[5152]_  | ~\new_[1578]_ ;
  assign \new_[4894]_  = \new_[5150]_  & \new_[5951]_ ;
  assign \new_[4895]_  = ~\new_[5152]_  | ~\new_[4560]_ ;
  assign \new_[4896]_  = ~\new_[5390]_  | ~\new_[5521]_  | ~\new_[5673]_  | ~\new_[5334]_ ;
  assign \new_[4897]_  = ~\new_[5666]_  | ~\new_[5804]_  | ~\new_[5285]_  | ~\new_[5408]_ ;
  assign \new_[4898]_  = ~\new_[5120]_ ;
  assign \new_[4899]_  = ~\new_[5778]_  | ~\new_[5595]_ ;
  assign \new_[4900]_  = ~\new_[5763]_  | ~\new_[5342]_  | ~\new_[5314]_ ;
  assign \new_[4901]_  = ~\new_[5774]_  | ~\new_[5437]_  | ~\new_[5363]_ ;
  assign \new_[4902]_  = ~\new_[5762]_  | ~\new_[5436]_  | ~\new_[5364]_ ;
  assign \new_[4903]_  = ~\new_[5180]_  | ~\new_[5599]_ ;
  assign \new_[4904]_  = ~\new_[5709]_  | ~\new_[5343]_  | ~\new_[5315]_ ;
  assign \new_[4905]_  = ~\new_[6128]_  | (~\new_[5303]_  & ~\new_[6032]_ );
  assign \new_[4906]_  = ~\new_[5711]_  | ~\new_[5440]_  | ~\new_[5313]_ ;
  assign \new_[4907]_  = ~\new_[5171]_  & ~\new_[5172]_ ;
  assign \new_[4908]_  = ~\new_[5171]_  | ~\new_[6084]_ ;
  assign \new_[4909]_  = ~\new_[5267]_  & (~\new_[2254]_  | ~\new_[7501]_ );
  assign \new_[4910]_  = \new_[5155]_  | \new_[6731]_ ;
  assign \new_[4911]_  = ~\new_[5466]_  & (~\new_[7561]_  | ~\new_[5257]_ );
  assign \new_[4912]_  = ~\new_[5756]_  | ~\new_[5664]_  | ~\new_[5190]_  | ~\new_[5433]_ ;
  assign \new_[4913]_  = ~\new_[5412]_  & (~\new_[5519]_  | ~\new_[5601]_ );
  assign \new_[4914]_  = ~\new_[5289]_  & (~\new_[5305]_  | ~\new_[5889]_ );
  assign \new_[4915]_  = ~\new_[5704]_  | ~\new_[6133]_  | ~\new_[5190]_  | ~\new_[5804]_ ;
  assign \new_[4916]_  = ~\new_[5633]_  & (~\new_[5860]_  | ~\new_[5331]_ );
  assign \new_[4917]_  = (~\new_[7376]_  & ~\new_[5428]_ ) | (~\new_[5872]_  & ~\new_[5298]_ );
  assign \new_[4918]_  = ~\new_[5673]_  | ~\new_[5418]_ ;
  assign \new_[4919]_  = ~\new_[5441]_  | ~\new_[5814]_ ;
  assign \new_[4920]_  = \new_[5398]_  | \new_[6495]_ ;
  assign \new_[4921]_  = \new_[5197]_  & \new_[6348]_ ;
  assign \new_[4922]_  = ~\new_[5206]_  | ~\new_[5760]_ ;
  assign \new_[4923]_  = ~\new_[5220]_  & ~\new_[6340]_ ;
  assign \new_[4924]_  = ~\new_[5045]_ ;
  assign \new_[4925]_  = ~\new_[5725]_  & ~\new_[5399]_ ;
  assign \new_[4926]_  = ~\new_[6013]_  | ~\new_[5185]_  | ~\new_[5742]_ ;
  assign \new_[4927]_  = ~\new_[5220]_  | ~\new_[6011]_ ;
  assign \new_[4928]_  = ~\new_[5196]_  & ~\new_[5200]_ ;
  assign \new_[4929]_  = ~\new_[5199]_  | ~\new_[1545]_ ;
  assign \new_[4930]_  = ~\new_[7466]_  & ~\new_[5295]_ ;
  assign \new_[4931]_  = \new_[5807]_  | \new_[5187]_ ;
  assign \new_[4932]_  = \new_[6216]_  | \new_[5188]_ ;
  assign \new_[4933]_  = ~\new_[5519]_  | ~\new_[6961]_ ;
  assign \new_[4934]_  = ~\new_[5138]_  | ~\new_[5895]_ ;
  assign \new_[4935]_  = ~\new_[5200]_  & ~\new_[5236]_ ;
  assign \new_[4936]_  = \new_[5201]_  & \new_[5636]_ ;
  assign \new_[4937]_  = \new_[5201]_  & \new_[5193]_ ;
  assign \new_[4938]_  = ~\new_[5198]_  & ~\new_[6675]_ ;
  assign \new_[4939]_  = ~\new_[6374]_  & (~\new_[5349]_  | ~\new_[6034]_ );
  assign \new_[4940]_  = ~\new_[5223]_  & ~\new_[6661]_ ;
  assign \new_[4941]_  = ~\new_[5223]_  & ~\new_[6582]_ ;
  assign \new_[4942]_  = ~\new_[5223]_  & ~\new_[6578]_ ;
  assign \new_[4943]_  = ~\new_[5223]_  & ~\new_[6575]_ ;
  assign \new_[4944]_  = ~\new_[5223]_  & ~\new_[6662]_ ;
  assign \new_[4945]_  = ~\new_[5223]_  & ~\new_[6535]_ ;
  assign \new_[4946]_  = ~\new_[5223]_  & ~\new_[6653]_ ;
  assign \new_[4947]_  = ~\new_[5223]_  & ~\new_[6568]_ ;
  assign \new_[4948]_  = ~\new_[5223]_  & ~\new_[6626]_ ;
  assign \new_[4949]_  = ~\new_[5223]_  & ~\new_[6676]_ ;
  assign \new_[4950]_  = ~\new_[5223]_  & ~\new_[6613]_ ;
  assign \new_[4951]_  = ~\new_[5234]_  & ~\new_[7159]_ ;
  assign \new_[4952]_  = ~\new_[5223]_  & ~\new_[6677]_ ;
  assign \new_[4953]_  = ~\new_[5223]_  & ~\new_[6646]_ ;
  assign \new_[4954]_  = ~\new_[5223]_  & ~\new_[6604]_ ;
  assign \new_[4955]_  = ~\new_[5223]_  & ~\new_[6550]_ ;
  assign \new_[4956]_  = ~\new_[7163]_  & ~\new_[5688]_ ;
  assign \new_[4957]_  = ~\new_[7172]_  & ~\new_[6271]_ ;
  assign \new_[4958]_  = ~\new_[5219]_  & ~\new_[5859]_ ;
  assign \new_[4959]_  = ~\new_[7315]_  | ~\new_[5428]_ ;
  assign \new_[4960]_  = \new_[5219]_  | \new_[5947]_ ;
  assign \new_[4961]_  = ~\new_[5239]_  | ~\new_[5862]_ ;
  assign \new_[4962]_  = \new_[7378]_  | \new_[5994]_ ;
  assign \new_[4963]_  = \new_[6016]_  | \new_[7017]_ ;
  assign \new_[4964]_  = \new_[5598]_  | \new_[5768]_ ;
  assign \new_[4965]_  = ~\new_[5211]_  | ~\new_[6106]_ ;
  assign \new_[4966]_  = ~\new_[6465]_  | ~\new_[5211]_  | ~\new_[6891]_ ;
  assign \new_[4967]_  = ~\new_[5221]_  & ~\new_[758]_ ;
  assign \new_[4968]_  = ~\new_[5598]_  | ~\new_[5752]_ ;
  assign \new_[4969]_  = ~\new_[5084]_ ;
  assign \new_[4970]_  = ~\new_[7008]_  & ~\new_[7200]_ ;
  assign \new_[4971]_  = ~\new_[5635]_  & ~\new_[5570]_ ;
  assign \new_[4972]_  = ~\new_[5239]_  | ~\new_[5767]_ ;
  assign \new_[4973]_  = ~\new_[5234]_  | ~\new_[6060]_ ;
  assign \new_[4974]_  = ~\new_[7378]_  | ~\new_[6405]_ ;
  assign \new_[4975]_  = ~\new_[5710]_  | ~\new_[5231]_ ;
  assign \new_[4976]_  = ~\new_[7006]_  & ~\new_[5234]_ ;
  assign \new_[4977]_  = ~\new_[7017]_  | ~\new_[6113]_ ;
  assign \new_[4978]_  = ~\new_[5215]_  | ~\new_[5831]_ ;
  assign \new_[4979]_  = ~\new_[5234]_  | ~\new_[7070]_ ;
  assign \new_[4980]_  = ~\new_[5426]_  | ~\new_[5598]_ ;
  assign \new_[4981]_  = ~\new_[5221]_  & ~\new_[759]_ ;
  assign \new_[4982]_  = ~\new_[5083]_ ;
  assign \new_[4983]_  = \new_[5212]_  & \new_[5776]_ ;
  assign \new_[4984]_  = ~\new_[5223]_  & ~\new_[6557]_ ;
  assign \new_[4985]_  = ~\new_[5443]_  | ~\new_[5772]_ ;
  assign \new_[4986]_  = ~\new_[5455]_  & (~\new_[5859]_  | ~\new_[6175]_ );
  assign \new_[4987]_  = ~\new_[7116]_  | ~\new_[5595]_ ;
  assign \new_[4988]_  = ~\new_[6397]_  | ~\new_[7550]_ ;
  assign \new_[4989]_  = ~\new_[5947]_  & ~\new_[6400]_ ;
  assign \new_[4990]_  = ~\new_[5875]_  & ~\new_[5601]_ ;
  assign \new_[4991]_  = \new_[5232]_  & \new_[5772]_ ;
  assign \new_[4992]_  = ~\new_[5458]_  & (~\new_[5350]_  | ~\new_[6593]_ );
  assign \new_[4993]_  = ~\new_[5915]_  & ~\new_[5688]_ ;
  assign \new_[4994]_  = ~\new_[6084]_  | ~\new_[6113]_  | ~\new_[5141]_  | ~\new_[6267]_ ;
  assign \new_[4995]_  = ~\new_[5675]_  | (~\new_[6461]_  & ~\new_[6080]_ );
  assign \new_[4996]_  = ~\new_[5125]_ ;
  assign \new_[4997]_  = ~\new_[6462]_  | ~\new_[5969]_  | ~\new_[5229]_  | ~\new_[5823]_ ;
  assign \new_[4998]_  = ~\new_[5220]_  & ~\new_[6310]_ ;
  assign \new_[4999]_  = ~\new_[5238]_  & ~\new_[2016]_ ;
  assign \new_[5000]_  = ~\new_[5238]_  | ~\new_[2016]_ ;
  assign \new_[5001]_  = ~\new_[2430]_  & ~\new_[7505]_ ;
  assign \new_[5002]_  = ~\new_[5692]_  & ~\new_[5772]_ ;
  assign \new_[5003]_  = ~\new_[7163]_  | ~\new_[5192]_ ;
  assign \new_[5004]_  = ~\new_[5581]_  & (~\new_[7549]_  | ~\new_[7253]_ );
  assign \new_[5005]_  = \new_[5232]_  | \new_[7550]_ ;
  assign \new_[5006]_  = \new_[5358]_  ? \new_[5696]_  : \new_[5718]_ ;
  assign \new_[5007]_  = \new_[5232]_  & \new_[5884]_ ;
  assign \new_[5008]_  = ~\new_[6084]_  & ~\new_[6227]_ ;
  assign \new_[5009]_  = ~\new_[5243]_  & ~\new_[5877]_ ;
  assign \new_[5010]_  = ~\new_[5113]_ ;
  assign \new_[5011]_  = ~\new_[5240]_  | (~\new_[5613]_  & ~\new_[5454]_ );
  assign \new_[5012]_  = ~\new_[5134]_ ;
  assign \new_[5013]_  = ~\new_[5228]_  | ~\new_[5958]_ ;
  assign \new_[5014]_  = ~\new_[5133]_ ;
  assign \new_[5015]_  = ~\new_[5219]_  & ~\new_[5896]_ ;
  assign \new_[5016]_  = \new_[5643]_  ? \new_[5250]_  : \new_[5735]_ ;
  assign \new_[5017]_  = \new_[5451]_  | \new_[5116]_ ;
  assign \new_[5018]_  = ~\new_[5221]_ ;
  assign \new_[5019]_  = ~\new_[5137]_ ;
  assign \new_[5020]_  = \new_[3264]_  ? \new_[5439]_  : \new_[6521]_ ;
  assign \new_[5021]_  = ~\new_[5310]_  | ~\new_[6004]_ ;
  assign \new_[5022]_  = ~\new_[5893]_  | ~\new_[5381]_  | ~\new_[5512]_  | ~\new_[7163]_ ;
  assign \new_[5023]_  = ~\new_[6457]_  & (~\new_[5598]_  | ~\new_[5380]_ );
  assign \new_[5024]_  = ~\new_[5376]_  | (~\new_[6083]_  & ~\new_[6316]_ );
  assign \new_[5025]_  = \new_[5384]_  ^ \new_[5662]_ ;
  assign \new_[5026]_  = \new_[5758]_  | \new_[5331]_ ;
  assign \new_[5027]_  = ~\new_[5955]_  | ~\new_[5817]_  | ~\new_[5599]_  | ~\new_[5461]_ ;
  assign \new_[5028]_  = ~\new_[5265]_  & ~\new_[5723]_ ;
  assign \new_[5029]_  = ~\new_[5259]_  | ~\new_[7180]_ ;
  assign \new_[5030]_  = ~\new_[5470]_  | ~\new_[5386]_  | ~\new_[5391]_ ;
  assign \new_[5031]_  = \new_[5288]_  | \new_[7563]_ ;
  assign \new_[5032]_  = ~\new_[5391]_  | ~\new_[5512]_  | ~\new_[6003]_ ;
  assign \new_[5033]_  = \new_[5260]_  & \new_[5764]_ ;
  assign \new_[5034]_  = ~\new_[5281]_  & ~\new_[6961]_ ;
  assign \new_[5035]_  = ~\new_[5334]_  | (~\new_[7376]_  & ~\new_[5802]_ );
  assign \new_[5036]_  = ~\new_[5898]_  | ~\new_[5658]_  | ~\new_[5655]_  | ~\new_[5419]_ ;
  assign \new_[5037]_  = \new_[7013]_  & \new_[7238]_ ;
  assign \new_[5038]_  = ~\new_[5556]_  | ~\new_[5285]_  | ~\new_[5408]_ ;
  assign \new_[5039]_  = ~\new_[6118]_  | ~\new_[5533]_  | ~\new_[5564]_  | ~\new_[5473]_ ;
  assign \new_[5040]_  = ~\new_[5406]_  & (~\new_[5407]_  | ~\new_[6128]_ );
  assign \new_[5041]_  = ~\new_[5151]_ ;
  assign \new_[5042]_  = (~\new_[5988]_  & ~\new_[5455]_ ) | (~\new_[5399]_  & ~\new_[5981]_ );
  assign \new_[5043]_  = ~\new_[5462]_  | ~\new_[5693]_  | ~\new_[5880]_  | ~\new_[5898]_ ;
  assign \new_[5044]_  = ~\new_[5257]_  | ~\new_[6006]_ ;
  assign \new_[5045]_  = ~\new_[2431]_  | ~\new_[7501]_ ;
  assign \new_[5046]_  = ~\new_[5561]_  & (~\new_[5456]_  | ~\new_[5786]_ );
  assign \new_[5047]_  = ~\new_[5307]_  | ~\new_[5984]_ ;
  assign \new_[5048]_  = ~\new_[5168]_ ;
  assign \new_[5049]_  = ~\new_[2780]_  | ~\new_[5546]_ ;
  assign \new_[5050]_  = ~\new_[5807]_  & ~\new_[5399]_ ;
  assign \new_[5051]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5424]_ );
  assign \new_[5052]_  = ~\new_[6041]_  & (~\new_[5538]_  | ~\new_[5434]_ );
  assign \new_[5053]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5422]_ );
  assign \new_[5054]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5423]_ );
  assign \new_[5055]_  = ~\new_[5545]_  | ~\new_[5556]_  | ~\new_[5541]_  | ~\new_[5553]_ ;
  assign \new_[5056]_  = ~\new_[5452]_  & (~\new_[5438]_  | ~\new_[6015]_ );
  assign \new_[5057]_  = ~\new_[7016]_ ;
  assign \new_[5058]_  = (~\new_[5555]_  | ~\new_[7378]_ ) & (~\new_[5592]_  | ~\new_[5438]_ );
  assign \new_[5059]_  = \new_[753]_  ? \new_[5439]_  : \new_[3271]_ ;
  assign \new_[5060]_  = \new_[740]_  ? \new_[5439]_  : \new_[3261]_ ;
  assign \new_[5061]_  = \new_[736]_  ? \new_[5439]_  : \new_[3267]_ ;
  assign \new_[5062]_  = \new_[6520]_  ? \new_[5439]_  : \new_[3263]_ ;
  assign \new_[5063]_  = \new_[6606]_  ? \new_[5439]_  : \new_[3262]_ ;
  assign \new_[5064]_  = \new_[6591]_  ? \new_[5439]_  : \new_[3251]_ ;
  assign \new_[5065]_  = \new_[6472]_  ? \new_[5439]_  : \new_[3266]_ ;
  assign \new_[5066]_  = \new_[844]_  ? \new_[5439]_  : \new_[3259]_ ;
  assign \new_[5067]_  = \new_[850]_  ? \new_[5439]_  : \new_[3265]_ ;
  assign \new_[5068]_  = \new_[762]_  ? \new_[5439]_  : \new_[3260]_ ;
  assign \new_[5069]_  = \new_[761]_  ? \new_[5439]_  : \new_[3268]_ ;
  assign \new_[5070]_  = \new_[758]_  ? \new_[5439]_  : \new_[3254]_ ;
  assign \new_[5071]_  = \new_[763]_  ? \new_[5439]_  : \new_[3269]_ ;
  assign \new_[5072]_  = \new_[759]_  ? \new_[5439]_  : \new_[3257]_ ;
  assign \new_[5073]_  = \new_[760]_  ? \new_[5439]_  : \new_[3270]_ ;
  assign \new_[5074]_  = \new_[6521]_  ? \new_[5439]_  : \new_[3264]_ ;
  assign \new_[5075]_  = \new_[3266]_  ? \new_[5439]_  : \new_[6472]_ ;
  assign \new_[5076]_  = \new_[3259]_  ? \new_[5439]_  : \new_[844]_ ;
  assign \new_[5077]_  = ~\new_[5860]_  | ~\new_[7209]_ ;
  assign \new_[5078]_  = ~\new_[6571]_  | ~\new_[6284]_  | ~\new_[6523]_  | ~\new_[5894]_ ;
  assign \new_[5079]_  = ~\new_[5799]_  | ~\new_[5598]_ ;
  assign \new_[5080]_  = ~\new_[5236]_ ;
  assign \new_[5081]_  = ~\new_[5189]_ ;
  assign \new_[5082]_  = \new_[5429]_  | \new_[6961]_ ;
  assign \new_[5083]_  = ~\new_[6107]_  | ~\new_[7209]_  | ~\new_[6233]_ ;
  assign \new_[5084]_  = \new_[5910]_  & \new_[7201]_ ;
  assign \new_[5085]_  = ~\new_[5193]_ ;
  assign \new_[5086]_  = ~\new_[7379]_  | ~\new_[5598]_ ;
  assign \new_[5087]_  = ~\new_[7377]_  | ~\new_[5758]_ ;
  assign \new_[5088]_  = \new_[5429]_  & \new_[6315]_ ;
  assign \new_[5089]_  = \new_[5598]_  & \new_[5635]_ ;
  assign \new_[5090]_  = ~\new_[5739]_  | ~\new_[6084]_ ;
  assign \new_[5091]_  = \new_[5443]_  & \new_[6128]_ ;
  assign \new_[5092]_  = ~\new_[5220]_ ;
  assign \new_[5093]_  = ~\new_[5233]_ ;
  assign \new_[5094]_  = ~\new_[5896]_  | ~\new_[5669]_ ;
  assign \new_[5095]_  = ~\new_[5209]_ ;
  assign \new_[5096]_  = ~\new_[5669]_  & ~\new_[6071]_ ;
  assign \new_[5097]_  = ~\new_[5353]_  | ~\new_[6995]_ ;
  assign \new_[5098]_  = ~\new_[5353]_  | ~\new_[6075]_ ;
  assign \new_[5099]_  = ~\new_[4554]_  | ~\new_[5724]_ ;
  assign \new_[5100]_  = ~\new_[4549]_  | ~\new_[5724]_ ;
  assign \new_[5101]_  = ~\new_[5530]_  | ~\new_[7209]_ ;
  assign \new_[5102]_  = ~\new_[4560]_  | ~\new_[5724]_ ;
  assign \new_[5103]_  = ~\new_[5689]_  & ~\new_[5357]_ ;
  assign \new_[5104]_  = ~\new_[5767]_  | ~\new_[6284]_ ;
  assign \new_[5105]_  = ~\new_[4557]_  | ~\new_[5724]_ ;
  assign \new_[5106]_  = ~\new_[5571]_  & (~\new_[6084]_  | ~\new_[5972]_ );
  assign \new_[5107]_  = (~\new_[6462]_  | ~\new_[6397]_ ) & (~\new_[6394]_  | ~\new_[6113]_ );
  assign \new_[5108]_  = (~\new_[6478]_  | ~\new_[7050]_ ) & (~\new_[1324]_  | ~\new_[5705]_ );
  assign \new_[5109]_  = ~\new_[5225]_ ;
  assign \new_[5110]_  = ~\new_[4559]_  | ~\new_[5724]_ ;
  assign \new_[5111]_  = ~\new_[5459]_  | ~\new_[740]_ ;
  assign \new_[5112]_  = \new_[5352]_  & \new_[6465]_ ;
  assign \new_[5113]_  = \new_[5350]_  | \new_[6593]_ ;
  assign \new_[5114]_  = ~\new_[5231]_ ;
  assign \new_[5115]_  = ~\new_[5238]_ ;
  assign \new_[5116]_  = ~\new_[5688]_ ;
  assign \new_[5117]_  = ~\new_[6325]_  & ~\new_[5356]_ ;
  assign \new_[5118]_  = ~\new_[6049]_  & ~\new_[5884]_ ;
  assign \new_[5119]_  = ~\new_[5347]_  | ~\new_[5884]_ ;
  assign \new_[5120]_  = ~\new_[5769]_  | ~\new_[6013]_  | ~\new_[7120]_  | ~\new_[7159]_ ;
  assign \new_[5121]_  = ~\new_[4556]_  | ~\new_[5724]_ ;
  assign \new_[5122]_  = ~\new_[6227]_  | ~\new_[6307]_  | ~\new_[6445]_ ;
  assign \new_[5123]_  = \new_[5823]_  & \new_[6193]_ ;
  assign \new_[5124]_  = i_tv80_core_NMI_s_reg;
  assign \new_[5125]_  = ~\new_[6216]_  | (~\new_[5641]_  & ~\new_[6272]_ );
  assign \new_[5126]_  = ~\new_[5613]_  | ~\new_[5361]_ ;
  assign \new_[5127]_  = ~\new_[5994]_  | ~\new_[6084]_ ;
  assign \new_[5128]_  = ~\new_[4553]_  | ~\new_[5724]_ ;
  assign \new_[5129]_  = (~\new_[5369]_  | ~\new_[6953]_ ) & (~\new_[6352]_  | ~\new_[5959]_ );
  assign \new_[5130]_  = (~\new_[6344]_  | ~\new_[6037]_ ) & (~\new_[5369]_  | ~\new_[6952]_ );
  assign \new_[5131]_  = ~\new_[4558]_  | ~\new_[5724]_ ;
  assign \new_[5132]_  = \new_[5370]_  ^ \new_[5464]_ ;
  assign \new_[5133]_  = ~\new_[5475]_  | ~\new_[5815]_  | ~\new_[5367]_  | ~\new_[5745]_ ;
  assign \new_[5134]_  = \new_[5347]_  & \new_[5772]_ ;
  assign \new_[5135]_  = \new_[5374]_  ? \new_[6625]_  : \new_[5372]_ ;
  assign \new_[5136]_  = ~\new_[5403]_  | ~\new_[6518]_ ;
  assign \new_[5137]_  = ~\new_[5388]_  & (~\new_[5820]_  | ~\new_[5729]_ );
  assign \new_[5138]_  = ~\new_[5257]_ ;
  assign \new_[5139]_  = \new_[6223]_  ^ \new_[5479]_ ;
  assign \new_[5140]_  = \new_[5375]_  & \new_[5951]_ ;
  assign \new_[5141]_  = ~\new_[5776]_  & ~\new_[6031]_ ;
  assign \new_[5142]_  = ~\new_[850]_  | ~\new_[6565]_  | ~\new_[6436]_  | ~\new_[6173]_ ;
  assign \new_[5143]_  = \new_[5504]_  | \new_[5387]_ ;
  assign \new_[5144]_  = \new_[6933]_  & \new_[7564]_ ;
  assign \new_[5145]_  = ~\new_[5435]_  & (~\new_[5906]_  | ~\new_[7116]_ );
  assign \new_[5146]_  = \new_[6926]_  ? \new_[6264]_  : \new_[845]_ ;
  assign \new_[5147]_  = ~\new_[5970]_  & ~\new_[5443]_ ;
  assign \new_[5148]_  = ~\new_[5259]_ ;
  assign \new_[5149]_  = \new_[6227]_  ? \new_[5680]_  : \di[1] ;
  assign \new_[5150]_  = ~\new_[7158]_  | ~\new_[7201]_  | ~\new_[5519]_ ;
  assign \new_[5151]_  = ~\new_[6168]_  | ~\new_[5880]_  | ~\new_[7024]_  | ~\new_[5532]_ ;
  assign \new_[5152]_  = (~\new_[5583]_  | ~\new_[6313]_ ) & (~\new_[5522]_  | ~\new_[6315]_ );
  assign \new_[5153]_  = ~\new_[5409]_  & (~\new_[5608]_  | ~\new_[6128]_ );
  assign \new_[5154]_  = ~\new_[6251]_  | ~\new_[5413]_ ;
  assign \new_[5155]_  = \new_[2928]_  & \new_[5397]_ ;
  assign \new_[5156]_  = ~\new_[2930]_  | ~\new_[5397]_ ;
  assign \new_[5157]_  = ~\new_[5268]_ ;
  assign \new_[5158]_  = ~\new_[5403]_  | ~\new_[6478]_ ;
  assign \new_[5159]_  = ~\new_[5279]_ ;
  assign \new_[5160]_  = ~\new_[6193]_  | ~\new_[5522]_  | ~\new_[6284]_ ;
  assign \new_[5161]_  = ~\new_[5403]_  | ~\new_[6548]_ ;
  assign \new_[5162]_  = \new_[5951]_  & \new_[5413]_ ;
  assign \new_[5163]_  = ~\new_[5866]_  | ~\new_[5385]_ ;
  assign \new_[5164]_  = ~\new_[5403]_  | ~\new_[6528]_ ;
  assign \new_[5165]_  = ~\new_[5403]_  | ~\new_[6542]_ ;
  assign \new_[5166]_  = ~\new_[5403]_  | ~\new_[6515]_ ;
  assign \new_[5167]_  = ~\new_[5536]_  | ~\new_[5928]_ ;
  assign \new_[5168]_  = ~\new_[5620]_  & ~\new_[6495]_ ;
  assign \new_[5169]_  = \new_[5994]_  | \new_[5404]_ ;
  assign \new_[5170]_  = \new_[7238]_  & \new_[7239]_ ;
  assign \new_[5171]_  = ~\new_[5462]_  | ~\new_[5366]_ ;
  assign \new_[5172]_  = ~\new_[5373]_  | ~\new_[5880]_ ;
  assign \new_[5173]_  = ~\new_[5287]_ ;
  assign \new_[5174]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5537]_ );
  assign \new_[5175]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5539]_ );
  assign \new_[5176]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5585]_ );
  assign \new_[5177]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5589]_ );
  assign \new_[5178]_  = ~\new_[5450]_  | (~\new_[5616]_  & ~\new_[5540]_ );
  assign \new_[5179]_  = (~\new_[5710]_  | ~\new_[5592]_ ) & (~\new_[5543]_  | ~\new_[6128]_ );
  assign \new_[5180]_  = ~\new_[5291]_ ;
  assign \new_[5181]_  = ~\new_[5396]_  | ~\new_[7120]_ ;
  assign \new_[5182]_  = ~\new_[5248]_ ;
  assign \new_[5183]_  = ~\new_[5247]_ ;
  assign \new_[5184]_  = ~\new_[5295]_ ;
  assign \new_[5185]_  = ~\new_[5296]_ ;
  assign \new_[5186]_  = ~\new_[5807]_  & ~\new_[6071]_ ;
  assign \new_[5187]_  = ~\new_[5399]_ ;
  assign \new_[5188]_  = \new_[5434]_  & \new_[5995]_ ;
  assign \new_[5189]_  = ~\new_[5985]_  | ~\new_[5805]_ ;
  assign \new_[5190]_  = \new_[5807]_  & \new_[6175]_ ;
  assign \new_[5191]_  = ~\new_[7200]_  & ~\new_[6803]_ ;
  assign \new_[5192]_  = ~\new_[5300]_ ;
  assign \new_[5193]_  = ~\new_[6961]_  | ~\new_[5595]_ ;
  assign \new_[5194]_  = ~\new_[5805]_  | ~\new_[5927]_ ;
  assign \new_[5195]_  = ~\new_[5994]_  | ~\new_[5428]_ ;
  assign \new_[5196]_  = ~\new_[5891]_  & ~\new_[5455]_ ;
  assign \new_[5197]_  = ~\new_[7440]_  & ~\new_[7335]_ ;
  assign \new_[5198]_  = ~\new_[5432]_  & ~\new_[6365]_ ;
  assign \new_[5199]_  = ~\new_[5304]_ ;
  assign \new_[5200]_  = ~\new_[7200]_  & ~\new_[5950]_ ;
  assign \new_[5201]_  = ~\new_[5429]_  | ~\new_[5595]_ ;
  assign \new_[5202]_  = ~\new_[7378]_  | ~\new_[6124]_ ;
  assign \new_[5203]_  = ~\new_[6133]_  | ~\new_[5554]_  | ~\new_[5915]_ ;
  assign \new_[5204]_  = ~\new_[5371]_  & (~\new_[1324]_  | ~\new_[6819]_ );
  assign \new_[5205]_  = ~\new_[5894]_  | ~\new_[6378]_  | ~\new_[6305]_ ;
  assign \new_[5206]_  = \new_[5617]_  | \new_[5897]_  | \new_[5864]_  | \new_[5786]_ ;
  assign \new_[5207]_  = \new_[5720]_  | \new_[5928]_ ;
  assign \new_[5208]_  = ~\new_[5705]_  | ~\new_[5823]_ ;
  assign \new_[5209]_  = ~\new_[5966]_  & ~\new_[5443]_ ;
  assign \new_[5210]_  = ~\new_[5443]_  & ~\new_[6400]_ ;
  assign \new_[5211]_  = ~\new_[5442]_  & ~\new_[6031]_ ;
  assign \new_[5212]_  = \new_[5442]_  | \new_[6484]_ ;
  assign \new_[5213]_  = ~\new_[5674]_  | ~\new_[5595]_ ;
  assign \new_[5214]_  = \new_[5417]_  | \new_[5552]_ ;
  assign \new_[5215]_  = ~\new_[5443]_  & ~\new_[5859]_ ;
  assign \new_[5216]_  = ~\new_[5988]_  & ~\new_[6394]_ ;
  assign \new_[5217]_  = ~\new_[6284]_  | ~\new_[5894]_  | ~\new_[6519]_ ;
  assign \new_[5218]_  = \new_[5394]_  | \new_[6227]_ ;
  assign \new_[5219]_  = ~\new_[5451]_  & (~\new_[6394]_  | ~\new_[5927]_ );
  assign \new_[5220]_  = ~\new_[1624]_  | ~\new_[1810]_  | ~\new_[5587]_ ;
  assign \new_[5221]_  = ~\new_[6465]_  | ~\new_[6400]_  | ~\new_[5445]_  | ~\new_[6267]_ ;
  assign \new_[5222]_  = ~\new_[5403]_  | ~\new_[2007]_ ;
  assign \new_[5223]_  = ~\new_[6523]_  | ~\new_[5889]_  | ~\new_[6603]_  | ~\new_[3281]_ ;
  assign \new_[5224]_  = ~\new_[5403]_  | ~\new_[2005]_ ;
  assign \new_[5225]_  = ~\new_[5775]_  & ~\new_[6400]_ ;
  assign \new_[5226]_  = ~\new_[5428]_  | ~\new_[5889]_ ;
  assign \new_[5227]_  = ~\new_[5357]_ ;
  assign \new_[5228]_  = ~\new_[5688]_  & ~\new_[7550]_ ;
  assign \new_[5229]_  = \new_[5446]_  & \new_[6039]_ ;
  assign \new_[5230]_  = ~\new_[6457]_  & ~\new_[5380]_ ;
  assign \new_[5231]_  = ~\new_[6400]_  & ~\new_[5688]_ ;
  assign \new_[5232]_  = ~\new_[6084]_  & ~\new_[6143]_ ;
  assign \new_[5233]_  = \new_[6986]_  | \new_[5688]_ ;
  assign \new_[5234]_  = ~\new_[7201]_ ;
  assign \new_[5235]_  = ~\new_[5695]_  | ~\new_[5443]_ ;
  assign \new_[5236]_  = ~\new_[6986]_  & ~\new_[7017]_ ;
  assign \new_[5237]_  = \new_[5460]_  ? \new_[5696]_  : \new_[5811]_ ;
  assign \new_[5238]_  = \new_[6462]_  & \new_[5772]_ ;
  assign \new_[5239]_  = ~\new_[5443]_  & ~\new_[6394]_ ;
  assign \new_[5240]_  = ~\new_[5613]_  | ~\new_[5454]_ ;
  assign \new_[5241]_  = ~\new_[5718]_  & (~\new_[5603]_  | ~\new_[5811]_ );
  assign \new_[5242]_  = ~\new_[5442]_  & ~\new_[7049]_ ;
  assign \new_[5243]_  = (~\new_[5457]_  | ~\new_[6625]_ ) & (~\new_[5707]_  | ~\new_[740]_ );
  assign \new_[5244]_  = ~\new_[5370]_  & ~\new_[5464]_ ;
  assign \new_[5245]_  = \new_[5365]_  | \new_[5877]_ ;
  assign \new_[5246]_  = ~\new_[5362]_ ;
  assign \new_[5247]_  = ~\new_[5486]_  & ~\new_[6264]_ ;
  assign \new_[5248]_  = ~\new_[5598]_  & ~\new_[6523]_ ;
  assign \new_[5249]_  = ~\new_[5467]_  & ~\new_[5877]_ ;
  assign \new_[5250]_  = ~\new_[6087]_  | (~\new_[5619]_  & ~\new_[6026]_ );
  assign \new_[5251]_  = \new_[3606]_  ? \new_[6271]_  : \A[12] ;
  assign \new_[5252]_  = \new_[3638]_  ? \new_[5724]_  : \A[9] ;
  assign \new_[5253]_  = ~\new_[5479]_  & ~\new_[6223]_ ;
  assign \new_[5254]_  = \new_[3626]_  ? \new_[5724]_  : \A[8] ;
  assign \new_[5255]_  = ~\new_[5864]_  & ~\new_[5617]_ ;
  assign \new_[5256]_  = (~\new_[5835]_  | ~\new_[6047]_ ) & (~\new_[799]_  | ~\new_[6264]_ );
  assign \new_[5257]_  = ~\new_[6107]_  | ~\new_[5598]_  | ~\new_[6006]_ ;
  assign \new_[5258]_  = (~\new_[7188]_  | ~\new_[6047]_ ) & (~\new_[849]_  | ~\new_[6264]_ );
  assign \new_[5259]_  = ~\new_[5511]_  | ~\new_[6234]_ ;
  assign \new_[5260]_  = \new_[5736]_  & \new_[5512]_ ;
  assign \new_[5261]_  = ~\new_[5234]_  | ~\new_[5630]_ ;
  assign \new_[5262]_  = ~\new_[5883]_  | ~\new_[5621]_  | ~\new_[5804]_ ;
  assign \new_[5263]_  = ~\new_[5383]_ ;
  assign \new_[5264]_  = ~\new_[6003]_  | ~\new_[5544]_  | ~\new_[5801]_ ;
  assign \new_[5265]_  = ~\new_[5557]_  | ~\new_[5932]_ ;
  assign \new_[5266]_  = \new_[2633]_  ? \new_[6271]_  : \A[0] ;
  assign \new_[5267]_  = \new_[2780]_  & \new_[6731]_ ;
  assign \new_[5268]_  = ~\new_[5520]_  & ~\new_[5525]_ ;
  assign \new_[5269]_  = ~\new_[5503]_  | ~\new_[6528]_ ;
  assign \new_[5270]_  = ~\new_[6481]_  | ~\new_[5588]_  | ~\new_[5672]_ ;
  assign \new_[5271]_  = ~\new_[5503]_  | ~\new_[6548]_ ;
  assign \new_[5272]_  = ~\new_[5503]_  | ~\new_[2007]_ ;
  assign \new_[5273]_  = ~\new_[5503]_  | ~\new_[2005]_ ;
  assign \new_[5274]_  = ~\new_[5503]_  | ~\new_[2003]_ ;
  assign \new_[5275]_  = ~\new_[5503]_  | ~\new_[2006]_ ;
  assign \new_[5276]_  = ~\new_[5503]_  | ~\new_[2002]_ ;
  assign \new_[5277]_  = ~\new_[5503]_  | ~\new_[2016]_ ;
  assign \new_[5278]_  = ~\new_[5532]_  | ~\new_[5634]_ ;
  assign \new_[5279]_  = \new_[5521]_  & \new_[5548]_ ;
  assign \new_[5280]_  = \new_[5523]_  & \new_[5639]_ ;
  assign \new_[5281]_  = ~\new_[5390]_ ;
  assign \new_[5282]_  = ~\new_[5575]_  | ~\new_[6113]_ ;
  assign \new_[5283]_  = \new_[5536]_  | \new_[5864]_ ;
  assign \new_[5284]_  = \new_[5994]_  | \new_[5522]_ ;
  assign \new_[5285]_  = \new_[5476]_  & \new_[5468]_ ;
  assign \new_[5286]_  = \new_[5551]_  & \new_[7153]_ ;
  assign \new_[5287]_  = ~\new_[6102]_  & (~\new_[7163]_  | ~\new_[5893]_ );
  assign \new_[5288]_  = ~\new_[5513]_  | ~\new_[6933]_ ;
  assign \new_[5289]_  = ~\new_[5787]_  & (~\new_[5612]_  | ~\new_[5826]_ );
  assign \new_[5290]_  = \new_[3600]_  ? \new_[6271]_  : \A[13] ;
  assign \new_[5291]_  = ~\new_[5741]_  | ~\new_[5948]_  | ~\new_[5903]_  | ~\new_[5987]_ ;
  assign \new_[5292]_  = ~\new_[5627]_  | ~\new_[6128]_ ;
  assign \new_[5293]_  = ~\new_[5430]_ ;
  assign \new_[5294]_  = ~\new_[5395]_ ;
  assign \new_[5295]_  = ~\new_[5397]_ ;
  assign \new_[5296]_  = \new_[7005]_  | \new_[7116]_ ;
  assign \new_[5297]_  = ~\new_[5406]_ ;
  assign \new_[5298]_  = \new_[7201]_  & \new_[6006]_ ;
  assign \new_[5299]_  = \new_[7163]_  | \new_[5234]_ ;
  assign \new_[5300]_  = \new_[5710]_  | \new_[5958]_ ;
  assign \new_[5301]_  = ~\new_[5765]_  | ~\new_[5554]_  | ~\new_[6168]_ ;
  assign \new_[5302]_  = ~\new_[6325]_  | ~\new_[7378]_  | ~\new_[6305]_ ;
  assign \new_[5303]_  = ~\new_[5441]_ ;
  assign \new_[5304]_  = ~\new_[5641]_  & ~\new_[6264]_ ;
  assign \new_[5305]_  = ~\new_[5640]_  | ~\new_[5863]_  | ~\new_[5901]_ ;
  assign \new_[5306]_  = ~\new_[6266]_  | ~\new_[7201]_ ;
  assign \new_[5307]_  = ~\new_[5234]_  | ~\new_[5787]_ ;
  assign \new_[5308]_  = (~\new_[5674]_  | ~\new_[6359]_ ) & (~\new_[7116]_  | ~\new_[6405]_ );
  assign n1869 = ~\new_[6441]_  & ~\new_[5754]_  & ~\new_[6519]_ ;
  assign \new_[5310]_  = ~\new_[5511]_  | ~\new_[5234]_ ;
  assign \new_[5311]_  = ~\new_[5712]_  & (~\new_[5862]_  | ~\new_[5927]_ );
  assign \new_[5312]_  = ~\new_[6284]_  | (~\new_[5674]_  & ~\new_[6064]_ );
  assign \new_[5313]_  = (~\new_[5679]_  | ~\new_[6518]_ ) & (~\new_[5861]_  | ~\new_[6478]_ );
  assign \new_[5314]_  = (~\new_[5679]_  | ~\new_[1247]_ ) & (~\new_[5861]_  | ~\new_[6518]_ );
  assign \new_[5315]_  = (~\new_[5679]_  | ~\new_[1248]_ ) & (~\new_[5861]_  | ~\new_[1247]_ );
  assign \new_[5316]_  = \new_[2661]_  ? \new_[6271]_  : \A[1] ;
  assign \new_[5317]_  = \new_[3615]_  ? \new_[6271]_  : \A[15] ;
  assign \new_[5318]_  = \new_[5733]_  ^ \new_[5606]_ ;
  assign \new_[5319]_  = \new_[2553]_  ? \new_[6271]_  : \A[3] ;
  assign \new_[5320]_  = \new_[2551]_  ? \new_[6271]_  : \A[6] ;
  assign \new_[5321]_  = \new_[3285]_  ? \new_[5724]_  : \A[7] ;
  assign \new_[5322]_  = \new_[2552]_  ? \new_[6271]_  : \A[5] ;
  assign \new_[5323]_  = \new_[2555]_  ? \new_[6271]_  : \A[4] ;
  assign \new_[5324]_  = \new_[3621]_  ? \new_[5724]_  : \A[14] ;
  assign \new_[5325]_  = \new_[3603]_  ? \new_[6271]_  : \A[10] ;
  assign \new_[5326]_  = \new_[6152]_  ? \new_[5680]_  : \di[6] ;
  assign \new_[5327]_  = \new_[6120]_  ? \new_[5680]_  : \di[7] ;
  assign \new_[5328]_  = \new_[2554]_  ? \new_[6271]_  : \A[2] ;
  assign \new_[5329]_  = \new_[3639]_  ? \new_[6271]_  : \A[11] ;
  assign \new_[5330]_  = \new_[5786]_  | \new_[5617]_ ;
  assign \new_[5331]_  = ~\new_[5428]_ ;
  assign \new_[5332]_  = ~\new_[5458]_  & (~\new_[5885]_  | ~\new_[6679]_ );
  assign \new_[5333]_  = ~\new_[5567]_  & ~\new_[6011]_ ;
  assign \new_[5334]_  = ~\new_[5527]_  & (~\new_[6054]_  | ~\new_[6085]_ );
  assign \new_[5335]_  = ~\new_[6995]_  | ~\new_[5116]_ ;
  assign \new_[5336]_  = ~\new_[5559]_  & ~\new_[6011]_ ;
  assign \new_[5337]_  = ~\new_[5573]_  | ~\new_[1126]_ ;
  assign \new_[5338]_  = ~\new_[6427]_  | ~\new_[5672]_  | ~\new_[6504]_ ;
  assign \new_[5339]_  = ~\new_[5816]_  | ~\new_[5823]_  | ~\new_[6492]_ ;
  assign \new_[5340]_  = ~reset_n | ~\new_[5672]_  | ~\new_[6452]_ ;
  assign \new_[5341]_  = ~\new_[5728]_  | (~\new_[5776]_  & ~\new_[6400]_ );
  assign \new_[5342]_  = (~\new_[6518]_  | ~\new_[5705]_ ) & (~\new_[1247]_  | ~\new_[7050]_ );
  assign \new_[5343]_  = (~\new_[1247]_  | ~\new_[5705]_ ) & (~\new_[1248]_  | ~\new_[7050]_ );
  assign \new_[5344]_  = ~\new_[6001]_  & ~\new_[5458]_ ;
  assign \new_[5345]_  = ~\new_[6076]_  & (~\new_[5679]_  | ~\new_[6478]_ );
  assign \new_[5346]_  = ~\new_[6648]_  | ~\new_[5459]_ ;
  assign \new_[5347]_  = ~\new_[6400]_  & ~\new_[6128]_ ;
  assign \new_[5348]_  = ~\new_[5866]_  | ~\new_[5116]_ ;
  assign \new_[5349]_  = ~\new_[7550]_  | ~\new_[5590]_  | ~\new_[6400]_ ;
  assign \new_[5350]_  = ~\new_[5996]_  | ~\new_[5884]_ ;
  assign \new_[5351]_  = ~\new_[7162]_  & ~\new_[6227]_ ;
  assign \new_[5352]_  = \new_[7231]_  & \new_[6084]_ ;
  assign \new_[5353]_  = \new_[5116]_  & \new_[6227]_ ;
  assign \new_[5354]_  = ~\new_[5860]_  & (~\new_[5895]_  | ~\new_[7201]_ );
  assign \new_[5355]_  = \new_[5696]_  ^ \new_[5812]_ ;
  assign \new_[5356]_  = ~\new_[5595]_ ;
  assign \new_[5357]_  = ~\new_[6143]_  | ~\new_[5823]_  | ~\new_[6465]_ ;
  assign \new_[5358]_  = \new_[5718]_  ^ \new_[5659]_ ;
  assign \new_[5359]_  = \new_[5569]_  & \new_[6138]_ ;
  assign \new_[5360]_  = ~\new_[5432]_ ;
  assign \new_[5361]_  = ~\new_[5454]_ ;
  assign \new_[5362]_  = \new_[6128]_  & \new_[6137]_ ;
  assign \new_[5363]_  = (~\new_[5679]_  | ~\new_[6542]_ ) & (~\new_[5861]_  | ~\new_[6515]_ );
  assign \new_[5364]_  = (~\new_[5679]_  | ~\new_[1126]_ ) & (~\new_[5861]_  | ~\new_[6542]_ );
  assign \new_[5365]_  = (~\new_[5716]_  | ~\new_[6625]_ ) & (~\new_[5784]_  | ~\new_[740]_ );
  assign \new_[5366]_  = ~\new_[5543]_ ;
  assign \new_[5367]_  = (~\new_[5726]_  | ~\new_[6952]_ ) & (~\new_[6422]_  | ~\new_[5959]_ );
  assign \new_[5368]_  = ~\new_[7170]_  | ~\new_[2002]_  | ~\new_[5779]_ ;
  assign \new_[5369]_  = \new_[5825]_  ^ \new_[5730]_ ;
  assign \new_[5370]_  = \new_[5975]_  ? \new_[5729]_  : \new_[5853]_ ;
  assign \new_[5371]_  = ~\new_[5465]_ ;
  assign \new_[5372]_  = ~\new_[5618]_  & ~\new_[5615]_ ;
  assign \new_[5373]_  = ~\new_[5608]_ ;
  assign \new_[5374]_  = ~\new_[5615]_  & (~\new_[6112]_  | ~\new_[6173]_ );
  assign \new_[5375]_  = ~\new_[5469]_ ;
  assign \new_[5376]_  = ~\new_[6083]_  | ~\new_[850]_ ;
  assign \new_[5377]_  = ~\new_[6011]_  & ~\new_[5685]_ ;
  assign \new_[5378]_  = ~\new_[5472]_ ;
  assign \new_[5379]_  = ~\new_[6457]_  & ~\new_[5949]_ ;
  assign \new_[5380]_  = ~\new_[7201]_  | ~\new_[5630]_ ;
  assign \new_[5381]_  = ~\new_[5642]_  & ~\new_[5626]_ ;
  assign \new_[5382]_  = ~\new_[5672]_  & ~\new_[6055]_ ;
  assign \new_[5383]_  = ~\new_[5701]_  & (~\new_[5781]_  | ~\new_[5904]_ );
  assign \new_[5384]_  = ~\new_[5632]_  | ~\new_[6036]_ ;
  assign \new_[5385]_  = \new_[7315]_  & \new_[5802]_ ;
  assign \new_[5386]_  = (~\new_[5928]_  | ~\new_[5924]_ ) & (~\new_[7201]_  | ~\new_[7117]_ );
  assign \new_[5387]_  = (~\new_[5793]_  & ~\new_[5879]_ ) | (~\new_[5720]_  & ~\new_[5946]_ );
  assign \new_[5388]_  = ~\new_[5649]_  & (~\new_[6030]_  | ~\new_[6565]_ );
  assign \new_[5389]_  = \new_[5636]_  & \new_[5637]_ ;
  assign \new_[5390]_  = \new_[5650]_  & \new_[5977]_ ;
  assign \new_[5391]_  = ~\new_[5608]_  | ~\new_[7201]_ ;
  assign \new_[5392]_  = ~\new_[5623]_  | ~\new_[6365]_ ;
  assign \new_[5393]_  = ~\new_[5511]_ ;
  assign \new_[5394]_  = ~\new_[5686]_  & ~\new_[6120]_ ;
  assign \new_[5395]_  = ~\new_[5627]_  | ~\new_[6084]_ ;
  assign \new_[5396]_  = ~\new_[5624]_  & (~\new_[5771]_  | ~\new_[6107]_ );
  assign \new_[5397]_  = ~\new_[5546]_ ;
  assign \new_[5398]_  = \new_[5850]_  & \new_[5663]_ ;
  assign \new_[5399]_  = ~\new_[5519]_ ;
  assign \new_[5400]_  = ~\new_[5614]_  | ~\new_[596]_ ;
  assign \new_[5401]_  = ~\new_[5753]_  | ~\new_[5804]_ ;
  assign \new_[5402]_  = ~\new_[5520]_ ;
  assign \new_[5403]_  = ~\new_[5503]_ ;
  assign \new_[5404]_  = ~\new_[5523]_ ;
  assign \new_[5405]_  = ~\new_[5660]_  & ~\new_[6284]_ ;
  assign \new_[5406]_  = ~\new_[5898]_  | ~\new_[5693]_ ;
  assign \new_[5407]_  = ~\new_[5462]_ ;
  assign \new_[5408]_  = ~\new_[5805]_  & ~\new_[5910]_ ;
  assign \new_[5409]_  = ~\new_[7163]_  & ~\new_[5629]_ ;
  assign \new_[5410]_  = \new_[5807]_  | \new_[7180]_ ;
  assign \new_[5411]_  = \new_[7008]_  & \new_[5704]_ ;
  assign \new_[5412]_  = ~\new_[5470]_ ;
  assign \new_[5413]_  = ~\new_[5710]_  | ~\new_[7201]_ ;
  assign \new_[5414]_  = \new_[5655]_  & \new_[5742]_ ;
  assign \new_[5415]_  = ~\new_[5657]_  | ~\new_[6359]_ ;
  assign \new_[5416]_  = ~\new_[5874]_  | ~\new_[5817]_  | ~\new_[5929]_  | ~\new_[5955]_ ;
  assign \new_[5417]_  = \new_[7315]_  | \new_[5607]_ ;
  assign \new_[5418]_  = ~\new_[5530]_ ;
  assign \new_[5419]_  = (~\new_[5954]_  | ~\new_[5906]_ ) & (~\new_[5934]_  | ~\new_[5787]_ );
  assign \new_[5420]_  = ~\new_[5549]_ ;
  assign \new_[5421]_  = ~\new_[7008]_  | ~\new_[7159]_ ;
  assign \new_[5422]_  = ~\di[5]  | ~\new_[6156]_ ;
  assign \new_[5423]_  = ~\di[3]  | ~\new_[6156]_ ;
  assign \new_[5424]_  = ~\di[4]  | ~\new_[6156]_ ;
  assign \new_[5425]_  = ~\new_[5909]_  | ~\new_[6452]_ ;
  assign \new_[5426]_  = ~\new_[5898]_  | ~\new_[5915]_ ;
  assign \new_[5427]_  = ~\new_[5909]_  | ~\new_[6504]_ ;
  assign \new_[5428]_  = \new_[7201]_ ;
  assign \new_[5429]_  = ~\new_[5660]_ ;
  assign \new_[5430]_  = ~\new_[5627]_  | ~\new_[5772]_ ;
  assign \new_[5431]_  = ~\new_[5987]_  | ~\new_[5929]_  | ~\new_[5748]_ ;
  assign \new_[5432]_  = \new_[5682]_  | \new_[7132]_ ;
  assign \new_[5433]_  = ~\new_[6075]_  & ~\new_[7058]_ ;
  assign \new_[5434]_  = ~\new_[5884]_  | ~\new_[5972]_  | ~\new_[6325]_  | ~\new_[5816]_ ;
  assign \new_[5435]_  = ~\new_[6003]_  | ~\new_[5901]_  | ~\new_[5801]_  | ~\new_[5968]_ ;
  assign \new_[5436]_  = (~\new_[6542]_  | ~\new_[5705]_ ) & (~\new_[1126]_  | ~\new_[7050]_ );
  assign \new_[5437]_  = (~\new_[6515]_  | ~\new_[5705]_ ) & (~\new_[6542]_  | ~\new_[7050]_ );
  assign \new_[5438]_  = \new_[5686]_  & \new_[6032]_ ;
  assign \new_[5439]_  = ~\new_[5972]_  | ~\new_[6397]_  | ~\new_[5678]_  | ~\new_[6313]_ ;
  assign \new_[5440]_  = (~\new_[6478]_  | ~\new_[5705]_ ) & (~\new_[6518]_  | ~\new_[7050]_ );
  assign \new_[5441]_  = ~\new_[7015]_  | ~\new_[7193]_ ;
  assign \new_[5442]_  = \new_[5692]_  | \new_[6400]_ ;
  assign \new_[5443]_  = ~\new_[5927]_  & ~\new_[5889]_ ;
  assign \new_[5444]_  = ~\new_[5991]_  | ~\new_[596]_ ;
  assign \new_[5445]_  = ~\new_[5692]_  & ~\new_[6031]_ ;
  assign \new_[5446]_  = ~\new_[5772]_  & ~\new_[6113]_ ;
  assign \new_[5447]_  = ~\new_[7155]_ ;
  assign \new_[5448]_  = ~\new_[5463]_ ;
  assign \new_[5449]_  = ~\new_[5909]_  | ~\new_[6442]_ ;
  assign \new_[5450]_  = ~\new_[6156]_  | ~\new_[6523]_  | ~\new_[3321]_  | ~\new_[6554]_ ;
  assign \new_[5451]_  = ~\new_[6394]_  & ~\new_[6107]_ ;
  assign \new_[5452]_  = ~\new_[6046]_  & ~\new_[7377]_ ;
  assign \new_[5453]_  = ~\new_[5779]_  | ~\new_[5885]_  | ~\new_[6548]_ ;
  assign \new_[5454]_  = ~\new_[5714]_  & ~\new_[5702]_ ;
  assign \new_[5455]_  = ~\new_[5598]_ ;
  assign \new_[5456]_  = \new_[5830]_  | \new_[5889]_ ;
  assign \new_[5457]_  = ~\new_[5971]_  | (~\new_[6043]_  & ~\new_[6083]_ );
  assign \new_[5458]_  = ~\new_[6534]_  | ~\new_[6440]_  | ~\new_[6429]_ ;
  assign \new_[5459]_  = ~\new_[5877]_ ;
  assign \new_[5460]_  = \new_[5812]_  ^ \new_[5811]_ ;
  assign \new_[5461]_  = ~\new_[5752]_  & ~\new_[5731]_ ;
  assign \new_[5462]_  = ~\new_[7121]_  | ~\new_[5927]_ ;
  assign \new_[5463]_  = \new_[5772]_  & \new_[6137]_ ;
  assign \new_[5464]_  = ~\new_[5730]_  | ~\new_[5825]_ ;
  assign \new_[5465]_  = (~\new_[5873]_  | ~\new_[1324]_ ) & (~\new_[1126]_  | ~\new_[6318]_ );
  assign \new_[5466]_  = ~\new_[5694]_ ;
  assign \new_[5467]_  = \new_[6515]_  ^ \new_[6083]_ ;
  assign \new_[5468]_  = ~\new_[7005]_  & ~\new_[5984]_ ;
  assign \new_[5469]_  = ~\new_[6800]_  | ~\new_[5926]_ ;
  assign \new_[5470]_  = ~\new_[7201]_  | ~\new_[5958]_ ;
  assign \new_[5471]_  = \new_[5719]_  | \new_[6523]_ ;
  assign \new_[5472]_  = ~\new_[7549]_  | ~\new_[6272]_ ;
  assign \new_[5473]_  = ~\new_[5705]_ ;
  assign \new_[5474]_  = \new_[1394]_  ^ \new_[5829]_ ;
  assign \new_[5475]_  = ~\new_[5726]_  | ~\new_[6953]_ ;
  assign \new_[5476]_  = \new_[5753]_  & \new_[7006]_ ;
  assign \new_[5477]_  = (~\new_[7223]_  | ~\new_[6047]_ ) & (~\new_[848]_  | ~\new_[6264]_ );
  assign \new_[5478]_  = (~\new_[5837]_  | ~\new_[6215]_ ) & (~\new_[792]_  | ~\new_[6264]_ );
  assign \new_[5479]_  = (~\new_[5833]_  | ~\new_[6384]_ ) & (~\new_[794]_  | ~\new_[6264]_ );
  assign \new_[5480]_  = (~\new_[5841]_  | ~\new_[6384]_ ) & (~\new_[742]_  | ~\new_[6264]_ );
  assign \new_[5481]_  = (~\new_[5832]_  | ~\new_[6215]_ ) & (~\new_[766]_  | ~\new_[6264]_ );
  assign \new_[5482]_  = (~\new_[5839]_  | ~\new_[6215]_ ) & (~\new_[764]_  | ~\new_[6264]_ );
  assign \new_[5483]_  = (~\new_[5834]_  | ~\new_[6215]_ ) & (~\new_[757]_  | ~\new_[6264]_ );
  assign \new_[5484]_  = (~\new_[5836]_  | ~\new_[6047]_ ) & (~\new_[853]_  | ~\new_[6264]_ );
  assign \new_[5485]_  = (~\new_[5840]_  | ~\new_[6047]_ ) & (~\new_[851]_  | ~\new_[6264]_ );
  assign \new_[5486]_  = ~\new_[6465]_  | ~\new_[6193]_  | ~\new_[5823]_  | ~\new_[6312]_ ;
  assign \new_[5487]_  = \new_[7339]_  & \new_[7440]_ ;
  assign \new_[5488]_  = \new_[7188]_  & \new_[7440]_ ;
  assign \new_[5489]_  = \new_[5832]_  & \new_[7440]_ ;
  assign \new_[5490]_  = \new_[5833]_  & \new_[7440]_ ;
  assign \new_[5491]_  = \new_[7223]_  & \new_[7440]_ ;
  assign \new_[5492]_  = \new_[5835]_  & \new_[7440]_ ;
  assign \new_[5493]_  = \new_[5834]_  & \new_[7440]_ ;
  assign \new_[5494]_  = \new_[6940]_  & \new_[7440]_ ;
  assign \new_[5495]_  = \new_[5841]_  & \new_[7440]_ ;
  assign \new_[5496]_  = \new_[5839]_  & \new_[7440]_ ;
  assign \new_[5497]_  = \new_[5837]_  & \new_[7440]_ ;
  assign \new_[5498]_  = \new_[5822]_  & \new_[7440]_ ;
  assign \new_[5499]_  = \new_[5838]_  & \new_[7440]_ ;
  assign \new_[5500]_  = ~\new_[7175]_  | ~\new_[5926]_ ;
  assign \new_[5501]_  = \new_[5840]_  & \new_[7440]_ ;
  assign \new_[5502]_  = \new_[5836]_  & \new_[7440]_ ;
  assign \new_[5503]_  = ~\new_[6315]_  | ~\new_[6961]_ ;
  assign \new_[5504]_  = ~\new_[7210]_  & (~\new_[5946]_  | ~\new_[5879]_ );
  assign \new_[5505]_  = ~\new_[5623]_ ;
  assign \new_[5506]_  = \new_[5904]_  ^ \new_[5819]_ ;
  assign \new_[5507]_  = \new_[5896]_  | \new_[6004]_ ;
  assign \new_[5508]_  = \new_[5855]_  | \new_[5723]_ ;
  assign \new_[5509]_  = ~\new_[6175]_  | ~\new_[5859]_  | ~\new_[5880]_ ;
  assign \new_[5510]_  = \new_[6926]_  & \new_[7440]_ ;
  assign \new_[5511]_  = \new_[7011]_ ;
  assign \new_[5512]_  = \new_[5843]_  & \new_[5715]_ ;
  assign \new_[5513]_  = ~\new_[5717]_  | ~\new_[6296]_ ;
  assign \new_[5514]_  = ~\new_[5666]_ ;
  assign \new_[5515]_  = ~\new_[5929]_  | ~\new_[5748]_ ;
  assign \new_[5516]_  = ~\new_[5848]_  | ~\new_[5795]_ ;
  assign \new_[5517]_  = \new_[5717]_  & \new_[6439]_ ;
  assign \new_[5518]_  = ~\new_[5634]_ ;
  assign \new_[5519]_  = ~\new_[7200]_  & ~\new_[6234]_ ;
  assign \new_[5520]_  = ~\new_[5744]_  | ~\new_[5792]_ ;
  assign \new_[5521]_  = \new_[5911]_  & \new_[5758]_ ;
  assign \new_[5522]_  = \new_[7379]_  | \new_[7315]_ ;
  assign \new_[5523]_  = ~\new_[7379]_  & ~\new_[5759]_ ;
  assign \new_[5524]_  = ~\new_[7121]_  & ~\new_[5924]_ ;
  assign \new_[5525]_  = ~\new_[5882]_  | ~\new_[5768]_ ;
  assign \new_[5526]_  = ~\new_[5882]_  | ~\new_[5792]_ ;
  assign \new_[5527]_  = \new_[6962]_  & \new_[6071]_ ;
  assign \new_[5528]_  = ~\new_[7005]_  & ~\new_[5894]_ ;
  assign \new_[5529]_  = ~\new_[5755]_  | ~\new_[5968]_ ;
  assign \new_[5530]_  = ~\new_[5650]_ ;
  assign \new_[5531]_  = ~\new_[5725]_  | ~\new_[5804]_ ;
  assign \new_[5532]_  = ~\new_[6085]_  | ~\new_[7121]_ ;
  assign \new_[5533]_  = ~\new_[6076]_  & (~\new_[5878]_  | ~\new_[6515]_ );
  assign \new_[5534]_  = \new_[5862]_  | \new_[7121]_ ;
  assign \new_[5535]_  = \new_[2633]_  ^ \new_[6156]_ ;
  assign \new_[5536]_  = \new_[5786]_  | \new_[5897]_ ;
  assign \new_[5537]_  = ~\di[2]  | ~\new_[6156]_ ;
  assign \new_[5538]_  = ~\new_[6009]_  | ~\new_[6067]_  | ~\new_[5887]_  | ~\new_[5996]_ ;
  assign \new_[5539]_  = ~\di[6]  | ~\new_[6156]_ ;
  assign \new_[5540]_  = ~\di[7]  | ~\new_[6156]_ ;
  assign \new_[5541]_  = ~\new_[5624]_ ;
  assign \new_[5542]_  = \new_[5766]_  | \new_[5933]_ ;
  assign \new_[5543]_  = \new_[5924]_  & \new_[5927]_ ;
  assign \new_[5544]_  = ~\new_[5601]_  & ~\new_[7116]_ ;
  assign \new_[5545]_  = ~\new_[5631]_ ;
  assign \new_[5546]_  = \new_[7129]_  & \new_[6458]_ ;
  assign \new_[5547]_  = ~\new_[7006]_  | ~\new_[5988]_  | ~\new_[5868]_ ;
  assign \new_[5548]_  = \new_[5796]_  & \new_[5721]_ ;
  assign \new_[5549]_  = ~\new_[5896]_  & ~\new_[6071]_ ;
  assign \new_[5550]_  = ~\new_[1624]_  | ~\new_[5925]_  | ~\new_[5877]_ ;
  assign \new_[5551]_  = ~\new_[5766]_  & ~\new_[6060]_ ;
  assign \new_[5552]_  = ~\new_[5911]_  | ~\new_[6016]_ ;
  assign \new_[5553]_  = ~\new_[5937]_  & ~\new_[6050]_ ;
  assign \new_[5554]_  = ~\new_[5954]_  & ~\new_[5794]_ ;
  assign \new_[5555]_  = ~\new_[5967]_  & ~\new_[5966]_ ;
  assign \new_[5556]_  = \new_[5988]_  & \new_[5883]_ ;
  assign \new_[5557]_  = ~\new_[7562]_  | ~\new_[7047]_ ;
  assign \new_[5558]_  = ~\new_[5612]_ ;
  assign \new_[5559]_  = ~\new_[2005]_  | ~\new_[5773]_ ;
  assign \new_[5560]_  = ~\new_[5693]_ ;
  assign \new_[5561]_  = ~\new_[5703]_  & (~\new_[6114]_  | ~\new_[6442]_ );
  assign \new_[5562]_  = \new_[5979]_  | \new_[595]_ ;
  assign \new_[5563]_  = (~\new_[5838]_  | ~\new_[6047]_ ) & (~\new_[755]_  | ~\new_[6264]_ );
  assign \new_[5564]_  = (~\new_[5873]_  | ~\new_[6515]_ ) & (~\new_[6014]_  | ~\new_[6520]_ );
  assign \new_[5565]_  = ~\new_[7175]_  | ~\new_[5824]_ ;
  assign \new_[5566]_  = ~\new_[5669]_ ;
  assign \new_[5567]_  = ~\new_[2006]_  | ~\new_[5773]_ ;
  assign \new_[5568]_  = ~\new_[5685]_ ;
  assign \new_[5569]_  = ~\new_[1248]_  | ~\new_[5705]_ ;
  assign \new_[5570]_  = ~\new_[5640]_ ;
  assign \new_[5571]_  = ~\new_[5775]_  & ~\new_[6084]_ ;
  assign \new_[5572]_  = ~\new_[1624]_  & ~\new_[5708]_ ;
  assign \new_[5573]_  = \new_[6268]_  | \new_[5705]_ ;
  assign \new_[5574]_  = ~\new_[5636]_ ;
  assign \new_[5575]_  = ~\new_[5741]_  | ~\new_[7159]_ ;
  assign \new_[5576]_  = ~\new_[5938]_  | ~\new_[5758]_ ;
  assign \new_[5577]_  = ~\new_[5744]_  | ~\new_[5768]_ ;
  assign \new_[5578]_  = ~\new_[6325]_  & ~\new_[6128]_ ;
  assign \new_[5579]_  = \new_[6528]_  & \new_[5779]_ ;
  assign \new_[5580]_  = ~\new_[6284]_  | (~\new_[5954]_  & ~\new_[6002]_ );
  assign \new_[5581]_  = ~\new_[6049]_  & ~\new_[6120]_ ;
  assign \new_[5582]_  = \new_[6039]_  & \new_[6067]_ ;
  assign \new_[5583]_  = ~\new_[5886]_  | ~\new_[5749]_ ;
  assign \new_[5584]_  = ~\new_[6120]_  & ~\new_[6227]_ ;
  assign \new_[5585]_  = ~\di[0]  | ~\new_[6156]_ ;
  assign \new_[5586]_  = (~\new_[5822]_  | ~\new_[6215]_ ) & (~\new_[793]_  | ~\new_[6264]_ );
  assign \new_[5587]_  = ~\new_[5722]_  | (~\new_[1811]_  & ~\new_[6460]_ );
  assign \new_[5588]_  = ~\new_[5605]_ ;
  assign \new_[5589]_  = ~\di[1]  | ~\new_[6156]_ ;
  assign \new_[5590]_  = ~\new_[5692]_ ;
  assign \new_[5591]_  = \new_[6940]_  ? \new_[6264]_  : \new_[684]_ ;
  assign \new_[5592]_  = ~\new_[5629]_ ;
  assign \new_[5593]_  = (~\new_[7339]_  | ~\new_[6047]_ ) & (~\new_[852]_  | ~\new_[6264]_ );
  assign \new_[5594]_  = \new_[6580]_  ^ \new_[5900]_ ;
  assign \new_[5595]_  = ~\new_[6107]_ ;
  assign \new_[5596]_  = ~\new_[7059]_  | ~\new_[5947]_  | ~\new_[5898]_  | ~\new_[6175]_ ;
  assign \new_[5597]_  = ~\new_[5775]_  & ~\new_[6959]_ ;
  assign \new_[5598]_  = ~\new_[7017]_ ;
  assign \new_[5599]_  = \new_[5748]_  & \new_[5874]_ ;
  assign \new_[5600]_  = \new_[1379]_  ^ \new_[5803]_ ;
  assign \new_[5601]_  = ~\new_[5901]_ ;
  assign \new_[5602]_  = ~\new_[5895]_ ;
  assign \new_[5603]_  = \new_[5707]_  & \new_[5812]_ ;
  assign \new_[5604]_  = \new_[1453]_  ^ \new_[5917]_ ;
  assign \new_[5605]_  = ~\new_[6632]_  | ~\new_[6637]_  | ~\new_[6571]_ ;
  assign \new_[5606]_  = \new_[5945]_  ^ \new_[5943]_ ;
  assign \new_[5607]_  = ~\new_[5796]_ ;
  assign \new_[5608]_  = ~\new_[5801]_ ;
  assign \new_[5609]_  = \new_[6084]_  & \new_[6137]_ ;
  assign \new_[5610]_  = ~\new_[5714]_ ;
  assign \new_[5611]_  = ~\new_[5722]_ ;
  assign \new_[5612]_  = ~\new_[6050]_  & ~\new_[7158]_ ;
  assign \new_[5613]_  = ~\new_[6072]_  | (~\new_[5963]_  & ~\new_[6280]_ );
  assign \new_[5614]_  = ~\new_[5847]_  | ~\new_[6055]_ ;
  assign \new_[5615]_  = \new_[6083]_  & \new_[6518]_ ;
  assign \new_[5616]_  = ~\new_[6571]_  | ~halt_n | ~\new_[5944]_ ;
  assign \new_[5617]_  = ~\new_[5703]_ ;
  assign \new_[5618]_  = ~\new_[6083]_  & (~\new_[6436]_  | ~\new_[6451]_ );
  assign \new_[5619]_  = ~\new_[5729]_ ;
  assign \new_[5620]_  = ~\new_[5723]_ ;
  assign \new_[5621]_  = ~\new_[5743]_ ;
  assign \new_[5622]_  = \new_[6055]_  & \new_[6504]_ ;
  assign \new_[5623]_  = ~\new_[5734]_ ;
  assign \new_[5624]_  = ~\new_[7159]_  | ~\new_[5949]_ ;
  assign \new_[5625]_  = \new_[6055]_  & \new_[6452]_ ;
  assign \new_[5626]_  = ~\new_[5923]_  | ~\new_[5801]_ ;
  assign \new_[5627]_  = ~\new_[5741]_ ;
  assign \new_[5628]_  = \new_[5862]_  | \new_[7070]_ ;
  assign \new_[5629]_  = ~\new_[6128]_  | ~\new_[5927]_ ;
  assign \new_[5630]_  = ~\new_[6004]_  & ~\new_[5889]_ ;
  assign \new_[5631]_  = \new_[5740]_ ;
  assign \new_[5632]_  = ~\new_[5904]_  | ~\new_[5999]_ ;
  assign \new_[5633]_  = ~\new_[5896]_  & ~\new_[5928]_ ;
  assign \new_[5634]_  = \new_[5807]_  & \new_[6133]_ ;
  assign \new_[5635]_  = ~\new_[5955]_  | ~\new_[5817]_ ;
  assign \new_[5636]_  = ~\new_[5892]_  | ~\new_[6140]_ ;
  assign \new_[5637]_  = ~\new_[7015]_  | ~\new_[6140]_ ;
  assign \new_[5638]_  = ~\new_[7024]_ ;
  assign \new_[5639]_  = ~\new_[7315]_  & ~\new_[5961]_ ;
  assign \new_[5640]_  = ~\new_[5731]_ ;
  assign \new_[5641]_  = ~\new_[5962]_ ;
  assign \new_[5642]_  = \new_[5854]_  | \new_[7056]_ ;
  assign \new_[5643]_  = ~\new_[5735]_ ;
  assign \new_[5644]_  = ~\new_[5848]_  | ~\new_[7157]_ ;
  assign \new_[5645]_  = ~\new_[5851]_  | ~\new_[5890]_ ;
  assign \new_[5646]_  = ~\new_[5891]_  | ~\new_[7163]_ ;
  assign \new_[5647]_  = ~\new_[5948]_  | ~\new_[5931]_  | ~\new_[5987]_ ;
  assign \new_[5648]_  = ~\new_[5805]_  | ~\new_[6305]_ ;
  assign \new_[5649]_  = ~\new_[5810]_  | ~\new_[5846]_ ;
  assign \new_[5650]_  = ~\new_[6317]_  | ~\new_[6044]_  | ~\new_[5908]_ ;
  assign \new_[5651]_  = (~\new_[7248]_  | ~\new_[6085]_ ) & (~\new_[6054]_  | ~\new_[7193]_ );
  assign \new_[5652]_  = \new_[6475]_  ? \new_[6271]_  : \new_[2661]_ ;
  assign \new_[5653]_  = \new_[5808]_  | \new_[6380]_ ;
  assign \new_[5654]_  = \new_[6055]_  & \new_[6442]_ ;
  assign \new_[5655]_  = \new_[5902]_  & \new_[6168]_ ;
  assign \new_[5656]_  = \new_[5864]_  | \new_[5897]_ ;
  assign \new_[5657]_  = ~\new_[5720]_ ;
  assign \new_[5658]_  = ~\new_[5809]_  | ~\new_[7193]_ ;
  assign \new_[5659]_  = ~\new_[5811]_  | ~\new_[5812]_ ;
  assign \new_[5660]_  = \new_[5888]_  | \new_[6969]_ ;
  assign \new_[5661]_  = ~\new_[5753]_ ;
  assign \new_[5662]_  = ~\new_[5867]_  & ~\new_[5953]_ ;
  assign \new_[5663]_  = ~\new_[5895]_  | ~\new_[6234]_ ;
  assign \new_[5664]_  = ~\new_[5952]_  & ~\new_[5934]_ ;
  assign \new_[5665]_  = ~\new_[5827]_  | ~\new_[1248]_ ;
  assign \new_[5666]_  = ~\new_[7349]_ ;
  assign \new_[5667]_  = ~\new_[6521]_  | (~\new_[5930]_  & ~\new_[6037]_ );
  assign \new_[5668]_  = ~\new_[5950]_  | ~\new_[6986]_  | ~\new_[6251]_ ;
  assign \new_[5669]_  = ~\new_[5789]_ ;
  assign \new_[5670]_  = ~\new_[5991]_  | ~\new_[597]_ ;
  assign \new_[5671]_  = ~\new_[5991]_  | ~\new_[6452]_ ;
  assign \new_[5672]_  = ~\new_[5847]_ ;
  assign \new_[5673]_  = ~\new_[5860]_ ;
  assign \new_[5674]_  = ~\new_[5765]_ ;
  assign \new_[5675]_  = ~\new_[5823]_  | ~\new_[6167]_ ;
  assign \new_[5676]_  = ~\new_[6041]_  | ~\new_[6216]_ ;
  assign \new_[5677]_  = ~\new_[5991]_  | ~\new_[6504]_ ;
  assign \new_[5678]_  = ~\new_[5885]_  & ~\new_[6484]_ ;
  assign \new_[5679]_  = \new_[5873]_  | \new_[6819]_ ;
  assign \new_[5680]_  = ~\new_[6216]_  & ~\new_[5995]_ ;
  assign \new_[5681]_  = ~\new_[6663]_  & ~\new_[5991]_ ;
  assign \new_[5682]_  = ~\new_[6084]_  | ~\new_[6104]_  | ~\new_[6171]_ ;
  assign \new_[5683]_  = ~\new_[6416]_  & ~\new_[6120]_ ;
  assign \new_[5684]_  = \new_[5823]_  & \new_[6039]_ ;
  assign \new_[5685]_  = \new_[5885]_  | \new_[6679]_ ;
  assign \new_[5686]_  = ~\new_[6325]_  | ~\new_[5884]_ ;
  assign \new_[5687]_  = \new_[5881]_  & \new_[1810]_ ;
  assign \new_[5688]_  = ~\new_[5927]_ ;
  assign \new_[5689]_  = ~\new_[5800]_  | ~\new_[6400]_ ;
  assign \new_[5690]_  = \new_[5903]_  & \new_[7159]_ ;
  assign \new_[5691]_  = ~\new_[5991]_  | ~\new_[6442]_ ;
  assign \new_[5692]_  = ~\new_[6128]_  | ~\new_[5972]_ ;
  assign \new_[5693]_  = ~\new_[5862]_  | ~\new_[6284]_ ;
  assign \new_[5694]_  = \new_[5814]_  & \new_[5851]_ ;
  assign \new_[5695]_  = ~\new_[5896]_ ;
  assign \new_[5696]_  = ~\new_[6520]_  & (~\new_[5989]_  | ~\new_[1324]_ );
  assign \new_[5697]_  = ~\new_[5793]_ ;
  assign \new_[5698]_  = ~\new_[6085]_  | ~\new_[5895]_ ;
  assign \new_[5699]_  = ~\new_[5827]_  | ~\new_[1324]_ ;
  assign \new_[5700]_  = ~\new_[6075]_  | ~\new_[5927]_ ;
  assign \new_[5701]_  = (~\new_[5978]_  | ~\new_[5953]_ ) & (~\new_[6036]_  | ~\new_[5978]_ );
  assign \new_[5702]_  = ~\new_[6073]_  | (~\new_[5976]_  & ~\new_[6280]_ );
  assign \new_[5703]_  = ~\new_[5973]_  | ~\new_[7324]_ ;
  assign \new_[5704]_  = ~\new_[5871]_ ;
  assign \new_[5705]_  = \new_[7557]_  & \new_[6128]_ ;
  assign \new_[5706]_  = ~\new_[6227]_  | ~\new_[6272]_ ;
  assign \new_[5707]_  = ~\new_[5971]_  | (~\new_[6089]_  & ~\new_[6083]_ );
  assign \new_[5708]_  = ~\new_[5982]_  | ~\new_[1810]_ ;
  assign \new_[5709]_  = (~\new_[6268]_  | ~\new_[1247]_ ) & (~\new_[1248]_  | ~\new_[6782]_ );
  assign \new_[5710]_  = ~\new_[5893]_ ;
  assign \new_[5711]_  = (~\new_[6268]_  | ~\new_[6478]_ ) & (~\new_[6518]_  | ~\new_[6782]_ );
  assign \new_[5712]_  = ~\new_[5898]_ ;
  assign \new_[5713]_  = ~\new_[5882]_ ;
  assign \new_[5714]_  = ~\new_[6122]_  | (~\new_[6059]_  & ~\new_[6280]_ );
  assign \new_[5715]_  = \new_[5234]_  | \new_[5968]_ ;
  assign \new_[5716]_  = ~\new_[5920]_  | (~\new_[6012]_  & ~\new_[6083]_ );
  assign \new_[5717]_  = ~\new_[7559]_ ;
  assign \new_[5718]_  = ~\new_[6072]_  | (~\new_[6021]_  & ~\new_[6083]_ );
  assign \new_[5719]_  = ~\new_[5844]_ ;
  assign \new_[5720]_  = ~\new_[6054]_  & ~\new_[5919]_ ;
  assign \new_[5721]_  = ~\new_[5974]_  | ~\new_[6228]_ ;
  assign \new_[5722]_  = ~\new_[1811]_  | ~\new_[6460]_ ;
  assign \new_[5723]_  = ~\new_[7210]_  & ~\new_[6309]_ ;
  assign \new_[5724]_  = ~\new_[6156]_ ;
  assign \new_[5725]_  = ~\new_[5984]_  & ~\new_[5937]_ ;
  assign \new_[5726]_  = \new_[6068]_  ^ \new_[6027]_ ;
  assign \new_[5727]_  = ~\new_[5824]_ ;
  assign \new_[5728]_  = \new_[6065]_  | \new_[6227]_ ;
  assign \new_[5729]_  = ~\new_[5939]_  | ~\new_[6212]_ ;
  assign \new_[5730]_  = \new_[5993]_  ? \new_[5998]_  : \new_[6081]_ ;
  assign \new_[5731]_  = ~\new_[7118]_  & ~\new_[6078]_ ;
  assign \new_[5732]_  = ~\new_[1248]_  | ~\new_[5930]_  | ~\new_[2002]_ ;
  assign \new_[5733]_  = \new_[6024]_  ^ \new_[6025]_ ;
  assign \new_[5734]_  = \new_[7200]_  & \new_[7134]_ ;
  assign \new_[5735]_  = ~\new_[6029]_  | ~\new_[5922]_ ;
  assign \new_[5736]_  = ~\new_[6085]_  | ~\new_[5924]_ ;
  assign \new_[5737]_  = ~\new_[6542]_  | ~\new_[5930]_  | ~\new_[2005]_ ;
  assign \new_[5738]_  = ~\new_[1126]_  | ~\new_[5930]_  | ~\new_[2006]_ ;
  assign \new_[5739]_  = ~\new_[7157]_ ;
  assign \new_[5740]_  = ~\new_[5942]_  | ~\new_[6205]_ ;
  assign \new_[5741]_  = ~\new_[6152]_  | ~\new_[7166]_  | ~\new_[7160]_ ;
  assign \new_[5742]_  = ~\new_[5934]_  & ~\new_[5954]_ ;
  assign \new_[5743]_  = ~\new_[5988]_  | ~\new_[6982]_ ;
  assign \new_[5744]_  = ~\new_[5845]_ ;
  assign \new_[5745]_  = ~\new_[6478]_  | ~\new_[5930]_  | ~\new_[6528]_ ;
  assign \new_[5746]_  = ~\new_[6156]_ ;
  assign \new_[5747]_  = ~\new_[6515]_  | ~\new_[5930]_  | ~\new_[6548]_ ;
  assign \new_[5748]_  = ~\new_[6916]_  | ~\new_[6465]_ ;
  assign \new_[5749]_  = ~\new_[5954]_  | ~\new_[6359]_ ;
  assign \new_[5750]_  = ~\new_[6518]_  | ~\new_[5930]_  | ~\new_[2007]_ ;
  assign \new_[5751]_  = ~\new_[5880]_ ;
  assign \new_[5752]_  = ~\new_[5931]_  | ~\new_[5929]_ ;
  assign \new_[5753]_  = ~\new_[6281]_  | ~\new_[6891]_  | ~\new_[6010]_ ;
  assign \new_[5754]_  = ~\new_[5124]_  & (~\new_[6017]_  | ~\new_[6619]_ );
  assign \new_[5755]_  = ~\new_[7116]_  & ~\new_[5958]_ ;
  assign \new_[5756]_  = ~\new_[5933]_  & ~\new_[7070]_ ;
  assign \new_[5757]_  = ~\new_[5967]_  & ~\new_[5970]_ ;
  assign \new_[5758]_  = ~\new_[7297]_  | ~\new_[6397]_  | ~\new_[5960]_  | ~\new_[7318]_ ;
  assign \new_[5759]_  = ~\new_[5869]_ ;
  assign \new_[5760]_  = ~\new_[5928]_ ;
  assign \new_[5761]_  = (~\new_[6014]_  | ~\new_[1126]_ ) & (~\new_[1324]_  | ~\new_[6782]_ );
  assign \new_[5762]_  = (~\new_[6268]_  | ~\new_[6542]_ ) & (~\new_[1126]_  | ~\new_[6782]_ );
  assign \new_[5763]_  = (~\new_[6268]_  | ~\new_[6518]_ ) & (~\new_[1247]_  | ~\new_[6782]_ );
  assign \new_[5764]_  = ~\new_[5958]_  | ~\new_[7193]_ ;
  assign \new_[5765]_  = ~\new_[5934]_ ;
  assign \new_[5766]_  = ~\new_[5968]_ ;
  assign \new_[5767]_  = ~\new_[5859]_ ;
  assign \new_[5768]_  = ~\new_[5956]_  | ~\new_[6152]_ ;
  assign \new_[5769]_  = ~\new_[5805]_ ;
  assign \new_[5770]_  = ~\new_[6394]_  | ~\new_[6400]_ ;
  assign \new_[5771]_  = ~\new_[5804]_ ;
  assign \new_[5772]_  = ~\new_[5884]_ ;
  assign \new_[5773]_  = ~\new_[5816]_ ;
  assign \new_[5774]_  = (~\new_[6268]_  | ~\new_[6515]_ ) & (~\new_[6542]_  | ~\new_[6782]_ );
  assign \new_[5775]_  = ~\new_[6989]_  | ~\new_[6120]_ ;
  assign \new_[5776]_  = ~\new_[6067]_  | ~\new_[7253]_ ;
  assign \new_[5777]_  = ~\new_[5931]_  | ~\new_[5987]_ ;
  assign \new_[5778]_  = ~\new_[5807]_ ;
  assign \new_[5779]_  = \new_[6351]_  & \new_[5982]_ ;
  assign \new_[5780]_  = ~\new_[6113]_  | ~\new_[6272]_ ;
  assign \new_[5781]_  = ~\new_[5957]_  & ~\new_[5953]_ ;
  assign \new_[5782]_  = ~\new_[5872]_ ;
  assign \new_[5783]_  = \new_[6953]_  | \new_[6952]_ ;
  assign \new_[5784]_  = ~\new_[5920]_  | (~\new_[6098]_  & ~\new_[6083]_ );
  assign \new_[5785]_  = \new_[1104]_  ^ \new_[6057]_ ;
  assign \new_[5786]_  = ~\new_[5914]_  & ~\new_[7169]_ ;
  assign \new_[5787]_  = ~\new_[5889]_ ;
  assign \new_[5788]_  = ~\new_[5954]_  | ~\new_[6405]_ ;
  assign \new_[5789]_  = \new_[5941]_  & \new_[6093]_ ;
  assign \new_[5790]_  = \new_[6061]_  | \new_[5942]_ ;
  assign \new_[5791]_  = \new_[5936]_  | \new_[5949]_ ;
  assign \new_[5792]_  = ~\new_[5980]_  | ~\new_[6152]_ ;
  assign \new_[5793]_  = ~\new_[5892]_ ;
  assign \new_[5794]_  = ~\new_[5902]_ ;
  assign \new_[5795]_  = ~\new_[5924]_  & ~\new_[5958]_ ;
  assign \new_[5796]_  = ~\new_[6009]_  | ~\new_[5960]_  | ~\new_[6125]_ ;
  assign \new_[5797]_  = ~\new_[1247]_  | ~\new_[5930]_  | ~\new_[2003]_ ;
  assign \new_[5798]_  = \new_[6062]_  | \new_[7325]_ ;
  assign \new_[5799]_  = ~\new_[5911]_ ;
  assign \new_[5800]_  = ~\new_[7550]_  & ~\new_[6495]_ ;
  assign \new_[5801]_  = ~\new_[6450]_  | ~\new_[7551]_  | ~\new_[7166]_  | ~\new_[7215]_ ;
  assign \new_[5802]_  = ~\new_[5906]_ ;
  assign \new_[5803]_  = ~\new_[1308]_  | ~\new_[1453]_  | ~\new_[6005]_  | ~\new_[6530]_ ;
  assign \new_[5804]_  = ~\new_[5990]_  | ~\new_[6010]_ ;
  assign \new_[5805]_  = \new_[5921]_ ;
  assign \new_[5806]_  = \new_[1610]_  ^ \new_[6074]_ ;
  assign \new_[5807]_  = ~\new_[7176]_ ;
  assign \new_[5808]_  = \new_[6045]_  | \new_[6094]_ ;
  assign \new_[5809]_  = ~\new_[5915]_ ;
  assign \new_[5810]_  = ~\new_[6087]_  | ~\new_[6029]_ ;
  assign \new_[5811]_  = ~\new_[6073]_  | (~\new_[6082]_  & ~\new_[6280]_ );
  assign \new_[5812]_  = ~\new_[6122]_  | (~\new_[6095]_  & ~\new_[6280]_ );
  assign \new_[5813]_  = ~\new_[5997]_  & ~\new_[6236]_ ;
  assign \new_[5814]_  = ~\new_[6121]_  | ~\new_[6228]_  | ~\new_[6096]_ ;
  assign \new_[5815]_  = ~\new_[6037]_  | (~\new_[6528]_  & ~\new_[1125]_ );
  assign \new_[5816]_  = \new_[6039]_  & \new_[6397]_ ;
  assign \new_[5817]_  = ~\new_[6053]_  | ~\new_[6109]_ ;
  assign \new_[5818]_  = ~\new_[6173]_  | ~\new_[1248]_  | ~\new_[6134]_  | ~\new_[1324]_ ;
  assign \new_[5819]_  = ~\new_[6036]_  | ~\new_[5999]_ ;
  assign \new_[5820]_  = ~\new_[6026]_  & ~\new_[6030]_ ;
  assign \new_[5821]_  = ~\new_[5930]_ ;
  assign \new_[5822]_  = ~\new_[6183]_  | ~\new_[6172]_  | ~\new_[6191]_  | ~\new_[6270]_ ;
  assign \new_[5823]_  = ~\new_[6120]_  & ~\new_[7298]_ ;
  assign \new_[5824]_  = ~\new_[7047]_  | ~\new_[7064]_ ;
  assign \new_[5825]_  = \new_[6027]_  & \new_[6068]_ ;
  assign \new_[5826]_  = ~\new_[5937]_ ;
  assign \new_[5827]_  = \new_[6811]_  | \new_[6014]_ ;
  assign \new_[5828]_  = ~\new_[6037]_  | (~\new_[2006]_  & ~\new_[1126]_ );
  assign \new_[5829]_  = ~\new_[1379]_  | ~\new_[1545]_  | ~\new_[6028]_  | ~\new_[1453]_ ;
  assign \new_[5830]_  = \new_[6048]_  | \new_[6405]_ ;
  assign \new_[5831]_  = ~\new_[5970]_ ;
  assign \new_[5832]_  = ~\new_[6146]_  | ~\new_[6260]_  | ~\new_[6182]_  | ~\new_[6184]_ ;
  assign \new_[5833]_  = ~\new_[6185]_  | ~\new_[6259]_  | ~\new_[6200]_  | ~\new_[6159]_ ;
  assign \new_[5834]_  = ~\new_[6187]_  | ~\new_[6273]_  | ~\new_[6235]_  | ~\new_[6241]_ ;
  assign \new_[5835]_  = ~\new_[6199]_  | ~\new_[6308]_  | ~\new_[6197]_  | ~\new_[6221]_ ;
  assign \new_[5836]_  = ~\new_[6195]_  | ~\new_[6288]_  | ~\new_[6214]_  | ~\new_[6208]_ ;
  assign \new_[5837]_  = ~\new_[6178]_  | ~\new_[6276]_  | ~\new_[6192]_  | ~\new_[6186]_ ;
  assign \new_[5838]_  = ~\new_[6179]_  | ~\new_[6303]_  | ~\new_[6176]_  | ~\new_[6238]_ ;
  assign \new_[5839]_  = ~\new_[6151]_  | ~\new_[6311]_  | ~\new_[6174]_  | ~\new_[6237]_ ;
  assign \new_[5840]_  = ~\new_[6201]_  | ~\new_[6289]_  | ~\new_[6157]_  | ~\new_[6155]_ ;
  assign \new_[5841]_  = ~\new_[6194]_  | ~\new_[6319]_  | ~\new_[6177]_  | ~\new_[6218]_ ;
  assign \new_[5842]_  = ~\new_[6953]_ ;
  assign \new_[5843]_  = ~\new_[7201]_  | ~\new_[6060]_ ;
  assign \new_[5844]_  = ~\new_[6055]_  | ~\new_[6401]_ ;
  assign \new_[5845]_  = ~\new_[6152]_  & ~\new_[6007]_ ;
  assign \new_[5846]_  = ~\new_[6088]_  | ~\new_[6030]_ ;
  assign \new_[5847]_  = ~\new_[5991]_  | ~\new_[1690]_ ;
  assign \new_[5848]_  = ~\new_[6995]_  & ~\new_[7116]_ ;
  assign \new_[5849]_  = \new_[5997]_  | \new_[6163]_ ;
  assign \new_[5850]_  = ~\new_[6054]_  | ~\new_[6234]_ ;
  assign \new_[5851]_  = ~\new_[6096]_  | ~\new_[6967]_  | ~\new_[6228]_ ;
  assign \new_[5852]_  = ~\new_[6011]_  & ~\new_[6000]_ ;
  assign \new_[5853]_  = ~\new_[5975]_ ;
  assign \new_[5854]_  = ~\new_[6140]_  & ~\new_[6986]_ ;
  assign \new_[5855]_  = ~\new_[5932]_ ;
  assign \new_[5856]_  = ~\new_[6037]_  | (~\new_[2003]_  & ~\new_[1247]_ );
  assign \new_[5857]_  = ~\new_[6018]_  & (~\new_[1248]_  | ~\new_[6318]_ );
  assign \new_[5858]_  = ~\new_[6037]_  | (~\new_[2002]_  & ~\new_[1248]_ );
  assign \new_[5859]_  = ~\new_[5952]_ ;
  assign \new_[5860]_  = ~\new_[6080]_  | ~\new_[6008]_  | ~\new_[6298]_ ;
  assign \new_[5861]_  = \new_[6014]_  | \new_[6318]_ ;
  assign \new_[5862]_  = ~\new_[5947]_ ;
  assign \new_[5863]_  = ~\new_[5984]_ ;
  assign \new_[5864]_  = ~\new_[7160]_  & ~\new_[6080]_ ;
  assign \new_[5865]_  = ~\new_[5988]_ ;
  assign \new_[5866]_  = ~\new_[5966]_ ;
  assign \new_[5867]_  = ~\new_[5978]_ ;
  assign \new_[5868]_  = ~\new_[5910]_ ;
  assign \new_[5869]_  = ~\new_[6963]_  | ~\new_[6228]_ ;
  assign \new_[5870]_  = ~\new_[6478]_  | ~\new_[6782]_ ;
  assign \new_[5871]_  = ~\new_[5942]_ ;
  assign \new_[5872]_  = ~\new_[6054]_ ;
  assign \new_[5873]_  = ~\new_[6492]_  & ~\new_[6143]_ ;
  assign \new_[5874]_  = ~\new_[6053]_  | ~\new_[6987]_ ;
  assign \new_[5875]_  = ~\new_[5951]_ ;
  assign \new_[5876]_  = ~\new_[6361]_  & ~\new_[6034]_ ;
  assign \new_[5877]_  = ~\new_[6058]_  | ~\new_[6440]_ ;
  assign \new_[5878]_  = \new_[7050]_  | \new_[6782]_ ;
  assign \new_[5879]_  = ~\new_[5234]_  & ~\new_[6015]_ ;
  assign \new_[5880]_  = ~\new_[7164]_  | ~\new_[7166]_  | ~\new_[7215]_ ;
  assign \new_[5881]_  = ~\new_[5982]_ ;
  assign \new_[5882]_  = \new_[6119]_  | \new_[6080]_ ;
  assign \new_[5883]_  = ~\new_[6053]_  | ~\new_[6164]_ ;
  assign \new_[5884]_  = ~\new_[6009]_ ;
  assign \new_[5885]_  = ~\new_[5996]_  | ~\new_[6009]_ ;
  assign \new_[5886]_  = ~\new_[7116]_  | ~\new_[6359]_ ;
  assign \new_[5887]_  = ~\new_[6049]_  & ~\new_[6397]_ ;
  assign \new_[5888]_  = ~\new_[5974]_ ;
  assign \new_[5889]_  = ~\new_[6107]_ ;
  assign \new_[5890]_  = ~\new_[6032]_ ;
  assign \new_[5891]_  = ~\new_[6125]_  | ~\new_[6267]_  | ~\new_[6109]_ ;
  assign \new_[5892]_  = ~\new_[5986]_ ;
  assign \new_[5893]_  = ~\new_[6115]_  | ~\new_[7166]_ ;
  assign \new_[5894]_  = ~\new_[5949]_ ;
  assign \new_[5895]_  = \new_[5919]_ ;
  assign \new_[5896]_  = \new_[5977]_ ;
  assign \new_[5897]_  = ~\new_[6298]_  & ~\new_[7160]_ ;
  assign \new_[5898]_  = ~\new_[6042]_  | ~\new_[6312]_ ;
  assign \new_[5899]_  = ~\new_[6037]_  | (~\new_[2007]_  & ~\new_[6518]_ );
  assign \new_[5900]_  = ~\new_[6529]_  | ~\new_[1379]_  | ~\new_[6019]_  | ~\new_[1453]_ ;
  assign \new_[5901]_  = ~\new_[5990]_  | ~\new_[6038]_ ;
  assign \new_[5902]_  = ~\new_[6053]_  | ~\new_[7061]_ ;
  assign \new_[5903]_  = ~\new_[6283]_  | ~\new_[6056]_ ;
  assign \new_[5904]_  = \new_[6210]_  & \new_[1247]_ ;
  assign \new_[5905]_  = \new_[6210]_  ^ \new_[1247]_ ;
  assign \new_[5906]_  = ~\new_[7180]_ ;
  assign \new_[5907]_  = \new_[1308]_  ^ \new_[6255]_ ;
  assign \new_[5908]_  = ~\new_[6111]_  & ~\new_[6232]_ ;
  assign \new_[5909]_  = ~\new_[6055]_ ;
  assign \new_[5910]_  = ~\new_[6982]_ ;
  assign \new_[5911]_  = ~\new_[7324]_  | ~\new_[6397]_  | ~\new_[6262]_  | ~\new_[6400]_ ;
  assign \new_[5912]_  = \new_[1646]_  ^ \new_[6219]_ ;
  assign \new_[5913]_  = \new_[2551]_  ^ \new_[6222]_ ;
  assign \new_[5914]_  = ~\new_[6120]_  | ~\new_[7164]_ ;
  assign \new_[5915]_  = ~\new_[7240]_  | ~\new_[6987]_ ;
  assign \new_[5916]_  = \new_[6203]_  ^ \new_[6355]_ ;
  assign \new_[5917]_  = ~\new_[6019]_ ;
  assign \new_[5918]_  = \new_[2552]_  ^ \new_[6250]_ ;
  assign \new_[5919]_  = ~\new_[6079]_  & ~\new_[7214]_ ;
  assign \new_[5920]_  = ~\new_[6083]_  | ~\new_[6542]_ ;
  assign \new_[5921]_  = ~\new_[6091]_  & ~\new_[6343]_ ;
  assign \new_[5922]_  = ~\new_[6030]_ ;
  assign \new_[5923]_  = ~\new_[6266]_  | ~\new_[6085]_ ;
  assign \new_[5924]_  = ~\new_[6078]_  & ~\new_[6918]_ ;
  assign \new_[5925]_  = ~\new_[6040]_ ;
  assign \new_[5926]_  = ~\new_[6266]_  | ~\new_[7047]_ ;
  assign \new_[5927]_  = ~\new_[7193]_ ;
  assign \new_[5928]_  = ~\new_[6004]_ ;
  assign \new_[5929]_  = ~\new_[7124]_  | ~\new_[6106]_  | ~\new_[7125]_ ;
  assign \new_[5930]_  = \new_[6447]_  & \new_[6460]_ ;
  assign \new_[5931]_  = ~\new_[6267]_  | ~\new_[6283]_  | ~\new_[7125]_ ;
  assign \new_[5932]_  = ~\new_[7248]_  | ~\new_[6284]_ ;
  assign \new_[5933]_  = ~\new_[6077]_  & ~\new_[7119]_ ;
  assign \new_[5934]_  = ~\new_[7118]_  & ~\new_[7071]_ ;
  assign \new_[5935]_  = \new_[1324]_  | \new_[1248]_  | \new_[6278]_  | \new_[6532]_ ;
  assign \new_[5936]_  = ~\new_[6085]_  & ~\new_[6457]_ ;
  assign \new_[5937]_  = ~\new_[6108]_  & ~\new_[6804]_ ;
  assign \new_[5938]_  = ~\new_[5994]_ ;
  assign \new_[5939]_  = ~\new_[6081]_  | ~\new_[6248]_ ;
  assign \new_[5940]_  = \new_[1545]_  ^ \new_[6148]_ ;
  assign \new_[5941]_  = \new_[7324]_  & \new_[7318]_ ;
  assign \new_[5942]_  = ~\new_[7240]_  | ~\new_[6109]_ ;
  assign \new_[5943]_  = \new_[6536]_  ^ \new_[6161]_ ;
  assign \new_[5944]_  = ~\new_[6523]_  | ~\new_[6603]_  | ~\new_[3281]_ ;
  assign \new_[5945]_  = ~\new_[6097]_  | (~\new_[6310]_  & ~\new_[1126]_ );
  assign \new_[5946]_  = \new_[7318]_  | \new_[6107]_ ;
  assign \new_[5947]_  = ~\new_[6123]_  | ~\new_[6103]_ ;
  assign \new_[5948]_  = \new_[6077]_  | \new_[6804]_ ;
  assign \new_[5949]_  = ~\new_[6801]_ ;
  assign \new_[5950]_  = ~\new_[7240]_  | ~\new_[7061]_ ;
  assign \new_[5951]_  = ~\new_[7056]_ ;
  assign \new_[5952]_  = \new_[6069]_  & \new_[6103]_ ;
  assign \new_[5953]_  = ~\new_[6117]_  & ~\new_[1248]_ ;
  assign \new_[5954]_  = ~\new_[7119]_  & ~\new_[6108]_ ;
  assign \new_[5955]_  = ~\new_[6009]_  | ~\new_[6164]_  | ~\new_[6445]_ ;
  assign \new_[5956]_  = ~\new_[6119]_  & ~\new_[7161]_ ;
  assign \new_[5957]_  = ~\new_[5999]_ ;
  assign \new_[5958]_  = ~\new_[6918]_  & ~\new_[7071]_ ;
  assign \new_[5959]_  = ~\new_[6127]_  & ~\new_[6620]_ ;
  assign \new_[5960]_  = \new_[6262]_  & \new_[6096]_ ;
  assign \new_[5961]_  = ~\new_[6016]_ ;
  assign \new_[5962]_  = ~\new_[6041]_ ;
  assign \new_[5963]_  = \new_[6169]_  ^ \new_[1324]_ ;
  assign \new_[5964]_  = ~\new_[6396]_  | (~\new_[6419]_  & ~\new_[6442]_ );
  assign \new_[5965]_  = \new_[2016]_  ^ \new_[6429]_ ;
  assign \new_[5966]_  = ~\new_[6394]_  | ~\new_[6128]_ ;
  assign \new_[5967]_  = ~\new_[6305]_  & ~\new_[6359]_ ;
  assign \new_[5968]_  = \new_[6077]_  | \new_[7071]_ ;
  assign \new_[5969]_  = ~\new_[6031]_ ;
  assign \new_[5970]_  = ~\new_[6394]_  | ~\new_[6084]_ ;
  assign \new_[5971]_  = ~\new_[6280]_  | ~\new_[1247]_ ;
  assign \new_[5972]_  = ~\new_[6080]_ ;
  assign \new_[5973]_  = ~\new_[6120]_  & ~\new_[7162]_ ;
  assign \new_[5974]_  = \new_[6121]_  & \new_[6965]_ ;
  assign \new_[5975]_  = ~\new_[6087]_  | ~\new_[6090]_ ;
  assign \new_[5976]_  = \new_[1248]_  ^ \new_[6160]_ ;
  assign \new_[5977]_  = ~\new_[6066]_  | ~\new_[6093]_ ;
  assign \new_[5978]_  = ~\new_[6117]_  | ~\new_[1248]_ ;
  assign \new_[5979]_  = ~\new_[5991]_ ;
  assign \new_[5980]_  = ~\new_[6007]_ ;
  assign \new_[5981]_  = ~\new_[6050]_ ;
  assign \new_[5982]_  = ~\new_[6620]_  & ~\new_[6460]_ ;
  assign \new_[5983]_  = ~\new_[5992]_ ;
  assign \new_[5984]_  = ~\new_[6077]_  & ~\new_[6078]_ ;
  assign \new_[5985]_  = ~\new_[6114]_  & ~\new_[6442]_ ;
  assign \new_[5986]_  = ~\new_[6101]_  | ~\new_[7215]_ ;
  assign \new_[5987]_  = ~\new_[6164]_  | ~\new_[7240]_ ;
  assign \new_[5988]_  = ~\new_[7064]_ ;
  assign \new_[5989]_  = ~\new_[6130]_  | ~\new_[6536]_ ;
  assign \new_[5990]_  = ~\new_[6108]_ ;
  assign \new_[5991]_  = i_tv80_core_BusReq_s_reg;
  assign \new_[5992]_  = \new_[6378]_  & \new_[6359]_ ;
  assign \new_[5993]_  = ~\new_[6081]_ ;
  assign \new_[5994]_  = \new_[7248]_ ;
  assign \new_[5995]_  = ~\new_[6272]_ ;
  assign \new_[5996]_  = \new_[6400]_  & \new_[6143]_ ;
  assign \new_[5997]_  = ~\new_[6236]_  & ~\new_[6163]_ ;
  assign \new_[5998]_  = ~\new_[6212]_  | ~\new_[6248]_ ;
  assign \new_[5999]_  = \new_[6158]_  | \new_[1126]_ ;
  assign \new_[6000]_  = ~\new_[2002]_  | ~\new_[6167]_ ;
  assign \new_[6001]_  = ~\new_[2002]_  & ~\new_[6167]_ ;
  assign \new_[6002]_  = ~\new_[6175]_ ;
  assign \new_[6003]_  = ~\new_[7201]_  | ~\new_[6995]_ ;
  assign \new_[6004]_  = \new_[7047]_ ;
  assign \new_[6005]_  = ~\new_[6074]_ ;
  assign \new_[6006]_  = ~\new_[6141]_  | ~\new_[6419]_ ;
  assign \new_[6007]_  = ~\new_[6244]_  | ~\new_[7161]_ ;
  assign \new_[6008]_  = ~\new_[7028]_  & (~\new_[7298]_  | ~\new_[7549]_ );
  assign \new_[6009]_  = ~\new_[7318]_ ;
  assign \new_[6010]_  = ~\new_[7071]_ ;
  assign \new_[6011]_  = ~\new_[1811]_  | ~\new_[6952]_  | ~\new_[1624]_ ;
  assign \new_[6012]_  = \new_[6451]_  ^ \new_[6565]_ ;
  assign \new_[6013]_  = ~\new_[6116]_ ;
  assign \new_[6014]_  = \new_[7557]_  & \new_[6143]_ ;
  assign \new_[6015]_  = ~\new_[6102]_ ;
  assign \new_[6016]_  = ~\new_[6139]_  | ~\new_[6307]_ ;
  assign \new_[6017]_  = i_tv80_core_Oldnmi_n_reg;
  assign \new_[6018]_  = ~\new_[6818]_ ;
  assign \new_[6019]_  = \new_[6353]_  & \new_[6219]_ ;
  assign \new_[6020]_  = ~\new_[6635]_  | ~\new_[6365]_ ;
  assign \new_[6021]_  = \new_[1324]_  ^ \new_[6274]_ ;
  assign \new_[6022]_  = \new_[6142]_  & \new_[7190]_ ;
  assign \new_[6023]_  = ~\new_[2135]_  | ~\new_[6190]_ ;
  assign \new_[6024]_  = \new_[1247]_  ^ \new_[6278]_ ;
  assign \new_[6025]_  = ~\new_[6256]_  | (~\new_[6340]_  & ~\new_[1324]_ );
  assign \new_[6026]_  = ~\new_[6090]_ ;
  assign \new_[6027]_  = ~\new_[6207]_  | (~\new_[6335]_  & ~\new_[6648]_ );
  assign \new_[6028]_  = ~\new_[6204]_  & ~\new_[6373]_ ;
  assign \new_[6029]_  = ~\new_[6135]_  | ~\new_[1231]_ ;
  assign \new_[6030]_  = ~\new_[6135]_  & ~\new_[1231]_ ;
  assign \new_[6031]_  = ~\new_[6313]_ ;
  assign \new_[6032]_  = ~\new_[6985]_  & ~\new_[6206]_ ;
  assign \new_[6033]_  = ~\A[2]  | ~\new_[6190]_ ;
  assign \new_[6034]_  = ~\new_[6067]_ ;
  assign \new_[6035]_  = i_tv80_core_INT_s_reg;
  assign \new_[6036]_  = ~\new_[6158]_  | ~\new_[1126]_ ;
  assign \new_[6037]_  = \new_[6447]_  & \new_[6429]_ ;
  assign \new_[6038]_  = ~\new_[6078]_ ;
  assign \new_[6039]_  = ~\new_[7550]_  & ~\new_[7253]_ ;
  assign \new_[6040]_  = \new_[6952]_  & \new_[6440]_ ;
  assign \new_[6041]_  = ~\new_[6141]_  | ~\new_[6452]_ ;
  assign \new_[6042]_  = ~\new_[6331]_  & ~\new_[7169]_ ;
  assign \new_[6043]_  = \new_[6316]_  ^ \new_[1247]_ ;
  assign \new_[6044]_  = \new_[7246]_  ^ \new_[7318]_ ;
  assign \new_[6045]_  = \new_[2863]_  ^ \new_[6442]_ ;
  assign \new_[6046]_  = ~\new_[6394]_  | ~\new_[6359]_ ;
  assign \new_[6047]_  = ~\new_[6264]_ ;
  assign \new_[6048]_  = ~\new_[6284]_  & ~\new_[6442]_ ;
  assign \new_[6049]_  = ~\new_[7550]_  | ~\new_[6227]_ ;
  assign \new_[6050]_  = ~\new_[7118]_  & ~\new_[6804]_ ;
  assign \new_[6051]_  = ~\A[6]  | ~\new_[6190]_ ;
  assign \new_[6052]_  = ~\A[5]  | ~\new_[6190]_ ;
  assign \new_[6053]_  = \new_[6171]_  & \new_[6281]_ ;
  assign \new_[6054]_  = ~\new_[6213]_  & ~\new_[7214]_ ;
  assign \new_[6055]_  = wait_n | \new_[6365]_ ;
  assign \new_[6056]_  = ~\new_[6918]_ ;
  assign \new_[6057]_  = ~\new_[6516]_  | ~\new_[1453]_  | ~\new_[6255]_  | ~\new_[1308]_ ;
  assign \new_[6058]_  = ~\new_[6127]_ ;
  assign \new_[6059]_  = ~\new_[6145]_  & (~\new_[6350]_  | ~\new_[1126]_ );
  assign \new_[6060]_  = ~\new_[7119]_  & ~\new_[7073]_ ;
  assign \new_[6061]_  = ~\new_[6085]_ ;
  assign \new_[6062]_  = ~\new_[6009]_  | ~\new_[7323]_ ;
  assign \new_[6063]_  = ~\A[1]  | ~\new_[6190]_ ;
  assign \new_[6064]_  = ~\new_[6133]_ ;
  assign \new_[6065]_  = ~\new_[6104]_ ;
  assign \new_[6066]_  = ~\new_[7325]_  & ~\new_[7318]_ ;
  assign \new_[6067]_  = ~\new_[6298]_ ;
  assign \new_[6068]_  = \new_[6460]_  ^ \new_[6362]_ ;
  assign \new_[6069]_  = ~\new_[7060]_ ;
  assign \new_[6070]_  = ~\new_[6251]_ ;
  assign \new_[6071]_  = ~\new_[6284]_ ;
  assign \new_[6072]_  = ~\new_[1324]_  | ~\new_[6280]_ ;
  assign \new_[6073]_  = ~\new_[6280]_  | ~\new_[1248]_ ;
  assign \new_[6074]_  = ~\new_[1578]_  | ~\new_[1646]_  | ~\new_[6320]_  | ~\new_[1689]_ ;
  assign \new_[6075]_  = ~\new_[6168]_ ;
  assign \new_[6076]_  = \new_[1324]_  & \new_[6318]_ ;
  assign \new_[6077]_  = ~\new_[6282]_  | ~\new_[7028]_ ;
  assign \new_[6078]_  = ~\new_[7124]_  | ~\new_[7030]_ ;
  assign \new_[6079]_  = ~\new_[7168]_  | ~\new_[6397]_ ;
  assign \new_[6080]_  = ~\new_[6229]_  | ~\new_[7298]_ ;
  assign \new_[6081]_  = ~\new_[6275]_  & ~\new_[6648]_ ;
  assign \new_[6082]_  = \new_[1248]_  ^ \new_[6368]_ ;
  assign \new_[6083]_  = ~\new_[6173]_ ;
  assign \new_[6084]_  = ~\new_[6400]_ ;
  assign \new_[6085]_  = \new_[6302]_  | \new_[6404]_ ;
  assign \new_[6086]_  = \new_[1689]_  ^ \new_[6373]_ ;
  assign \new_[6087]_  = \new_[6265]_  | \new_[6668]_ ;
  assign \new_[6088]_  = ~\new_[6135]_ ;
  assign \new_[6089]_  = \new_[6336]_  ^ \new_[1247]_ ;
  assign \new_[6090]_  = ~\new_[6265]_  | ~\new_[6668]_ ;
  assign \new_[6091]_  = ~\new_[7061]_  | ~\new_[7231]_ ;
  assign \new_[6092]_  = \new_[2555]_  ^ \new_[6345]_ ;
  assign \new_[6093]_  = \new_[6307]_  & \new_[7552]_ ;
  assign \new_[6094]_  = \new_[2929]_  ^ \new_[6452]_ ;
  assign \new_[6095]_  = \new_[6367]_  ^ \new_[1126]_ ;
  assign \new_[6096]_  = ~\new_[6400]_  & ~\new_[7253]_ ;
  assign \new_[6097]_  = ~\new_[6310]_  | ~\new_[1126]_ ;
  assign \new_[6098]_  = \new_[6292]_  & \new_[6336]_ ;
  assign \new_[6099]_  = ~\new_[1690]_ ;
  assign \new_[6100]_  = ~\new_[6279]_  & ~\new_[6523]_ ;
  assign \new_[6101]_  = ~\new_[7214]_  & ~\new_[7213]_ ;
  assign \new_[6102]_  = \new_[7319]_  | \new_[7193]_ ;
  assign \new_[6103]_  = \new_[6488]_  & \new_[7253]_ ;
  assign \new_[6104]_  = ~\new_[7246]_  & ~\new_[6298]_ ;
  assign \new_[6105]_  = \new_[2553]_  ^ \new_[6377]_ ;
  assign \new_[6106]_  = \new_[6267]_  & \new_[6465]_ ;
  assign \new_[6107]_  = ~\new_[6234]_ ;
  assign \new_[6108]_  = ~\new_[6282]_  | ~\new_[7125]_ ;
  assign \new_[6109]_  = ~\new_[6960]_ ;
  assign \new_[6110]_  = ~\new_[6161]_ ;
  assign \new_[6111]_  = \new_[7246]_  ^ \new_[6397]_ ;
  assign \new_[6112]_  = \new_[6586]_  ^ \new_[6668]_ ;
  assign \new_[6113]_  = ~\new_[6397]_ ;
  assign \new_[6114]_  = ~\new_[6142]_ ;
  assign \new_[6115]_  = ~\new_[7326]_  & ~\new_[7162]_ ;
  assign \new_[6116]_  = ~\new_[6205]_ ;
  assign \new_[6117]_  = \new_[2002]_  ^ \new_[6429]_ ;
  assign \new_[6118]_  = ~\new_[6515]_  | ~\new_[6819]_ ;
  assign \new_[6119]_  = ~\new_[6244]_ ;
  assign \new_[6120]_  = ~\new_[6229]_ ;
  assign \new_[6121]_  = ~\new_[7296]_ ;
  assign \new_[6122]_  = ~\new_[6280]_  | ~\new_[1126]_ ;
  assign \new_[6123]_  = ~\new_[7036]_ ;
  assign \new_[6124]_  = ~\new_[6394]_  & ~\new_[6293]_ ;
  assign \new_[6125]_  = ~\new_[6240]_ ;
  assign \new_[6126]_  = ~\new_[1690]_ ;
  assign \new_[6127]_  = ~\new_[6460]_  | ~\new_[1810]_ ;
  assign \new_[6128]_  = ~\new_[6143]_ ;
  assign \new_[6129]_  = ~\new_[1690]_ ;
  assign \new_[6130]_  = ~\new_[1126]_  & (~\new_[6423]_  | ~\new_[1247]_ );
  assign \new_[6131]_  = \new_[1578]_  ^ \new_[6349]_ ;
  assign \new_[6132]_  = ~\new_[1690]_ ;
  assign \new_[6133]_  = ~\new_[7145]_ ;
  assign \new_[6134]_  = ~\new_[6160]_ ;
  assign \new_[6135]_  = ~\new_[6395]_  | ~\new_[6366]_ ;
  assign \new_[6136]_  = ~\new_[1811]_  | ~\new_[6406]_ ;
  assign \new_[6137]_  = ~\new_[6985]_  & ~\new_[6331]_ ;
  assign \new_[6138]_  = ~\new_[1324]_  | ~\new_[7050]_ ;
  assign \new_[6139]_  = ~\new_[7067]_ ;
  assign \new_[6140]_  = ~\new_[7193]_ ;
  assign \new_[6141]_  = ~\new_[6895]_  & ~\new_[6442]_ ;
  assign \new_[6142]_  = ~\new_[6455]_  | ~\new_[6981]_ ;
  assign \new_[6143]_  = ~\new_[6296]_ ;
  assign \new_[6144]_  = (~\new_[6408]_  | ~\new_[6612]_ ) & (~\new_[6446]_  | ~\new_[6597]_ );
  assign \new_[6145]_  = ~\new_[6350]_  & ~\new_[1126]_ ;
  assign \new_[6146]_  = (~\new_[6463]_  | ~\new_[660]_ ) & (~\new_[6381]_  | ~\new_[661]_ );
  assign \new_[6147]_  = (~\new_[6404]_  & ~\new_[6895]_ ) | (~\new_[6399]_  & ~\new_[6452]_ );
  assign \new_[6148]_  = ~\new_[6373]_  & ~\new_[6421]_ ;
  assign \new_[6149]_  = ~\new_[6387]_ ;
  assign \new_[6150]_  = (~\new_[6389]_  | ~\new_[6583]_ ) & (~\new_[6386]_  | ~\new_[6639]_ );
  assign \new_[6151]_  = (~\new_[6463]_  | ~\new_[652]_ ) & (~\new_[6381]_  | ~\new_[653]_ );
  assign \new_[6152]_  = ~\new_[7298]_ ;
  assign \new_[6153]_  = (~\new_[6463]_  | ~\new_[429]_ ) & (~\new_[6381]_  | ~\new_[430]_ );
  assign n1879 = ~\new_[6619]_  & ~\new_[6371]_ ;
  assign \new_[6155]_  = (~\new_[6389]_  | ~\new_[539]_ ) & (~\new_[6386]_  | ~\new_[540]_ );
  assign \new_[6156]_  = ~\new_[6271]_ ;
  assign \new_[6157]_  = (~\new_[6408]_  | ~\new_[520]_ ) & (~\new_[6446]_  | ~\new_[542]_ );
  assign \new_[6158]_  = \new_[2006]_  ^ \new_[6429]_ ;
  assign \new_[6159]_  = (~\new_[6389]_  | ~\new_[788]_ ) & (~\new_[6386]_  | ~\new_[789]_ );
  assign \new_[6160]_  = ~\new_[1126]_  | ~\new_[6423]_  | ~\new_[1247]_ ;
  assign \new_[6161]_  = (~\new_[6548]_  | ~\new_[6620]_ ) & (~\new_[2006]_  | ~\new_[1811]_ );
  assign \new_[6162]_  = ~\new_[6258]_ ;
  assign \new_[6163]_  = ~\new_[6333]_  & ~\new_[1620]_ ;
  assign \new_[6164]_  = \new_[6341]_  & \new_[6917]_ ;
  assign \new_[6165]_  = ~\new_[6387]_ ;
  assign \new_[6166]_  = \new_[7252]_  | \new_[7553]_ ;
  assign \new_[6167]_  = ~\new_[7170]_ ;
  assign \new_[6168]_  = \new_[6996]_  | \new_[7326]_ ;
  assign \new_[6169]_  = \new_[6538]_  | \new_[6350]_ ;
  assign \new_[6170]_  = \new_[1861]_  ^ \new_[6409]_ ;
  assign \new_[6171]_  = \new_[6282]_ ;
  assign \new_[6172]_  = (~\new_[6463]_  | ~\new_[731]_ ) & (~\new_[6381]_  | ~\new_[735]_ );
  assign \new_[6173]_  = ~\new_[6280]_ ;
  assign \new_[6174]_  = (~\new_[6408]_  | ~\new_[656]_ ) & (~\new_[6446]_  | ~\new_[657]_ );
  assign \new_[6175]_  = ~\new_[6337]_  | ~\new_[7324]_ ;
  assign \new_[6176]_  = (~\new_[6408]_  | ~\new_[572]_ ) & (~\new_[6446]_  | ~\new_[573]_ );
  assign \new_[6177]_  = (~\new_[6408]_  | ~\new_[778]_ ) & (~\new_[6446]_  | ~\new_[779]_ );
  assign \new_[6178]_  = (~\new_[6463]_  | ~\new_[768]_ ) & (~\new_[6381]_  | ~\new_[769]_ );
  assign \new_[6179]_  = (~\new_[6463]_  | ~\new_[568]_ ) & (~\new_[6381]_  | ~\new_[569]_ );
  assign \new_[6180]_  = (~\new_[6408]_  | ~\new_[433]_ ) & (~\new_[6446]_  | ~\new_[434]_ );
  assign \new_[6181]_  = (~\new_[6408]_  | ~n324) & (~\new_[6446]_  | ~n329);
  assign \new_[6182]_  = (~\new_[6408]_  | ~\new_[665]_ ) & (~\new_[6446]_  | ~\new_[663]_ );
  assign \new_[6183]_  = (~\new_[6408]_  | ~\new_[685]_ ) & (~\new_[6446]_  | ~\new_[686]_ );
  assign \new_[6184]_  = (~\new_[6389]_  | ~\new_[662]_ ) & (~\new_[6386]_  | ~\new_[646]_ );
  assign \new_[6185]_  = (~\new_[6463]_  | ~\new_[786]_ ) & (~\new_[6381]_  | ~\new_[787]_ );
  assign \new_[6186]_  = (~\new_[6389]_  | ~\new_[770]_ ) & (~\new_[6386]_  | ~\new_[796]_ );
  assign \new_[6187]_  = (~\new_[6463]_  | ~\new_[529]_ ) & (~\new_[6381]_  | ~\new_[530]_ );
  assign \new_[6188]_  = (~\new_[6463]_  | ~\new_[6618]_ ) & (~\new_[6381]_  | ~\new_[6615]_ );
  assign \new_[6189]_  = (~\new_[6408]_  | ~\new_[6672]_ ) & (~\new_[6446]_  | ~\new_[7513]_ );
  assign \new_[6190]_  = ~\new_[6388]_ ;
  assign \new_[6191]_  = (~\new_[6389]_  | ~\new_[732]_ ) & (~\new_[6386]_  | ~\new_[733]_ );
  assign \new_[6192]_  = (~\new_[6408]_  | ~\new_[771]_ ) & (~\new_[6446]_  | ~\new_[772]_ );
  assign \new_[6193]_  = ~\new_[6495]_ ;
  assign \new_[6194]_  = (~\new_[6463]_  | ~\new_[775]_ ) & (~\new_[6381]_  | ~\new_[776]_ );
  assign \new_[6195]_  = (~\new_[6463]_  | ~\new_[575]_ ) & (~\new_[6381]_  | ~\new_[576]_ );
  assign \new_[6196]_  = (~\new_[6389]_  | ~\new_[6660]_ ) & (~\new_[6386]_  | ~\new_[6599]_ );
  assign \new_[6197]_  = (~\new_[6408]_  | ~\new_[6496]_ ) & (~\new_[6446]_  | ~\new_[6512]_ );
  assign \new_[6198]_  = (~\new_[6389]_  | ~n314) & (~\new_[6386]_  | ~n319);
  assign \new_[6199]_  = (~\new_[6463]_  | ~\new_[6627]_ ) & (~\new_[6381]_  | ~\new_[6645]_ );
  assign \new_[6200]_  = (~\new_[6408]_  | ~\new_[790]_ ) & (~\new_[6446]_  | ~\new_[797]_ );
  assign \new_[6201]_  = (~\new_[6463]_  | ~\new_[537]_ ) & (~\new_[6381]_  | ~\new_[538]_ );
  assign \new_[6202]_  = (~\new_[6463]_  | ~\new_[6566]_ ) & (~\new_[6381]_  | ~\new_[6642]_ );
  assign \new_[6203]_  = \new_[6392]_  ^ \new_[6485]_ ;
  assign \new_[6204]_  = ~\new_[6372]_  | ~\new_[1308]_ ;
  assign \new_[6205]_  = ~\new_[6337]_  | ~\new_[6369]_ ;
  assign \new_[6206]_  = ~\new_[6307]_ ;
  assign \new_[6207]_  = ~\new_[6335]_  | ~\new_[6648]_ ;
  assign \new_[6208]_  = (~\new_[6389]_  | ~\new_[577]_ ) & (~\new_[6386]_  | ~\new_[560]_ );
  assign \new_[6209]_  = \new_[6674]_  ^ \new_[6430]_ ;
  assign \new_[6210]_  = \new_[2003]_  ^ \new_[6429]_ ;
  assign \new_[6211]_  = ~\new_[1810]_  | ~\new_[6406]_ ;
  assign \new_[6212]_  = \new_[6346]_  | \new_[6586]_ ;
  assign \new_[6213]_  = \new_[7169]_  | \new_[6397]_ ;
  assign \new_[6214]_  = (~\new_[6408]_  | ~\new_[578]_ ) & (~\new_[6446]_  | ~\new_[579]_ );
  assign \new_[6215]_  = ~\new_[6264]_ ;
  assign \new_[6216]_  = ~\new_[6730]_ ;
  assign \new_[6217]_  = (~\new_[6389]_  | ~\new_[431]_ ) & (~\new_[6386]_  | ~\new_[432]_ );
  assign \new_[6218]_  = (~\new_[6389]_  | ~\new_[777]_ ) & (~\new_[6386]_  | ~\new_[737]_ );
  assign \new_[6219]_  = ~\new_[6321]_  & ~\new_[6543]_ ;
  assign \new_[6220]_  = ~\new_[1690]_ ;
  assign \new_[6221]_  = (~\new_[6389]_  | ~\new_[6641]_ ) & (~\new_[6386]_  | ~\new_[6587]_ );
  assign \new_[6222]_  = ~\new_[2552]_  | ~\new_[2553]_  | ~\new_[6377]_  | ~\new_[2555]_ ;
  assign \new_[6223]_  = ~\new_[4560]_  & ~\new_[6264]_ ;
  assign \new_[6224]_  = ~\new_[1690]_ ;
  assign \new_[6225]_  = ~\new_[6387]_ ;
  assign \new_[6226]_  = ~\new_[6388]_ ;
  assign \new_[6227]_  = ~\new_[7253]_ ;
  assign \new_[6228]_  = ~\new_[6358]_  & ~\new_[6331]_ ;
  assign \new_[6229]_  = ~\new_[7161]_ ;
  assign n1874 = ~busrq_n & ~\new_[6371]_ ;
  assign \new_[6231]_  = ~\new_[6473]_  | ~\new_[6917]_ ;
  assign \new_[6232]_  = ~\new_[6262]_ ;
  assign \new_[6233]_  = ~\new_[6305]_ ;
  assign \new_[6234]_  = ~\new_[6309]_ ;
  assign \new_[6235]_  = (~\new_[6389]_  | ~\new_[534]_ ) & (~\new_[6386]_  | ~\new_[535]_ );
  assign \new_[6236]_  = ~\new_[6333]_  & ~\new_[6634]_ ;
  assign \new_[6237]_  = (~\new_[6389]_  | ~\new_[654]_ ) & (~\new_[6386]_  | ~\new_[655]_ );
  assign \new_[6238]_  = (~\new_[6389]_  | ~\new_[570]_ ) & (~\new_[6386]_  | ~\new_[571]_ );
  assign \new_[6239]_  = ~\new_[6387]_ ;
  assign \new_[6240]_  = ~\new_[6281]_ ;
  assign \new_[6241]_  = (~\new_[6408]_  | ~\new_[531]_ ) & (~\new_[6446]_  | ~\new_[532]_ );
  assign \new_[6242]_  = (~\new_[6408]_  | ~\new_[6559]_ ) & (~\new_[6446]_  | ~\new_[6482]_ );
  assign \new_[6243]_  = ~\new_[1579]_  | ~\new_[6634]_  | ~\new_[6453]_  | ~\new_[6570]_ ;
  assign \new_[6244]_  = \new_[6420]_  | \new_[7553]_ ;
  assign \new_[6245]_  = \new_[6360]_  | \new_[6634]_ ;
  assign \new_[6246]_  = ~\new_[6379]_  & ~\new_[6634]_ ;
  assign \new_[6247]_  = (~\new_[6463]_  | ~\new_[6590]_ ) & (~\new_[6381]_  | ~\new_[6564]_ );
  assign \new_[6248]_  = ~\new_[6346]_  | ~\new_[6586]_ ;
  assign \new_[6249]_  = (~\new_[6463]_  | ~n304) & (~\new_[6381]_  | ~n309);
  assign \new_[6250]_  = \new_[6524]_  & \new_[6377]_ ;
  assign \new_[6251]_  = ~\new_[6266]_ ;
  assign \new_[6252]_  = ~\new_[6348]_ ;
  assign n1884 = ~int_n & ~\new_[6371]_ ;
  assign \new_[6254]_  = (~\new_[6389]_  | ~\new_[6556]_ ) & (~\new_[6386]_  | ~\new_[6657]_ );
  assign \new_[6255]_  = ~\new_[6354]_  & ~\new_[6349]_ ;
  assign \new_[6256]_  = ~\new_[6340]_  | ~\new_[1324]_ ;
  assign \new_[6257]_  = ~\new_[6379]_  & ~\new_[1620]_ ;
  assign \new_[6258]_  = ~\new_[6326]_ ;
  assign \new_[6259]_  = (~\new_[6464]_  | ~\new_[785]_ ) & (~\new_[6459]_  | ~\new_[791]_ );
  assign \new_[6260]_  = (~\new_[6464]_  | ~\new_[659]_ ) & (~\new_[6459]_  | ~\new_[664]_ );
  assign \new_[6261]_  = ~\new_[6714]_ ;
  assign \new_[6262]_  = ~\new_[6385]_  & ~\new_[7553]_ ;
  assign \new_[6263]_  = ~\new_[6347]_ ;
  assign \new_[6264]_  = ~\new_[6384]_ ;
  assign \new_[6265]_  = ~\new_[6493]_  & ~\new_[6390]_ ;
  assign \new_[6266]_  = \new_[6407]_  & \new_[6470]_ ;
  assign \new_[6267]_  = ~\new_[6959]_ ;
  assign \new_[6268]_  = \new_[6811]_ ;
  assign \new_[6269]_  = (~\new_[6464]_  | ~\new_[6598]_ ) & (~\new_[6459]_  | ~\new_[6652]_ );
  assign \new_[6270]_  = (~\new_[6464]_  | ~\new_[730]_ ) & (~\new_[6459]_  | ~\new_[734]_ );
  assign \new_[6271]_  = ~wait_n | ~\new_[7308]_ ;
  assign \new_[6272]_  = \new_[6364]_ ;
  assign \new_[6273]_  = (~\new_[6464]_  | ~\new_[528]_ ) & (~\new_[6459]_  | ~\new_[533]_ );
  assign \new_[6274]_  = ~\new_[6536]_  | ~\new_[6436]_  | ~\new_[6444]_ ;
  assign \new_[6275]_  = ~\new_[6335]_ ;
  assign \new_[6276]_  = (~\new_[6464]_  | ~\new_[767]_ ) & (~\new_[6459]_  | ~\new_[773]_ );
  assign \new_[6277]_  = ~\new_[6360]_ ;
  assign \new_[6278]_  = \new_[2007]_  ? \new_[1811]_  : \new_[2002]_ ;
  assign \new_[6279]_  = ~\new_[6571]_  | ~halt_n;
  assign \new_[6280]_  = ~\new_[6423]_  & ~\new_[850]_ ;
  assign \new_[6281]_  = ~\new_[6343]_ ;
  assign \new_[6282]_  = \new_[7245]_ ;
  assign \new_[6283]_  = \new_[6465]_  & \new_[7031]_ ;
  assign \new_[6284]_  = ~\new_[6981]_ ;
  assign \new_[6285]_  = \new_[2554]_  ^ \new_[6474]_ ;
  assign \new_[6286]_  = (~\new_[6464]_  | ~\new_[6644]_ ) & (~\new_[6459]_  | ~\new_[6673]_ );
  assign \new_[6287]_  = \new_[1892]_  ^ \new_[6456]_ ;
  assign \new_[6288]_  = (~\new_[6464]_  | ~\new_[574]_ ) & (~\new_[6459]_  | ~\new_[580]_ );
  assign \new_[6289]_  = (~\new_[6464]_  | ~\new_[536]_ ) & (~\new_[6459]_  | ~\new_[543]_ );
  assign \new_[6290]_  = \new_[6677]_  ^ \new_[6525]_ ;
  assign \new_[6291]_  = (~\new_[6464]_  | ~n299) & (~\new_[6459]_  | ~n334);
  assign \new_[6292]_  = \new_[6436]_  | \new_[6565]_ ;
  assign \new_[6293]_  = ~\new_[6359]_ ;
  assign \new_[6294]_  = (~\new_[6464]_  | ~\new_[6491]_ ) & (~\new_[6459]_  | ~\new_[6607]_ );
  assign \new_[6295]_  = ~\new_[6441]_ ;
  assign \new_[6296]_  = ~\new_[7246]_ ;
  assign \new_[6297]_  = ~\new_[6406]_  | ~\new_[2926]_ ;
  assign \new_[6298]_  = \new_[6651]_  | \new_[7298]_ ;
  assign \new_[6299]_  = ~\new_[6348]_ ;
  assign \new_[6300]_  = ~\new_[6664]_  | ~\new_[6565]_ ;
  assign \new_[6301]_  = (~\new_[6464]_  | ~\new_[428]_ ) & (~\new_[6459]_  | ~\new_[435]_ );
  assign \new_[6302]_  = ~\new_[6391]_  | ~\new_[6895]_ ;
  assign \new_[6303]_  = (~\new_[6464]_  | ~\new_[567]_ ) & (~\new_[6459]_  | ~\new_[562]_ );
  assign \new_[6304]_  = ~\new_[6441]_ ;
  assign \new_[6305]_  = \new_[6405]_  & \new_[6442]_ ;
  assign \new_[6306]_  = \new_[2005]_  ^ \new_[6542]_ ;
  assign \new_[6307]_  = \new_[6651]_  & \new_[6397]_ ;
  assign \new_[6308]_  = (~\new_[6464]_  | ~\new_[6633]_ ) & (~\new_[6459]_  | ~\new_[6665]_ );
  assign \new_[6309]_  = ~\new_[7127]_ ;
  assign \new_[6310]_  = (~\new_[2005]_  | ~\new_[6620]_ ) & (~\new_[2016]_  | ~\new_[1811]_ );
  assign \new_[6311]_  = (~\new_[6464]_  | ~\new_[650]_ ) & (~\new_[6459]_  | ~\new_[658]_ );
  assign \new_[6312]_  = ~\new_[6358]_ ;
  assign \new_[6313]_  = ~\new_[6935]_ ;
  assign \new_[6314]_  = ~\new_[1690]_ ;
  assign \new_[6315]_  = ~\new_[7128]_  & ~\new_[6495]_ ;
  assign \new_[6316]_  = ~\new_[6423]_ ;
  assign \new_[6317]_  = ~\new_[6400]_  & ~\new_[7325]_ ;
  assign \new_[6318]_  = \new_[6375]_ ;
  assign \new_[6319]_  = (~\new_[6464]_  | ~\new_[774]_ ) & (~\new_[6459]_  | ~\new_[780]_ );
  assign \new_[6320]_  = ~\new_[6409]_  & ~\new_[6661]_ ;
  assign \new_[6321]_  = ~\new_[6456]_  | ~\new_[6505]_ ;
  assign \new_[6322]_  = ~\new_[6387]_ ;
  assign \new_[6323]_  = ~reset_n;
  assign \new_[6324]_  = \new_[2002]_  ^ \new_[1248]_ ;
  assign \new_[6325]_  = ~\new_[6394]_ ;
  assign \new_[6326]_  = \new_[6714]_ ;
  assign \new_[6327]_  = ~reset_n;
  assign \new_[6328]_  = ~\new_[6437]_  & ~\new_[6704]_ ;
  assign \new_[6329]_  = ~reset_n;
  assign \new_[6330]_  = ~\new_[7134]_  & (~\new_[6517]_  | ~\new_[597]_ );
  assign \new_[6331]_  = ~\new_[7251]_ ;
  assign \new_[6332]_  = ~\new_[6539]_  & ~\new_[597]_ ;
  assign \new_[6333]_  = ~\new_[6453]_  | ~\new_[6511]_ ;
  assign \new_[6334]_  = ~\new_[6388]_ ;
  assign \new_[6335]_  = ~\new_[6487]_  | ~\new_[6443]_ ;
  assign \new_[6336]_  = ~\new_[6436]_  | ~\new_[6565]_ ;
  assign \new_[6337]_  = \new_[6435]_  & \new_[7552]_ ;
  assign \new_[6338]_  = ~\new_[6388]_ ;
  assign \new_[6339]_  = \new_[6654]_  ^ \new_[6668]_ ;
  assign \new_[6340]_  = (~\new_[6528]_  | ~\new_[6620]_ ) & (~\new_[2003]_  | ~\new_[1811]_ );
  assign \new_[6341]_  = ~\new_[6988]_ ;
  assign \new_[6342]_  = ~\new_[6623]_  & ~\new_[1690]_ ;
  assign \new_[6343]_  = \new_[7246]_  | \new_[7299]_ ;
  assign \new_[6344]_  = ~\new_[6679]_  | ~\new_[6586]_ ;
  assign \new_[6345]_  = \new_[6544]_  & \new_[6474]_ ;
  assign \new_[6346]_  = ~\new_[6479]_  & ~\new_[6469]_ ;
  assign \new_[6347]_  = ~busak_n;
  assign \new_[6348]_  = ~\new_[1690]_ ;
  assign \new_[6349]_  = ~\new_[1861]_  | ~\new_[1689]_  | ~\new_[6456]_  | ~\new_[1892]_ ;
  assign \new_[6350]_  = ~\new_[1247]_  | ~\new_[6451]_  | ~\new_[1231]_ ;
  assign \new_[6351]_  = ~\new_[6589]_  & ~\new_[1810]_ ;
  assign \new_[6352]_  = \new_[6679]_  ^ \new_[6586]_ ;
  assign \new_[6353]_  = ~\new_[6433]_  & ~\new_[6617]_ ;
  assign \new_[6354]_  = \new_[6433]_  | \new_[6557]_ ;
  assign \new_[6355]_  = \new_[6498]_  ^ \new_[6507]_ ;
  assign \new_[6356]_  = ~\new_[6406]_ ;
  assign \new_[6357]_  = ~\new_[6399]_ ;
  assign \new_[6358]_  = ~\new_[7246]_  | ~\new_[7554]_ ;
  assign \new_[6359]_  = ~\new_[7128]_ ;
  assign \new_[6360]_  = ~\new_[1739]_  | ~\new_[6649]_  | ~\new_[6489]_ ;
  assign \new_[6361]_  = ~\new_[6465]_ ;
  assign \new_[6362]_  = \new_[6467]_  | \new_[6620]_ ;
  assign \new_[6363]_  = ~\new_[6412]_ ;
  assign \new_[6364]_  = ~\new_[6411]_ ;
  assign \new_[6365]_  = ~\new_[7308]_ ;
  assign \new_[6366]_  = ~\new_[6664]_  | ~\new_[6526]_ ;
  assign \new_[6367]_  = ~\new_[6432]_  | ~\new_[6436]_ ;
  assign \new_[6368]_  = ~\new_[6436]_  | ~\new_[6444]_ ;
  assign \new_[6369]_  = ~\new_[6418]_ ;
  assign \new_[6370]_  = ~\new_[6427]_ ;
  assign \new_[6371]_  = ~\new_[6427]_ ;
  assign \new_[6372]_  = ~\new_[6421]_ ;
  assign \new_[6373]_  = ~\new_[1925]_  | ~\new_[6503]_  | ~\new_[6483]_ ;
  assign \new_[6374]_  = ~\new_[7030]_ ;
  assign \new_[6375]_  = ~\new_[6414]_ ;
  assign \new_[6376]_  = ~\new_[6412]_ ;
  assign \new_[6377]_  = \new_[6474]_  & \new_[2554]_ ;
  assign \new_[6378]_  = ~\new_[6637]_  & ~\new_[6519]_ ;
  assign \new_[6379]_  = ~\new_[6649]_  | ~\new_[6454]_  | ~\new_[1739]_ ;
  assign \new_[6380]_  = \new_[2926]_  ^ \new_[6504]_ ;
  assign \new_[6381]_  = \new_[6499]_  & \new_[6608]_ ;
  assign \new_[6382]_  = ~reset_n;
  assign busak_n = ~\new_[6438]_ ;
  assign \new_[6384]_  = \new_[7134]_ ;
  assign \new_[6385]_  = ~\new_[6651]_ ;
  assign \new_[6386]_  = \new_[6502]_  & \new_[6608]_ ;
  assign \new_[6387]_  = ~\new_[6438]_ ;
  assign \new_[6388]_  = ~\new_[6438]_ ;
  assign \new_[6389]_  = \new_[6499]_  & \new_[2550]_ ;
  assign \new_[6390]_  = ~\new_[2007]_  & ~\new_[6647]_ ;
  assign \new_[6391]_  = \new_[7182]_  | \new_[7048]_ ;
  assign \new_[6392]_  = \new_[4559]_  ^ \new_[4553]_ ;
  assign \new_[6393]_  = ~\new_[6441]_ ;
  assign \new_[6394]_  = \new_[6437]_ ;
  assign \new_[6395]_  = ~\new_[2005]_  | ~\new_[6501]_ ;
  assign \new_[6396]_  = ~\new_[6894]_ ;
  assign \new_[6397]_  = ~\new_[6450]_ ;
  assign \new_[6398]_  = ~\new_[7052]_ ;
  assign \new_[6399]_  = ~\new_[6895]_  | ~\new_[7048]_ ;
  assign \new_[6400]_  = ~\new_[6439]_ ;
  assign \new_[6401]_  = \new_[6497]_  | \new_[597]_ ;
  assign \new_[6402]_  = ~reset_n;
  assign \new_[6403]_  = ~reset_n;
  assign \new_[6404]_  = \new_[7182]_  & \new_[7048]_ ;
  assign \new_[6405]_  = ~\new_[6455]_ ;
  assign \new_[6406]_  = ~\new_[6623]_  & ~\new_[6348]_ ;
  assign \new_[6407]_  = ~\new_[7326]_  & ~\new_[7213]_ ;
  assign \new_[6408]_  = \new_[6502]_  & \new_[2550]_ ;
  assign \new_[6409]_  = ~\new_[1892]_  | ~\new_[6503]_  | ~\new_[1925]_ ;
  assign \new_[6410]_  = ~\new_[2135]_  | ~\new_[6513]_ ;
  assign \new_[6411]_  = ~\new_[6495]_  | ~\new_[2660]_ ;
  assign \new_[6412]_  = ~reset_n;
  assign \new_[6413]_  = ~\new_[6481]_ ;
  assign \new_[6414]_  = ~\new_[6812]_  | ~\new_[7365]_ ;
  assign \new_[6415]_  = ~\new_[6470]_ ;
  assign \new_[6416]_  = ~\new_[6462]_ ;
  assign \new_[6417]_  = ~reset_n;
  assign \new_[6418]_  = ~\new_[2665]_  | ~\new_[7253]_ ;
  assign \new_[6419]_  = ~\new_[6452]_ ;
  assign \new_[6420]_  = ~\new_[7072]_ ;
  assign \new_[6421]_  = ~\new_[1610]_  | ~\new_[6505]_  | ~\new_[1646]_ ;
  assign \new_[6422]_  = \new_[6593]_  ^ \new_[6648]_ ;
  assign \new_[6423]_  = ~\new_[6506]_  & ~\new_[6565]_ ;
  assign \new_[6424]_  = ~reset_n;
  assign \new_[6425]_  = ~\new_[7063]_  | ~\new_[6704]_ ;
  assign \new_[6426]_  = \new_[6424]_ ;
  assign \new_[6427]_  = ~\new_[6424]_ ;
  assign \new_[6428]_  = ~\new_[7115]_  & ~\new_[2826]_ ;
  assign \new_[6429]_  = ~\new_[6460]_ ;
  assign \new_[6430]_  = \new_[6663]_  & \new_[6667]_ ;
  assign \new_[6431]_  = \new_[6663]_  ^ \new_[6667]_ ;
  assign \new_[6432]_  = ~\new_[6542]_  & ~\new_[1247]_ ;
  assign \new_[6433]_  = ~\new_[6530]_  | ~\new_[1646]_ ;
  assign \new_[6434]_  = ~\new_[7217]_ ;
  assign \new_[6435]_  = ~\new_[6508]_ ;
  assign \new_[6436]_  = ~\new_[6518]_  | ~\new_[6515]_ ;
  assign \new_[6437]_  = ~\new_[7363]_ ;
  assign \new_[6438]_  = ~\new_[6714]_ ;
  assign \new_[6439]_  = ~\new_[7035]_ ;
  assign \new_[6440]_  = ~\new_[6589]_  & ~\new_[1811]_ ;
  assign \new_[6441]_  = ~\new_[6481]_ ;
  assign \new_[6442]_  = ~\new_[7048]_ ;
  assign \new_[6443]_  = ~\new_[6486]_ ;
  assign \new_[6444]_  = ~\new_[6532]_  & ~\new_[6542]_ ;
  assign \new_[6445]_  = ~\new_[7249]_ ;
  assign \new_[6446]_  = \new_[6608]_  & \new_[6527]_ ;
  assign \new_[6447]_  = ~\new_[1811]_  & ~\new_[6534]_ ;
  assign \new_[6448]_  = ~\new_[6492]_ ;
  assign \new_[6449]_  = \new_[6613]_  ^ \new_[6676]_ ;
  assign \new_[6450]_  = ~\new_[7213]_ ;
  assign \new_[6451]_  = ~\new_[6506]_ ;
  assign \new_[6452]_  = ~\new_[7182]_ ;
  assign \new_[6453]_  = ~\new_[1739]_  & ~\new_[1481]_ ;
  assign \new_[6454]_  = ~\new_[6489]_ ;
  assign \new_[6455]_  = ~\new_[6480]_ ;
  assign \new_[6456]_  = ~\new_[6525]_  & ~\new_[6677]_ ;
  assign \new_[6457]_  = ~\new_[6803]_ ;
  assign \new_[6458]_  = ~\new_[6539]_  & ~\new_[6707]_ ;
  assign \new_[6459]_  = \new_[2550]_  & \new_[6527]_ ;
  assign \new_[6460]_  = \new_[6501]_ ;
  assign \new_[6461]_  = \new_[6484]_ ;
  assign \new_[6462]_  = \new_[6892]_ ;
  assign \new_[6463]_  = ~\new_[6514]_  & ~\new_[6608]_ ;
  assign \new_[6464]_  = ~\new_[6514]_  & ~\new_[2550]_ ;
  assign \new_[6465]_  = ~\new_[7062]_ ;
  assign \new_[6466]_  = \new_[7115]_ ;
  assign \new_[6467]_  = ~\new_[6490]_ ;
  assign \new_[6468]_  = ~\new_[6488]_ ;
  assign \new_[6469]_  = \new_[6679]_  & \new_[6526]_ ;
  assign \new_[6470]_  = ~\new_[7552]_  & ~\new_[6651]_ ;
  assign \new_[6471]_  = ~\new_[6495]_ ;
  assign \new_[6472]_  = ~\new_[6513]_ ;
  assign \new_[6473]_  = ~\new_[6935]_ ;
  assign \new_[6474]_  = \new_[2633]_  & \new_[2661]_ ;
  assign \new_[6475]_  = \new_[2633]_  ^ \new_[2661]_ ;
  assign \new_[6476]_  = \new_[2006]_  ^ \new_[1126]_ ;
  assign \new_[6477]_  = ~\new_[506]_ ;
  assign \new_[6478]_  = ~\new_[6648]_ ;
  assign \new_[6479]_  = \new_[2004]_  & \new_[6647]_ ;
  assign \new_[6480]_  = \new_[1032]_  & \new_[7182]_ ;
  assign \new_[6481]_  = ~\new_[6623]_ ;
  assign \new_[6482]_  = ~\new_[418]_ ;
  assign \new_[6483]_  = ~\new_[6543]_ ;
  assign \new_[6484]_  = ~\new_[7552]_  | ~\new_[6997]_ ;
  assign \new_[6485]_  = \new_[4549]_  ^ \new_[4554]_ ;
  assign \new_[6486]_  = ~\new_[1866]_  & ~\new_[6601]_ ;
  assign \new_[6487]_  = ~\new_[1866]_  | ~\new_[6647]_ ;
  assign \new_[6488]_  = \new_[7299]_  & \new_[7552]_ ;
  assign \new_[6489]_  = ~\new_[6570]_  | ~\new_[6622]_ ;
  assign \new_[6490]_  = ~\new_[1810]_  & ~\new_[6584]_ ;
  assign \new_[6491]_  = ~\new_[505]_ ;
  assign \new_[6492]_  = \new_[6581]_  | \new_[6705]_ ;
  assign \new_[6493]_  = \new_[2007]_  & \new_[6647]_ ;
  assign \new_[6494]_  = \new_[595]_  | \new_[6666]_ ;
  assign \new_[6495]_  = ~\new_[2716]_ ;
  assign \new_[6496]_  = ~\new_[425]_ ;
  assign \new_[6497]_  = ~\new_[595]_  | ~\new_[6666]_ ;
  assign \new_[6498]_  = \new_[4558]_  ^ \new_[4557]_ ;
  assign \new_[6499]_  = ~\new_[6574]_  & ~\new_[4126]_ ;
  assign \new_[6500]_  = ~\new_[7247]_ ;
  assign \new_[6501]_  = ~\new_[6526]_ ;
  assign \new_[6502]_  = \new_[6574]_  & \new_[4126]_ ;
  assign \new_[6503]_  = ~\new_[6525]_ ;
  assign \new_[6504]_  = ~\new_[6895]_ ;
  assign \new_[6505]_  = ~\new_[6646]_  & ~\new_[6557]_ ;
  assign \new_[6506]_  = \new_[6668]_  & \new_[6586]_ ;
  assign \new_[6507]_  = \new_[4560]_  ^ \new_[4556]_ ;
  assign \new_[6508]_  = ~\new_[2666]_  | ~\new_[6621]_ ;
  assign \new_[6509]_  = \new_[2003]_  ^ \new_[1247]_ ;
  assign \new_[6510]_  = \new_[2016]_  ^ \new_[1324]_ ;
  assign \new_[6511]_  = ~\new_[6570]_  & ~\new_[6622]_ ;
  assign \new_[6512]_  = ~\new_[426]_ ;
  assign \new_[6513]_  = ~\new_[751]_ ;
  assign \new_[6514]_  = \new_[2134]_  | \new_[4126]_ ;
  assign \new_[6515]_  = ~\new_[6586]_ ;
  assign \new_[6516]_  = \new_[1379]_  & \new_[1394]_ ;
  assign \new_[6517]_  = ~\new_[595]_  | ~\new_[596]_ ;
  assign \new_[6518]_  = ~\new_[6668]_ ;
  assign \new_[6519]_  = ~\new_[6571]_ ;
  assign \new_[6520]_  = ~\new_[6584]_ ;
  assign \new_[6521]_  = ~\new_[6659]_ ;
  assign \new_[6522]_  = ~\new_[7299]_ ;
  assign \new_[6523]_  = ~\new_[6637]_ ;
  assign \new_[6524]_  = \new_[2555]_  & \new_[2553]_ ;
  assign \new_[6525]_  = ~\new_[2429]_  | ~\new_[2034]_ ;
  assign \new_[6526]_  = ~\new_[6647]_ ;
  assign \new_[6527]_  = \new_[2134]_  & \new_[4126]_ ;
  assign \new_[6528]_  = ~\new_[6593]_ ;
  assign \new_[6529]_  = \new_[1394]_  & \new_[1104]_ ;
  assign \new_[6530]_  = \new_[1610]_  & \new_[1545]_ ;
  assign \new_[6531]_  = ~\new_[4560]_  & ~\new_[4558]_ ;
  assign \new_[6532]_  = \new_[1247]_  | \new_[1126]_ ;
  assign \new_[6533]_  = ~\new_[7216]_ ;
  assign \new_[6534]_  = ~\new_[1810]_ ;
  assign \new_[6535]_  = ~\new_[1892]_ ;
  assign \new_[6536]_  = ~\new_[1248]_ ;
  assign \new_[6537]_  = ~\new_[774]_ ;
  assign \new_[6538]_  = ~\new_[1126]_  | ~\new_[1248]_ ;
  assign \new_[6539]_  = \new_[595]_  | \new_[596]_ ;
  assign \new_[6540]_  = ~\new_[4549]_  & ~\new_[4556]_ ;
  assign \new_[6541]_  = ~\new_[4557]_  & ~\new_[4553]_ ;
  assign \new_[6542]_  = ~\new_[6565]_ ;
  assign \new_[6543]_  = ~\new_[1892]_  | ~\new_[1861]_ ;
  assign \new_[6544]_  = \new_[2554]_  & \new_[2553]_ ;
  assign \new_[6545]_  = ~\new_[785]_ ;
  assign \new_[6546]_  = ~\new_[6614]_ ;
  assign \new_[6547]_  = ~\new_[6588]_ ;
  assign \new_[6548]_  = ~\new_[6679]_ ;
  assign \new_[6549]_  = ~\new_[775]_ ;
  assign \new_[6550]_  = ~\new_[1646]_ ;
  assign \new_[6551]_  = ~\new_[1692]_ ;
  assign \new_[6552]_  = ~\new_[1863]_ ;
  assign \new_[6553]_  = ~\new_[560]_ ;
  assign \new_[6554]_  = ~\new_[3281]_ ;
  assign \new_[6555]_  = ~\new_[579]_ ;
  assign \new_[6556]_  = ~\new_[467]_ ;
  assign \new_[6557]_  = ~\new_[1578]_ ;
  assign \new_[6558]_  = ~\new_[1581]_ ;
  assign \new_[6559]_  = ~\new_[417]_ ;
  assign \new_[6560]_  = ~\new_[1860]_ ;
  assign \new_[6561]_  = ~\new_[776]_ ;
  assign \new_[6563]_  = ~\new_[686]_ ;
  assign \new_[6564]_  = ~\new_[414]_ ;
  assign \new_[6565]_  = ~\new_[1231]_ ;
  assign \new_[6566]_  = ~\new_[465]_ ;
  assign \new_[6567]_  = ~\new_[2664]_ ;
  assign \new_[6568]_  = ~\new_[3626]_ ;
  assign \new_[6569]_  = ~\new_[1787]_ ;
  assign \new_[6570]_  = ~\new_[1621]_ ;
  assign \new_[6571]_  = ~\new_[1124]_ ;
  assign \new_[6572]_  = ~\new_[4559]_ ;
  assign \new_[6573]_  = ~\new_[1809]_ ;
  assign \new_[6574]_  = ~\new_[2134]_ ;
  assign \new_[6575]_  = ~\new_[3603]_ ;
  assign \new_[6576]_  = ~\new_[1862]_ ;
  assign \new_[6577]_  = ~\new_[3029]_ ;
  assign \new_[6578]_  = ~\new_[3638]_ ;
  assign \new_[6580]_  = ~\new_[1337]_ ;
  assign \new_[6581]_  = ~\new_[2727]_ ;
  assign \new_[6582]_  = ~\new_[3639]_ ;
  assign \new_[6583]_  = ~\new_[508]_ ;
  assign \new_[6584]_  = ~\new_[752]_ ;
  assign \new_[6586]_  = ~\new_[1338]_ ;
  assign \new_[6587]_  = ~\new_[424]_ ;
  assign \new_[6588]_  = ~\new_[537]_ ;
  assign \new_[6589]_  = ~\new_[1624]_ ;
  assign \new_[6590]_  = ~\new_[413]_ ;
  assign \new_[6591]_  = ~\new_[847]_ ;
  assign \new_[6592]_  = ~\new_[1236]_ ;
  assign \new_[6593]_  = ~\new_[1866]_ ;
  assign \new_[6595]_  = ~\new_[1580]_ ;
  assign \new_[6596]_  = ~\new_[1808]_ ;
  assign \new_[6597]_  = ~\new_[511]_ ;
  assign \new_[6598]_  = ~\new_[412]_ ;
  assign \new_[6599]_  = ~\new_[416]_ ;
  assign \new_[6600]_  = ~\new_[787]_ ;
  assign \new_[6601]_  = ~\new_[1622]_ ;
  assign \new_[6602]_  = \new_[685]_ ;
  assign \new_[6603]_  = ~\new_[3321]_ ;
  assign \new_[6604]_  = ~\new_[3600]_ ;
  assign \new_[6605]_  = ~\new_[1865]_ ;
  assign \new_[6606]_  = ~\new_[846]_ ;
  assign \new_[6607]_  = ~\new_[512]_ ;
  assign \new_[6608]_  = ~\new_[2550]_ ;
  assign \new_[6609]_  = ~\new_[731]_ ;
  assign \new_[6610]_  = ~\new_[786]_ ;
  assign \new_[6611]_  = ~\new_[577]_ ;
  assign \new_[6612]_  = ~\new_[510]_ ;
  assign \new_[6613]_  = ~\new_[2429]_ ;
  assign \new_[6614]_  = ~\new_[562]_ ;
  assign \new_[6615]_  = ~\new_[507]_ ;
  assign \new_[6616]_  = ~\new_[1052]_ ;
  assign \new_[6617]_  = ~\new_[1308]_ ;
  assign \new_[6618]_  = ~\new_[506]_ ;
  assign \new_[6619]_  = ~nmi_n;
  assign \new_[6620]_  = ~\new_[1811]_ ;
  assign \new_[6621]_  = ~\new_[2662]_ ;
  assign \new_[6622]_  = ~\new_[1579]_ ;
  assign \new_[6623]_  = ~reset_n;
  assign \new_[6624]_  = ~\new_[1909]_ ;
  assign \new_[6625]_  = ~\new_[740]_ ;
  assign \new_[6626]_  = ~\new_[3615]_ ;
  assign \new_[6627]_  = ~\new_[421]_ ;
  assign \new_[6629]_  = ~\new_[1292]_ ;
  assign \new_[6630]_  = ~\new_[733]_ ;
  assign \new_[6631]_  = ~\new_[1293]_ ;
  assign \new_[6632]_  = ~halt_n;
  assign \new_[6633]_  = ~\new_[420]_ ;
  assign \new_[6634]_  = ~\new_[1620]_ ;
  assign \new_[6635]_  = ~\new_[1110]_ ;
  assign \new_[6637]_  = ~\new_[1123]_ ;
  assign \new_[6638]_  = ~\new_[575]_ ;
  assign \new_[6639]_  = ~\new_[509]_ ;
  assign \new_[6640]_  = ~\new_[2660]_ ;
  assign \new_[6641]_  = ~\new_[423]_ ;
  assign \new_[6642]_  = ~\new_[466]_ ;
  assign \new_[6643]_  = ~\new_[1691]_ ;
  assign \new_[6644]_  = ~\new_[464]_ ;
  assign \new_[6645]_  = ~\new_[422]_ ;
  assign \new_[6646]_  = ~\new_[1689]_ ;
  assign \new_[6647]_  = ~\new_[1622]_ ;
  assign \new_[6648]_  = ~\new_[1125]_ ;
  assign \new_[6649]_  = ~\new_[1481]_ ;
  assign \new_[6651]_  = ~\new_[2666]_ ;
  assign \new_[6652]_  = ~\new_[419]_ ;
  assign \new_[6653]_  = ~\new_[3621]_ ;
  assign \new_[6654]_  = ~\new_[2007]_ ;
  assign \new_[6655]_  = ~\new_[3841]_ ;
  assign \new_[6656]_  = ~\new_[1647]_ ;
  assign \new_[6657]_  = ~\new_[468]_ ;
  assign \new_[6658]_  = ~\new_[1864]_ ;
  assign \new_[6659]_  = ~\new_[651]_ ;
  assign \new_[6660]_  = ~\new_[415]_ ;
  assign \new_[6661]_  = ~\new_[1861]_ ;
  assign \new_[6662]_  = ~\new_[3606]_ ;
  assign \new_[6663]_  = ~\new_[1244]_ ;
  assign \new_[6664]_  = ~\new_[2005]_ ;
  assign \new_[6665]_  = ~\new_[427]_ ;
  assign \new_[6666]_  = ~\new_[596]_ ;
  assign \new_[6667]_  = ~\new_[1245]_ ;
  assign \new_[6668]_  = ~\new_[1246]_ ;
  assign \new_[6669]_  = ~\new_[3002]_ ;
  assign \new_[6670]_  = ~\new_[2826]_ ;
  assign \new_[6671]_  = ~\new_[1693]_ ;
  assign \new_[6672]_  = ~\new_[470]_ ;
  assign \new_[6673]_  = ~\new_[469]_ ;
  assign \new_[6674]_  = ~\new_[1228]_ ;
  assign \new_[6675]_  = ~\new_[1111]_ ;
  assign \new_[6676]_  = ~\new_[2034]_ ;
  assign \new_[6677]_  = ~\new_[1925]_ ;
  assign \new_[6678]_  = ~\new_[1908]_ ;
  assign \new_[6679]_  = ~\new_[2004]_ ;
  assign \new_[6680]_  = \new_[6681]_ ;
  assign \new_[6681]_  = \new_[2121]_ ;
  assign \new_[6682]_  = ~\new_[6683]_ ;
  assign \new_[6683]_  = ~\new_[7460]_ ;
  assign \new_[6684]_  = ~\new_[6975]_ ;
  assign \new_[6685]_  = ~\new_[6686]_ ;
  assign \new_[6686]_  = \new_[7394]_ ;
  assign \new_[6687]_  = ~\new_[6688]_ ;
  assign \new_[6688]_  = ~\new_[7078]_ ;
  assign \new_[6689]_  = \new_[2448]_ ;
  assign \new_[6690]_  = \new_[6691]_ ;
  assign \new_[6691]_  = \new_[2039]_ ;
  assign \new_[6692]_  = ~\new_[2039]_ ;
  assign \new_[6693]_  = \new_[2064]_ ;
  assign \new_[6694]_  = \new_[2066]_ ;
  assign \new_[6695]_  = \new_[1574]_ ;
  assign \new_[6696]_  = ~\new_[6697]_  | ~\new_[2780]_ ;
  assign \new_[6697]_  = \new_[6698]_ ;
  assign \new_[6698]_  = ~\new_[7268]_ ;
  assign \new_[6699]_  = ~\new_[3305]_  | ~\new_[6700]_ ;
  assign \new_[6700]_  = \new_[7266]_  & \new_[3029]_ ;
  assign \new_[6701]_  = ~\new_[4482]_  | ~\new_[3304]_  | ~\new_[3362]_ ;
  assign \new_[6702]_  = ~\new_[6927]_  | ~\new_[6703]_ ;
  assign \new_[6703]_  = \new_[6495]_  | \new_[5028]_ ;
  assign \new_[6704]_  = ~\new_[7322]_ ;
  assign \new_[6705]_  = ~\new_[2779]_ ;
  assign \new_[6706]_  = \new_[7194]_ ;
  assign \new_[6707]_  = ~\new_[597]_ ;
  assign \new_[6708]_  = ~\new_[6715]_  | (~\new_[6709]_  & ~\new_[6710]_ );
  assign \new_[6709]_  = (~\new_[5724]_  | ~\new_[2106]_ ) & (~\new_[1850]_  | ~\new_[6156]_ );
  assign \new_[6710]_  = ~\new_[6711]_  | ~\new_[6714]_ ;
  assign \new_[6711]_  = ~\new_[6712]_ ;
  assign \new_[6712]_  = \new_[6713]_ ;
  assign \new_[6713]_  = ~\new_[597]_  & ~\new_[7209]_ ;
  assign \new_[6714]_  = ~\new_[1690]_ ;
  assign \new_[6715]_  = \new_[1235]_  ? \new_[6714]_  : \new_[6716]_ ;
  assign \new_[6716]_  = ~\new_[2323]_  | ~\new_[6712]_ ;
  assign \new_[6717]_  = ~\new_[6718]_ ;
  assign \new_[6718]_  = \new_[6458]_  & \new_[7208]_ ;
  assign \new_[6719]_  = ~\new_[684]_  & ~\new_[6156]_ ;
  assign \new_[6720]_  = (~\new_[3509]_  | ~\new_[2136]_ ) & (~\new_[6721]_  | ~\new_[684]_ );
  assign \new_[6721]_  = \new_[3563]_  | \new_[6722]_ ;
  assign \new_[6722]_  = ~\new_[6156]_  & ~\new_[6718]_ ;
  assign \new_[6723]_  = \new_[6722]_ ;
  assign \new_[6724]_  = \new_[6725]_  & \new_[6726]_ ;
  assign \new_[6725]_  = ~\new_[6825]_  & ~\new_[6826]_ ;
  assign \new_[6726]_  = ~\new_[7539]_ ;
  assign \new_[6727]_  = \new_[6728]_  & \new_[6041]_ ;
  assign \new_[6728]_  = \new_[6895]_  | \new_[6729]_ ;
  assign \new_[6729]_  = \new_[6391]_  | \new_[6272]_ ;
  assign \new_[6730]_  = ~\new_[6391]_  & ~\new_[6895]_ ;
  assign \new_[6731]_  = ~\new_[7502]_ ;
  assign \new_[6732]_  = ~\new_[6733]_  & ~\new_[7111]_ ;
  assign \new_[6733]_  = ~\new_[6734]_  | ~\new_[7331]_ ;
  assign \new_[6734]_  = ~\new_[1887]_  | ~\new_[7332]_ ;
  assign \new_[6735]_  = ~\new_[7482]_ ;
  assign \new_[6736]_  = ~\new_[7110]_  | ~\new_[7112]_ ;
  assign \new_[6737]_  = ~\new_[7107]_  | ~\new_[7331]_ ;
  assign \new_[6738]_  = ~\new_[6734]_ ;
  assign \new_[6739]_  = \new_[6738]_  ^ \new_[7104]_ ;
  assign \new_[6745]_  = ~\new_[7501]_ ;
  assign \new_[6747]_  = \new_[4137]_  | \new_[4068]_ ;
  assign \new_[6753]_  = ~\new_[1691]_  & ~\new_[5184]_ ;
  assign \new_[6754]_  = ~\new_[7468]_  | ~\new_[7464]_ ;
  assign n159 = ~\new_[6758]_  | (~\new_[6756]_  & ~\new_[6757]_ );
  assign \new_[6756]_  = ~\new_[7397]_  & ~\new_[6769]_ ;
  assign \new_[6757]_  = ~\new_[7515]_  | (~\new_[7398]_  & ~\new_[6633]_ );
  assign \new_[6758]_  = ~\new_[1187]_  | ~\new_[6633]_ ;
  assign n184 = ~\new_[6762]_  | (~\new_[6760]_  & ~\new_[6761]_ );
  assign \new_[6760]_  = ~\new_[7432]_  & ~\new_[6769]_ ;
  assign \new_[6761]_  = ~\new_[7515]_  | (~\new_[7426]_  & ~\new_[6496]_ );
  assign \new_[6762]_  = ~\new_[1183]_  | ~\new_[6496]_ ;
  assign n169 = ~\new_[6766]_  | (~\new_[6764]_  & ~\new_[6765]_ );
  assign \new_[6764]_  = ~\new_[6830]_  & ~\new_[6769]_ ;
  assign \new_[6765]_  = ~\new_[7515]_  | (~\new_[7389]_  & ~\new_[6645]_ );
  assign \new_[6766]_  = ~\new_[1183]_  | ~\new_[6645]_ ;
  assign n189 = ~\new_[6772]_  | (~\new_[6768]_  & ~\new_[6771]_ );
  assign \new_[6768]_  = ~\new_[6853]_  & ~\new_[6769]_ ;
  assign \new_[6769]_  = ~\new_[6770]_ ;
  assign \new_[6770]_  = ~\new_[6773]_ ;
  assign \new_[6771]_  = ~\new_[7515]_  | (~\new_[7514]_  & ~\new_[6512]_ );
  assign \new_[6772]_  = ~\new_[1183]_  | ~\new_[6512]_ ;
  assign \new_[6773]_  = ~\new_[6779]_  | ~\new_[6774]_  | ~\new_[6777]_ ;
  assign \new_[6774]_  = ~\new_[6775]_  | ~\new_[7469]_ ;
  assign \new_[6775]_  = ~\new_[6776]_ ;
  assign \new_[6776]_  = ~\new_[7501]_  | ~\new_[3571]_  | ~\new_[5184]_ ;
  assign \new_[6777]_  = ~\new_[6778]_  | ~\new_[7501]_ ;
  assign \new_[6778]_  = ~\new_[2897]_  | ~\new_[4613]_ ;
  assign \new_[6779]_  = ~\new_[3934]_  | ~\new_[7466]_ ;
  assign \new_[6780]_  = ~\new_[6375]_  | ~\new_[6513]_ ;
  assign \new_[6781]_  = ~\new_[751]_  | ~\new_[6398]_  | ~\new_[6815]_ ;
  assign \new_[6782]_  = \new_[6398]_  & \new_[6815]_ ;
  assign \new_[6783]_  = ~\new_[7440]_  & (~\new_[6784]_  | ~\new_[6785]_ );
  assign \new_[6784]_  = ~\new_[5223]_  | ~\new_[1510]_  | ~\new_[6796]_ ;
  assign \new_[6785]_  = \new_[6786]_  & \new_[6787]_ ;
  assign \new_[6786]_  = ~\new_[6796]_  | (~\new_[4952]_  & ~\new_[6792]_ );
  assign \new_[6787]_  = ~\new_[7174]_  | ~\new_[1925]_ ;
  assign \new_[6788]_  = ~\new_[7440]_  & (~\new_[6789]_  | ~\new_[6790]_ );
  assign \new_[6789]_  = ~\new_[5223]_  | ~\new_[1513]_  | ~\new_[6796]_ ;
  assign \new_[6790]_  = \new_[6791]_  & \new_[6793]_ ;
  assign \new_[6791]_  = ~\new_[6796]_  | (~\new_[4953]_  & ~\new_[6792]_ );
  assign \new_[6792]_  = ~\new_[7171]_ ;
  assign \new_[6793]_  = ~\new_[7174]_  | ~\new_[1689]_ ;
  assign \new_[6794]_  = ~\new_[7440]_  & (~\new_[6795]_  | ~\new_[6797]_ );
  assign \new_[6795]_  = ~\new_[5223]_  | ~\new_[1514]_  | ~\new_[6796]_ ;
  assign \new_[6796]_  = ~\new_[7174]_ ;
  assign \new_[6797]_  = \new_[6798]_  & \new_[6799]_ ;
  assign \new_[6798]_  = ~\new_[6796]_  | (~\new_[4984]_  & ~\new_[6792]_ );
  assign \new_[6799]_  = ~\new_[7174]_  | ~\new_[1578]_ ;
  assign \new_[6800]_  = ~\new_[6801]_  | ~\new_[6802]_ ;
  assign \new_[6801]_  = ~\new_[7027]_ ;
  assign \new_[6802]_  = \new_[7047]_  & \new_[6803]_ ;
  assign \new_[6803]_  = ~\new_[6571]_  | ~\new_[6637]_ ;
  assign \new_[6804]_  = ~\new_[7031]_  | ~\new_[7030]_ ;
  assign \new_[6805]_  = ~\new_[7440]_  & (~\new_[6806]_  | ~\new_[6807]_ );
  assign \new_[6806]_  = ~\new_[5223]_  | ~\new_[1509]_  | ~\new_[6796]_ ;
  assign \new_[6807]_  = \new_[6808]_  & \new_[6809]_ ;
  assign \new_[6808]_  = ~\new_[6796]_  | (~\new_[4949]_  & ~\new_[6792]_ );
  assign \new_[6809]_  = ~\new_[7174]_  | ~\new_[2034]_ ;
  assign \new_[6810]_  = ~\new_[7073]_ ;
  assign \new_[6811]_  = \new_[6812]_  & \new_[2664]_ ;
  assign \new_[6812]_  = ~\new_[2727]_  & ~\new_[2779]_ ;
  assign \new_[6813]_  = ~\new_[651]_  | ~\new_[7051]_ ;
  assign \new_[6814]_  = ~\new_[6584]_  | ~\new_[7558]_  | ~\new_[6815]_ ;
  assign \new_[6815]_  = \new_[7365]_ ;
  assign \new_[6816]_  = ~\new_[6328]_  | ~\new_[844]_ ;
  assign \new_[6817]_  = ~\new_[752]_  | ~\new_[6448]_  | ~\new_[6815]_ ;
  assign \new_[6818]_  = ~\new_[6819]_  | ~\new_[752]_ ;
  assign \new_[6819]_  = \new_[6448]_  & \new_[6815]_ ;
  assign \new_[6820]_  = \new_[2842]_  & \new_[7540]_ ;
  assign \new_[6821]_  = ~\new_[6822]_  | ~\new_[6824]_ ;
  assign \new_[6822]_  = ~\new_[6823]_ ;
  assign \new_[6823]_  = ~\new_[5052]_  & (~\new_[6041]_  | ~\new_[3560]_ );
  assign \new_[6824]_  = ~\new_[6825]_ ;
  assign \new_[6825]_  = ~\new_[6272]_  & ~\new_[6216]_ ;
  assign \new_[6826]_  = ~\new_[5052]_  & (~\new_[3560]_  | ~\new_[6041]_ );
  assign \new_[6827]_  = ~\new_[595]_ ;
  assign n129 = ~\new_[6832]_  | (~\new_[6829]_  & ~\new_[6831]_ );
  assign \new_[6829]_  = ~\new_[6830]_  & ~\new_[6847]_ ;
  assign \new_[6830]_  = ~\new_[7389]_ ;
  assign \new_[6831]_  = ~\new_[7515]_  | (~\new_[7389]_  & ~\new_[6564]_ );
  assign \new_[6832]_  = ~\new_[1192]_  | ~\new_[6564]_ ;
  assign n144 = ~\new_[6836]_  | (~\new_[6834]_  & ~\new_[6835]_ );
  assign \new_[6834]_  = ~\new_[6847]_  & ~\new_[7432]_ ;
  assign \new_[6835]_  = ~\new_[7515]_  | (~\new_[7426]_  & ~\new_[6559]_ );
  assign \new_[6836]_  = ~\new_[1185]_  | ~\new_[6559]_ ;
  assign \new_[6837]_  = ~\new_[6839]_  | (~\new_[1356]_  & ~\new_[6838]_ );
  assign \new_[6838]_  = ~\new_[1635]_  | (~\new_[1407]_  & ~\new_[1703]_ );
  assign \new_[6839]_  = ~\new_[6840]_ ;
  assign \new_[6840]_  = \new_[7535]_  & \new_[7331]_ ;
  assign \new_[6841]_  = \new_[6842]_  & \new_[6840]_ ;
  assign \new_[6842]_  = ~\new_[1704]_  | ~\new_[1639]_  | ~\new_[1472]_ ;
  assign \new_[6843]_  = ~\new_[6838]_ ;
  assign n124 = ~\new_[6849]_  | (~\new_[6845]_  & ~\new_[6848]_ );
  assign \new_[6845]_  = ~\new_[6846]_  & ~\new_[6847]_ ;
  assign \new_[6846]_  = ~\new_[7383]_ ;
  assign \new_[6847]_  = ~\new_[6852]_ ;
  assign \new_[6848]_  = ~\new_[7515]_  | (~\new_[7383]_  & ~\new_[6590]_ );
  assign \new_[6849]_  = ~\new_[1185]_  | ~\new_[6590]_ ;
  assign n149 = ~\new_[6855]_  | (~\new_[6851]_  & ~\new_[6854]_ );
  assign \new_[6851]_  = ~\new_[6847]_  & ~\new_[6853]_ ;
  assign \new_[6852]_  = ~\new_[6882]_ ;
  assign \new_[6853]_  = ~\new_[7514]_ ;
  assign \new_[6854]_  = ~\new_[7515]_  | (~\new_[7514]_  & ~\new_[6482]_ );
  assign \new_[6855]_  = ~\new_[1184]_  | ~\new_[6482]_ ;
  assign \new_[6856]_  = ~\new_[7515]_ ;
  assign n204 = ~\new_[6860]_  | (~\new_[6858]_  & ~\new_[6859]_ );
  assign \new_[6858]_  = ~\new_[7382]_  & ~\new_[6910]_ ;
  assign \new_[6859]_  = ~\new_[7515]_  | (~\new_[7383]_  & ~\new_[429]_ );
  assign \new_[6860]_  = ~\new_[1185]_  | ~\new_[429]_ ;
  assign n544 = ~\new_[6862]_  | ~\new_[6867]_ ;
  assign \new_[6862]_  = ~\new_[6866]_  | ~\new_[6863]_  | ~\new_[7515]_ ;
  assign \new_[6863]_  = ~\new_[6864]_  | ~\new_[7398]_  | ~\new_[3767]_ ;
  assign \new_[6864]_  = ~\new_[6865]_  | ~\new_[7501]_ ;
  assign \new_[6865]_  = ~\new_[1113]_ ;
  assign \new_[6866]_  = \new_[574]_  | \new_[7398]_ ;
  assign \new_[6867]_  = ~\new_[1187]_  | ~\new_[574]_ ;
  assign \new_[6868]_  = ~\new_[6864]_  | ~\new_[3767]_ ;
  assign n229 = ~\new_[6872]_  | (~\new_[6870]_  & ~\new_[6871]_ );
  assign \new_[6870]_  = ~\new_[7419]_  & ~\new_[6910]_ ;
  assign \new_[6871]_  = ~\new_[7515]_  | (~\new_[7514]_  & ~\new_[434]_ );
  assign \new_[6872]_  = ~\new_[1185]_  | ~\new_[434]_ ;
  assign \new_[6873]_  = \new_[6874]_ ;
  assign \new_[6874]_  = ~\new_[6876]_  | ~\new_[6944]_  | ~\new_[6875]_ ;
  assign \new_[6875]_  = ~\new_[2016]_  | ~\new_[5930]_  | ~\new_[1324]_ ;
  assign \new_[6876]_  = (~\new_[6510]_  | ~\new_[5959]_ ) & (~\new_[6037]_  | ~\new_[6877]_ );
  assign \new_[6877]_  = \new_[2016]_  | \new_[1324]_ ;
  assign n209 = ~\new_[6881]_  | (~\new_[6879]_  & ~\new_[6880]_ );
  assign \new_[6879]_  = ~\new_[2711]_  & ~\new_[6910]_ ;
  assign \new_[6880]_  = ~\new_[7515]_  | (~\new_[7389]_  & ~\new_[430]_ );
  assign \new_[6881]_  = ~\new_[1192]_  | ~\new_[430]_ ;
  assign \new_[6882]_  = ~\new_[6888]_  | ~\new_[6883]_  | ~\new_[6887]_ ;
  assign \new_[6883]_  = ~\new_[7501]_  | ~\new_[6886]_  | ~\new_[6885]_  | ~\new_[6884]_ ;
  assign \new_[6884]_  = ~\new_[7109]_  | ~\new_[6732]_ ;
  assign \new_[6885]_  = ~\new_[6738]_  | (~\new_[6736]_  & ~\new_[6737]_ );
  assign \new_[6886]_  = ~\new_[6735]_ ;
  assign \new_[6887]_  = ~\new_[7501]_  | (~\new_[2720]_  & ~\new_[4530]_ );
  assign \new_[6888]_  = ~\new_[3944]_  | ~\new_[7466]_ ;
  assign \new_[6889]_  = \new_[6080]_  | \new_[7209]_  | \new_[6890]_  | \new_[6420]_ ;
  assign \new_[6890]_  = ~\new_[6891]_  | ~\new_[6892]_ ;
  assign \new_[6891]_  = ~\new_[7049]_ ;
  assign \new_[6892]_  = ~\new_[6567]_  & ~\new_[7364]_ ;
  assign \new_[6893]_  = \new_[1032]_  | \new_[6616]_ ;
  assign \new_[6894]_  = ~\new_[6616]_  & ~\new_[6452]_ ;
  assign \new_[6895]_  = ~\new_[1032]_ ;
  assign n344 = ~\new_[6902]_  | (~\new_[6897]_  & ~\new_[6901]_ );
  assign \new_[6897]_  = ~\new_[6898]_  & ~\new_[6899]_ ;
  assign \new_[6898]_  = \new_[7382]_  | \new_[6972]_ ;
  assign \new_[6899]_  = ~\new_[6900]_ ;
  assign \new_[6900]_  = ~\new_[7086]_ ;
  assign \new_[6901]_  = ~\new_[7515]_  | (~\new_[7383]_  & ~\new_[6566]_ );
  assign \new_[6902]_  = ~\new_[1192]_  | ~\new_[6566]_ ;
  assign \new_[6903]_  = ~\new_[7515]_ ;
  assign \new_[6904]_  = ~\new_[6972]_ ;
  assign n224 = ~\new_[6909]_  | (~\new_[6906]_  & ~\new_[6908]_ );
  assign \new_[6906]_  = ~\new_[6910]_  & ~\new_[6907]_ ;
  assign \new_[6907]_  = ~\new_[7426]_ ;
  assign \new_[6908]_  = ~\new_[7515]_  | (~\new_[7426]_  & ~\new_[433]_ );
  assign \new_[6909]_  = ~\new_[1182]_  | ~\new_[433]_ ;
  assign \new_[6910]_  = ~\new_[7461]_  | ~\new_[6911]_ ;
  assign \new_[6911]_  = (~\new_[7466]_  | ~\new_[3938]_ ) & (~\new_[6912]_  | ~\new_[7501]_ );
  assign \new_[6912]_  = \new_[6753]_  | \new_[3231]_ ;
  assign \new_[6913]_  = ~\new_[6915]_  | (~\new_[6133]_  & ~\new_[6914]_ );
  assign \new_[6914]_  = ~\new_[6920]_ ;
  assign \new_[6915]_  = ~\new_[7145]_  | ~\new_[6919]_ ;
  assign \new_[6916]_  = ~\new_[7122]_ ;
  assign \new_[6917]_  = ~\new_[7181]_ ;
  assign \new_[6918]_  = ~\new_[7123]_  | ~\new_[7125]_ ;
  assign \new_[6919]_  = ~\new_[7012]_  & ~\new_[7011]_ ;
  assign \new_[6920]_  = ~\new_[7128]_ ;
  assign \new_[6921]_  = ~\new_[6924]_  | (~\new_[6922]_  & ~\new_[2143]_ );
  assign \new_[6922]_  = \new_[7335]_  | \new_[6923]_ ;
  assign \new_[6923]_  = \new_[6723]_  & \new_[845]_ ;
  assign \new_[6924]_  = \new_[6925]_  | \new_[5682]_ ;
  assign \new_[6925]_  = \new_[6231]_  | \new_[6926]_ ;
  assign \new_[6926]_  = ~\new_[6181]_  | ~\new_[6249]_  | ~\new_[6291]_  | ~\new_[6198]_ ;
  assign \new_[6927]_  = ~\new_[6928]_  | ~\new_[6934]_ ;
  assign \new_[6928]_  = ~\new_[6933]_  | ~\new_[6929]_  | ~\new_[7143]_ ;
  assign \new_[6929]_  = ~\new_[6930]_ ;
  assign \new_[6930]_  = ~\new_[5375]_  | ~\new_[7565]_ ;
  assign \new_[6931]_  = ~\new_[5921]_  | ~\new_[6022]_ ;
  assign \new_[6932]_  = ~\new_[6980]_ ;
  assign \new_[6933]_  = ~\new_[5740]_  | ~\new_[6284]_ ;
  assign \new_[6934]_  = ~\new_[6935]_ ;
  assign \new_[6935]_  = ~\new_[6495]_  | ~\new_[6640]_ ;
  assign \new_[6936]_  = ~\new_[6980]_  & ~\new_[7147]_ ;
  assign \new_[6937]_  = \new_[6931]_ ;
  assign \new_[6938]_  = ~\new_[6939]_  & ~\new_[6941]_ ;
  assign \new_[6939]_  = \new_[7335]_  & \new_[6940]_ ;
  assign \new_[6940]_  = ~\new_[6242]_  | ~\new_[6269]_  | ~\new_[6247]_  | ~\new_[6196]_ ;
  assign \new_[6941]_  = ~\new_[6942]_  & ~\new_[6720]_ ;
  assign \new_[6942]_  = ~\new_[6943]_ ;
  assign \new_[6943]_  = ~\new_[7335]_  & (~\new_[6717]_  | ~\new_[6719]_ );
  assign \new_[6944]_  = ~\new_[6954]_  | (~\new_[6945]_  & ~\new_[6948]_ );
  assign \new_[6945]_  = ~\new_[6946]_ ;
  assign \new_[6946]_  = ~\new_[6947]_ ;
  assign \new_[6947]_  = ~\new_[3987]_ ;
  assign \new_[6948]_  = ~\new_[6950]_  & (~\new_[5383]_  | ~\new_[7293]_ );
  assign \new_[6949]_  = ~\new_[5965]_  | ~\new_[1324]_ ;
  assign \new_[6950]_  = ~\new_[6951]_  | (~\new_[5383]_  & ~\new_[7293]_ );
  assign \new_[6951]_  = \new_[6952]_  | \new_[6953]_ ;
  assign \new_[6952]_  = ~\new_[1810]_  & ~\new_[6429]_ ;
  assign \new_[6953]_  = ~\new_[6447]_  & ~\new_[6460]_ ;
  assign \new_[6954]_  = \new_[6955]_  | \new_[6946]_ ;
  assign \new_[6955]_  = ~\new_[6956]_  & (~\new_[5263]_  | ~\new_[7293]_ );
  assign \new_[6956]_  = ~\new_[6951]_  | (~\new_[5263]_  & ~\new_[7293]_ );
  assign \new_[6957]_  = ~\new_[5263]_ ;
  assign \new_[6958]_  = ~\new_[5383]_  & ~\new_[6947]_ ;
  assign \new_[6959]_  = \new_[7552]_  | \new_[7321]_ ;
  assign \new_[6960]_  = ~\new_[7179]_  | ~\new_[7178]_ ;
  assign \new_[6961]_  = \new_[6962]_ ;
  assign \new_[6962]_  = \new_[6963]_  & \new_[6968]_ ;
  assign \new_[6963]_  = ~\new_[6964]_ ;
  assign \new_[6964]_  = ~\new_[6965]_  | ~\new_[6967]_ ;
  assign \new_[6965]_  = ~\new_[6966]_ ;
  assign \new_[6966]_  = ~\new_[7254]_  | ~\new_[7035]_ ;
  assign \new_[6967]_  = ~\new_[7299]_  & ~\new_[7319]_ ;
  assign \new_[6968]_  = ~\new_[7246]_  & ~\new_[6166]_ ;
  assign \new_[6969]_  = ~\new_[6968]_ ;
  assign \new_[6970]_  = ~\new_[3942]_  | ~\new_[7466]_ ;
  assign \new_[6971]_  = ~\new_[7088]_  | ~\new_[7501]_ ;
  assign \new_[6972]_  = ~\new_[6970]_ ;
  assign \new_[6973]_  = ~\new_[6979]_  | ~\new_[6974]_  | ~\new_[6978]_ ;
  assign \new_[6974]_  = (~\new_[6627]_  | ~\new_[2706]_ ) & (~\new_[6975]_  | ~\new_[6512]_ );
  assign \new_[6975]_  = \new_[6976]_ ;
  assign \new_[6976]_  = \new_[6977]_ ;
  assign \new_[6977]_  = ~\new_[7460]_ ;
  assign \new_[6978]_  = ~\new_[7489]_  | ~\new_[6633]_ ;
  assign \new_[6979]_  = ~\new_[7442]_  | ~\new_[6496]_ ;
  assign \new_[6980]_  = ~\new_[6981]_  & ~\new_[6982]_ ;
  assign \new_[6981]_  = \new_[7191]_ ;
  assign \new_[6982]_  = ~\new_[7066]_  | ~\new_[6984]_  | ~\new_[7320]_  | ~\new_[6983]_ ;
  assign \new_[6983]_  = ~\new_[6500]_ ;
  assign \new_[6984]_  = ~\new_[6484]_ ;
  assign \new_[6985]_  = ~\new_[6983]_  | ~\new_[6984]_ ;
  assign \new_[6986]_  = ~\new_[7231]_  | ~\new_[6987]_  | ~\new_[6989]_ ;
  assign \new_[6987]_  = ~\new_[7062]_  & ~\new_[6988]_ ;
  assign \new_[6988]_  = \new_[7035]_  | \new_[6651]_ ;
  assign \new_[6989]_  = ~\new_[7241]_ ;
  assign \new_[6990]_  = ~\new_[6991]_  | ~\new_[2716]_ ;
  assign \new_[6991]_  = ~\new_[5398]_  | ~\new_[6992]_ ;
  assign \new_[6992]_  = \new_[5389]_  & \new_[5932]_ ;
  assign \new_[6993]_  = ~\new_[6473]_  | (~\new_[5031]_  & ~\new_[4445]_ );
  assign \new_[6994]_  = \new_[7301]_ ;
  assign \new_[6995]_  = ~\new_[7169]_  & ~\new_[6996]_ ;
  assign \new_[6996]_  = \new_[7552]_  | \new_[6508]_ ;
  assign \new_[6997]_  = ~\new_[2663]_ ;
  assign \new_[6998]_  = ~\new_[6999]_  | ~\new_[7007]_ ;
  assign \new_[6999]_  = ~\new_[7000]_  & ~\new_[5027]_ ;
  assign \new_[7000]_  = ~\new_[7006]_  | ~\new_[7004]_  | ~\new_[7001]_  | ~\new_[7002]_ ;
  assign \new_[7001]_  = ~\new_[5291]_  & (~\new_[5805]_  | ~\new_[6147]_ );
  assign \new_[7002]_  = \new_[7003]_  & \new_[7159]_ ;
  assign \new_[7003]_  = \new_[5883]_  & \new_[5981]_ ;
  assign \new_[7004]_  = ~\new_[7005]_  & (~\new_[6085]_  | ~\new_[5743]_ );
  assign \new_[7005]_  = ~\new_[6091]_  & ~\new_[7241]_ ;
  assign \new_[7006]_  = ~\new_[7231]_  | ~\new_[6125]_  | ~\new_[6987]_ ;
  assign \new_[7007]_  = ~\new_[4209]_ ;
  assign \new_[7008]_  = ~\new_[7005]_ ;
  assign \new_[7009]_  = ~\new_[6780]_  | ~\new_[6816]_ ;
  assign \new_[7010]_  = ~\new_[6814]_ ;
  assign \new_[7011]_  = ~\new_[7126]_ ;
  assign \new_[7012]_  = ~\new_[7127]_ ;
  assign \new_[7013]_  = \new_[5669]_  & \new_[7239]_ ;
  assign \new_[7014]_  = ~\new_[7015]_  | ~\new_[7201]_ ;
  assign \new_[7015]_  = ~\new_[7210]_ ;
  assign \new_[7016]_  = ~\new_[5405]_  & (~\new_[5697]_  | ~\new_[7201]_ );
  assign \new_[7017]_  = ~\new_[7201]_ ;
  assign \new_[7018]_  = ~\new_[7026]_  | ~\new_[4129]_  | ~\new_[7019]_ ;
  assign \new_[7019]_  = ~\new_[7020]_  & ~\new_[7025]_ ;
  assign \new_[7020]_  = ~\new_[7022]_  | ~\new_[7021]_  | ~\new_[7156]_ ;
  assign \new_[7021]_  = ~\new_[7058]_  & ~\new_[5509]_ ;
  assign \new_[7022]_  = \new_[7023]_  & \new_[7024]_ ;
  assign \new_[7023]_  = ~\new_[5933]_  | ~\new_[7201]_ ;
  assign \new_[7024]_  = ~\new_[7070]_  | ~\new_[7201]_ ;
  assign \new_[7025]_  = ~\new_[7153]_  | ~\new_[5901]_ ;
  assign \new_[7026]_  = ~\new_[5534]_ ;
  assign \new_[7027]_  = ~\new_[7031]_  | ~\new_[7030]_  | ~\new_[7028]_  | ~\new_[7231]_ ;
  assign \new_[7028]_  = ~\new_[7029]_ ;
  assign \new_[7029]_  = ~\new_[7242]_  | ~\new_[7299]_ ;
  assign \new_[7030]_  = \new_[6997]_  & \new_[7216]_ ;
  assign \new_[7031]_  = ~\new_[2666]_  & ~\new_[7063]_ ;
  assign \new_[7032]_  = ~\new_[7033]_  & ~\new_[7366]_ ;
  assign \new_[7033]_  = ~\new_[6781]_  | ~\new_[6813]_  | ~\new_[6817]_ ;
  assign \new_[7034]_  = ~\new_[7009]_  & ~\new_[7010]_ ;
  assign \new_[7035]_  = ~\new_[7063]_ ;
  assign \new_[7036]_  = \new_[7252]_  | \new_[7320]_ ;
  assign \new_[7037]_  = ~\new_[7043]_  | ~\new_[4563]_  | ~\new_[7038]_ ;
  assign \new_[7038]_  = ~\new_[7039]_  & ~\new_[5036]_ ;
  assign \new_[7039]_  = ~\new_[7040]_  | ~\new_[7042]_ ;
  assign \new_[7040]_  = ~\new_[7041]_  & ~\new_[5278]_ ;
  assign \new_[7041]_  = ~\new_[6251]_  | ~\new_[5891]_  | ~\new_[7163]_ ;
  assign \new_[7042]_  = ~\new_[5628]_  & ~\new_[5509]_ ;
  assign \new_[7043]_  = ~\new_[7044]_  & ~\new_[7046]_ ;
  assign \new_[7044]_  = ~\new_[5950]_  | ~\new_[7045]_  | ~\new_[7155]_ ;
  assign \new_[7045]_  = \new_[7059]_  & \new_[7023]_ ;
  assign \new_[7046]_  = ~\new_[5162]_ ;
  assign \new_[7047]_  = ~\new_[7189]_  | ~\new_[7202]_ ;
  assign \new_[7048]_  = ~\new_[7190]_ ;
  assign \new_[7049]_  = ~\new_[7123]_ ;
  assign \new_[7050]_  = \new_[7051]_ ;
  assign \new_[7051]_  = ~\new_[7365]_  & ~\new_[7052]_ ;
  assign \new_[7052]_  = ~\new_[7322]_  | ~\new_[7364]_ ;
  assign \new_[7053]_  = \new_[7054]_  & \new_[7251]_ ;
  assign \new_[7054]_  = ~\new_[7253]_  & ~\new_[6468]_ ;
  assign \new_[7055]_  = \new_[7319]_ ;
  assign \new_[7056]_  = ~\new_[7057]_  & ~\new_[7036]_ ;
  assign \new_[7057]_  = ~\new_[7054]_ ;
  assign \new_[7058]_  = ~\new_[7059]_ ;
  assign \new_[7059]_  = \new_[7057]_  | \new_[7060]_ ;
  assign \new_[7060]_  = ~\new_[7055]_  | ~\new_[7251]_ ;
  assign \new_[7061]_  = ~\new_[7137]_  & ~\new_[7062]_ ;
  assign \new_[7062]_  = \new_[6621]_  | \new_[6997]_ ;
  assign \new_[7063]_  = ~\new_[7364]_ ;
  assign \new_[7064]_  = ~\new_[7067]_  & ~\new_[7065]_ ;
  assign \new_[7065]_  = ~\new_[7066]_  | ~\new_[7320]_ ;
  assign \new_[7066]_  = ~\new_[7216]_  & ~\new_[6651]_ ;
  assign \new_[7067]_  = ~\new_[6445]_  | ~\new_[7253]_ ;
  assign \new_[7068]_  = \new_[7069]_ ;
  assign \new_[7069]_  = ~\new_[7282]_  | ~\new_[7340]_ ;
  assign \new_[7070]_  = ~\new_[7071]_  & ~\new_[7073]_ ;
  assign \new_[7071]_  = ~\new_[7124]_  | ~\new_[7072]_ ;
  assign \new_[7072]_  = \new_[7216]_  & \new_[2663]_ ;
  assign \new_[7073]_  = ~\new_[7028]_  | ~\new_[7231]_ ;
  assign \new_[7074]_  = ~\new_[7482]_ ;
  assign \new_[7075]_  = ~\new_[7371]_ ;
  assign \new_[7076]_  = \new_[5143]_  & \new_[2716]_ ;
  assign \new_[7077]_  = ~\new_[7358]_ ;
  assign \new_[7078]_  = ~\new_[7357]_  & ~\new_[7079]_ ;
  assign \new_[7079]_  = ~\new_[7084]_  | ~\new_[7080]_  | ~\new_[7083]_ ;
  assign \new_[7080]_  = ~\new_[7081]_  & ~\new_[7082]_ ;
  assign \new_[7081]_  = ~\new_[2598]_  | ~\new_[2691]_ ;
  assign \new_[7082]_  = ~\new_[2596]_  | ~\new_[2701]_ ;
  assign \new_[7083]_  = \new_[2689]_  & \new_[2610]_ ;
  assign \new_[7084]_  = \new_[2597]_  & \new_[2690]_ ;
  assign \new_[7085]_  = ~\new_[7084]_  | ~\new_[7080]_  | ~\new_[7083]_ ;
  assign \new_[7086]_  = \new_[7087]_  | \new_[7089]_ ;
  assign \new_[7087]_  = \new_[7088]_  & \new_[7501]_ ;
  assign \new_[7088]_  = ~\new_[2883]_  | ~\new_[4614]_ ;
  assign \new_[7089]_  = ~\new_[7090]_  & (~\new_[7570]_  | ~\new_[6837]_ );
  assign \new_[7090]_  = \new_[7466]_  | \new_[7074]_ ;
  assign \new_[7091]_  = ~\new_[7092]_ ;
  assign \new_[7092]_  = ~\new_[7077]_  & ~\new_[2064]_ ;
  assign \new_[7093]_  = ~\new_[7094]_  & ~\new_[7095]_ ;
  assign \new_[7094]_  = \new_[7358]_ ;
  assign \new_[7095]_  = \new_[7096]_ ;
  assign \new_[7096]_  = ~\new_[7097]_ ;
  assign \new_[7097]_  = ~\new_[2231]_  | ~\new_[2230]_ ;
  assign \new_[7098]_  = ~\new_[7099]_ ;
  assign \new_[7099]_  = ~\new_[3926]_  | ~\new_[2064]_ ;
  assign \new_[7100]_  = ~\new_[7094]_  & ~\new_[7095]_ ;
  assign \new_[7101]_  = ~\new_[7100]_ ;
  assign \new_[7102]_  = ~\new_[7077]_  & ~\new_[2064]_ ;
  assign \new_[7103]_  = ~\new_[7095]_ ;
  assign \new_[7104]_  = ~\new_[7331]_  | ~\new_[7105]_  | ~\new_[7108]_ ;
  assign \new_[7105]_  = \new_[7106]_  & \new_[7107]_ ;
  assign \new_[7106]_  = ~\new_[7473]_  | ~\new_[1597]_ ;
  assign \new_[7107]_  = ~\new_[7532]_  | ~\new_[1405]_  | ~\new_[1698]_ ;
  assign \new_[7108]_  = ~\new_[1598]_  & (~\new_[1544]_  | ~\new_[7532]_ );
  assign \new_[7109]_  = \new_[7110]_  & \new_[7107]_ ;
  assign \new_[7110]_  = ~\new_[7473]_  | ~\new_[1597]_ ;
  assign \new_[7111]_  = ~\new_[7112]_ ;
  assign \new_[7112]_  = ~\new_[1598]_  & (~\new_[1544]_  | ~\new_[7532]_ );
  assign \new_[7113]_  = ~\new_[7501]_  | ~\new_[7267]_  | ~\new_[7114]_ ;
  assign \new_[7114]_  = \new_[2976]_  | \new_[5295]_ ;
  assign \new_[7115]_  = \new_[7269]_ ;
  assign \new_[7116]_  = \new_[7117]_ ;
  assign \new_[7117]_  = ~\new_[7118]_  & ~\new_[7119]_ ;
  assign \new_[7118]_  = ~\new_[7125]_  | ~\new_[7231]_ ;
  assign \new_[7119]_  = ~\new_[7031]_  | ~\new_[7072]_ ;
  assign \new_[7120]_  = ~\new_[7349]_  | ~\new_[7201]_ ;
  assign \new_[7121]_  = ~\new_[7181]_  & ~\new_[7122]_ ;
  assign \new_[7122]_  = ~\new_[7125]_  | ~\new_[7123]_  | ~\new_[7124]_ ;
  assign \new_[7123]_  = \new_[7554]_  & \new_[7321]_ ;
  assign \new_[7124]_  = ~\new_[2666]_  & ~\new_[7035]_ ;
  assign \new_[7125]_  = ~\new_[6522]_  & ~\new_[7242]_ ;
  assign \new_[7126]_  = ~\new_[7032]_  | ~\new_[7034]_ ;
  assign \new_[7127]_  = ~\new_[6616]_  & ~\new_[7191]_ ;
  assign \new_[7128]_  = ~\new_[6480]_  | ~\new_[7048]_ ;
  assign \new_[7129]_  = ~\new_[7130]_ ;
  assign \new_[7130]_  = ~\new_[7131]_  | ~\new_[6171]_ ;
  assign \new_[7131]_  = ~\new_[7132]_  & ~\new_[7133]_ ;
  assign \new_[7132]_  = ~\new_[6465]_  | ~\new_[6934]_ ;
  assign \new_[7133]_  = ~\new_[6400]_  | ~\new_[6104]_ ;
  assign \new_[7134]_  = ~\new_[597]_  & ~\new_[6517]_ ;
  assign \new_[7135]_  = ~\new_[7136]_  | ~\new_[6171]_ ;
  assign \new_[7136]_  = ~\new_[7133]_ ;
  assign \new_[7137]_  = ~\new_[7364]_  | ~\new_[2666]_ ;
  assign \new_[7138]_  = ~\new_[7556]_  | ~\new_[7246]_  | ~\new_[7322]_ ;
  assign \new_[7139]_  = ~\new_[7140]_  | ~\new_[7141]_ ;
  assign \new_[7140]_  = ~\new_[2118]_  | ~\new_[4002]_ ;
  assign \new_[7141]_  = ~\new_[7358]_  & ~\new_[2117]_ ;
  assign \new_[7142]_  = ~\new_[2066]_  | ~\new_[7077]_ ;
  assign \new_[7143]_  = ~\new_[7144]_  & ~\new_[7146]_ ;
  assign \new_[7144]_  = ~\new_[6133]_  & (~\new_[7541]_  | ~\new_[7128]_ );
  assign \new_[7145]_  = ~\new_[6418]_  & ~\new_[6996]_ ;
  assign \new_[7146]_  = ~\new_[6932]_  | ~\new_[7560]_  | ~\new_[6931]_ ;
  assign \new_[7147]_  = ~\new_[6133]_  & (~\new_[7128]_  | ~\new_[7542]_ );
  assign \new_[7148]_  = ~\new_[7150]_  | ~\new_[5033]_  | ~\new_[4306]_  | ~\new_[7149]_ ;
  assign \new_[7149]_  = ~\new_[5291]_  & ~\new_[5027]_ ;
  assign \new_[7150]_  = ~\new_[7151]_  & ~\new_[7046]_ ;
  assign \new_[7151]_  = \new_[7152]_  | \new_[7154]_ ;
  assign \new_[7152]_  = ~\new_[7153]_  | ~\new_[7163]_ ;
  assign \new_[7153]_  = \new_[5891]_  & \new_[5950]_ ;
  assign \new_[7154]_  = ~\new_[7155]_  | ~\new_[7157]_ ;
  assign \new_[7155]_  = \new_[7156]_ ;
  assign \new_[7156]_  = ~\new_[6810]_  | ~\new_[6038]_ ;
  assign \new_[7157]_  = \new_[6986]_  & \new_[6251]_ ;
  assign \new_[7158]_  = ~\new_[7156]_ ;
  assign \new_[7159]_  = ~\new_[7161]_  | ~\new_[7160]_  | ~\new_[7298]_ ;
  assign \new_[7160]_  = ~\new_[7350]_ ;
  assign \new_[7161]_  = \new_[2666]_ ;
  assign \new_[7162]_  = ~\new_[7164]_ ;
  assign \new_[7163]_  = ~\new_[7168]_  | ~\new_[7166]_  | ~\new_[7164]_ ;
  assign \new_[7164]_  = ~\new_[7165]_ ;
  assign \new_[7165]_  = \new_[6450]_  | \new_[7552]_ ;
  assign \new_[7166]_  = ~\new_[2666]_  & ~\new_[7167]_ ;
  assign \new_[7167]_  = \new_[7368]_ ;
  assign \new_[7168]_  = ~\new_[7169]_ ;
  assign \new_[7169]_  = ~\new_[7254]_  | ~\new_[7299]_ ;
  assign \new_[7170]_  = ~\new_[7167]_ ;
  assign \new_[7171]_  = \new_[6571]_  | \new_[5653]_ ;
  assign \new_[7172]_  = ~\new_[5595]_  | ~\new_[6313]_  | ~\new_[6070]_ ;
  assign \new_[7173]_  = ~\new_[6305]_  | ~\new_[5518]_  | ~\new_[6313]_ ;
  assign \new_[7174]_  = ~\new_[7172]_  | ~\new_[7173]_ ;
  assign \new_[7175]_  = ~\new_[7180]_  | ~\new_[7176]_ ;
  assign \new_[7176]_  = ~\new_[7177]_  & ~\new_[7138]_ ;
  assign \new_[7177]_  = ~\new_[7247]_  | ~\new_[7178]_  | ~\new_[7179]_ ;
  assign \new_[7178]_  = \new_[6533]_  & \new_[6997]_ ;
  assign \new_[7179]_  = ~\new_[7137]_ ;
  assign \new_[7180]_  = ~\new_[6309]_  | ~\new_[7128]_ ;
  assign \new_[7181]_  = ~\new_[7178]_ ;
  assign \new_[7182]_  = ~\new_[952]_ ;
  assign \new_[7183]_  = ~\new_[7186]_  | (~\new_[7184]_  & ~\new_[2261]_ );
  assign \new_[7184]_  = \new_[7335]_  | \new_[7185]_ ;
  assign \new_[7185]_  = \new_[6723]_  & \new_[849]_ ;
  assign \new_[7186]_  = \new_[7187]_  | \new_[5682]_ ;
  assign \new_[7187]_  = \new_[6231]_  | \new_[7188]_ ;
  assign \new_[7188]_  = ~\new_[6189]_  | ~\new_[6286]_  | ~\new_[6202]_  | ~\new_[6254]_ ;
  assign \new_[7189]_  = \new_[7190]_  | \new_[7191]_ ;
  assign \new_[7190]_  = \new_[1052]_ ;
  assign \new_[7191]_  = ~\new_[7192]_  | ~\new_[952]_ ;
  assign \new_[7192]_  = ~\new_[1032]_ ;
  assign \new_[7193]_  = \new_[7189]_ ;
  assign \new_[7194]_  = ~\new_[7198]_  | ~\new_[7195]_  | ~\new_[7196]_ ;
  assign \new_[7195]_  = \new_[595]_  ? \new_[3237]_  : \new_[6827]_ ;
  assign \new_[7196]_  = \new_[6707]_  ? \new_[7197]_  : \new_[597]_ ;
  assign \new_[7197]_  = ~\new_[7199]_  | ~\new_[6041]_ ;
  assign \new_[7198]_  = \new_[596]_  ? \new_[3087]_  : \new_[6666]_ ;
  assign \new_[7199]_  = ~\new_[7200]_  | ~\new_[7204]_ ;
  assign \new_[7200]_  = ~\new_[7201]_ ;
  assign \new_[7201]_  = \new_[7202]_ ;
  assign \new_[7202]_  = ~\new_[7203]_  | ~\new_[7182]_ ;
  assign \new_[7203]_  = ~\new_[6893]_ ;
  assign \new_[7204]_  = ~\new_[7206]_  | (~\new_[7205]_  & ~\new_[6031]_ );
  assign \new_[7205]_  = ~\new_[4011]_  & ~\new_[3624]_ ;
  assign \new_[7206]_  = ~\new_[7207]_  & (~\new_[6193]_  | ~\new_[4060]_ );
  assign \new_[7207]_  = \new_[4335]_  & \new_[6272]_ ;
  assign \new_[7208]_  = \new_[7200]_ ;
  assign \new_[7209]_  = ~\new_[7200]_ ;
  assign \new_[7210]_  = ~\new_[7555]_  | ~\new_[7253]_  | ~\new_[7211]_  | ~\new_[6500]_ ;
  assign \new_[7211]_  = \new_[7212]_  & \new_[7213]_ ;
  assign \new_[7212]_  = \new_[7243]_  & \new_[2666]_ ;
  assign \new_[7213]_  = ~\new_[2662]_ ;
  assign \new_[7214]_  = ~\new_[7555]_  | ~\new_[7212]_ ;
  assign \new_[7215]_  = \new_[7253]_  & \new_[6500]_ ;
  assign \new_[7216]_  = ~\new_[2662]_ ;
  assign \new_[7217]_  = ~\new_[7550]_  | ~\new_[2666]_ ;
  assign \new_[7218]_  = ~\new_[7221]_  | (~\new_[7219]_  & ~\new_[2137]_ );
  assign \new_[7219]_  = \new_[7335]_  | \new_[7220]_ ;
  assign \new_[7220]_  = \new_[6723]_  & \new_[848]_ ;
  assign \new_[7221]_  = \new_[7222]_  | \new_[5682]_ ;
  assign \new_[7222]_  = \new_[6231]_  | \new_[7223]_ ;
  assign \new_[7223]_  = ~\new_[6180]_  | ~\new_[6301]_  | ~\new_[6153]_  | ~\new_[6217]_ ;
  assign \new_[7224]_  = ~\new_[7227]_  | ~\new_[4798]_  | ~\new_[7225]_  | ~\new_[7013]_ ;
  assign \new_[7225]_  = ~\new_[7226]_ ;
  assign \new_[7226]_  = ~\new_[6016]_  | ~\new_[5279]_  | ~\new_[5390]_ ;
  assign \new_[7227]_  = ~\new_[7228]_  & ~\new_[7229]_ ;
  assign \new_[7228]_  = ~\new_[7014]_  | ~\new_[5869]_  | ~\new_[5673]_  | ~\new_[5698]_ ;
  assign \new_[7229]_  = ~\new_[7238]_  | ~\new_[7230]_  | ~\new_[7016]_  | ~\new_[5694]_ ;
  assign \new_[7230]_  = ~\new_[7316]_  | ~\new_[5906]_ ;
  assign \new_[7231]_  = ~\new_[2556]_  & ~\new_[7322]_ ;
  assign \new_[7232]_  = ~\new_[7233]_  | ~\new_[7234]_ ;
  assign \new_[7233]_  = ~\new_[5566]_  | ~\new_[5928]_ ;
  assign \new_[7234]_  = ~\new_[7235]_  & (~\new_[5138]_  | ~\new_[7562]_ );
  assign \new_[7235]_  = ~\new_[7236]_  | ~\new_[7237]_ ;
  assign \new_[7236]_  = \new_[5399]_  | \new_[5660]_ ;
  assign \new_[7237]_  = \new_[7238]_  & \new_[7239]_ ;
  assign \new_[7238]_  = ~\new_[6137]_  | ~\new_[7201]_ ;
  assign \new_[7239]_  = ~\new_[6032]_  | ~\new_[7201]_ ;
  assign \new_[7240]_  = ~\new_[7241]_  & ~\new_[7244]_ ;
  assign \new_[7241]_  = ~\new_[2665]_  | ~\new_[7242]_ ;
  assign \new_[7242]_  = ~\new_[7243]_ ;
  assign \new_[7243]_  = \new_[2664]_ ;
  assign \new_[7244]_  = ~\new_[7245]_ ;
  assign \new_[7245]_  = ~\new_[7556]_  & ~\new_[7321]_ ;
  assign \new_[7246]_  = \new_[7242]_ ;
  assign \new_[7247]_  = ~\new_[7299]_ ;
  assign \new_[7248]_  = ~\new_[7249]_  & ~\new_[7250]_ ;
  assign \new_[7249]_  = \new_[7299]_  | \new_[7552]_ ;
  assign \new_[7250]_  = ~\new_[7251]_  | ~\new_[7253]_ ;
  assign \new_[7251]_  = ~\new_[7252]_ ;
  assign \new_[7252]_  = ~\new_[6651]_  | ~\new_[2662]_ ;
  assign \new_[7253]_  = ~\new_[7254]_ ;
  assign \new_[7254]_  = \new_[2663]_ ;
  assign \new_[7255]_  = ~\new_[7260]_  | ~\new_[7257]_  | ~\new_[4003]_  | ~\new_[7256]_ ;
  assign \new_[7256]_  = ~\new_[4590]_  & ~\new_[4447]_ ;
  assign \new_[7257]_  = ~\new_[7258]_  & ~\new_[7259]_ ;
  assign \new_[7258]_  = ~\new_[5883]_  | ~\new_[4517]_  | ~\new_[4757]_ ;
  assign \new_[7259]_  = ~\new_[4969]_  | ~\new_[4591]_  | ~\new_[4685]_ ;
  assign \new_[7260]_  = ~\new_[7261]_ ;
  assign \new_[7261]_  = ~\new_[4845]_  | ~\new_[7262]_  | ~\new_[7263]_ ;
  assign \new_[7262]_  = ~\new_[4383]_  & (~\new_[5598]_  | ~\new_[5301]_ );
  assign \new_[7263]_  = ~\new_[4903]_  | ~\new_[5598]_ ;
  assign \new_[7264]_  = ~\new_[7393]_  | ~\new_[7075]_ ;
  assign \new_[7265]_  = ~\new_[7266]_  | ~\new_[7267]_ ;
  assign \new_[7266]_  = ~\new_[7300]_ ;
  assign \new_[7267]_  = \new_[7268]_ ;
  assign \new_[7268]_  = ~\new_[7303]_  | ~\new_[7269]_ ;
  assign \new_[7269]_  = \new_[6577]_  & \new_[6669]_ ;
  assign \new_[7270]_  = \new_[7271]_  & \new_[7274]_ ;
  assign \new_[7271]_  = ~\new_[7272]_  | ~\new_[732]_ ;
  assign \new_[7272]_  = ~\new_[7273]_ ;
  assign \new_[7273]_  = ~\new_[7451]_  | ~\new_[3008]_  | ~\new_[7446]_ ;
  assign \new_[7274]_  = ~\new_[7275]_  | ~\new_[735]_ ;
  assign \new_[7275]_  = ~\new_[7276]_ ;
  assign \new_[7276]_  = ~\new_[7448]_  | ~\new_[2952]_  | ~\new_[7451]_ ;
  assign \new_[7277]_  = ~\new_[732]_ ;
  assign \new_[7278]_  = ~\new_[7501]_  | ~\new_[5184]_  | ~\new_[7279]_  | ~\new_[3571]_ ;
  assign \new_[7279]_  = ~\new_[7569]_  | ~\new_[6837]_ ;
  assign \new_[7280]_  = \new_[6971]_  & \new_[6970]_ ;
  assign \new_[7281]_  = ~\new_[7501]_  | ~\new_[5184]_  | ~\new_[7279]_  | ~\new_[3571]_ ;
  assign \new_[7282]_  = ~\new_[7287]_  | ~\new_[7283]_  | ~\new_[7353]_ ;
  assign \new_[7283]_  = ~\new_[7284]_  | ~\new_[7286]_ ;
  assign \new_[7284]_  = ~\new_[7285]_ ;
  assign \new_[7285]_  = ~\new_[7139]_  | ~\new_[7142]_ ;
  assign \new_[7286]_  = ~\new_[2032]_  | ~\new_[1929]_  | ~\new_[2040]_ ;
  assign \new_[7287]_  = ~\new_[7348]_ ;
  assign \new_[7288]_  = \new_[7283]_ ;
  assign \new_[7289]_  = \new_[7290]_  ? \new_[7292]_  : \new_[7291]_ ;
  assign \new_[7290]_  = ~\new_[5965]_  | ~\new_[1324]_ ;
  assign \new_[7291]_  = ~\new_[7290]_ ;
  assign \new_[7292]_  = \new_[7293]_  | \new_[7294]_ ;
  assign \new_[7293]_  = ~\new_[6949]_  | (~\new_[5965]_  & ~\new_[1324]_ );
  assign \new_[7294]_  = ~\new_[6958]_  & (~\new_[6947]_  | ~\new_[6957]_ );
  assign \new_[7295]_  = ~\new_[7294]_ ;
  assign \new_[7296]_  = ~\new_[7297]_  | ~\new_[7321]_ ;
  assign \new_[7297]_  = ~\new_[7298]_ ;
  assign \new_[7298]_  = \new_[7299]_ ;
  assign \new_[7299]_  = ~\new_[2665]_ ;
  assign \new_[7300]_  = ~\new_[7301]_  | ~\new_[7303]_  | ~\new_[7302]_ ;
  assign \new_[7301]_  = ~\new_[6990]_  | ~\new_[6993]_ ;
  assign \new_[7302]_  = ~\new_[4058]_  & (~\new_[5508]_  | ~\new_[2716]_ );
  assign \new_[7303]_  = ~\new_[7304]_  | ~\new_[7305]_ ;
  assign \new_[7304]_  = ~\new_[6702]_  | ~\new_[5734]_ ;
  assign \new_[7305]_  = ~\new_[7306]_  | ~\new_[7307]_ ;
  assign \new_[7306]_  = ~\new_[6494]_ ;
  assign \new_[7307]_  = ~\new_[597]_ ;
  assign \new_[7308]_  = ~\new_[7305]_ ;
  assign \new_[7309]_  = ~\new_[7310]_  & ~\new_[7312]_ ;
  assign \new_[7310]_  = ~\new_[7567]_  & ~\new_[7311]_ ;
  assign \new_[7311]_  = ~\new_[7075]_  | ~\new_[7393]_ ;
  assign \new_[7312]_  = ~\new_[7314]_  | ~\new_[7313]_ ;
  assign \new_[7313]_  = ~\new_[7393]_  | ~\new_[1886]_ ;
  assign \new_[7314]_  = ~\new_[1942]_  | ~\new_[3854]_ ;
  assign \new_[7315]_  = \new_[7316]_ ;
  assign \new_[7316]_  = \new_[7317]_  & \new_[7324]_ ;
  assign \new_[7317]_  = \new_[7318]_  & \new_[7323]_ ;
  assign \new_[7318]_  = \new_[7319]_ ;
  assign \new_[7319]_  = \new_[7320]_ ;
  assign \new_[7320]_  = \new_[7321]_ ;
  assign \new_[7321]_  = ~\new_[7322]_ ;
  assign \new_[7322]_  = \new_[2779]_ ;
  assign \new_[7323]_  = ~\new_[6331]_  & ~\new_[7551]_ ;
  assign \new_[7324]_  = ~\new_[7325]_ ;
  assign \new_[7325]_  = \new_[7326]_ ;
  assign \new_[7326]_  = \new_[6997]_  | \new_[7299]_ ;
  assign \new_[7327]_  = ~\new_[3854]_  | ~\new_[7328]_  | ~\new_[7329]_ ;
  assign \new_[7328]_  = ~\new_[7375]_  | ~\new_[3705]_ ;
  assign \new_[7329]_  = ~\new_[7330]_ ;
  assign \new_[7330]_  = ~\new_[1944]_  & (~\new_[1837]_  | ~\new_[1887]_ );
  assign \new_[7331]_  = ~\new_[1837]_  | ~\new_[3854]_ ;
  assign \new_[7332]_  = ~\new_[1944]_  | ~\new_[3854]_ ;
  assign \new_[7333]_  = ~\new_[7337]_  | (~\new_[7334]_  & ~\new_[2311]_ );
  assign \new_[7334]_  = \new_[7335]_  | \new_[7336]_ ;
  assign \new_[7335]_  = ~\new_[6231]_  & ~\new_[5682]_ ;
  assign \new_[7336]_  = \new_[6723]_  & \new_[852]_ ;
  assign \new_[7337]_  = \new_[7338]_  | \new_[5682]_ ;
  assign \new_[7338]_  = \new_[6231]_  | \new_[7339]_ ;
  assign \new_[7339]_  = ~\new_[6144]_  | ~\new_[6294]_  | ~\new_[6188]_  | ~\new_[6150]_ ;
  assign \new_[7340]_  = ~\new_[7341]_  & ~\new_[7345]_ ;
  assign \new_[7341]_  = ~\new_[7344]_  & (~\new_[7342]_  | ~\new_[7373]_ );
  assign \new_[7342]_  = ~\new_[7343]_ ;
  assign \new_[7343]_  = ~\new_[7362]_  & ~\new_[4002]_ ;
  assign \new_[7344]_  = ~\new_[7360]_  | ~\new_[2031]_  | ~\new_[6688]_ ;
  assign \new_[7345]_  = ~\new_[1825]_  | ~\new_[1991]_ ;
  assign \new_[7346]_  = ~\new_[7342]_  | (~\new_[7374]_  & ~\new_[7347]_ );
  assign \new_[7347]_  = ~\new_[7360]_ ;
  assign \new_[7348]_  = ~\new_[2031]_  | ~\new_[6688]_ ;
  assign \new_[7349]_  = ~\new_[7350]_  & ~\new_[7351]_ ;
  assign \new_[7350]_  = ~\new_[7253]_  & ~\new_[7165]_ ;
  assign \new_[7351]_  = \new_[7296]_  | \new_[6400]_  | \new_[2666]_  | \new_[7352]_ ;
  assign \new_[7352]_  = \new_[7246]_ ;
  assign \new_[7353]_  = ~\new_[7354]_ ;
  assign \new_[7354]_  = ~\new_[7355]_  | ~\new_[7360]_ ;
  assign \new_[7355]_  = ~\new_[7356]_ ;
  assign \new_[7356]_  = ~\new_[7357]_  & ~\new_[2121]_ ;
  assign \new_[7357]_  = ~\new_[7358]_ ;
  assign \new_[7358]_  = \new_[7359]_ ;
  assign \new_[7359]_  = ~\new_[7076]_  & (~\new_[4448]_  | ~\new_[6473]_ );
  assign \new_[7360]_  = ~\new_[7358]_  | ~\new_[7361]_ ;
  assign \new_[7361]_  = ~\new_[2322]_  & ~\new_[2321]_ ;
  assign \new_[7362]_  = ~\new_[2322]_  & ~\new_[2321]_ ;
  assign \new_[7363]_  = ~\new_[6567]_  & ~\new_[7364]_ ;
  assign \new_[7364]_  = ~\new_[2727]_ ;
  assign \new_[7365]_  = ~\new_[2664]_ ;
  assign \new_[7366]_  = ~\new_[7367]_  | ~\new_[7370]_ ;
  assign \new_[7367]_  = ~\new_[7368]_  | ~\new_[7369]_ ;
  assign \new_[7368]_  = \new_[6892]_  & \new_[6704]_ ;
  assign \new_[7369]_  = ~\new_[844]_ ;
  assign \new_[7370]_  = ~\new_[6811]_  | ~\new_[6659]_ ;
  assign \new_[7371]_  = ~\new_[7357]_  & ~\new_[7538]_ ;
  assign \new_[7372]_  = ~\new_[7357]_  & ~\new_[7538]_ ;
  assign \new_[7373]_  = ~\new_[6681]_  | ~\new_[3927]_ ;
  assign \new_[7374]_  = ~\new_[6681]_  | ~\new_[3927]_ ;
  assign \new_[7375]_  = ~\new_[1887]_ ;
  assign \new_[7376]_  = ~\new_[7379]_ ;
  assign \new_[7377]_  = ~\new_[7378]_ ;
  assign \new_[7378]_  = \new_[7379]_ ;
  assign \new_[7379]_  = ~\new_[5798]_ ;
  assign n469 = ~\new_[7385]_  | (~\new_[7381]_  & ~\new_[7384]_ );
  assign \new_[7381]_  = ~\new_[7382]_  & ~\new_[7474]_ ;
  assign \new_[7382]_  = ~\new_[7383]_ ;
  assign \new_[7383]_  = ~\new_[2849]_  & ~\new_[2809]_ ;
  assign \new_[7384]_  = ~\new_[7515]_  | (~\new_[7383]_  & ~\new_[537]_ );
  assign \new_[7385]_  = ~\new_[1192]_  | ~\new_[537]_ ;
  assign n349 = ~\new_[7387]_  | ~\new_[7391]_ ;
  assign \new_[7387]_  = ~\new_[7515]_  | ~\new_[7388]_  | ~\new_[7390]_ ;
  assign \new_[7388]_  = ~\new_[7389]_  | ~\new_[7278]_  | ~\new_[7280]_ ;
  assign \new_[7389]_  = ~\new_[2899]_  & ~\new_[2845]_ ;
  assign \new_[7390]_  = \new_[6642]_  | \new_[7389]_ ;
  assign \new_[7391]_  = ~\new_[1184]_  | ~\new_[6642]_ ;
  assign \new_[7392]_  = ~\new_[7278]_  | ~\new_[7280]_ ;
  assign \new_[7393]_  = ~\new_[1996]_  | ~\new_[4001]_ ;
  assign \new_[7394]_  = ~\new_[6692]_  | ~\new_[3853]_ ;
  assign n464 = ~\new_[7400]_  | (~\new_[7396]_  & ~\new_[7399]_ );
  assign \new_[7396]_  = ~\new_[7397]_  & ~\new_[7474]_ ;
  assign \new_[7397]_  = ~\new_[7398]_ ;
  assign \new_[7398]_  = \new_[2758]_  & \new_[2814]_ ;
  assign \new_[7399]_  = ~\new_[7515]_  | (~\new_[7398]_  & ~\new_[536]_ );
  assign \new_[7400]_  = ~\new_[1187]_  | ~\new_[536]_ ;
  assign \new_[7401]_  = ~\new_[7415]_  | (~\new_[7402]_  & ~\new_[7410]_ );
  assign \new_[7402]_  = ~\new_[886]_  | ~\new_[729]_  | ~\new_[7403]_ ;
  assign \new_[7403]_  = ~\new_[7404]_ ;
  assign \new_[7404]_  = ~\new_[7407]_  | ~\new_[937]_  | ~\new_[7405]_ ;
  assign \new_[7405]_  = ~\new_[7406]_ ;
  assign \new_[7406]_  = \new_[1757]_  ^ \new_[7288]_ ;
  assign \new_[7407]_  = \new_[7408]_  & \new_[7409]_ ;
  assign \new_[7408]_  = ~\new_[1625]_ ;
  assign \new_[7409]_  = ~\new_[1747]_ ;
  assign \new_[7410]_  = ~\new_[7413]_  | ~\new_[887]_  | ~\new_[7411]_ ;
  assign \new_[7411]_  = ~\new_[7412]_ ;
  assign \new_[7412]_  = ~\new_[1945]_  | ~\new_[1215]_  | ~\new_[1153]_ ;
  assign \new_[7413]_  = ~\new_[7414]_ ;
  assign \new_[7414]_  = ~\new_[5392]_  | ~\new_[3842]_  | ~\new_[3998]_  | ~\new_[3754]_ ;
  assign \new_[7415]_  = \new_[7413]_  | \new_[7416]_ ;
  assign \new_[7416]_  = \new_[2078]_  ? \new_[4511]_  : \new_[407]_ ;
  assign n489 = ~\new_[7421]_  | (~\new_[7418]_  & ~\new_[7420]_ );
  assign \new_[7418]_  = ~\new_[7419]_  & ~\new_[7474]_ ;
  assign \new_[7419]_  = ~\new_[7514]_ ;
  assign \new_[7420]_  = ~\new_[7515]_  | (~\new_[7514]_  & ~\new_[542]_ );
  assign \new_[7421]_  = ~\new_[1181]_  | ~\new_[542]_ ;
  assign n369 = ~\new_[7423]_  | ~\new_[7429]_ ;
  assign \new_[7423]_  = ~\new_[7428]_  | ~\new_[7424]_  | ~\new_[7427]_ ;
  assign \new_[7424]_  = ~\new_[6900]_  | ~\new_[7425]_  | ~\new_[6904]_ ;
  assign \new_[7425]_  = \new_[7426]_ ;
  assign \new_[7426]_  = ~\new_[2809]_  & ~\new_[2814]_ ;
  assign \new_[7427]_  = \new_[6672]_  | \new_[7425]_ ;
  assign \new_[7428]_  = \new_[7515]_ ;
  assign \new_[7429]_  = ~\new_[1184]_  | ~\new_[6672]_ ;
  assign \new_[7430]_  = ~\new_[7428]_ ;
  assign \new_[7431]_  = ~\new_[6900]_  | ~\new_[6904]_ ;
  assign \new_[7432]_  = ~\new_[7425]_ ;
  assign \new_[7433]_  = ~\new_[7440]_  & (~\new_[7434]_  | ~\new_[7437]_ );
  assign \new_[7434]_  = ~\new_[5223]_  | ~\new_[1502]_  | ~\new_[7435]_ ;
  assign \new_[7435]_  = ~\new_[7436]_ ;
  assign \new_[7436]_  = ~\new_[7173]_  | ~\new_[7172]_  | ~\new_[7171]_ ;
  assign \new_[7437]_  = ~\new_[7438]_  & (~\new_[7435]_  | ~\new_[4950]_ );
  assign \new_[7438]_  = ~\new_[7439]_ ;
  assign \new_[7439]_  = ~\new_[7174]_  | ~\new_[2429]_ ;
  assign \new_[7440]_  = ~\new_[6231]_  & ~\new_[7135]_ ;
  assign \new_[7441]_  = ~\new_[7442]_  | ~\new_[433]_ ;
  assign \new_[7442]_  = \new_[7443]_ ;
  assign \new_[7443]_  = \new_[7444]_ ;
  assign \new_[7444]_  = ~\new_[7445]_ ;
  assign \new_[7445]_  = ~\new_[7450]_  | ~\new_[7447]_  | ~\new_[7543]_ ;
  assign \new_[7446]_  = ~\new_[7543]_ ;
  assign \new_[7447]_  = ~\new_[7448]_ ;
  assign \new_[7448]_  = ~\new_[7449]_ ;
  assign \new_[7449]_  = ~\new_[7265]_  | ~\new_[3248]_  | ~\new_[7113]_ ;
  assign \new_[7450]_  = ~\new_[7451]_ ;
  assign \new_[7451]_  = ~\new_[7452]_ ;
  assign \new_[7452]_  = ~\new_[3193]_  & ~\new_[3241]_ ;
  assign \new_[7453]_  = ~\new_[7456]_  | ~\new_[7454]_  | ~\new_[7455]_ ;
  assign \new_[7454]_  = ~\new_[7442]_  | ~\new_[6559]_ ;
  assign \new_[7455]_  = ~\new_[7489]_  | ~\new_[6598]_ ;
  assign \new_[7456]_  = (~\new_[6590]_  | ~\new_[2706]_ ) & (~\new_[7457]_  | ~\new_[6482]_ );
  assign \new_[7457]_  = ~\new_[7458]_ ;
  assign \new_[7458]_  = ~\new_[7459]_ ;
  assign \new_[7459]_  = ~\new_[7460]_ ;
  assign \new_[7460]_  = ~\new_[2894]_  | ~\new_[2898]_ ;
  assign \new_[7461]_  = ~\new_[7462]_  | ~\new_[7465]_ ;
  assign \new_[7462]_  = ~\new_[7463]_  | ~\new_[7464]_ ;
  assign \new_[7463]_  = ~\new_[1214]_  | ~\new_[1706]_ ;
  assign \new_[7464]_  = ~\new_[1213]_  | ~\new_[1641]_ ;
  assign \new_[7465]_  = ~\new_[7466]_  & ~\new_[7467]_ ;
  assign \new_[7466]_  = ~\new_[7501]_ ;
  assign \new_[7467]_  = ~\new_[7482]_ ;
  assign \new_[7468]_  = ~\new_[1706]_  | ~\new_[1214]_ ;
  assign \new_[7469]_  = \new_[7470]_  ^ \new_[7471]_ ;
  assign \new_[7470]_  = \new_[1834]_  & \new_[1836]_ ;
  assign \new_[7471]_  = ~\new_[7472]_  | ~\new_[7517]_  | ~\new_[7490]_ ;
  assign \new_[7472]_  = ~\new_[7473]_ ;
  assign \new_[7473]_  = ~\new_[1715]_  | (~\new_[6685]_  & ~\new_[7314]_ );
  assign \new_[7474]_  = ~\new_[7480]_  | ~\new_[7475]_  | ~\new_[7479]_ ;
  assign \new_[7475]_  = ~\new_[7476]_  | ~\new_[7477]_ ;
  assign \new_[7476]_  = \new_[1705]_  ? \new_[1355]_  : \new_[1754]_ ;
  assign \new_[7477]_  = ~\new_[7478]_ ;
  assign \new_[7478]_  = ~\new_[7501]_  | ~\new_[3571]_  | ~\new_[5184]_ ;
  assign \new_[7479]_  = ~\new_[3932]_  | ~\new_[7466]_ ;
  assign \new_[7480]_  = ~\new_[7481]_  | ~\new_[7501]_ ;
  assign \new_[7481]_  = ~\new_[3235]_  | (~\new_[5184]_  & ~\new_[1809]_ );
  assign \new_[7482]_  = \new_[3571]_  & \new_[5184]_ ;
  assign \new_[7483]_  = ~\new_[7488]_  | (~\new_[7484]_  & ~\new_[505]_ );
  assign \new_[7484]_  = ~\new_[7485]_ ;
  assign \new_[7485]_  = \new_[7486]_ ;
  assign \new_[7486]_  = ~\new_[7487]_ ;
  assign \new_[7487]_  = ~\new_[2952]_  | ~\new_[3015]_  | ~\new_[3009]_ ;
  assign \new_[7488]_  = ~\new_[2706]_  | ~\new_[6477]_ ;
  assign \new_[7489]_  = ~\new_[7484]_ ;
  assign \new_[7490]_  = ~\new_[7520]_  | ~\new_[7494]_  | ~\new_[7491]_  | ~\new_[7522]_ ;
  assign \new_[7491]_  = \new_[7492]_  & \new_[7493]_ ;
  assign \new_[7492]_  = ~\new_[1742]_  | ~\new_[1701]_ ;
  assign \new_[7493]_  = \new_[7360]_  & \new_[2031]_ ;
  assign \new_[7494]_  = ~\new_[7495]_ ;
  assign \new_[7495]_  = ~\new_[7496]_ ;
  assign \new_[7496]_  = ~\new_[1927]_  & ~\new_[6687]_ ;
  assign \new_[7497]_  = ~\new_[7498]_  | ~\new_[7499]_ ;
  assign \new_[7498]_  = \new_[2808]_  & \new_[2849]_ ;
  assign \new_[7499]_  = ~\new_[7503]_  & (~\new_[1320]_  | ~\new_[7500]_ );
  assign \new_[7500]_  = \new_[7482]_  & \new_[7501]_ ;
  assign \new_[7501]_  = \new_[7502]_ ;
  assign \new_[7502]_  = ~\new_[7129]_  | ~\new_[7134]_ ;
  assign \new_[7503]_  = ~\new_[7504]_ ;
  assign \new_[7504]_  = (~\new_[6745]_  | ~\new_[3933]_ ) & (~\new_[2170]_  | ~\new_[7501]_ );
  assign \new_[7505]_  = ~\new_[7501]_ ;
  assign n374 = ~\new_[7507]_  | ~\new_[7516]_ ;
  assign \new_[7507]_  = ~\new_[7508]_  | ~\new_[7511]_ ;
  assign \new_[7508]_  = ~\new_[7509]_  | ~\new_[7281]_ ;
  assign \new_[7509]_  = \new_[7510]_  & \new_[6971]_ ;
  assign \new_[7510]_  = ~\new_[6972]_  & ~\new_[6853]_ ;
  assign \new_[7511]_  = \new_[7512]_  & \new_[7515]_ ;
  assign \new_[7512]_  = \new_[7513]_  | \new_[7514]_ ;
  assign \new_[7513]_  = ~\new_[471]_ ;
  assign \new_[7514]_  = ~\new_[2845]_  & ~\new_[2814]_ ;
  assign \new_[7515]_  = ~\new_[1690]_  & (~\new_[1370]_  | ~\new_[4930]_ );
  assign \new_[7516]_  = \new_[471]_  | \new_[7515]_ ;
  assign \new_[7517]_  = ~\new_[7522]_  | (~\new_[7518]_  & ~\new_[7521]_ );
  assign \new_[7518]_  = ~\new_[7519]_  & (~\new_[1700]_  | ~\new_[1741]_ );
  assign \new_[7519]_  = ~\new_[7520]_ ;
  assign \new_[7520]_  = ~\new_[7102]_  & ~\new_[7372]_ ;
  assign \new_[7521]_  = ~\new_[1932]_  | (~\new_[7371]_  & ~\new_[7099]_ );
  assign \new_[7522]_  = ~\new_[7533]_ ;
  assign \new_[7523]_  = ~\new_[7521]_ ;
  assign \new_[7524]_  = ~\new_[1700]_  | ~\new_[1741]_ ;
  assign \new_[7525]_  = ~\new_[7526]_  | ~\new_[7529]_  | ~\new_[7531]_  | ~\new_[7528]_ ;
  assign \new_[7526]_  = ~\new_[7527]_  & (~\new_[6975]_  | ~\new_[7513]_ );
  assign \new_[7527]_  = \new_[2712]_  & \new_[6556]_ ;
  assign \new_[7528]_  = ~\new_[2236]_ ;
  assign \new_[7529]_  = ~\new_[7530]_  & (~\new_[7442]_  | ~\new_[6672]_ );
  assign \new_[7530]_  = \new_[2713]_  & \new_[6642]_ ;
  assign \new_[7531]_  = ~\new_[2327]_ ;
  assign \new_[7532]_  = ~\new_[7533]_  & ~\new_[7534]_ ;
  assign \new_[7533]_  = ~\new_[7394]_  | ~\new_[7393]_ ;
  assign \new_[7534]_  = ~\new_[7535]_  | ~\new_[7536]_ ;
  assign \new_[7535]_  = ~\new_[1894]_  | ~\new_[3853]_ ;
  assign \new_[7536]_  = ~\new_[1997]_  | ~\new_[4001]_ ;
  assign \new_[7537]_  = ~\new_[2160]_  | ~\new_[2124]_ ;
  assign \new_[7538]_  = ~\new_[2160]_  | ~\new_[2124]_ ;
  assign \new_[7539]_  = \new_[3088]_  & \new_[6727]_ ;
  assign \new_[7540]_  = \new_[3088]_  & \new_[6727]_ ;
  assign \new_[7541]_  = ~\new_[7126]_  | ~\new_[7127]_ ;
  assign \new_[7542]_  = ~\new_[7126]_  | ~\new_[7127]_ ;
  assign \new_[7543]_  = ~\new_[6701]_  | ~\new_[6696]_  | ~\new_[6699]_ ;
  assign \new_[7544]_  = ~\new_[6701]_  | ~\new_[6696]_  | ~\new_[6699]_ ;
  assign \new_[7545]_  = ~\new_[7359]_  & ~\new_[6384]_ ;
  assign \new_[7546]_  = ~\new_[7359]_  & ~\new_[6384]_ ;
  assign \new_[7547]_  = ~\new_[1408]_  | ~\new_[7309]_ ;
  assign \new_[7548]_  = ~\new_[1408]_  | ~\new_[7309]_ ;
  assign \new_[7549]_  = ~\new_[7550]_ ;
  assign \new_[7550]_  = \new_[7552]_ ;
  assign \new_[7551]_  = ~\new_[7552]_ ;
  assign \new_[7552]_  = ~\new_[2556]_ ;
  assign \new_[7553]_  = ~\new_[7554]_ ;
  assign \new_[7554]_  = \new_[7556]_ ;
  assign \new_[7555]_  = ~\new_[7556]_ ;
  assign \new_[7556]_  = \new_[2556]_ ;
  assign \new_[7557]_  = \new_[7558]_ ;
  assign \new_[7558]_  = ~\new_[6425]_ ;
  assign \new_[7559]_  = ~\new_[7056]_  & (~\new_[7055]_  | ~\new_[7053]_ );
  assign \new_[7560]_  = ~\new_[7056]_  & (~\new_[7055]_  | ~\new_[7053]_ );
  assign \new_[7561]_  = ~\new_[7210]_  | ~\new_[5986]_ ;
  assign \new_[7562]_  = ~\new_[7210]_  | ~\new_[5986]_ ;
  assign \new_[7563]_  = ~\new_[7564]_ ;
  assign \new_[7564]_  = \new_[7565]_ ;
  assign \new_[7565]_  = ~\new_[5565]_ ;
  assign \new_[7566]_  = ~\new_[1824]_ ;
  assign \new_[7567]_  = ~\new_[7098]_  & (~\new_[7093]_  | ~\new_[7091]_ );
  assign \new_[7568]_  = ~\new_[7098]_  & (~\new_[7093]_  | ~\new_[7091]_ );
  assign \new_[7569]_  = ~\new_[6841]_  | ~\new_[6843]_ ;
  assign \new_[7570]_  = ~\new_[6841]_  | ~\new_[6843]_ ;
  always @ (posedge clock) begin
    i_tv80_core_IncDecZ_reg <= n94;
    \\i_tv80_core_A_reg[1]  <= n99;
    \\i_tv80_core_A_reg[2]  <= n104;
    \\i_tv80_core_A_reg[5]  <= n109;
    \\i_tv80_core_A_reg[6]  <= n114;
    \\i_tv80_core_i_reg_RegsH_reg[0][6]  <= n119;
    \\i_tv80_core_i_reg_RegsH_reg[1][6]  <= n124;
    \\i_tv80_core_i_reg_RegsH_reg[2][6]  <= n129;
    \\i_tv80_core_i_reg_RegsH_reg[3][6]  <= n134;
    \\i_tv80_core_i_reg_RegsH_reg[4][6]  <= n139;
    \\i_tv80_core_i_reg_RegsH_reg[5][6]  <= n144;
    \\i_tv80_core_i_reg_RegsH_reg[6][6]  <= n149;
    \\i_tv80_core_i_reg_RegsH_reg[7][6]  <= n154;
    \\i_tv80_core_i_reg_RegsH_reg[0][4]  <= n159;
    \\i_tv80_core_i_reg_RegsH_reg[1][4]  <= n164;
    \\i_tv80_core_i_reg_RegsH_reg[2][4]  <= n169;
    \\i_tv80_core_i_reg_RegsH_reg[3][4]  <= n174;
    \\i_tv80_core_i_reg_RegsH_reg[4][4]  <= n179;
    \\i_tv80_core_i_reg_RegsH_reg[5][4]  <= n184;
    \\i_tv80_core_i_reg_RegsH_reg[6][4]  <= n189;
    \\i_tv80_core_i_reg_RegsH_reg[7][4]  <= n194;
    \\i_tv80_core_i_reg_RegsH_reg[0][2]  <= n199;
    \\i_tv80_core_i_reg_RegsH_reg[1][2]  <= n204;
    \\i_tv80_core_i_reg_RegsH_reg[2][2]  <= n209;
    \\i_tv80_core_i_reg_RegsH_reg[3][2]  <= n214;
    \\i_tv80_core_i_reg_RegsH_reg[4][2]  <= n219;
    \\i_tv80_core_i_reg_RegsH_reg[5][2]  <= n224;
    \\i_tv80_core_i_reg_RegsH_reg[6][2]  <= n229;
    \\i_tv80_core_i_reg_RegsH_reg[7][2]  <= n234;
    \\i_tv80_core_A_reg[11]  <= n239;
    \\i_tv80_core_A_reg[12]  <= n244;
    \\i_tv80_core_A_reg[13]  <= n249;
    \\i_tv80_core_A_reg[14]  <= n254;
    \\i_tv80_core_A_reg[10]  <= n259;
    \\i_tv80_core_A_reg[4]  <= n264;
    \\i_tv80_core_A_reg[0]  <= n269;
    \\i_tv80_core_A_reg[3]  <= n274;
    \\i_tv80_core_A_reg[15]  <= n279;
    \\i_tv80_core_A_reg[8]  <= n284;
    \\i_tv80_core_A_reg[7]  <= n289;
    \\i_tv80_core_A_reg[9]  <= n294;
    \\i_tv80_core_i_reg_RegsH_reg[0][7]  <= n299;
    \\i_tv80_core_i_reg_RegsH_reg[1][7]  <= n304;
    \\i_tv80_core_i_reg_RegsH_reg[2][7]  <= n309;
    \\i_tv80_core_i_reg_RegsH_reg[3][7]  <= n314;
    \\i_tv80_core_i_reg_RegsH_reg[4][7]  <= n319;
    \\i_tv80_core_i_reg_RegsH_reg[5][7]  <= n324;
    \\i_tv80_core_i_reg_RegsH_reg[6][7]  <= n329;
    \\i_tv80_core_i_reg_RegsH_reg[7][7]  <= n334;
    \\i_tv80_core_i_reg_RegsH_reg[0][5]  <= n339;
    \\i_tv80_core_i_reg_RegsH_reg[1][5]  <= n344;
    \\i_tv80_core_i_reg_RegsH_reg[2][5]  <= n349;
    \\i_tv80_core_i_reg_RegsH_reg[3][5]  <= n354;
    \\i_tv80_core_i_reg_RegsH_reg[4][5]  <= n359;
    \\i_tv80_core_i_reg_RegsH_reg[7][5]  <= n364;
    \\i_tv80_core_i_reg_RegsH_reg[5][5]  <= n369;
    \\i_tv80_core_i_reg_RegsH_reg[6][5]  <= n374;
    \\i_tv80_core_i_reg_RegsH_reg[0][3]  <= n379;
    \\i_tv80_core_i_reg_RegsH_reg[1][3]  <= n384;
    \\i_tv80_core_i_reg_RegsH_reg[2][3]  <= n389;
    \\i_tv80_core_i_reg_RegsH_reg[3][3]  <= n394;
    \\i_tv80_core_i_reg_RegsH_reg[4][3]  <= n399;
    \\i_tv80_core_i_reg_RegsH_reg[5][3]  <= n404;
    \\i_tv80_core_i_reg_RegsH_reg[6][3]  <= n409;
    \\i_tv80_core_i_reg_RegsH_reg[7][3]  <= n414;
    \\i_tv80_core_i_reg_RegsH_reg[5][1]  <= n419;
    \\i_tv80_core_i_reg_RegsL_reg[0][6]  <= n424;
    \\i_tv80_core_i_reg_RegsL_reg[1][6]  <= n429;
    \\i_tv80_core_i_reg_RegsL_reg[2][6]  <= n434;
    \\i_tv80_core_i_reg_RegsL_reg[5][6]  <= n439;
    \\i_tv80_core_i_reg_RegsL_reg[6][6]  <= n444;
    \\i_tv80_core_i_reg_RegsL_reg[7][6]  <= n449;
    \\i_tv80_core_i_reg_RegsL_reg[3][6]  <= n454;
    \\i_tv80_core_i_reg_RegsL_reg[4][6]  <= n459;
    \\i_tv80_core_i_reg_RegsH_reg[0][1]  <= n464;
    \\i_tv80_core_i_reg_RegsH_reg[1][1]  <= n469;
    \\i_tv80_core_i_reg_RegsH_reg[2][1]  <= n474;
    \\i_tv80_core_i_reg_RegsH_reg[3][1]  <= n479;
    \\i_tv80_core_i_reg_RegsH_reg[4][1]  <= n484;
    \\i_tv80_core_i_reg_RegsH_reg[6][1]  <= n489;
    \\i_tv80_core_i_reg_RegsH_reg[7][1]  <= n494;
    \\i_tv80_core_i_reg_RegsH_reg[4][0]  <= n499;
    \\i_tv80_core_i_reg_RegsL_reg[7][7]  <= n504;
    \\i_tv80_core_i_reg_RegsL_reg[0][7]  <= n509;
    \\i_tv80_core_i_reg_RegsL_reg[1][7]  <= n514;
    \\i_tv80_core_i_reg_RegsL_reg[2][7]  <= n519;
    \\i_tv80_core_i_reg_RegsL_reg[3][7]  <= n524;
    \\i_tv80_core_i_reg_RegsL_reg[4][7]  <= n529;
    \\i_tv80_core_i_reg_RegsL_reg[5][7]  <= n534;
    \\i_tv80_core_i_reg_RegsL_reg[6][7]  <= n539;
    \\i_tv80_core_i_reg_RegsH_reg[0][0]  <= n544;
    \\i_tv80_core_i_reg_RegsH_reg[1][0]  <= n549;
    \\i_tv80_core_i_reg_RegsH_reg[2][0]  <= n554;
    \\i_tv80_core_i_reg_RegsH_reg[3][0]  <= n559;
    \\i_tv80_core_i_reg_RegsH_reg[5][0]  <= n564;
    \\i_tv80_core_i_reg_RegsH_reg[6][0]  <= n569;
    \\i_tv80_core_i_reg_RegsH_reg[7][0]  <= n574;
    \\i_tv80_core_tstate_reg[0]  <= n579;
    \\i_tv80_core_tstate_reg[1]  <= n584;
    \\i_tv80_core_tstate_reg[2]  <= n589;
    \\i_tv80_core_i_reg_RegsL_reg[4][4]  <= n594;
    \\i_tv80_core_i_reg_RegsL_reg[0][5]  <= n599;
    \\i_tv80_core_F_reg[2]  <= n604;
    \\i_tv80_core_i_reg_RegsL_reg[1][5]  <= n609;
    \\i_tv80_core_i_reg_RegsL_reg[2][5]  <= n614;
    \\i_tv80_core_i_reg_RegsL_reg[3][5]  <= n619;
    \\i_tv80_core_i_reg_RegsL_reg[4][5]  <= n624;
    \\i_tv80_core_i_reg_RegsL_reg[5][5]  <= n629;
    \\i_tv80_core_i_reg_RegsL_reg[6][5]  <= n634;
    \\i_tv80_core_i_reg_RegsL_reg[7][5]  <= n639;
    \\i_tv80_core_i_reg_RegsL_reg[0][4]  <= n644;
    \\i_tv80_core_i_reg_RegsL_reg[1][4]  <= n649;
    \\i_tv80_core_i_reg_RegsL_reg[2][4]  <= n654;
    \\i_tv80_core_i_reg_RegsL_reg[3][4]  <= n659;
    \\i_tv80_core_i_reg_RegsL_reg[6][4]  <= n664;
    \\i_tv80_core_i_reg_RegsL_reg[7][4]  <= n669;
    \\i_tv80_core_i_reg_RegsL_reg[5][4]  <= n674;
    \\i_tv80_core_SP_reg[14]  <= n679;
    \\i_tv80_core_i_reg_RegsL_reg[5][3]  <= n684;
    \\i_tv80_core_i_reg_RegsL_reg[6][3]  <= n689;
    \\i_tv80_core_i_reg_RegsL_reg[0][3]  <= n694;
    \\i_tv80_core_i_reg_RegsL_reg[1][3]  <= n699;
    \\i_tv80_core_i_reg_RegsL_reg[3][3]  <= n704;
    \\i_tv80_core_i_reg_RegsL_reg[4][3]  <= n709;
    \\i_tv80_core_i_reg_RegsL_reg[7][3]  <= n714;
    \\i_tv80_core_i_reg_RegsL_reg[2][3]  <= n719;
    \\i_tv80_core_ACC_reg[0]  <= n724;
    \\i_tv80_core_i_reg_RegsL_reg[4][1]  <= n729;
    \\i_tv80_core_do_reg[5]  <= n734;
    \\i_tv80_core_F_reg[1]  <= n739;
    \\i_tv80_core_SP_reg[1]  <= n744;
    \\i_tv80_core_F_reg[6]  <= n749;
    \\i_tv80_core_F_reg[0]  <= n754;
    \\i_tv80_core_ACC_reg[7]  <= n759;
    \\i_tv80_core_do_reg[7]  <= n764;
    \\i_tv80_core_SP_reg[7]  <= n769;
    \\i_tv80_core_do_reg[6]  <= n774;
    \\i_tv80_core_SP_reg[6]  <= n779;
    \\i_tv80_core_ACC_reg[3]  <= n784;
    \\i_tv80_core_ACC_reg[5]  <= n789;
    \\i_tv80_core_ACC_reg[6]  <= n794;
    \\i_tv80_core_ACC_reg[2]  <= n799;
    \\i_tv80_core_ACC_reg[1]  <= n804;
    \\i_tv80_core_ACC_reg[4]  <= n809;
    \\i_tv80_core_SP_reg[5]  <= n814;
    \\i_tv80_core_do_reg[4]  <= n819;
    \\i_tv80_core_SP_reg[4]  <= n824;
    \\i_tv80_core_i_reg_RegsL_reg[0][2]  <= n829;
    \\i_tv80_core_i_reg_RegsL_reg[1][2]  <= n834;
    \\i_tv80_core_i_reg_RegsL_reg[2][2]  <= n839;
    \\i_tv80_core_i_reg_RegsL_reg[3][2]  <= n844;
    \\i_tv80_core_i_reg_RegsL_reg[5][2]  <= n849;
    \\i_tv80_core_i_reg_RegsL_reg[6][2]  <= n854;
    \\i_tv80_core_i_reg_RegsL_reg[7][2]  <= n859;
    \\i_tv80_core_i_reg_RegsL_reg[0][1]  <= n864;
    \\i_tv80_core_i_reg_RegsL_reg[1][1]  <= n869;
    \\i_tv80_core_i_reg_RegsL_reg[2][1]  <= n874;
    \\i_tv80_core_i_reg_RegsL_reg[3][1]  <= n879;
    \\i_tv80_core_i_reg_RegsL_reg[5][1]  <= n884;
    \\i_tv80_core_i_reg_RegsL_reg[6][1]  <= n889;
    \\i_tv80_core_i_reg_RegsL_reg[7][1]  <= n894;
    \\i_tv80_core_do_reg[0]  <= n899;
    \\i_tv80_core_do_reg[1]  <= n904;
    \\i_tv80_core_do_reg[2]  <= n909;
    \\i_tv80_core_do_reg[3]  <= n914;
    \\i_tv80_core_i_reg_RegsL_reg[0][0]  <= n919;
    \\i_tv80_core_i_reg_RegsL_reg[1][0]  <= n924;
    \\i_tv80_core_i_reg_RegsL_reg[2][0]  <= n929;
    \\i_tv80_core_i_reg_RegsL_reg[3][0]  <= n934;
    \\i_tv80_core_i_reg_RegsL_reg[4][0]  <= n939;
    \\i_tv80_core_i_reg_RegsL_reg[5][0]  <= n944;
    \\i_tv80_core_i_reg_RegsL_reg[7][0]  <= n949;
    \\i_tv80_core_SP_reg[2]  <= n954;
    \\i_tv80_core_SP_reg[3]  <= n959;
    \\i_tv80_core_SP_reg[0]  <= n964;
    \\i_tv80_core_i_reg_RegsL_reg[4][2]  <= n969;
    \\i_tv80_core_i_reg_RegsL_reg[6][0]  <= n974;
    \\i_tv80_core_SP_reg[12]  <= n979;
    \\i_tv80_core_F_reg[7]  <= n984;
    \\i_tv80_core_SP_reg[15]  <= n989;
    \\i_tv80_core_F_reg[3]  <= n994;
    \\i_tv80_core_F_reg[5]  <= n999;
    \\i_tv80_core_SP_reg[10]  <= n1004;
    \\i_tv80_core_SP_reg[13]  <= n1009;
    \\i_tv80_core_F_reg[4]  <= n1014;
    \\i_tv80_core_SP_reg[9]  <= n1019;
    \\i_tv80_core_SP_reg[11]  <= n1024;
    \\i_tv80_core_SP_reg[8]  <= n1029;
    \\i_tv80_core_mcycle_reg[1]  <= n1034;
    \\i_tv80_core_mcycle_reg[2]  <= n1039;
    \\i_tv80_core_mcycle_reg[0]  <= n1044;
    \\i_tv80_core_TmpAddr_reg[14]  <= n1049;
    i_tv80_core_IntE_FF1_reg <= n1054;
    i_tv80_core_IntE_FF2_reg <= n1059;
    i_tv80_core_m1_n_reg <= n1064;
    i_tv80_core_IntCycle_reg <= n1069;
    i_tv80_core_NMICycle_reg <= n1074;
    \\i_tv80_core_BusA_reg[0]  <= n1079;
    \\i_tv80_core_BusA_reg[5]  <= n1084;
    \\i_tv80_core_PC_reg[9]  <= n1089;
    \\i_tv80_core_PC_reg[7]  <= n1094;
    \\i_tv80_core_Pre_XY_F_M_reg[2]  <= n1099;
    \\i_tv80_core_BusA_reg[3]  <= n1104;
    \\i_tv80_core_PC_reg[11]  <= n1109;
    \\i_tv80_core_PC_reg[12]  <= n1114;
    \\i_tv80_core_PC_reg[13]  <= n1119;
    \\i_tv80_core_PC_reg[1]  <= n1124;
    \\i_tv80_core_PC_reg[2]  <= n1129;
    \\i_tv80_core_PC_reg[3]  <= n1134;
    \\i_tv80_core_PC_reg[4]  <= n1139;
    \\i_tv80_core_PC_reg[5]  <= n1144;
    \\i_tv80_core_PC_reg[6]  <= n1149;
    \\i_tv80_core_PC_reg[8]  <= n1154;
    \\i_tv80_core_Pre_XY_F_M_reg[0]  <= n1159;
    \\i_tv80_core_Pre_XY_F_M_reg[1]  <= n1164;
    \\i_tv80_core_BusA_reg[2]  <= n1169;
    \\i_tv80_core_BusA_reg[4]  <= n1174;
    \\i_tv80_core_BusA_reg[6]  <= n1179;
    \\i_tv80_core_PC_reg[15]  <= n1184;
    \\i_tv80_core_PC_reg[14]  <= n1189;
    \\i_tv80_core_PC_reg[0]  <= n1194;
    \\i_tv80_core_PC_reg[10]  <= n1199;
    \\i_tv80_core_TmpAddr_reg[10]  <= n1204;
    \\i_tv80_core_BusA_reg[7]  <= n1209;
    \\i_tv80_core_TmpAddr_reg[15]  <= n1214;
    \\i_tv80_core_BusA_reg[1]  <= n1219;
    \\i_tv80_core_TmpAddr_reg[12]  <= n1224;
    \\i_tv80_core_TmpAddr_reg[13]  <= n1229;
    i_tv80_core_BTR_r_reg <= n1234;
    \\i_tv80_core_TmpAddr_reg[11]  <= n1239;
    i_tv80_core_Halt_FF_reg <= n1244;
    \\i_tv80_core_Read_To_Reg_r_reg[4]  <= n1249;
    \\i_tv80_core_TmpAddr_reg[9]  <= n1254;
    \\i_tv80_core_TmpAddr_reg[6]  <= n1259;
    \\i_tv80_core_Read_To_Reg_r_reg[2]  <= n1264;
    \\i_tv80_core_RegBusA_r_reg[0]  <= n1269;
    \\i_tv80_core_RegBusA_r_reg[13]  <= n1274;
    i_tv80_core_Auto_Wait_t2_reg <= n1279;
    \\i_tv80_core_TmpAddr_reg[8]  <= n1284;
    \\i_tv80_core_Read_To_Reg_r_reg[0]  <= n1289;
    \\i_tv80_core_Read_To_Reg_r_reg[1]  <= n1294;
    \\i_tv80_core_ALU_Op_r_reg[1]  <= n1299;
    i_tv80_core_Save_ALU_r_reg <= n1304;
    \\i_tv80_core_ALU_Op_r_reg[3]  <= n1309;
    \\i_tv80_core_TmpAddr_reg[7]  <= n1314;
    \\i_tv80_core_RegBusA_r_reg[11]  <= n1319;
    \\i_tv80_core_TmpAddr_reg[5]  <= n1324;
    i_tv80_core_BusAck_reg <= n1329;
    \\i_tv80_core_RegBusA_r_reg[10]  <= n1334;
    \\i_tv80_core_RegBusA_r_reg[12]  <= n1339;
    \\i_tv80_core_RegBusA_r_reg[14]  <= n1344;
    \\i_tv80_core_Read_To_Reg_r_reg[3]  <= n1349;
    i_tv80_core_Auto_Wait_t1_reg <= n1354;
    \\i_tv80_core_RegBusA_r_reg[15]  <= n1359;
    \\i_tv80_core_RegBusA_r_reg[7]  <= n1364;
    \\i_tv80_core_RegBusA_r_reg[9]  <= n1369;
    \\i_tv80_core_ALU_Op_r_reg[2]  <= n1374;
    \\i_tv80_core_ALU_Op_r_reg[0]  <= n1379;
    \\i_tv80_core_RegBusA_r_reg[8]  <= n1384;
    \\i_tv80_core_TmpAddr_reg[4]  <= n1389;
    \\i_tv80_core_RegBusA_r_reg[1]  <= n1394;
    \\i_tv80_core_RegBusA_r_reg[2]  <= n1399;
    \\i_tv80_core_RegBusA_r_reg[5]  <= n1404;
    \\i_tv80_core_RegBusA_r_reg[6]  <= n1409;
    \\i_tv80_core_BusB_reg[0]  <= n1414;
    \\i_tv80_core_TmpAddr_reg[3]  <= n1419;
    \\i_tv80_core_RegBusA_r_reg[4]  <= n1424;
    \\i_tv80_core_RegBusA_r_reg[3]  <= n1429;
    \\i_tv80_core_TmpAddr_reg[2]  <= n1434;
    \\i_tv80_core_BusB_reg[6]  <= n1439;
    \\i_tv80_core_BusB_reg[4]  <= n1444;
    \\i_tv80_core_BusB_reg[1]  <= n1449;
    \\i_tv80_core_BusB_reg[3]  <= n1454;
    \\i_tv80_core_BusB_reg[5]  <= n1459;
    \\i_tv80_core_BusB_reg[2]  <= n1464;
    \\i_tv80_core_BusB_reg[7]  <= n1469;
    \\i_tv80_core_TmpAddr_reg[1]  <= n1474;
    \\i_tv80_core_RegAddrC_reg[1]  <= n1479;
    i_tv80_core_Z16_r_reg <= n1484;
    iorq_n_reg <= n1489;
    \\i_tv80_core_RegAddrB_r_reg[2]  <= n1494;
    mreq_n_reg <= n1499;
    \\i_tv80_core_TmpAddr_reg[0]  <= n1504;
    \\i_tv80_core_RegAddrB_r_reg[0]  <= n1509;
    \\i_tv80_core_RegAddrB_r_reg[1]  <= n1514;
    \\i_tv80_core_RegAddrC_reg[0]  <= n1519;
    \\i_tv80_core_R_reg[6]  <= n1524;
    \\i_tv80_core_R_reg[5]  <= n1529;
    \\i_tv80_core_R_reg[3]  <= n1534;
    \\i_tv80_core_R_reg[2]  <= n1539;
    \\i_tv80_core_R_reg[4]  <= n1544;
    \\i_tv80_core_IR_reg[2]  <= n1549;
    \\i_tv80_core_R_reg[0]  <= n1554;
    rd_n_reg <= n1559;
    \\i_tv80_core_ISet_reg[0]  <= n1564;
    \\i_tv80_core_R_reg[1]  <= n1569;
    \\i_tv80_core_IR_reg[0]  <= n1574;
    \\i_tv80_core_IR_reg[1]  <= n1579;
    \\i_tv80_core_IR_reg[5]  <= n1584;
    \\i_tv80_core_IR_reg[6]  <= n1589;
    \\i_tv80_core_IR_reg[7]  <= n1594;
    \\i_tv80_core_ISet_reg[1]  <= n1599;
    \\i_tv80_core_IR_reg[4]  <= n1604;
    \\i_tv80_core_IR_reg[3]  <= n1609;
    i_tv80_core_Alternate_reg <= n1614;
    i_tv80_core_XY_Ind_reg <= n1619;
    wr_n_reg <= n1624;
    \\i_tv80_core_mcycles_reg[0]  <= n1629;
    \\i_tv80_core_mcycles_reg[2]  <= n1634;
    \\i_tv80_core_RegAddrA_r_reg[1]  <= n1639;
    \\i_tv80_core_mcycles_reg[1]  <= n1644;
    \\i_tv80_core_RegAddrA_r_reg[2]  <= n1649;
    \\i_tv80_core_RegAddrA_r_reg[0]  <= n1654;
    \\i_tv80_core_XY_State_reg[0]  <= n1659;
    \\i_tv80_core_XY_State_reg[1]  <= n1664;
    \\i_tv80_core_Fp_reg[5]  <= n1669;
    \\i_tv80_core_Ap_reg[3]  <= n1674;
    \\i_tv80_core_Ap_reg[5]  <= n1679;
    \\i_tv80_core_Fp_reg[7]  <= n1684;
    \\i_tv80_core_Ap_reg[1]  <= n1689;
    \\i_tv80_core_Fp_reg[1]  <= n1694;
    \\i_tv80_core_Fp_reg[3]  <= n1699;
    \\i_tv80_core_Fp_reg[0]  <= n1704;
    \\i_tv80_core_Fp_reg[2]  <= n1709;
    \\i_tv80_core_Fp_reg[4]  <= n1714;
    \\i_tv80_core_Fp_reg[6]  <= n1719;
    \\i_tv80_core_Ap_reg[0]  <= n1724;
    \\i_tv80_core_Ap_reg[2]  <= n1729;
    \\i_tv80_core_Ap_reg[4]  <= n1734;
    \\i_tv80_core_Ap_reg[6]  <= n1739;
    \\i_tv80_core_Ap_reg[7]  <= n1744;
    \\i_tv80_core_IStatus_reg[1]  <= n1749;
    \\i_tv80_core_R_reg[7]  <= n1754;
    \\i_tv80_core_IStatus_reg[0]  <= n1759;
    i_tv80_core_rfsh_n_reg <= n1764;
    i_tv80_core_PreserveC_r_reg <= n1769;
    \\i_tv80_core_I_reg[5]  <= n1774;
    \\i_tv80_core_I_reg[2]  <= n1779;
    \\i_tv80_core_I_reg[4]  <= n1784;
    \\i_tv80_core_I_reg[7]  <= n1789;
    \\i_tv80_core_I_reg[6]  <= n1794;
    \\i_tv80_core_I_reg[0]  <= n1799;
    \\i_tv80_core_I_reg[1]  <= n1804;
    \\i_tv80_core_I_reg[3]  <= n1809;
    i_tv80_core_Arith16_r_reg <= n1814;
    i_tv80_core_No_BTR_reg <= n1819;
    \\i_tv80_core_RegAddrC_reg[2]  <= n1824;
    \\di_reg_reg[6]  <= n1829;
    \\di_reg_reg[3]  <= n1834;
    \\di_reg_reg[1]  <= n1839;
    \\di_reg_reg[7]  <= n1844;
    \\di_reg_reg[2]  <= n1849;
    \\di_reg_reg[4]  <= n1854;
    \\di_reg_reg[5]  <= n1859;
    \\di_reg_reg[0]  <= n1864;
    i_tv80_core_NMI_s_reg <= n1869;
    i_tv80_core_BusReq_s_reg <= n1874;
    i_tv80_core_Oldnmi_n_reg <= n1879;
    i_tv80_core_INT_s_reg <= n1884;
  end
endmodule


