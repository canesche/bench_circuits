module top ( 
    pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv56_13_, pv56_22_, pv88_7_,
    pv88_29_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_, pv56_15_,
    pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv9_5_, pv56_30_, pv88_2_,
    pv88_15_, pv88_26_, pv9_6_, pv24_10_, pv56_31_, pv88_3_, pv88_16_,
    pv88_25_, pv9_7_, pv9_10_, pv56_10_, pv56_21_, pv88_4_, pv88_13_,
    pv88_24_, pv9_8_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_,
    pv56_5_, pv88_11_, pv88_22_, pv56_4_, pv88_12_, pv88_21_, pv56_7_,
    pv88_20_, pv56_6_, pv88_10_, pv24_8_, pv56_9_, pv24_9_, pv56_8_,
    pv24_6_, pv24_7_, pv24_4_, pv24_5_, pv24_2_, pv24_3_, pv24_0_, pv56_1_,
    pv24_1_, pv56_0_, pv88_30_, pv56_3_, pv88_31_, pv56_2_, pv9_1_,
    pv24_13_, pv9_2_, pv24_14_, pv9_3_, pv24_11_, pv88_0_, pv24_12_,
    pv88_1_, pv56_16_, pv56_27_, pv56_17_, pv56_26_, pv56_18_, pv56_29_,
    pv9_0_, pv56_19_, pv56_28_,
    pv119_1_, pv119_0_, pv119_3_, pv119_30_, pv119_2_, pv151_1_, pv151_18_,
    pv151_0_, pv151_19_, pv119_21_, pv151_3_, pv151_16_, pv119_20_,
    pv151_2_, pv151_17_, pv119_9_, pv119_23_, pv151_27_, pv119_8_,
    pv119_22_, pv151_26_, pv119_25_, pv151_29_, pv119_24_, pv151_28_,
    pv119_5_, pv119_27_, pv119_4_, pv119_26_, pv119_7_, pv119_29_,
    pv119_6_, pv119_28_, pv119_18_, pv119_19_, pv119_16_, pv151_21_,
    pv119_17_, pv151_20_, pv119_14_, pv151_23_, pv119_15_, pv151_22_,
    pv119_12_, pv151_25_, pv151_30_, pv119_13_, pv151_24_, pv151_31_,
    pv119_10_, pv151_5_, pv151_14_, pv119_11_, pv151_4_, pv151_15_,
    pv151_7_, pv151_12_, pv151_6_, pv151_13_, pv151_9_, pv151_10_,
    pv151_8_, pv151_11_  );
  input  pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv56_13_, pv56_22_,
    pv88_7_, pv88_29_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_,
    pv56_15_, pv56_24_, pv88_9_, pv88_18_, pv88_27_, pv9_5_, pv56_30_,
    pv88_2_, pv88_15_, pv88_26_, pv9_6_, pv24_10_, pv56_31_, pv88_3_,
    pv88_16_, pv88_25_, pv9_7_, pv9_10_, pv56_10_, pv56_21_, pv88_4_,
    pv88_13_, pv88_24_, pv9_8_, pv56_11_, pv56_20_, pv88_5_, pv88_14_,
    pv88_23_, pv56_5_, pv88_11_, pv88_22_, pv56_4_, pv88_12_, pv88_21_,
    pv56_7_, pv88_20_, pv56_6_, pv88_10_, pv24_8_, pv56_9_, pv24_9_,
    pv56_8_, pv24_6_, pv24_7_, pv24_4_, pv24_5_, pv24_2_, pv24_3_, pv24_0_,
    pv56_1_, pv24_1_, pv56_0_, pv88_30_, pv56_3_, pv88_31_, pv56_2_,
    pv9_1_, pv24_13_, pv9_2_, pv24_14_, pv9_3_, pv24_11_, pv88_0_,
    pv24_12_, pv88_1_, pv56_16_, pv56_27_, pv56_17_, pv56_26_, pv56_18_,
    pv56_29_, pv9_0_, pv56_19_, pv56_28_;
  output pv119_1_, pv119_0_, pv119_3_, pv119_30_, pv119_2_, pv151_1_,
    pv151_18_, pv151_0_, pv151_19_, pv119_21_, pv151_3_, pv151_16_,
    pv119_20_, pv151_2_, pv151_17_, pv119_9_, pv119_23_, pv151_27_,
    pv119_8_, pv119_22_, pv151_26_, pv119_25_, pv151_29_, pv119_24_,
    pv151_28_, pv119_5_, pv119_27_, pv119_4_, pv119_26_, pv119_7_,
    pv119_29_, pv119_6_, pv119_28_, pv119_18_, pv119_19_, pv119_16_,
    pv151_21_, pv119_17_, pv151_20_, pv119_14_, pv151_23_, pv119_15_,
    pv151_22_, pv119_12_, pv151_25_, pv151_30_, pv119_13_, pv151_24_,
    pv151_31_, pv119_10_, pv151_5_, pv151_14_, pv119_11_, pv151_4_,
    pv151_15_, pv151_7_, pv151_12_, pv151_6_, pv151_13_, pv151_9_,
    pv151_10_, pv151_8_, pv151_11_;
  wire new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_,
    new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_;
  assign new_n152_ = pv9_8_ & pv9_1_;
  assign new_n153_ = ~pv9_10_ & new_n152_;
  assign new_n154_ = ~pv9_6_ & ~pv9_2_;
  assign new_n155_ = ~pv9_5_ & new_n154_;
  assign new_n156_ = pv9_1_ & new_n155_;
  assign new_n157_ = ~pv9_10_ & new_n156_;
  assign new_n158_ = pv9_2_ & pv9_0_;
  assign new_n159_ = ~pv9_5_ & new_n158_;
  assign new_n160_ = ~pv9_1_ & new_n159_;
  assign new_n161_ = ~pv9_10_ & new_n160_;
  assign new_n162_ = ~pv9_6_ & new_n161_;
  assign new_n163_ = pv9_2_ & ~pv9_3_;
  assign new_n164_ = pv9_1_ & new_n163_;
  assign new_n165_ = ~pv9_10_ & new_n164_;
  assign new_n166_ = pv9_8_ & pv9_2_;
  assign new_n167_ = ~pv9_1_ & new_n166_;
  assign new_n168_ = ~pv9_10_ & new_n167_;
  assign new_n169_ = ~pv9_1_ & ~pv9_2_;
  assign new_n170_ = pv9_10_ & new_n169_;
  assign new_n171_ = ~pv9_5_ & ~pv9_2_;
  assign new_n172_ = ~pv9_1_ & new_n171_;
  assign new_n173_ = ~pv9_6_ & new_n172_;
  assign new_n174_ = pv9_7_ & new_n169_;
  assign new_n175_ = pv9_10_ & pv9_2_;
  assign new_n176_ = pv9_1_ & pv9_2_;
  assign new_n177_ = pv9_3_ & new_n176_;
  assign new_n178_ = pv9_10_ & pv9_1_;
  assign new_n179_ = ~pv9_5_ & ~pv9_0_;
  assign new_n180_ = ~pv9_10_ & new_n179_;
  assign new_n181_ = pv9_7_ & ~pv9_0_;
  assign new_n182_ = ~pv9_10_ & new_n181_;
  assign new_n183_ = ~new_n153_ & ~new_n157_;
  assign new_n184_ = ~new_n162_ & ~new_n165_;
  assign new_n185_ = new_n183_ & new_n184_;
  assign new_n186_ = ~new_n168_ & ~new_n170_;
  assign new_n187_ = ~new_n173_ & new_n186_;
  assign new_n188_ = new_n185_ & new_n187_;
  assign new_n189_ = ~new_n178_ & ~new_n180_;
  assign new_n190_ = ~new_n182_ & new_n189_;
  assign new_n191_ = ~new_n174_ & ~new_n175_;
  assign new_n192_ = ~new_n177_ & new_n191_;
  assign new_n193_ = new_n190_ & new_n192_;
  assign new_n194_ = new_n188_ & new_n193_;
  assign new_n195_ = ~new_n157_ & ~new_n180_;
  assign new_n196_ = ~new_n173_ & ~new_n174_;
  assign new_n197_ = new_n195_ & new_n196_;
  assign new_n198_ = ~new_n170_ & ~new_n182_;
  assign new_n199_ = ~new_n153_ & new_n198_;
  assign new_n200_ = new_n197_ & new_n199_;
  assign new_n201_ = ~new_n170_ & ~new_n174_;
  assign new_n202_ = ~new_n168_ & new_n201_;
  assign new_n203_ = ~new_n173_ & new_n184_;
  assign new_n204_ = new_n202_ & new_n203_;
  assign new_n205_ = ~new_n194_ & new_n200_;
  assign new_n206_ = new_n204_ & new_n205_;
  assign new_n207_ = pv56_2_ & new_n206_;
  assign new_n208_ = ~new_n204_ & new_n205_;
  assign new_n209_ = pv88_2_ & new_n208_;
  assign new_n210_ = ~new_n200_ & new_n204_;
  assign new_n211_ = ~new_n194_ & new_n210_;
  assign new_n212_ = ~new_n194_ & ~new_n200_;
  assign new_n213_ = ~new_n204_ & new_n212_;
  assign new_n214_ = pv24_1_ & new_n213_;
  assign new_n215_ = ~new_n211_ & ~new_n214_;
  assign new_n216_ = ~new_n194_ & ~new_n207_;
  assign new_n217_ = ~new_n209_ & new_n216_;
  assign pv119_1_ = ~new_n215_ | ~new_n217_;
  assign new_n219_ = pv56_1_ & new_n206_;
  assign new_n220_ = pv88_1_ & new_n208_;
  assign new_n221_ = pv24_0_ & new_n213_;
  assign new_n222_ = ~new_n211_ & ~new_n221_;
  assign new_n223_ = ~new_n194_ & ~new_n219_;
  assign new_n224_ = ~new_n220_ & new_n223_;
  assign pv119_0_ = ~new_n222_ | ~new_n224_;
  assign new_n226_ = pv56_4_ & new_n206_;
  assign new_n227_ = pv88_4_ & new_n208_;
  assign new_n228_ = pv24_3_ & new_n213_;
  assign new_n229_ = ~new_n211_ & ~new_n228_;
  assign new_n230_ = ~new_n194_ & ~new_n226_;
  assign new_n231_ = ~new_n227_ & new_n230_;
  assign pv119_3_ = ~new_n229_ | ~new_n231_;
  assign new_n233_ = pv56_31_ & new_n206_;
  assign new_n234_ = pv56_20_ & new_n208_;
  assign new_n235_ = pv56_23_ & new_n211_;
  assign new_n236_ = pv56_16_ & new_n213_;
  assign new_n237_ = ~new_n235_ & ~new_n236_;
  assign new_n238_ = ~new_n194_ & ~new_n233_;
  assign new_n239_ = ~new_n234_ & new_n238_;
  assign pv119_30_ = ~new_n237_ | ~new_n239_;
  assign new_n241_ = pv56_3_ & new_n206_;
  assign new_n242_ = pv88_3_ & new_n208_;
  assign new_n243_ = pv24_2_ & new_n213_;
  assign new_n244_ = ~new_n211_ & ~new_n243_;
  assign new_n245_ = ~new_n194_ & ~new_n241_;
  assign new_n246_ = ~new_n242_ & new_n245_;
  assign pv119_2_ = ~new_n244_ | ~new_n246_;
  assign new_n248_ = pv88_1_ & new_n206_;
  assign new_n249_ = ~new_n200_ & ~new_n204_;
  assign new_n250_ = new_n194_ & new_n249_;
  assign new_n251_ = pv56_22_ & new_n208_;
  assign new_n252_ = new_n204_ & new_n212_;
  assign new_n253_ = pv56_25_ & new_n252_;
  assign new_n254_ = pv56_18_ & new_n213_;
  assign new_n255_ = new_n200_ & new_n204_;
  assign new_n256_ = new_n194_ & new_n255_;
  assign new_n257_ = new_n200_ & ~new_n204_;
  assign new_n258_ = new_n194_ & new_n257_;
  assign new_n259_ = new_n194_ & new_n210_;
  assign new_n260_ = ~new_n258_ & ~new_n259_;
  assign new_n261_ = ~new_n254_ & ~new_n256_;
  assign new_n262_ = new_n260_ & new_n261_;
  assign new_n263_ = ~new_n248_ & ~new_n250_;
  assign new_n264_ = ~new_n251_ & ~new_n253_;
  assign new_n265_ = new_n263_ & new_n264_;
  assign pv151_1_ = ~new_n262_ | ~new_n265_;
  assign new_n267_ = pv88_18_ & new_n206_;
  assign new_n268_ = pv88_7_ & new_n208_;
  assign new_n269_ = pv88_10_ & new_n252_;
  assign new_n270_ = pv88_3_ & new_n213_;
  assign new_n271_ = ~new_n256_ & ~new_n270_;
  assign new_n272_ = new_n260_ & new_n271_;
  assign new_n273_ = ~new_n250_ & ~new_n267_;
  assign new_n274_ = ~new_n268_ & ~new_n269_;
  assign new_n275_ = new_n273_ & new_n274_;
  assign pv151_18_ = ~new_n272_ | ~new_n275_;
  assign new_n277_ = pv88_0_ & new_n206_;
  assign new_n278_ = pv56_21_ & new_n208_;
  assign new_n279_ = pv56_24_ & new_n252_;
  assign new_n280_ = pv56_17_ & new_n213_;
  assign new_n281_ = ~new_n256_ & ~new_n280_;
  assign new_n282_ = new_n260_ & new_n281_;
  assign new_n283_ = ~new_n250_ & ~new_n277_;
  assign new_n284_ = ~new_n278_ & ~new_n279_;
  assign new_n285_ = new_n283_ & new_n284_;
  assign pv151_0_ = ~new_n282_ | ~new_n285_;
  assign new_n287_ = pv88_19_ & new_n206_;
  assign new_n288_ = pv88_8_ & new_n208_;
  assign new_n289_ = pv88_11_ & new_n252_;
  assign new_n290_ = pv88_4_ & new_n213_;
  assign new_n291_ = ~new_n256_ & ~new_n290_;
  assign new_n292_ = new_n260_ & new_n291_;
  assign new_n293_ = ~new_n250_ & ~new_n287_;
  assign new_n294_ = ~new_n288_ & ~new_n289_;
  assign new_n295_ = new_n293_ & new_n294_;
  assign pv151_19_ = ~new_n292_ | ~new_n295_;
  assign new_n297_ = pv56_22_ & new_n206_;
  assign new_n298_ = pv56_11_ & new_n208_;
  assign new_n299_ = pv56_14_ & new_n211_;
  assign new_n300_ = pv56_7_ & new_n213_;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = ~new_n194_ & ~new_n297_;
  assign new_n303_ = ~new_n298_ & new_n302_;
  assign pv119_21_ = ~new_n301_ | ~new_n303_;
  assign new_n305_ = pv88_3_ & new_n206_;
  assign new_n306_ = pv56_24_ & new_n208_;
  assign new_n307_ = pv56_27_ & new_n252_;
  assign new_n308_ = pv56_20_ & new_n213_;
  assign new_n309_ = ~new_n256_ & ~new_n308_;
  assign new_n310_ = new_n260_ & new_n309_;
  assign new_n311_ = ~new_n250_ & ~new_n305_;
  assign new_n312_ = ~new_n306_ & ~new_n307_;
  assign new_n313_ = new_n311_ & new_n312_;
  assign pv151_3_ = ~new_n310_ | ~new_n313_;
  assign new_n315_ = pv88_16_ & new_n206_;
  assign new_n316_ = pv88_5_ & new_n208_;
  assign new_n317_ = pv88_8_ & new_n252_;
  assign new_n318_ = pv88_1_ & new_n213_;
  assign new_n319_ = ~new_n256_ & ~new_n318_;
  assign new_n320_ = new_n260_ & new_n319_;
  assign new_n321_ = ~new_n250_ & ~new_n315_;
  assign new_n322_ = ~new_n316_ & ~new_n317_;
  assign new_n323_ = new_n321_ & new_n322_;
  assign pv151_16_ = ~new_n320_ | ~new_n323_;
  assign new_n325_ = pv56_21_ & new_n206_;
  assign new_n326_ = pv56_10_ & new_n208_;
  assign new_n327_ = pv56_13_ & new_n211_;
  assign new_n328_ = pv56_6_ & new_n213_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~new_n194_ & ~new_n325_;
  assign new_n331_ = ~new_n326_ & new_n330_;
  assign pv119_20_ = ~new_n329_ | ~new_n331_;
  assign new_n333_ = pv88_2_ & new_n206_;
  assign new_n334_ = pv56_23_ & new_n208_;
  assign new_n335_ = pv56_26_ & new_n252_;
  assign new_n336_ = pv56_19_ & new_n213_;
  assign new_n337_ = ~new_n256_ & ~new_n336_;
  assign new_n338_ = new_n260_ & new_n337_;
  assign new_n339_ = ~new_n250_ & ~new_n333_;
  assign new_n340_ = ~new_n334_ & ~new_n335_;
  assign new_n341_ = new_n339_ & new_n340_;
  assign pv151_2_ = ~new_n338_ | ~new_n341_;
  assign new_n343_ = pv88_17_ & new_n206_;
  assign new_n344_ = pv88_6_ & new_n208_;
  assign new_n345_ = pv88_9_ & new_n252_;
  assign new_n346_ = pv88_2_ & new_n213_;
  assign new_n347_ = ~new_n256_ & ~new_n346_;
  assign new_n348_ = new_n260_ & new_n347_;
  assign new_n349_ = ~new_n250_ & ~new_n343_;
  assign new_n350_ = ~new_n344_ & ~new_n345_;
  assign new_n351_ = new_n349_ & new_n350_;
  assign pv151_17_ = ~new_n348_ | ~new_n351_;
  assign new_n353_ = pv56_10_ & new_n206_;
  assign new_n354_ = pv88_10_ & new_n208_;
  assign new_n355_ = pv56_2_ & new_n211_;
  assign new_n356_ = pv24_9_ & new_n213_;
  assign new_n357_ = ~new_n355_ & ~new_n356_;
  assign new_n358_ = ~new_n194_ & ~new_n353_;
  assign new_n359_ = ~new_n354_ & new_n358_;
  assign pv119_9_ = ~new_n357_ | ~new_n359_;
  assign new_n361_ = pv56_24_ & new_n206_;
  assign new_n362_ = pv56_13_ & new_n208_;
  assign new_n363_ = pv56_16_ & new_n211_;
  assign new_n364_ = pv56_9_ & new_n213_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = ~new_n194_ & ~new_n361_;
  assign new_n367_ = ~new_n362_ & new_n366_;
  assign pv119_23_ = ~new_n365_ | ~new_n367_;
  assign new_n369_ = pv88_27_ & new_n206_;
  assign new_n370_ = pv88_16_ & new_n208_;
  assign new_n371_ = pv88_19_ & new_n252_;
  assign new_n372_ = pv88_12_ & new_n213_;
  assign new_n373_ = ~new_n256_ & ~new_n372_;
  assign new_n374_ = new_n260_ & new_n373_;
  assign new_n375_ = ~new_n250_ & ~new_n369_;
  assign new_n376_ = ~new_n370_ & ~new_n371_;
  assign new_n377_ = new_n375_ & new_n376_;
  assign pv151_27_ = ~new_n374_ | ~new_n377_;
  assign new_n379_ = pv56_9_ & new_n206_;
  assign new_n380_ = pv88_9_ & new_n208_;
  assign new_n381_ = pv56_1_ & new_n211_;
  assign new_n382_ = pv24_8_ & new_n213_;
  assign new_n383_ = ~new_n381_ & ~new_n382_;
  assign new_n384_ = ~new_n194_ & ~new_n379_;
  assign new_n385_ = ~new_n380_ & new_n384_;
  assign pv119_8_ = ~new_n383_ | ~new_n385_;
  assign new_n387_ = pv56_23_ & new_n206_;
  assign new_n388_ = pv56_12_ & new_n208_;
  assign new_n389_ = pv56_15_ & new_n211_;
  assign new_n390_ = pv56_8_ & new_n213_;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = ~new_n194_ & ~new_n387_;
  assign new_n393_ = ~new_n388_ & new_n392_;
  assign pv119_22_ = ~new_n391_ | ~new_n393_;
  assign new_n395_ = pv88_26_ & new_n206_;
  assign new_n396_ = pv88_15_ & new_n208_;
  assign new_n397_ = pv88_18_ & new_n252_;
  assign new_n398_ = pv88_11_ & new_n213_;
  assign new_n399_ = ~new_n256_ & ~new_n398_;
  assign new_n400_ = new_n260_ & new_n399_;
  assign new_n401_ = ~new_n250_ & ~new_n395_;
  assign new_n402_ = ~new_n396_ & ~new_n397_;
  assign new_n403_ = new_n401_ & new_n402_;
  assign pv151_26_ = ~new_n400_ | ~new_n403_;
  assign new_n405_ = pv56_26_ & new_n206_;
  assign new_n406_ = pv56_15_ & new_n208_;
  assign new_n407_ = pv56_18_ & new_n211_;
  assign new_n408_ = pv56_11_ & new_n213_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = ~new_n194_ & ~new_n405_;
  assign new_n411_ = ~new_n406_ & new_n410_;
  assign pv119_25_ = ~new_n409_ | ~new_n411_;
  assign new_n413_ = pv88_29_ & new_n206_;
  assign new_n414_ = pv88_18_ & new_n208_;
  assign new_n415_ = pv88_21_ & new_n252_;
  assign new_n416_ = pv88_14_ & new_n213_;
  assign new_n417_ = ~new_n256_ & ~new_n416_;
  assign new_n418_ = new_n260_ & new_n417_;
  assign new_n419_ = ~new_n250_ & ~new_n413_;
  assign new_n420_ = ~new_n414_ & ~new_n415_;
  assign new_n421_ = new_n419_ & new_n420_;
  assign pv151_29_ = ~new_n418_ | ~new_n421_;
  assign new_n423_ = pv56_25_ & new_n206_;
  assign new_n424_ = pv56_14_ & new_n208_;
  assign new_n425_ = pv56_17_ & new_n211_;
  assign new_n426_ = pv56_10_ & new_n213_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = ~new_n194_ & ~new_n423_;
  assign new_n429_ = ~new_n424_ & new_n428_;
  assign pv119_24_ = ~new_n427_ | ~new_n429_;
  assign new_n431_ = pv88_28_ & new_n206_;
  assign new_n432_ = pv88_17_ & new_n208_;
  assign new_n433_ = pv88_20_ & new_n252_;
  assign new_n434_ = pv88_13_ & new_n213_;
  assign new_n435_ = ~new_n256_ & ~new_n434_;
  assign new_n436_ = new_n260_ & new_n435_;
  assign new_n437_ = ~new_n250_ & ~new_n431_;
  assign new_n438_ = ~new_n432_ & ~new_n433_;
  assign new_n439_ = new_n437_ & new_n438_;
  assign pv151_28_ = ~new_n436_ | ~new_n439_;
  assign new_n441_ = pv56_6_ & new_n206_;
  assign new_n442_ = pv24_5_ & new_n213_;
  assign new_n443_ = ~new_n211_ & ~new_n442_;
  assign new_n444_ = ~new_n194_ & ~new_n441_;
  assign new_n445_ = ~new_n344_ & new_n444_;
  assign pv119_5_ = ~new_n443_ | ~new_n445_;
  assign new_n447_ = pv56_28_ & new_n206_;
  assign new_n448_ = pv56_17_ & new_n208_;
  assign new_n449_ = pv56_20_ & new_n211_;
  assign new_n450_ = pv56_13_ & new_n213_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = ~new_n194_ & ~new_n447_;
  assign new_n453_ = ~new_n448_ & new_n452_;
  assign pv119_27_ = ~new_n451_ | ~new_n453_;
  assign new_n455_ = pv56_5_ & new_n206_;
  assign new_n456_ = pv24_4_ & new_n213_;
  assign new_n457_ = ~new_n211_ & ~new_n456_;
  assign new_n458_ = ~new_n194_ & ~new_n455_;
  assign new_n459_ = ~new_n316_ & new_n458_;
  assign pv119_4_ = ~new_n457_ | ~new_n459_;
  assign new_n461_ = pv56_27_ & new_n206_;
  assign new_n462_ = pv56_16_ & new_n208_;
  assign new_n463_ = pv56_19_ & new_n211_;
  assign new_n464_ = pv56_12_ & new_n213_;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign new_n466_ = ~new_n194_ & ~new_n461_;
  assign new_n467_ = ~new_n462_ & new_n466_;
  assign pv119_26_ = ~new_n465_ | ~new_n467_;
  assign new_n469_ = pv56_8_ & new_n206_;
  assign new_n470_ = pv56_0_ & new_n211_;
  assign new_n471_ = pv24_7_ & new_n213_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = ~new_n194_ & ~new_n469_;
  assign new_n474_ = ~new_n288_ & new_n473_;
  assign pv119_7_ = ~new_n472_ | ~new_n474_;
  assign new_n476_ = pv56_30_ & new_n206_;
  assign new_n477_ = pv56_19_ & new_n208_;
  assign new_n478_ = pv56_22_ & new_n211_;
  assign new_n479_ = pv56_15_ & new_n213_;
  assign new_n480_ = ~new_n478_ & ~new_n479_;
  assign new_n481_ = ~new_n194_ & ~new_n476_;
  assign new_n482_ = ~new_n477_ & new_n481_;
  assign pv119_29_ = ~new_n480_ | ~new_n482_;
  assign new_n484_ = pv56_7_ & new_n206_;
  assign new_n485_ = pv24_6_ & new_n213_;
  assign new_n486_ = ~new_n211_ & ~new_n485_;
  assign new_n487_ = ~new_n194_ & ~new_n484_;
  assign new_n488_ = ~new_n268_ & new_n487_;
  assign pv119_6_ = ~new_n486_ | ~new_n488_;
  assign new_n490_ = pv56_29_ & new_n206_;
  assign new_n491_ = pv56_18_ & new_n208_;
  assign new_n492_ = pv56_21_ & new_n211_;
  assign new_n493_ = pv56_14_ & new_n213_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = ~new_n194_ & ~new_n490_;
  assign new_n496_ = ~new_n491_ & new_n495_;
  assign pv119_28_ = ~new_n494_ | ~new_n496_;
  assign new_n498_ = pv56_19_ & new_n206_;
  assign new_n499_ = pv56_8_ & new_n208_;
  assign new_n500_ = pv56_11_ & new_n211_;
  assign new_n501_ = pv56_4_ & new_n213_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~new_n194_ & ~new_n498_;
  assign new_n504_ = ~new_n499_ & new_n503_;
  assign pv119_18_ = ~new_n502_ | ~new_n504_;
  assign new_n506_ = pv56_20_ & new_n206_;
  assign new_n507_ = pv56_9_ & new_n208_;
  assign new_n508_ = pv56_12_ & new_n211_;
  assign new_n509_ = pv56_5_ & new_n213_;
  assign new_n510_ = ~new_n508_ & ~new_n509_;
  assign new_n511_ = ~new_n194_ & ~new_n506_;
  assign new_n512_ = ~new_n507_ & new_n511_;
  assign pv119_19_ = ~new_n510_ | ~new_n512_;
  assign new_n514_ = pv56_17_ & new_n206_;
  assign new_n515_ = pv56_6_ & new_n208_;
  assign new_n516_ = pv56_9_ & new_n211_;
  assign new_n517_ = pv56_2_ & new_n213_;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign new_n519_ = ~new_n194_ & ~new_n514_;
  assign new_n520_ = ~new_n515_ & new_n519_;
  assign pv119_16_ = ~new_n518_ | ~new_n520_;
  assign new_n522_ = pv88_21_ & new_n206_;
  assign new_n523_ = pv88_13_ & new_n252_;
  assign new_n524_ = pv88_6_ & new_n213_;
  assign new_n525_ = ~new_n256_ & ~new_n524_;
  assign new_n526_ = new_n260_ & new_n525_;
  assign new_n527_ = ~new_n250_ & ~new_n522_;
  assign new_n528_ = ~new_n354_ & ~new_n523_;
  assign new_n529_ = new_n527_ & new_n528_;
  assign pv151_21_ = ~new_n526_ | ~new_n529_;
  assign new_n531_ = pv56_18_ & new_n206_;
  assign new_n532_ = pv56_7_ & new_n208_;
  assign new_n533_ = pv56_10_ & new_n211_;
  assign new_n534_ = pv56_3_ & new_n213_;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~new_n194_ & ~new_n531_;
  assign new_n537_ = ~new_n532_ & new_n536_;
  assign pv119_17_ = ~new_n535_ | ~new_n537_;
  assign new_n539_ = pv88_20_ & new_n206_;
  assign new_n540_ = pv88_12_ & new_n252_;
  assign new_n541_ = pv88_5_ & new_n213_;
  assign new_n542_ = ~new_n256_ & ~new_n541_;
  assign new_n543_ = new_n260_ & new_n542_;
  assign new_n544_ = ~new_n250_ & ~new_n539_;
  assign new_n545_ = ~new_n380_ & ~new_n540_;
  assign new_n546_ = new_n544_ & new_n545_;
  assign pv151_20_ = ~new_n543_ | ~new_n546_;
  assign new_n548_ = pv56_15_ & new_n206_;
  assign new_n549_ = pv56_4_ & new_n208_;
  assign new_n550_ = pv56_7_ & new_n211_;
  assign new_n551_ = pv24_14_ & new_n213_;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~new_n194_ & ~new_n548_;
  assign new_n554_ = ~new_n549_ & new_n553_;
  assign pv119_14_ = ~new_n552_ | ~new_n554_;
  assign new_n556_ = pv88_23_ & new_n206_;
  assign new_n557_ = pv88_12_ & new_n208_;
  assign new_n558_ = pv88_15_ & new_n252_;
  assign new_n559_ = pv88_8_ & new_n213_;
  assign new_n560_ = ~new_n256_ & ~new_n559_;
  assign new_n561_ = new_n260_ & new_n560_;
  assign new_n562_ = ~new_n250_ & ~new_n556_;
  assign new_n563_ = ~new_n557_ & ~new_n558_;
  assign new_n564_ = new_n562_ & new_n563_;
  assign pv151_23_ = ~new_n561_ | ~new_n564_;
  assign new_n566_ = pv56_16_ & new_n206_;
  assign new_n567_ = pv56_5_ & new_n208_;
  assign new_n568_ = pv56_8_ & new_n211_;
  assign new_n569_ = pv56_1_ & new_n213_;
  assign new_n570_ = ~new_n568_ & ~new_n569_;
  assign new_n571_ = ~new_n194_ & ~new_n566_;
  assign new_n572_ = ~new_n567_ & new_n571_;
  assign pv119_15_ = ~new_n570_ | ~new_n572_;
  assign new_n574_ = pv88_22_ & new_n206_;
  assign new_n575_ = pv88_11_ & new_n208_;
  assign new_n576_ = pv88_14_ & new_n252_;
  assign new_n577_ = pv88_7_ & new_n213_;
  assign new_n578_ = ~new_n256_ & ~new_n577_;
  assign new_n579_ = new_n260_ & new_n578_;
  assign new_n580_ = ~new_n250_ & ~new_n574_;
  assign new_n581_ = ~new_n575_ & ~new_n576_;
  assign new_n582_ = new_n580_ & new_n581_;
  assign pv151_22_ = ~new_n579_ | ~new_n582_;
  assign new_n584_ = pv56_13_ & new_n206_;
  assign new_n585_ = pv56_2_ & new_n208_;
  assign new_n586_ = pv56_5_ & new_n211_;
  assign new_n587_ = pv24_12_ & new_n213_;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = ~new_n194_ & ~new_n584_;
  assign new_n590_ = ~new_n585_ & new_n589_;
  assign pv119_12_ = ~new_n588_ | ~new_n590_;
  assign new_n592_ = pv88_25_ & new_n206_;
  assign new_n593_ = pv88_14_ & new_n208_;
  assign new_n594_ = pv88_17_ & new_n252_;
  assign new_n595_ = pv88_10_ & new_n213_;
  assign new_n596_ = ~new_n256_ & ~new_n595_;
  assign new_n597_ = new_n260_ & new_n596_;
  assign new_n598_ = ~new_n250_ & ~new_n592_;
  assign new_n599_ = ~new_n593_ & ~new_n594_;
  assign new_n600_ = new_n598_ & new_n599_;
  assign pv151_25_ = ~new_n597_ | ~new_n600_;
  assign new_n602_ = pv88_30_ & new_n206_;
  assign new_n603_ = pv88_19_ & new_n208_;
  assign new_n604_ = pv88_22_ & new_n252_;
  assign new_n605_ = pv88_15_ & new_n213_;
  assign new_n606_ = ~new_n256_ & ~new_n605_;
  assign new_n607_ = new_n260_ & new_n606_;
  assign new_n608_ = ~new_n250_ & ~new_n602_;
  assign new_n609_ = ~new_n603_ & ~new_n604_;
  assign new_n610_ = new_n608_ & new_n609_;
  assign pv151_30_ = ~new_n607_ | ~new_n610_;
  assign new_n612_ = pv56_14_ & new_n206_;
  assign new_n613_ = pv56_3_ & new_n208_;
  assign new_n614_ = pv56_6_ & new_n211_;
  assign new_n615_ = pv24_13_ & new_n213_;
  assign new_n616_ = ~new_n614_ & ~new_n615_;
  assign new_n617_ = ~new_n194_ & ~new_n612_;
  assign new_n618_ = ~new_n613_ & new_n617_;
  assign pv119_13_ = ~new_n616_ | ~new_n618_;
  assign new_n620_ = pv88_24_ & new_n206_;
  assign new_n621_ = pv88_13_ & new_n208_;
  assign new_n622_ = pv88_16_ & new_n252_;
  assign new_n623_ = pv88_9_ & new_n213_;
  assign new_n624_ = ~new_n256_ & ~new_n623_;
  assign new_n625_ = new_n260_ & new_n624_;
  assign new_n626_ = ~new_n250_ & ~new_n620_;
  assign new_n627_ = ~new_n621_ & ~new_n622_;
  assign new_n628_ = new_n626_ & new_n627_;
  assign pv151_24_ = ~new_n625_ | ~new_n628_;
  assign new_n630_ = pv88_31_ & new_n206_;
  assign new_n631_ = pv88_20_ & new_n208_;
  assign new_n632_ = pv88_23_ & new_n252_;
  assign new_n633_ = pv88_16_ & new_n213_;
  assign new_n634_ = ~new_n256_ & ~new_n633_;
  assign new_n635_ = new_n260_ & new_n634_;
  assign new_n636_ = ~new_n250_ & ~new_n630_;
  assign new_n637_ = ~new_n631_ & ~new_n632_;
  assign new_n638_ = new_n636_ & new_n637_;
  assign pv151_31_ = ~new_n635_ | ~new_n638_;
  assign new_n640_ = pv56_11_ & new_n206_;
  assign new_n641_ = pv56_3_ & new_n211_;
  assign new_n642_ = pv24_10_ & new_n213_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = ~new_n194_ & ~new_n640_;
  assign new_n645_ = ~new_n575_ & new_n644_;
  assign pv119_10_ = ~new_n643_ | ~new_n645_;
  assign new_n647_ = pv88_5_ & new_n206_;
  assign new_n648_ = pv56_26_ & new_n208_;
  assign new_n649_ = pv56_29_ & new_n252_;
  assign new_n650_ = pv56_22_ & new_n213_;
  assign new_n651_ = ~new_n256_ & ~new_n650_;
  assign new_n652_ = new_n260_ & new_n651_;
  assign new_n653_ = ~new_n250_ & ~new_n647_;
  assign new_n654_ = ~new_n648_ & ~new_n649_;
  assign new_n655_ = new_n653_ & new_n654_;
  assign pv151_5_ = ~new_n652_ | ~new_n655_;
  assign new_n657_ = pv88_14_ & new_n206_;
  assign new_n658_ = pv88_6_ & new_n252_;
  assign new_n659_ = pv56_31_ & new_n213_;
  assign new_n660_ = ~new_n256_ & ~new_n659_;
  assign new_n661_ = new_n260_ & new_n660_;
  assign new_n662_ = ~new_n250_ & ~new_n657_;
  assign new_n663_ = ~new_n242_ & ~new_n658_;
  assign new_n664_ = new_n662_ & new_n663_;
  assign pv151_14_ = ~new_n661_ | ~new_n664_;
  assign new_n666_ = pv56_12_ & new_n206_;
  assign new_n667_ = pv56_1_ & new_n208_;
  assign new_n668_ = pv56_4_ & new_n211_;
  assign new_n669_ = pv24_11_ & new_n213_;
  assign new_n670_ = ~new_n668_ & ~new_n669_;
  assign new_n671_ = ~new_n194_ & ~new_n666_;
  assign new_n672_ = ~new_n667_ & new_n671_;
  assign pv119_11_ = ~new_n670_ | ~new_n672_;
  assign new_n674_ = pv88_4_ & new_n206_;
  assign new_n675_ = pv56_25_ & new_n208_;
  assign new_n676_ = pv56_28_ & new_n252_;
  assign new_n677_ = pv56_21_ & new_n213_;
  assign new_n678_ = ~new_n256_ & ~new_n677_;
  assign new_n679_ = new_n260_ & new_n678_;
  assign new_n680_ = ~new_n250_ & ~new_n674_;
  assign new_n681_ = ~new_n675_ & ~new_n676_;
  assign new_n682_ = new_n680_ & new_n681_;
  assign pv151_4_ = ~new_n679_ | ~new_n682_;
  assign new_n684_ = pv88_15_ & new_n206_;
  assign new_n685_ = pv88_7_ & new_n252_;
  assign new_n686_ = pv88_0_ & new_n213_;
  assign new_n687_ = ~new_n256_ & ~new_n686_;
  assign new_n688_ = new_n260_ & new_n687_;
  assign new_n689_ = ~new_n250_ & ~new_n684_;
  assign new_n690_ = ~new_n227_ & ~new_n685_;
  assign new_n691_ = new_n689_ & new_n690_;
  assign pv151_15_ = ~new_n688_ | ~new_n691_;
  assign new_n693_ = pv88_7_ & new_n206_;
  assign new_n694_ = pv56_28_ & new_n208_;
  assign new_n695_ = pv56_31_ & new_n252_;
  assign new_n696_ = pv56_24_ & new_n213_;
  assign new_n697_ = ~new_n256_ & ~new_n696_;
  assign new_n698_ = new_n260_ & new_n697_;
  assign new_n699_ = ~new_n250_ & ~new_n693_;
  assign new_n700_ = ~new_n694_ & ~new_n695_;
  assign new_n701_ = new_n699_ & new_n700_;
  assign pv151_7_ = ~new_n698_ | ~new_n701_;
  assign new_n703_ = pv88_12_ & new_n206_;
  assign new_n704_ = pv88_4_ & new_n252_;
  assign new_n705_ = pv56_29_ & new_n213_;
  assign new_n706_ = ~new_n256_ & ~new_n705_;
  assign new_n707_ = new_n260_ & new_n706_;
  assign new_n708_ = ~new_n250_ & ~new_n703_;
  assign new_n709_ = ~new_n220_ & ~new_n704_;
  assign new_n710_ = new_n708_ & new_n709_;
  assign pv151_12_ = ~new_n707_ | ~new_n710_;
  assign new_n712_ = pv88_6_ & new_n206_;
  assign new_n713_ = pv56_27_ & new_n208_;
  assign new_n714_ = pv56_30_ & new_n252_;
  assign new_n715_ = pv56_23_ & new_n213_;
  assign new_n716_ = ~new_n256_ & ~new_n715_;
  assign new_n717_ = new_n260_ & new_n716_;
  assign new_n718_ = ~new_n250_ & ~new_n712_;
  assign new_n719_ = ~new_n713_ & ~new_n714_;
  assign new_n720_ = new_n718_ & new_n719_;
  assign pv151_6_ = ~new_n717_ | ~new_n720_;
  assign new_n722_ = pv88_13_ & new_n206_;
  assign new_n723_ = pv88_5_ & new_n252_;
  assign new_n724_ = pv56_30_ & new_n213_;
  assign new_n725_ = ~new_n256_ & ~new_n724_;
  assign new_n726_ = new_n260_ & new_n725_;
  assign new_n727_ = ~new_n250_ & ~new_n722_;
  assign new_n728_ = ~new_n209_ & ~new_n723_;
  assign new_n729_ = new_n727_ & new_n728_;
  assign pv151_13_ = ~new_n726_ | ~new_n729_;
  assign new_n731_ = pv88_9_ & new_n206_;
  assign new_n732_ = pv56_30_ & new_n208_;
  assign new_n733_ = pv88_1_ & new_n252_;
  assign new_n734_ = pv56_26_ & new_n213_;
  assign new_n735_ = ~new_n256_ & ~new_n734_;
  assign new_n736_ = new_n260_ & new_n735_;
  assign new_n737_ = ~new_n250_ & ~new_n731_;
  assign new_n738_ = ~new_n732_ & ~new_n733_;
  assign new_n739_ = new_n737_ & new_n738_;
  assign pv151_9_ = ~new_n736_ | ~new_n739_;
  assign new_n741_ = pv88_10_ & new_n206_;
  assign new_n742_ = pv56_31_ & new_n208_;
  assign new_n743_ = pv88_2_ & new_n252_;
  assign new_n744_ = pv56_27_ & new_n213_;
  assign new_n745_ = ~new_n256_ & ~new_n744_;
  assign new_n746_ = new_n260_ & new_n745_;
  assign new_n747_ = ~new_n250_ & ~new_n741_;
  assign new_n748_ = ~new_n742_ & ~new_n743_;
  assign new_n749_ = new_n747_ & new_n748_;
  assign pv151_10_ = ~new_n746_ | ~new_n749_;
  assign new_n751_ = pv88_8_ & new_n206_;
  assign new_n752_ = pv56_29_ & new_n208_;
  assign new_n753_ = pv88_0_ & new_n252_;
  assign new_n754_ = pv56_25_ & new_n213_;
  assign new_n755_ = ~new_n256_ & ~new_n754_;
  assign new_n756_ = new_n260_ & new_n755_;
  assign new_n757_ = ~new_n250_ & ~new_n751_;
  assign new_n758_ = ~new_n752_ & ~new_n753_;
  assign new_n759_ = new_n757_ & new_n758_;
  assign pv151_8_ = ~new_n756_ | ~new_n759_;
  assign new_n761_ = pv88_11_ & new_n206_;
  assign new_n762_ = pv88_0_ & new_n208_;
  assign new_n763_ = pv88_3_ & new_n252_;
  assign new_n764_ = pv56_28_ & new_n213_;
  assign new_n765_ = ~new_n256_ & ~new_n764_;
  assign new_n766_ = new_n260_ & new_n765_;
  assign new_n767_ = ~new_n250_ & ~new_n761_;
  assign new_n768_ = ~new_n762_ & ~new_n763_;
  assign new_n769_ = new_n767_ & new_n768_;
  assign pv151_11_ = ~new_n766_ | ~new_n769_;
endmodule

