module count ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, u, v, w, x, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0,
    k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, u, v,
    w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0;
  output k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0;
  wire new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n59_,
    new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n83_,
    new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_;
  assign new_n52_ = ~r & u;
  assign new_n53_ = r & ~u;
  assign new_n54_ = ~new_n52_ & ~new_n53_;
  assign new_n55_ = q & new_n54_;
  assign new_n56_ = ~p & ~q;
  assign new_n57_ = ~new_n55_ & ~new_n56_;
  assign k0 = s | ~new_n57_;
  assign new_n59_ = ~r & ~u;
  assign new_n60_ = ~v & ~new_n59_;
  assign new_n61_ = v & new_n59_;
  assign new_n62_ = ~new_n60_ & ~new_n61_;
  assign new_n63_ = q & new_n62_;
  assign new_n64_ = ~o & ~q;
  assign new_n65_ = ~new_n63_ & ~new_n64_;
  assign l0 = s | ~new_n65_;
  assign new_n67_ = ~v & new_n59_;
  assign new_n68_ = w & new_n67_;
  assign new_n69_ = ~w & ~new_n67_;
  assign new_n70_ = ~new_n68_ & ~new_n69_;
  assign new_n71_ = q & new_n70_;
  assign new_n72_ = ~n & ~q;
  assign new_n73_ = ~new_n71_ & ~new_n72_;
  assign m0 = s | ~new_n73_;
  assign new_n75_ = ~w & new_n67_;
  assign new_n76_ = ~x & ~new_n75_;
  assign new_n77_ = x & new_n75_;
  assign new_n78_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = q & new_n78_;
  assign new_n80_ = ~m & ~q;
  assign new_n81_ = ~new_n79_ & ~new_n80_;
  assign n0 = s | ~new_n81_;
  assign new_n83_ = ~x & new_n75_;
  assign new_n84_ = y & new_n83_;
  assign new_n85_ = ~y & ~new_n83_;
  assign new_n86_ = ~new_n84_ & ~new_n85_;
  assign new_n87_ = q & new_n86_;
  assign new_n88_ = ~l & ~q;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign o0 = s | ~new_n89_;
  assign new_n91_ = ~y & new_n83_;
  assign new_n92_ = ~z & ~new_n91_;
  assign new_n93_ = z & new_n91_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = q & new_n94_;
  assign new_n96_ = ~k & ~q;
  assign new_n97_ = ~new_n95_ & ~new_n96_;
  assign p0 = s | ~new_n97_;
  assign new_n99_ = ~z & new_n91_;
  assign new_n100_ = a0 & new_n99_;
  assign new_n101_ = ~a0 & ~new_n99_;
  assign new_n102_ = ~new_n100_ & ~new_n101_;
  assign new_n103_ = q & new_n102_;
  assign new_n104_ = ~j & ~q;
  assign new_n105_ = ~new_n103_ & ~new_n104_;
  assign q0 = s | ~new_n105_;
  assign new_n107_ = ~a0 & new_n99_;
  assign new_n108_ = ~b0 & ~new_n107_;
  assign new_n109_ = b0 & new_n107_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = q & new_n110_;
  assign new_n112_ = ~i & ~q;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign r0 = s | ~new_n113_;
  assign new_n115_ = ~b0 & new_n107_;
  assign new_n116_ = c0 & new_n115_;
  assign new_n117_ = ~c0 & ~new_n115_;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = q & new_n118_;
  assign new_n120_ = ~h & ~q;
  assign new_n121_ = ~new_n119_ & ~new_n120_;
  assign s0 = s | ~new_n121_;
  assign new_n123_ = ~c0 & new_n115_;
  assign new_n124_ = ~d0 & ~new_n123_;
  assign new_n125_ = d0 & new_n123_;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign new_n127_ = q & new_n126_;
  assign new_n128_ = ~g & ~q;
  assign new_n129_ = ~new_n127_ & ~new_n128_;
  assign t0 = s | ~new_n129_;
  assign new_n131_ = ~d0 & new_n123_;
  assign new_n132_ = e0 & new_n131_;
  assign new_n133_ = ~e0 & ~new_n131_;
  assign new_n134_ = ~new_n132_ & ~new_n133_;
  assign new_n135_ = q & new_n134_;
  assign new_n136_ = ~f & ~q;
  assign new_n137_ = ~new_n135_ & ~new_n136_;
  assign u0 = s | ~new_n137_;
  assign new_n139_ = ~e0 & new_n131_;
  assign new_n140_ = ~f0 & ~new_n139_;
  assign new_n141_ = f0 & new_n139_;
  assign new_n142_ = ~new_n140_ & ~new_n141_;
  assign new_n143_ = q & new_n142_;
  assign new_n144_ = ~e & ~q;
  assign new_n145_ = ~new_n143_ & ~new_n144_;
  assign v0 = s | ~new_n145_;
  assign new_n147_ = ~f0 & new_n139_;
  assign new_n148_ = g0 & new_n147_;
  assign new_n149_ = ~g0 & ~new_n147_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = q & new_n150_;
  assign new_n152_ = ~d & ~q;
  assign new_n153_ = ~new_n151_ & ~new_n152_;
  assign w0 = s | ~new_n153_;
  assign new_n155_ = ~g0 & new_n147_;
  assign new_n156_ = ~h0 & ~new_n155_;
  assign new_n157_ = h0 & new_n155_;
  assign new_n158_ = ~new_n156_ & ~new_n157_;
  assign new_n159_ = q & new_n158_;
  assign new_n160_ = ~c & ~q;
  assign new_n161_ = ~new_n159_ & ~new_n160_;
  assign x0 = s | ~new_n161_;
  assign new_n163_ = ~h0 & new_n155_;
  assign new_n164_ = i0 & new_n163_;
  assign new_n165_ = ~i0 & ~new_n163_;
  assign new_n166_ = ~new_n164_ & ~new_n165_;
  assign new_n167_ = q & new_n166_;
  assign new_n168_ = ~b & ~q;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign y0 = s | ~new_n169_;
  assign new_n171_ = ~i0 & new_n163_;
  assign new_n172_ = ~j0 & ~new_n171_;
  assign new_n173_ = j0 & new_n171_;
  assign new_n174_ = ~new_n172_ & ~new_n173_;
  assign new_n175_ = q & new_n174_;
  assign new_n176_ = ~a & ~q;
  assign new_n177_ = ~new_n175_ & ~new_n176_;
  assign z0 = s | ~new_n177_;
endmodule

