module top ( 
    pv144_18_, pv126_20_, pv126_31_, pv94_30_, pv126_9_, pv129_0_,
    pv94_31_, pv144_19_, pv94_10_, pv94_21_, pv126_7_, pv126_10_,
    pv144_27_, pv176_31_, pv190_0_, pv94_11_, pv94_20_, pv126_8_,
    pv144_28_, pv176_30_, pv30_18_, pv30_29_, pv126_5_, pv144_29_,
    pv30_19_, pv30_28_, pv126_6_, pv128_0_, pv190_1_, pv30_9_, pv62_2_,
    pv64_0_, pv126_14_, pv126_27_, pv176_8_, pv176_22_, pv188_23_, pv30_8_,
    pv62_3_, pv126_13_, pv126_28_, pv176_7_, pv176_23_, pv178_1_,
    pv188_24_, pv30_7_, pv62_0_, pv126_12_, pv126_25_, pv176_6_, pv176_20_,
    pv178_0_, pv188_25_, pv30_6_, pv62_1_, pv63_0_, pv126_11_, pv126_26_,
    pv176_5_, pv176_21_, pv188_26_, pv30_5_, pv62_6_, pv94_7_, pv126_18_,
    pv126_23_, pv176_13_, pv188_27_, pv30_4_, pv62_7_, pv94_6_, pv126_17_,
    pv126_24_, pv176_12_, pv188_28_, pv30_3_, pv62_4_, pv94_9_, pv126_16_,
    pv126_21_, pv126_30_, pv130_0_, pv176_11_, pv188_29_, pv30_2_, pv62_5_,
    pv94_8_, pv126_15_, pv126_22_, pv176_9_, pv176_10_, pv30_30_, pv62_15_,
    pv62_26_, pv94_3_, pv176_0_, pv176_17_, pv30_31_, pv62_16_, pv62_25_,
    pv94_2_, pv176_16_, pv201_0_, pv62_8_, pv62_17_, pv62_28_, pv94_5_,
    pv176_15_, pv176_28_, pv201_1_, pv62_9_, pv62_18_, pv62_27_, pv94_4_,
    pv126_19_, pv176_14_, pv176_29_, pv191_31_, pv201_2_, pv62_19_,
    pv176_4_, pv176_26_, pv62_29_, pv176_3_, pv176_27_, pv188_31_,
    pv126_29_, pv176_2_, pv176_19_, pv176_24_, pv188_30_, pv176_1_,
    pv176_18_, pv176_25_, pv188_22_, pv30_16_, pv30_27_, pv94_14_,
    pv94_25_, pv126_3_, pv127_0_, pv144_23_, pv201_7_, pv30_17_, pv30_26_,
    pv62_30_, pv94_15_, pv94_24_, pv126_4_, pv144_24_, pv30_14_, pv30_25_,
    pv62_20_, pv94_12_, pv94_23_, pv126_1_, pv144_25_, pv30_15_, pv30_24_,
    pv62_10_, pv94_13_, pv94_22_, pv126_2_, pv144_26_, pv30_12_, pv30_23_,
    pv62_11_, pv62_22_, pv94_18_, pv94_29_, pv201_3_, pv30_13_, pv30_22_,
    pv62_12_, pv62_21_, pv94_19_, pv94_28_, pv126_0_, pv144_20_, pv144_31_,
    pv201_4_, pv30_10_, pv30_21_, pv62_13_, pv62_24_, pv62_31_, pv94_16_,
    pv94_27_, pv144_21_, pv144_30_, pv193_1_, pv201_5_, pv30_11_, pv30_20_,
    pv62_14_, pv62_23_, pv94_17_, pv94_26_, pv144_22_, pv193_0_, pv201_6_,
    pv202_0_  );
  input  pv144_18_, pv126_20_, pv126_31_, pv94_30_, pv126_9_, pv129_0_,
    pv94_31_, pv144_19_, pv94_10_, pv94_21_, pv126_7_, pv126_10_,
    pv144_27_, pv176_31_, pv190_0_, pv94_11_, pv94_20_, pv126_8_,
    pv144_28_, pv176_30_, pv30_18_, pv30_29_, pv126_5_, pv144_29_,
    pv30_19_, pv30_28_, pv126_6_, pv128_0_, pv190_1_, pv30_9_, pv62_2_,
    pv64_0_, pv126_14_, pv126_27_, pv176_8_, pv176_22_, pv188_23_, pv30_8_,
    pv62_3_, pv126_13_, pv126_28_, pv176_7_, pv176_23_, pv178_1_,
    pv188_24_, pv30_7_, pv62_0_, pv126_12_, pv126_25_, pv176_6_, pv176_20_,
    pv178_0_, pv188_25_, pv30_6_, pv62_1_, pv63_0_, pv126_11_, pv126_26_,
    pv176_5_, pv176_21_, pv188_26_, pv30_5_, pv62_6_, pv94_7_, pv126_18_,
    pv126_23_, pv176_13_, pv188_27_, pv30_4_, pv62_7_, pv94_6_, pv126_17_,
    pv126_24_, pv176_12_, pv188_28_, pv30_3_, pv62_4_, pv94_9_, pv126_16_,
    pv126_21_, pv126_30_, pv130_0_, pv176_11_, pv188_29_, pv30_2_, pv62_5_,
    pv94_8_, pv126_15_, pv126_22_, pv176_9_, pv176_10_, pv30_30_, pv62_15_,
    pv62_26_, pv94_3_, pv176_0_, pv176_17_, pv30_31_, pv62_16_, pv62_25_,
    pv94_2_, pv176_16_, pv201_0_, pv62_8_, pv62_17_, pv62_28_, pv94_5_,
    pv176_15_, pv176_28_, pv201_1_, pv62_9_, pv62_18_, pv62_27_, pv94_4_,
    pv126_19_, pv176_14_, pv176_29_, pv191_31_, pv201_2_, pv62_19_,
    pv176_4_, pv176_26_, pv62_29_, pv176_3_, pv176_27_, pv188_31_,
    pv126_29_, pv176_2_, pv176_19_, pv176_24_, pv188_30_, pv176_1_,
    pv176_18_, pv176_25_, pv188_22_, pv30_16_, pv30_27_, pv94_14_,
    pv94_25_, pv126_3_, pv127_0_, pv144_23_, pv201_7_, pv30_17_, pv30_26_,
    pv62_30_, pv94_15_, pv94_24_, pv126_4_, pv144_24_, pv30_14_, pv30_25_,
    pv62_20_, pv94_12_, pv94_23_, pv126_1_, pv144_25_, pv30_15_, pv30_24_,
    pv62_10_, pv94_13_, pv94_22_, pv126_2_, pv144_26_, pv30_12_, pv30_23_,
    pv62_11_, pv62_22_, pv94_18_, pv94_29_, pv201_3_, pv30_13_, pv30_22_,
    pv62_12_, pv62_21_, pv94_19_, pv94_28_, pv126_0_, pv144_20_, pv144_31_,
    pv201_4_, pv30_10_, pv30_21_, pv62_13_, pv62_24_, pv62_31_, pv94_16_,
    pv94_27_, pv144_21_, pv144_30_, pv193_1_, pv201_5_, pv30_11_, pv30_20_,
    pv62_14_, pv62_23_, pv94_17_, pv94_26_, pv144_22_, pv193_0_, pv201_6_;
  output pv202_0_;
  wire new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_;
  assign new_n203_ = ~pv190_1_ & ~pv188_30_;
  assign new_n204_ = ~pv190_0_ & ~pv188_31_;
  assign new_n205_ = new_n203_ & new_n204_;
  assign new_n206_ = pv201_4_ & ~new_n205_;
  assign new_n207_ = pv201_5_ & new_n206_;
  assign new_n208_ = pv193_1_ & pv201_6_;
  assign new_n209_ = pv201_7_ & new_n208_;
  assign new_n210_ = pv191_31_ & pv201_6_;
  assign new_n211_ = pv201_7_ & new_n210_;
  assign new_n212_ = ~pv176_3_ & ~pv176_2_;
  assign new_n213_ = ~pv176_6_ & ~pv176_4_;
  assign new_n214_ = new_n212_ & new_n213_;
  assign new_n215_ = ~pv176_5_ & ~pv176_9_;
  assign new_n216_ = ~pv176_7_ & ~pv176_17_;
  assign new_n217_ = new_n215_ & new_n216_;
  assign new_n218_ = new_n214_ & new_n217_;
  assign new_n219_ = ~pv176_13_ & ~pv176_15_;
  assign new_n220_ = ~pv176_11_ & ~pv176_16_;
  assign new_n221_ = new_n219_ & new_n220_;
  assign new_n222_ = ~pv176_8_ & ~pv176_10_;
  assign new_n223_ = ~pv176_12_ & ~pv176_14_;
  assign new_n224_ = new_n222_ & new_n223_;
  assign new_n225_ = new_n221_ & new_n224_;
  assign new_n226_ = new_n218_ & new_n225_;
  assign new_n227_ = pv201_2_ & ~new_n226_;
  assign new_n228_ = ~pv176_19_ & ~pv176_18_;
  assign new_n229_ = ~pv176_22_ & ~pv176_20_;
  assign new_n230_ = new_n228_ & new_n229_;
  assign new_n231_ = ~pv176_21_ & ~pv176_25_;
  assign new_n232_ = ~pv176_23_ & ~pv178_1_;
  assign new_n233_ = new_n231_ & new_n232_;
  assign new_n234_ = new_n230_ & new_n233_;
  assign new_n235_ = ~pv176_31_ & ~pv176_29_;
  assign new_n236_ = ~pv178_0_ & ~pv176_27_;
  assign new_n237_ = new_n235_ & new_n236_;
  assign new_n238_ = ~pv176_26_ & ~pv176_24_;
  assign new_n239_ = ~pv176_30_ & ~pv176_28_;
  assign new_n240_ = new_n238_ & new_n239_;
  assign new_n241_ = new_n237_ & new_n240_;
  assign new_n242_ = new_n234_ & new_n241_;
  assign new_n243_ = pv201_3_ & ~new_n242_;
  assign new_n244_ = ~pv188_26_ & ~pv188_29_;
  assign new_n245_ = ~pv188_27_ & ~pv188_28_;
  assign new_n246_ = new_n244_ & new_n245_;
  assign new_n247_ = pv201_4_ & ~new_n246_;
  assign new_n248_ = pv201_5_ & new_n247_;
  assign new_n249_ = pv201_7_ & pv193_1_;
  assign new_n250_ = ~pv30_22_ & ~pv30_20_;
  assign new_n251_ = ~pv30_18_ & ~pv30_16_;
  assign new_n252_ = new_n250_ & new_n251_;
  assign new_n253_ = ~pv30_14_ & ~pv30_10_;
  assign new_n254_ = ~pv30_12_ & ~pv30_11_;
  assign new_n255_ = new_n253_ & new_n254_;
  assign new_n256_ = new_n252_ & new_n255_;
  assign new_n257_ = ~pv62_1_ & ~pv30_13_;
  assign new_n258_ = ~pv30_2_ & ~pv30_31_;
  assign new_n259_ = new_n257_ & new_n258_;
  assign new_n260_ = ~pv30_19_ & ~pv30_4_;
  assign new_n261_ = ~pv30_6_ & ~pv30_21_;
  assign new_n262_ = new_n260_ & new_n261_;
  assign new_n263_ = new_n259_ & new_n262_;
  assign new_n264_ = new_n256_ & new_n263_;
  assign new_n265_ = ~pv30_9_ & ~pv30_17_;
  assign new_n266_ = ~pv30_8_ & ~pv30_15_;
  assign new_n267_ = new_n265_ & new_n266_;
  assign new_n268_ = ~pv30_7_ & ~pv30_27_;
  assign new_n269_ = ~pv30_29_ & ~pv30_5_;
  assign new_n270_ = new_n268_ & new_n269_;
  assign new_n271_ = new_n267_ & new_n270_;
  assign new_n272_ = ~pv30_3_ & ~pv30_23_;
  assign new_n273_ = ~pv62_0_ & ~pv30_25_;
  assign new_n274_ = new_n272_ & new_n273_;
  assign new_n275_ = ~pv30_26_ & ~pv30_24_;
  assign new_n276_ = ~pv30_28_ & ~pv30_30_;
  assign new_n277_ = new_n275_ & new_n276_;
  assign new_n278_ = new_n274_ & new_n277_;
  assign new_n279_ = new_n271_ & new_n278_;
  assign new_n280_ = new_n264_ & new_n279_;
  assign new_n281_ = ~pv201_0_ & ~new_n280_;
  assign new_n282_ = pv201_1_ & new_n281_;
  assign new_n283_ = pv193_0_ & pv201_6_;
  assign new_n284_ = pv130_0_ & pv201_0_;
  assign new_n285_ = ~pv126_20_ & ~pv126_22_;
  assign new_n286_ = ~pv126_18_ & ~pv126_16_;
  assign new_n287_ = new_n285_ & new_n286_;
  assign new_n288_ = ~pv126_10_ & ~pv126_14_;
  assign new_n289_ = ~pv126_12_ & ~pv126_11_;
  assign new_n290_ = new_n288_ & new_n289_;
  assign new_n291_ = new_n287_ & new_n290_;
  assign new_n292_ = ~pv128_0_ & ~pv126_13_;
  assign new_n293_ = ~pv126_31_ & ~pv126_2_;
  assign new_n294_ = new_n292_ & new_n293_;
  assign new_n295_ = ~pv126_19_ & ~pv126_4_;
  assign new_n296_ = ~pv126_6_ & ~pv126_21_;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = new_n294_ & new_n297_;
  assign new_n299_ = new_n291_ & new_n298_;
  assign new_n300_ = ~pv126_9_ & ~pv126_17_;
  assign new_n301_ = ~pv126_8_ & ~pv126_15_;
  assign new_n302_ = new_n300_ & new_n301_;
  assign new_n303_ = ~pv126_7_ & ~pv126_27_;
  assign new_n304_ = ~pv126_5_ & ~pv126_29_;
  assign new_n305_ = new_n303_ & new_n304_;
  assign new_n306_ = new_n302_ & new_n305_;
  assign new_n307_ = ~pv126_23_ & ~pv126_3_;
  assign new_n308_ = ~pv126_25_ & ~pv127_0_;
  assign new_n309_ = new_n307_ & new_n308_;
  assign new_n310_ = ~pv126_26_ & ~pv126_24_;
  assign new_n311_ = ~pv126_28_ & ~pv126_30_;
  assign new_n312_ = new_n310_ & new_n311_;
  assign new_n313_ = new_n309_ & new_n312_;
  assign new_n314_ = new_n306_ & new_n313_;
  assign new_n315_ = new_n299_ & new_n314_;
  assign new_n316_ = pv201_0_ & ~new_n315_;
  assign new_n317_ = pv201_1_ & new_n316_;
  assign new_n318_ = pv201_3_ & new_n227_;
  assign new_n319_ = pv201_7_ & new_n283_;
  assign new_n320_ = ~pv62_20_ & ~pv62_22_;
  assign new_n321_ = ~pv62_16_ & ~pv62_18_;
  assign new_n322_ = new_n320_ & new_n321_;
  assign new_n323_ = ~pv62_10_ & ~pv62_14_;
  assign new_n324_ = ~pv62_11_ & ~pv62_12_;
  assign new_n325_ = new_n323_ & new_n324_;
  assign new_n326_ = new_n322_ & new_n325_;
  assign new_n327_ = ~pv64_0_ & ~pv62_13_;
  assign new_n328_ = ~pv62_2_ & ~pv62_31_;
  assign new_n329_ = new_n327_ & new_n328_;
  assign new_n330_ = ~pv62_4_ & ~pv62_19_;
  assign new_n331_ = ~pv62_6_ & ~pv62_21_;
  assign new_n332_ = new_n330_ & new_n331_;
  assign new_n333_ = new_n329_ & new_n332_;
  assign new_n334_ = new_n326_ & new_n333_;
  assign new_n335_ = ~pv62_17_ & ~pv62_9_;
  assign new_n336_ = ~pv62_15_ & ~pv62_8_;
  assign new_n337_ = new_n335_ & new_n336_;
  assign new_n338_ = ~pv62_7_ & ~pv62_27_;
  assign new_n339_ = ~pv62_5_ & ~pv62_29_;
  assign new_n340_ = new_n338_ & new_n339_;
  assign new_n341_ = new_n337_ & new_n340_;
  assign new_n342_ = ~pv62_3_ & ~pv62_23_;
  assign new_n343_ = ~pv63_0_ & ~pv62_25_;
  assign new_n344_ = new_n342_ & new_n343_;
  assign new_n345_ = ~pv62_26_ & ~pv62_24_;
  assign new_n346_ = ~pv62_28_ & ~pv62_30_;
  assign new_n347_ = new_n345_ & new_n346_;
  assign new_n348_ = new_n344_ & new_n347_;
  assign new_n349_ = new_n341_ & new_n348_;
  assign new_n350_ = new_n334_ & new_n349_;
  assign new_n351_ = ~pv201_0_ & ~new_n350_;
  assign new_n352_ = pv201_1_ & new_n351_;
  assign new_n353_ = pv201_5_ & ~new_n205_;
  assign new_n354_ = pv129_0_ & ~pv201_0_;
  assign new_n355_ = ~pv94_20_ & ~pv94_22_;
  assign new_n356_ = ~pv94_18_ & ~pv94_16_;
  assign new_n357_ = new_n355_ & new_n356_;
  assign new_n358_ = ~pv94_10_ & ~pv94_14_;
  assign new_n359_ = ~pv94_11_ & ~pv94_12_;
  assign new_n360_ = new_n358_ & new_n359_;
  assign new_n361_ = new_n357_ & new_n360_;
  assign new_n362_ = ~pv126_1_ & ~pv94_13_;
  assign new_n363_ = ~pv94_31_ & ~pv94_2_;
  assign new_n364_ = new_n362_ & new_n363_;
  assign new_n365_ = ~pv94_4_ & ~pv94_19_;
  assign new_n366_ = ~pv94_21_ & ~pv94_6_;
  assign new_n367_ = new_n365_ & new_n366_;
  assign new_n368_ = new_n364_ & new_n367_;
  assign new_n369_ = new_n361_ & new_n368_;
  assign new_n370_ = ~pv94_9_ & ~pv94_17_;
  assign new_n371_ = ~pv94_8_ & ~pv94_15_;
  assign new_n372_ = new_n370_ & new_n371_;
  assign new_n373_ = ~pv94_7_ & ~pv94_27_;
  assign new_n374_ = ~pv94_5_ & ~pv94_29_;
  assign new_n375_ = new_n373_ & new_n374_;
  assign new_n376_ = new_n372_ & new_n375_;
  assign new_n377_ = ~pv94_3_ & ~pv94_23_;
  assign new_n378_ = ~pv94_25_ & ~pv126_0_;
  assign new_n379_ = new_n377_ & new_n378_;
  assign new_n380_ = ~pv94_24_ & ~pv94_26_;
  assign new_n381_ = ~pv94_30_ & ~pv94_28_;
  assign new_n382_ = new_n380_ & new_n381_;
  assign new_n383_ = new_n379_ & new_n382_;
  assign new_n384_ = new_n376_ & new_n383_;
  assign new_n385_ = new_n369_ & new_n384_;
  assign new_n386_ = pv201_0_ & ~new_n385_;
  assign new_n387_ = pv201_1_ & new_n386_;
  assign new_n388_ = pv201_2_ & ~new_n242_;
  assign new_n389_ = pv201_3_ & new_n388_;
  assign new_n390_ = ~pv144_18_ & ~pv144_19_;
  assign new_n391_ = ~pv144_20_ & ~pv144_22_;
  assign new_n392_ = new_n390_ & new_n391_;
  assign new_n393_ = ~pv144_25_ & ~pv144_21_;
  assign new_n394_ = ~pv176_1_ & ~pv144_23_;
  assign new_n395_ = new_n393_ & new_n394_;
  assign new_n396_ = new_n392_ & new_n395_;
  assign new_n397_ = ~pv144_29_ & ~pv144_31_;
  assign new_n398_ = ~pv144_27_ & ~pv176_0_;
  assign new_n399_ = new_n397_ & new_n398_;
  assign new_n400_ = ~pv144_24_ & ~pv144_26_;
  assign new_n401_ = ~pv144_28_ & ~pv144_30_;
  assign new_n402_ = new_n400_ & new_n401_;
  assign new_n403_ = new_n399_ & new_n402_;
  assign new_n404_ = new_n396_ & new_n403_;
  assign new_n405_ = pv201_2_ & ~new_n404_;
  assign new_n406_ = pv201_3_ & new_n405_;
  assign new_n407_ = ~pv188_25_ & ~pv188_22_;
  assign new_n408_ = ~pv188_23_ & ~pv188_24_;
  assign new_n409_ = new_n407_ & new_n408_;
  assign new_n410_ = pv201_4_ & ~new_n409_;
  assign new_n411_ = pv201_5_ & new_n410_;
  assign new_n412_ = ~new_n406_ & ~new_n411_;
  assign new_n413_ = ~new_n388_ & new_n412_;
  assign new_n414_ = ~new_n354_ & ~new_n387_;
  assign new_n415_ = ~new_n389_ & new_n414_;
  assign new_n416_ = new_n413_ & new_n415_;
  assign new_n417_ = ~new_n319_ & ~new_n352_;
  assign new_n418_ = ~new_n353_ & new_n417_;
  assign new_n419_ = ~new_n284_ & ~new_n317_;
  assign new_n420_ = ~new_n318_ & new_n419_;
  assign new_n421_ = new_n418_ & new_n420_;
  assign new_n422_ = new_n416_ & new_n421_;
  assign new_n423_ = ~new_n249_ & ~new_n282_;
  assign new_n424_ = ~new_n283_ & new_n423_;
  assign new_n425_ = ~new_n243_ & ~new_n248_;
  assign new_n426_ = ~new_n247_ & new_n425_;
  assign new_n427_ = new_n424_ & new_n426_;
  assign new_n428_ = ~new_n208_ & ~new_n211_;
  assign new_n429_ = ~new_n227_ & new_n428_;
  assign new_n430_ = ~new_n206_ & ~new_n207_;
  assign new_n431_ = ~new_n209_ & new_n430_;
  assign new_n432_ = new_n429_ & new_n431_;
  assign new_n433_ = new_n427_ & new_n432_;
  assign pv202_0_ = ~new_n422_ | ~new_n433_;
endmodule

