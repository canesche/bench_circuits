module top ( 
    pv96_30_, pv128_5_, pv160_1_, pv160_12_, pv160_25_, pv96_31_, pv128_6_,
    pv160_2_, pv160_11_, pv160_26_, pv96_10_, pv96_21_, pv128_3_,
    pv160_14_, pv160_27_, pv192_0_, pv96_11_, pv96_20_, pv128_4_, pv160_0_,
    pv160_13_, pv160_28_, pv128_1_, pv160_5_, pv160_29_, pv128_2_,
    pv128_19_, pv160_6_, pv199_4_, pv160_3_, pv160_10_, pv128_0_, pv160_4_,
    pv32_7_, pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv128_29_, pv192_19_,
    pv199_1_, pv32_6_, pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv192_18_,
    pv199_0_, pv32_5_, pv192_17_, pv192_31_, pv199_3_, pv32_4_, pv192_16_,
    pv192_30_, pv32_3_, pv64_4_, pv96_5_, pv128_9_, pv192_15_, pv192_20_,
    pv32_2_, pv64_5_, pv96_4_, pv192_14_, pv192_21_, pv32_1_, pv64_2_,
    pv96_7_, pv128_7_, pv192_13_, pv32_0_, pv64_3_, pv96_6_, pv128_8_,
    pv192_12_, pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_,
    pv128_21_, pv192_11_, pv192_24_, pv32_11_, pv32_20_, pv64_9_, pv64_18_,
    pv64_27_, pv96_0_, pv128_22_, pv192_10_, pv192_25_, pv32_12_, pv32_23_,
    pv32_30_, pv64_6_, pv64_15_, pv64_26_, pv96_3_, pv128_10_, pv128_23_,
    pv192_22_, pv32_13_, pv32_22_, pv32_31_, pv64_7_, pv64_16_, pv64_25_,
    pv96_2_, pv128_24_, pv128_31_, pv192_23_, pv32_14_, pv32_25_,
    pv128_25_, pv192_28_, pv32_15_, pv32_24_, pv128_26_, pv192_9_,
    pv192_29_, pv195_0_, pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv128_27_,
    pv192_26_, pv32_8_, pv32_17_, pv32_26_, pv64_29_, pv128_28_, pv192_27_,
    pv64_20_, pv64_31_, pv96_16_, pv96_27_, pv128_16_, pv160_9_, pv160_30_,
    pv192_6_, pv194_0_, pv64_10_, pv96_17_, pv96_26_, pv128_15_, pv160_19_,
    pv192_5_, pv96_18_, pv96_29_, pv128_18_, pv160_7_, pv192_8_, pv96_19_,
    pv96_28_, pv128_17_, pv160_8_, pv160_20_, pv192_7_, pv194_1_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv128_12_, pv128_30_, pv160_16_,
    pv160_21_, pv192_2_, pv64_14_, pv64_23_, pv96_13_, pv96_22_, pv128_11_,
    pv160_15_, pv160_22_, pv192_1_, pv64_11_, pv64_22_, pv96_14_, pv96_25_,
    pv128_14_, pv160_18_, pv160_23_, pv192_4_, pv64_12_, pv64_21_,
    pv64_30_, pv96_15_, pv96_24_, pv128_13_, pv128_20_, pv160_17_,
    pv160_24_, pv160_31_, pv192_3_,
    pv227_10_, pv227_23_, pv266_6_, pv227_0_, pv227_24_, pv227_21_,
    pv266_4_, pv227_22_, pv266_5_, pv227_27_, pv259_0_, pv227_25_,
    pv259_2_, pv227_26_, pv259_1_, pv227_7_, pv227_18_, pv259_17_,
    pv227_8_, pv227_17_, pv259_16_, pv227_5_, pv227_16_, pv259_19_,
    pv227_6_, pv227_15_, pv259_18_, pv227_3_, pv227_14_, pv259_26_,
    pv266_2_, pv227_4_, pv227_13_, pv227_20_, pv259_27_, pv266_3_,
    pv227_1_, pv227_12_, pv259_28_, pv266_0_, pv227_2_, pv227_11_,
    pv259_29_, pv266_1_, pv259_22_, pv259_23_, pv259_11_, pv259_24_,
    pv259_10_, pv259_25_, pv259_13_, pv259_31_, pv259_12_, pv259_30_,
    pv227_9_, pv259_15_, pv259_20_, pv227_19_, pv259_14_, pv259_21_,
    pv259_4_, pv259_3_, pv259_6_, pv259_5_, pv259_8_, pv259_7_, pv259_9_  );
  input  pv96_30_, pv128_5_, pv160_1_, pv160_12_, pv160_25_, pv96_31_,
    pv128_6_, pv160_2_, pv160_11_, pv160_26_, pv96_10_, pv96_21_, pv128_3_,
    pv160_14_, pv160_27_, pv192_0_, pv96_11_, pv96_20_, pv128_4_, pv160_0_,
    pv160_13_, pv160_28_, pv128_1_, pv160_5_, pv160_29_, pv128_2_,
    pv128_19_, pv160_6_, pv199_4_, pv160_3_, pv160_10_, pv128_0_, pv160_4_,
    pv32_7_, pv32_18_, pv32_29_, pv64_0_, pv96_9_, pv128_29_, pv192_19_,
    pv199_1_, pv32_6_, pv32_19_, pv32_28_, pv64_1_, pv96_8_, pv192_18_,
    pv199_0_, pv32_5_, pv192_17_, pv192_31_, pv199_3_, pv32_4_, pv192_16_,
    pv192_30_, pv32_3_, pv64_4_, pv96_5_, pv128_9_, pv192_15_, pv192_20_,
    pv32_2_, pv64_5_, pv96_4_, pv192_14_, pv192_21_, pv32_1_, pv64_2_,
    pv96_7_, pv128_7_, pv192_13_, pv32_0_, pv64_3_, pv96_6_, pv128_8_,
    pv192_12_, pv32_10_, pv32_21_, pv64_8_, pv64_17_, pv64_28_, pv96_1_,
    pv128_21_, pv192_11_, pv192_24_, pv32_11_, pv32_20_, pv64_9_, pv64_18_,
    pv64_27_, pv96_0_, pv128_22_, pv192_10_, pv192_25_, pv32_12_, pv32_23_,
    pv32_30_, pv64_6_, pv64_15_, pv64_26_, pv96_3_, pv128_10_, pv128_23_,
    pv192_22_, pv32_13_, pv32_22_, pv32_31_, pv64_7_, pv64_16_, pv64_25_,
    pv96_2_, pv128_24_, pv128_31_, pv192_23_, pv32_14_, pv32_25_,
    pv128_25_, pv192_28_, pv32_15_, pv32_24_, pv128_26_, pv192_9_,
    pv192_29_, pv195_0_, pv32_9_, pv32_16_, pv32_27_, pv64_19_, pv128_27_,
    pv192_26_, pv32_8_, pv32_17_, pv32_26_, pv64_29_, pv128_28_, pv192_27_,
    pv64_20_, pv64_31_, pv96_16_, pv96_27_, pv128_16_, pv160_9_, pv160_30_,
    pv192_6_, pv194_0_, pv64_10_, pv96_17_, pv96_26_, pv128_15_, pv160_19_,
    pv192_5_, pv96_18_, pv96_29_, pv128_18_, pv160_7_, pv192_8_, pv96_19_,
    pv96_28_, pv128_17_, pv160_8_, pv160_20_, pv192_7_, pv194_1_, pv64_13_,
    pv64_24_, pv96_12_, pv96_23_, pv128_12_, pv128_30_, pv160_16_,
    pv160_21_, pv192_2_, pv64_14_, pv64_23_, pv96_13_, pv96_22_, pv128_11_,
    pv160_15_, pv160_22_, pv192_1_, pv64_11_, pv64_22_, pv96_14_, pv96_25_,
    pv128_14_, pv160_18_, pv160_23_, pv192_4_, pv64_12_, pv64_21_,
    pv64_30_, pv96_15_, pv96_24_, pv128_13_, pv128_20_, pv160_17_,
    pv160_24_, pv160_31_, pv192_3_;
  output pv227_10_, pv227_23_, pv266_6_, pv227_0_, pv227_24_, pv227_21_,
    pv266_4_, pv227_22_, pv266_5_, pv227_27_, pv259_0_, pv227_25_,
    pv259_2_, pv227_26_, pv259_1_, pv227_7_, pv227_18_, pv259_17_,
    pv227_8_, pv227_17_, pv259_16_, pv227_5_, pv227_16_, pv259_19_,
    pv227_6_, pv227_15_, pv259_18_, pv227_3_, pv227_14_, pv259_26_,
    pv266_2_, pv227_4_, pv227_13_, pv227_20_, pv259_27_, pv266_3_,
    pv227_1_, pv227_12_, pv259_28_, pv266_0_, pv227_2_, pv227_11_,
    pv259_29_, pv266_1_, pv259_22_, pv259_23_, pv259_11_, pv259_24_,
    pv259_10_, pv259_25_, pv259_13_, pv259_31_, pv259_12_, pv259_30_,
    pv227_9_, pv259_15_, pv259_20_, pv227_19_, pv259_14_, pv259_21_,
    pv259_4_, pv259_3_, pv259_6_, pv259_5_, pv259_8_, pv259_7_, pv259_9_;
  wire new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n326_, new_n327_, new_n328_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_;
  assign new_n267_ = ~pv199_1_ & pv199_0_;
  assign new_n268_ = pv32_10_ & new_n267_;
  assign new_n269_ = pv199_1_ & pv199_0_;
  assign new_n270_ = pv64_10_ & new_n269_;
  assign new_n271_ = ~pv199_1_ & ~pv199_0_;
  assign new_n272_ = pv96_10_ & new_n271_;
  assign new_n273_ = pv199_1_ & ~pv199_0_;
  assign new_n274_ = ~pv96_10_ & new_n273_;
  assign new_n275_ = ~new_n272_ & ~new_n274_;
  assign new_n276_ = ~new_n268_ & ~new_n270_;
  assign pv227_10_ = ~new_n275_ | ~new_n276_;
  assign new_n278_ = pv32_23_ & new_n267_;
  assign new_n279_ = pv64_23_ & new_n269_;
  assign new_n280_ = pv96_23_ & new_n271_;
  assign new_n281_ = ~pv96_23_ & new_n273_;
  assign new_n282_ = ~new_n280_ & ~new_n281_;
  assign new_n283_ = ~new_n278_ & ~new_n279_;
  assign pv227_23_ = ~new_n282_ | ~new_n283_;
  assign new_n285_ = ~pv199_0_ & pv199_3_;
  assign new_n286_ = pv199_1_ & new_n285_;
  assign new_n287_ = pv195_0_ & new_n286_;
  assign new_n288_ = ~pv199_1_ & new_n285_;
  assign new_n289_ = pv195_0_ & new_n288_;
  assign pv266_6_ = new_n287_ | new_n289_;
  assign new_n291_ = pv32_0_ & new_n267_;
  assign new_n292_ = pv64_0_ & new_n269_;
  assign new_n293_ = pv96_0_ & new_n271_;
  assign new_n294_ = ~pv96_0_ & new_n273_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = ~new_n291_ & ~new_n292_;
  assign pv227_0_ = ~new_n295_ | ~new_n296_;
  assign new_n298_ = pv32_24_ & new_n267_;
  assign new_n299_ = pv64_24_ & new_n269_;
  assign new_n300_ = pv96_24_ & new_n271_;
  assign new_n301_ = ~pv96_24_ & new_n273_;
  assign new_n302_ = ~new_n300_ & ~new_n301_;
  assign new_n303_ = ~new_n298_ & ~new_n299_;
  assign pv227_24_ = ~new_n302_ | ~new_n303_;
  assign new_n305_ = pv32_21_ & new_n267_;
  assign new_n306_ = pv64_21_ & new_n269_;
  assign new_n307_ = pv96_21_ & new_n271_;
  assign new_n308_ = ~pv96_21_ & new_n273_;
  assign new_n309_ = ~new_n307_ & ~new_n308_;
  assign new_n310_ = ~new_n305_ & ~new_n306_;
  assign pv227_21_ = ~new_n309_ | ~new_n310_;
  assign new_n312_ = pv199_1_ & ~pv199_3_;
  assign new_n313_ = pv199_3_ & new_n269_;
  assign new_n314_ = pv194_0_ & new_n288_;
  assign new_n315_ = ~pv194_0_ & new_n286_;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = ~new_n312_ & ~new_n313_;
  assign pv266_4_ = ~new_n316_ | ~new_n317_;
  assign new_n319_ = pv32_22_ & new_n267_;
  assign new_n320_ = pv64_22_ & new_n269_;
  assign new_n321_ = pv96_22_ & new_n271_;
  assign new_n322_ = ~pv96_22_ & new_n273_;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign new_n324_ = ~new_n319_ & ~new_n320_;
  assign pv227_22_ = ~new_n323_ | ~new_n324_;
  assign new_n326_ = pv194_1_ & new_n288_;
  assign new_n327_ = ~pv194_1_ & new_n286_;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign pv266_5_ = ~new_n317_ | ~new_n328_;
  assign new_n330_ = pv32_27_ & new_n267_;
  assign new_n331_ = pv64_27_ & new_n269_;
  assign new_n332_ = pv96_27_ & new_n271_;
  assign new_n333_ = ~pv96_27_ & new_n273_;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = ~new_n330_ & ~new_n331_;
  assign pv227_27_ = ~new_n334_ | ~new_n335_;
  assign new_n337_ = pv199_4_ & ~pv199_0_;
  assign new_n338_ = ~pv199_1_ & new_n337_;
  assign new_n339_ = pv96_28_ & new_n338_;
  assign new_n340_ = pv199_4_ & pv199_0_;
  assign new_n341_ = ~pv199_1_ & new_n340_;
  assign new_n342_ = pv32_28_ & new_n341_;
  assign new_n343_ = pv199_1_ & new_n337_;
  assign new_n344_ = ~pv96_28_ & new_n343_;
  assign new_n345_ = pv199_1_ & new_n340_;
  assign new_n346_ = pv64_28_ & new_n345_;
  assign new_n347_ = ~pv199_4_ & pv199_1_;
  assign new_n348_ = ~new_n346_ & ~new_n347_;
  assign new_n349_ = ~new_n339_ & ~new_n342_;
  assign new_n350_ = ~new_n344_ & new_n349_;
  assign pv259_0_ = ~new_n348_ | ~new_n350_;
  assign new_n352_ = pv32_25_ & new_n267_;
  assign new_n353_ = pv64_25_ & new_n269_;
  assign new_n354_ = pv96_25_ & new_n271_;
  assign new_n355_ = ~pv96_25_ & new_n273_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = ~new_n352_ & ~new_n353_;
  assign pv227_25_ = ~new_n356_ | ~new_n357_;
  assign new_n359_ = pv96_30_ & new_n338_;
  assign new_n360_ = pv32_30_ & new_n341_;
  assign new_n361_ = ~pv96_30_ & new_n343_;
  assign new_n362_ = pv64_30_ & new_n345_;
  assign new_n363_ = ~new_n347_ & ~new_n362_;
  assign new_n364_ = ~new_n359_ & ~new_n360_;
  assign new_n365_ = ~new_n361_ & new_n364_;
  assign pv259_2_ = ~new_n363_ | ~new_n365_;
  assign new_n367_ = pv32_26_ & new_n267_;
  assign new_n368_ = pv64_26_ & new_n269_;
  assign new_n369_ = pv96_26_ & new_n271_;
  assign new_n370_ = ~pv96_26_ & new_n273_;
  assign new_n371_ = ~new_n369_ & ~new_n370_;
  assign new_n372_ = ~new_n367_ & ~new_n368_;
  assign pv227_26_ = ~new_n371_ | ~new_n372_;
  assign new_n374_ = pv96_29_ & new_n338_;
  assign new_n375_ = pv32_29_ & new_n341_;
  assign new_n376_ = ~pv96_29_ & new_n343_;
  assign new_n377_ = pv64_29_ & new_n345_;
  assign new_n378_ = ~new_n347_ & ~new_n377_;
  assign new_n379_ = ~new_n374_ & ~new_n375_;
  assign new_n380_ = ~new_n376_ & new_n379_;
  assign pv259_1_ = ~new_n378_ | ~new_n380_;
  assign new_n382_ = pv32_7_ & new_n267_;
  assign new_n383_ = pv64_7_ & new_n269_;
  assign new_n384_ = pv96_7_ & new_n271_;
  assign new_n385_ = ~pv96_7_ & new_n273_;
  assign new_n386_ = ~new_n384_ & ~new_n385_;
  assign new_n387_ = ~new_n382_ & ~new_n383_;
  assign pv227_7_ = ~new_n386_ | ~new_n387_;
  assign new_n389_ = pv32_18_ & new_n267_;
  assign new_n390_ = pv64_18_ & new_n269_;
  assign new_n391_ = pv96_18_ & new_n271_;
  assign new_n392_ = ~pv96_18_ & new_n273_;
  assign new_n393_ = ~new_n391_ & ~new_n392_;
  assign new_n394_ = ~new_n389_ & ~new_n390_;
  assign pv227_18_ = ~new_n393_ | ~new_n394_;
  assign new_n396_ = pv192_13_ & new_n338_;
  assign new_n397_ = pv128_13_ & new_n341_;
  assign new_n398_ = ~pv192_13_ & new_n343_;
  assign new_n399_ = pv160_13_ & new_n345_;
  assign new_n400_ = ~new_n347_ & ~new_n399_;
  assign new_n401_ = ~new_n396_ & ~new_n397_;
  assign new_n402_ = ~new_n398_ & new_n401_;
  assign pv259_17_ = ~new_n400_ | ~new_n402_;
  assign new_n404_ = pv32_8_ & new_n267_;
  assign new_n405_ = pv64_8_ & new_n269_;
  assign new_n406_ = pv96_8_ & new_n271_;
  assign new_n407_ = ~pv96_8_ & new_n273_;
  assign new_n408_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = ~new_n404_ & ~new_n405_;
  assign pv227_8_ = ~new_n408_ | ~new_n409_;
  assign new_n411_ = pv32_17_ & new_n267_;
  assign new_n412_ = pv64_17_ & new_n269_;
  assign new_n413_ = pv96_17_ & new_n271_;
  assign new_n414_ = ~pv96_17_ & new_n273_;
  assign new_n415_ = ~new_n413_ & ~new_n414_;
  assign new_n416_ = ~new_n411_ & ~new_n412_;
  assign pv227_17_ = ~new_n415_ | ~new_n416_;
  assign new_n418_ = pv192_12_ & new_n338_;
  assign new_n419_ = pv128_12_ & new_n341_;
  assign new_n420_ = ~pv192_12_ & new_n343_;
  assign new_n421_ = pv160_12_ & new_n345_;
  assign new_n422_ = ~new_n347_ & ~new_n421_;
  assign new_n423_ = ~new_n418_ & ~new_n419_;
  assign new_n424_ = ~new_n420_ & new_n423_;
  assign pv259_16_ = ~new_n422_ | ~new_n424_;
  assign new_n426_ = pv32_5_ & new_n267_;
  assign new_n427_ = pv64_5_ & new_n269_;
  assign new_n428_ = pv96_5_ & new_n271_;
  assign new_n429_ = ~pv96_5_ & new_n273_;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = ~new_n426_ & ~new_n427_;
  assign pv227_5_ = ~new_n430_ | ~new_n431_;
  assign new_n433_ = pv32_16_ & new_n267_;
  assign new_n434_ = pv64_16_ & new_n269_;
  assign new_n435_ = pv96_16_ & new_n271_;
  assign new_n436_ = ~pv96_16_ & new_n273_;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = ~new_n433_ & ~new_n434_;
  assign pv227_16_ = ~new_n437_ | ~new_n438_;
  assign new_n440_ = pv192_15_ & new_n338_;
  assign new_n441_ = pv128_15_ & new_n341_;
  assign new_n442_ = ~pv192_15_ & new_n343_;
  assign new_n443_ = pv160_15_ & new_n345_;
  assign new_n444_ = ~new_n347_ & ~new_n443_;
  assign new_n445_ = ~new_n440_ & ~new_n441_;
  assign new_n446_ = ~new_n442_ & new_n445_;
  assign pv259_19_ = ~new_n444_ | ~new_n446_;
  assign new_n448_ = pv32_6_ & new_n267_;
  assign new_n449_ = pv64_6_ & new_n269_;
  assign new_n450_ = pv96_6_ & new_n271_;
  assign new_n451_ = ~pv96_6_ & new_n273_;
  assign new_n452_ = ~new_n450_ & ~new_n451_;
  assign new_n453_ = ~new_n448_ & ~new_n449_;
  assign pv227_6_ = ~new_n452_ | ~new_n453_;
  assign new_n455_ = pv32_15_ & new_n267_;
  assign new_n456_ = pv64_15_ & new_n269_;
  assign new_n457_ = pv96_15_ & new_n271_;
  assign new_n458_ = ~pv96_15_ & new_n273_;
  assign new_n459_ = ~new_n457_ & ~new_n458_;
  assign new_n460_ = ~new_n455_ & ~new_n456_;
  assign pv227_15_ = ~new_n459_ | ~new_n460_;
  assign new_n462_ = pv192_14_ & new_n338_;
  assign new_n463_ = pv128_14_ & new_n341_;
  assign new_n464_ = ~pv192_14_ & new_n343_;
  assign new_n465_ = pv160_14_ & new_n345_;
  assign new_n466_ = ~new_n347_ & ~new_n465_;
  assign new_n467_ = ~new_n462_ & ~new_n463_;
  assign new_n468_ = ~new_n464_ & new_n467_;
  assign pv259_18_ = ~new_n466_ | ~new_n468_;
  assign new_n470_ = pv32_3_ & new_n267_;
  assign new_n471_ = pv64_3_ & new_n269_;
  assign new_n472_ = pv96_3_ & new_n271_;
  assign new_n473_ = ~pv96_3_ & new_n273_;
  assign new_n474_ = ~new_n472_ & ~new_n473_;
  assign new_n475_ = ~new_n470_ & ~new_n471_;
  assign pv227_3_ = ~new_n474_ | ~new_n475_;
  assign new_n477_ = pv32_14_ & new_n267_;
  assign new_n478_ = pv64_14_ & new_n269_;
  assign new_n479_ = pv96_14_ & new_n271_;
  assign new_n480_ = ~pv96_14_ & new_n273_;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = ~new_n477_ & ~new_n478_;
  assign pv227_14_ = ~new_n481_ | ~new_n482_;
  assign new_n484_ = pv192_22_ & new_n338_;
  assign new_n485_ = pv128_22_ & new_n341_;
  assign new_n486_ = ~pv192_22_ & new_n343_;
  assign new_n487_ = pv160_22_ & new_n345_;
  assign new_n488_ = ~new_n347_ & ~new_n487_;
  assign new_n489_ = ~new_n484_ & ~new_n485_;
  assign new_n490_ = ~new_n486_ & new_n489_;
  assign pv259_26_ = ~new_n488_ | ~new_n490_;
  assign new_n492_ = pv192_30_ & new_n288_;
  assign new_n493_ = pv199_0_ & pv199_3_;
  assign new_n494_ = ~pv199_1_ & new_n493_;
  assign new_n495_ = pv128_30_ & new_n494_;
  assign new_n496_ = ~pv192_30_ & new_n286_;
  assign new_n497_ = pv160_30_ & new_n313_;
  assign new_n498_ = ~new_n312_ & ~new_n497_;
  assign new_n499_ = ~new_n492_ & ~new_n495_;
  assign new_n500_ = ~new_n496_ & new_n499_;
  assign pv266_2_ = ~new_n498_ | ~new_n500_;
  assign new_n502_ = pv32_4_ & new_n267_;
  assign new_n503_ = pv64_4_ & new_n269_;
  assign new_n504_ = pv96_4_ & new_n271_;
  assign new_n505_ = ~pv96_4_ & new_n273_;
  assign new_n506_ = ~new_n504_ & ~new_n505_;
  assign new_n507_ = ~new_n502_ & ~new_n503_;
  assign pv227_4_ = ~new_n506_ | ~new_n507_;
  assign new_n509_ = pv32_13_ & new_n267_;
  assign new_n510_ = pv64_13_ & new_n269_;
  assign new_n511_ = pv96_13_ & new_n271_;
  assign new_n512_ = ~pv96_13_ & new_n273_;
  assign new_n513_ = ~new_n511_ & ~new_n512_;
  assign new_n514_ = ~new_n509_ & ~new_n510_;
  assign pv227_13_ = ~new_n513_ | ~new_n514_;
  assign new_n516_ = pv32_20_ & new_n267_;
  assign new_n517_ = pv64_20_ & new_n269_;
  assign new_n518_ = pv96_20_ & new_n271_;
  assign new_n519_ = ~pv96_20_ & new_n273_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = ~new_n516_ & ~new_n517_;
  assign pv227_20_ = ~new_n520_ | ~new_n521_;
  assign new_n523_ = pv192_23_ & new_n338_;
  assign new_n524_ = pv128_23_ & new_n341_;
  assign new_n525_ = ~pv192_23_ & new_n343_;
  assign new_n526_ = pv160_23_ & new_n345_;
  assign new_n527_ = ~new_n347_ & ~new_n526_;
  assign new_n528_ = ~new_n523_ & ~new_n524_;
  assign new_n529_ = ~new_n525_ & new_n528_;
  assign pv259_27_ = ~new_n527_ | ~new_n529_;
  assign new_n531_ = pv192_31_ & new_n288_;
  assign new_n532_ = pv128_31_ & new_n494_;
  assign new_n533_ = ~pv192_31_ & new_n286_;
  assign new_n534_ = pv160_31_ & new_n313_;
  assign new_n535_ = ~new_n312_ & ~new_n534_;
  assign new_n536_ = ~new_n531_ & ~new_n532_;
  assign new_n537_ = ~new_n533_ & new_n536_;
  assign pv266_3_ = ~new_n535_ | ~new_n537_;
  assign new_n539_ = pv32_1_ & new_n267_;
  assign new_n540_ = pv64_1_ & new_n269_;
  assign new_n541_ = pv96_1_ & new_n271_;
  assign new_n542_ = ~pv96_1_ & new_n273_;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = ~new_n539_ & ~new_n540_;
  assign pv227_1_ = ~new_n543_ | ~new_n544_;
  assign new_n546_ = pv32_12_ & new_n267_;
  assign new_n547_ = pv64_12_ & new_n269_;
  assign new_n548_ = pv96_12_ & new_n271_;
  assign new_n549_ = ~pv96_12_ & new_n273_;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = ~new_n546_ & ~new_n547_;
  assign pv227_12_ = ~new_n550_ | ~new_n551_;
  assign new_n553_ = pv192_24_ & new_n338_;
  assign new_n554_ = pv128_24_ & new_n341_;
  assign new_n555_ = ~pv192_24_ & new_n343_;
  assign new_n556_ = pv160_24_ & new_n345_;
  assign new_n557_ = ~new_n347_ & ~new_n556_;
  assign new_n558_ = ~new_n553_ & ~new_n554_;
  assign new_n559_ = ~new_n555_ & new_n558_;
  assign pv259_28_ = ~new_n557_ | ~new_n559_;
  assign new_n561_ = pv192_28_ & new_n288_;
  assign new_n562_ = pv128_28_ & new_n494_;
  assign new_n563_ = ~pv192_28_ & new_n286_;
  assign new_n564_ = pv160_28_ & new_n313_;
  assign new_n565_ = ~new_n312_ & ~new_n564_;
  assign new_n566_ = ~new_n561_ & ~new_n562_;
  assign new_n567_ = ~new_n563_ & new_n566_;
  assign pv266_0_ = ~new_n565_ | ~new_n567_;
  assign new_n569_ = pv32_2_ & new_n267_;
  assign new_n570_ = pv64_2_ & new_n269_;
  assign new_n571_ = pv96_2_ & new_n271_;
  assign new_n572_ = ~pv96_2_ & new_n273_;
  assign new_n573_ = ~new_n571_ & ~new_n572_;
  assign new_n574_ = ~new_n569_ & ~new_n570_;
  assign pv227_2_ = ~new_n573_ | ~new_n574_;
  assign new_n576_ = pv32_11_ & new_n267_;
  assign new_n577_ = pv64_11_ & new_n269_;
  assign new_n578_ = pv96_11_ & new_n271_;
  assign new_n579_ = ~pv96_11_ & new_n273_;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = ~new_n576_ & ~new_n577_;
  assign pv227_11_ = ~new_n580_ | ~new_n581_;
  assign new_n583_ = pv192_25_ & new_n338_;
  assign new_n584_ = pv128_25_ & new_n341_;
  assign new_n585_ = ~pv192_25_ & new_n343_;
  assign new_n586_ = pv160_25_ & new_n345_;
  assign new_n587_ = ~new_n347_ & ~new_n586_;
  assign new_n588_ = ~new_n583_ & ~new_n584_;
  assign new_n589_ = ~new_n585_ & new_n588_;
  assign pv259_29_ = ~new_n587_ | ~new_n589_;
  assign new_n591_ = pv192_29_ & new_n288_;
  assign new_n592_ = pv128_29_ & new_n494_;
  assign new_n593_ = ~pv192_29_ & new_n286_;
  assign new_n594_ = pv160_29_ & new_n313_;
  assign new_n595_ = ~new_n312_ & ~new_n594_;
  assign new_n596_ = ~new_n591_ & ~new_n592_;
  assign new_n597_ = ~new_n593_ & new_n596_;
  assign pv266_1_ = ~new_n595_ | ~new_n597_;
  assign new_n599_ = pv192_18_ & new_n338_;
  assign new_n600_ = pv128_18_ & new_n341_;
  assign new_n601_ = ~pv192_18_ & new_n343_;
  assign new_n602_ = pv160_18_ & new_n345_;
  assign new_n603_ = ~new_n347_ & ~new_n602_;
  assign new_n604_ = ~new_n599_ & ~new_n600_;
  assign new_n605_ = ~new_n601_ & new_n604_;
  assign pv259_22_ = ~new_n603_ | ~new_n605_;
  assign new_n607_ = pv192_19_ & new_n338_;
  assign new_n608_ = pv128_19_ & new_n341_;
  assign new_n609_ = ~pv192_19_ & new_n343_;
  assign new_n610_ = pv160_19_ & new_n345_;
  assign new_n611_ = ~new_n347_ & ~new_n610_;
  assign new_n612_ = ~new_n607_ & ~new_n608_;
  assign new_n613_ = ~new_n609_ & new_n612_;
  assign pv259_23_ = ~new_n611_ | ~new_n613_;
  assign new_n615_ = pv192_7_ & new_n338_;
  assign new_n616_ = pv128_7_ & new_n341_;
  assign new_n617_ = ~pv192_7_ & new_n343_;
  assign new_n618_ = pv160_7_ & new_n345_;
  assign new_n619_ = ~new_n347_ & ~new_n618_;
  assign new_n620_ = ~new_n615_ & ~new_n616_;
  assign new_n621_ = ~new_n617_ & new_n620_;
  assign pv259_11_ = ~new_n619_ | ~new_n621_;
  assign new_n623_ = pv192_20_ & new_n338_;
  assign new_n624_ = pv128_20_ & new_n341_;
  assign new_n625_ = ~pv192_20_ & new_n343_;
  assign new_n626_ = pv160_20_ & new_n345_;
  assign new_n627_ = ~new_n347_ & ~new_n626_;
  assign new_n628_ = ~new_n623_ & ~new_n624_;
  assign new_n629_ = ~new_n625_ & new_n628_;
  assign pv259_24_ = ~new_n627_ | ~new_n629_;
  assign new_n631_ = pv192_6_ & new_n338_;
  assign new_n632_ = pv128_6_ & new_n341_;
  assign new_n633_ = ~pv192_6_ & new_n343_;
  assign new_n634_ = pv160_6_ & new_n345_;
  assign new_n635_ = ~new_n347_ & ~new_n634_;
  assign new_n636_ = ~new_n631_ & ~new_n632_;
  assign new_n637_ = ~new_n633_ & new_n636_;
  assign pv259_10_ = ~new_n635_ | ~new_n637_;
  assign new_n639_ = pv192_21_ & new_n338_;
  assign new_n640_ = pv128_21_ & new_n341_;
  assign new_n641_ = ~pv192_21_ & new_n343_;
  assign new_n642_ = pv160_21_ & new_n345_;
  assign new_n643_ = ~new_n347_ & ~new_n642_;
  assign new_n644_ = ~new_n639_ & ~new_n640_;
  assign new_n645_ = ~new_n641_ & new_n644_;
  assign pv259_25_ = ~new_n643_ | ~new_n645_;
  assign new_n647_ = pv192_9_ & new_n338_;
  assign new_n648_ = pv128_9_ & new_n341_;
  assign new_n649_ = ~pv192_9_ & new_n343_;
  assign new_n650_ = pv160_9_ & new_n345_;
  assign new_n651_ = ~new_n347_ & ~new_n650_;
  assign new_n652_ = ~new_n647_ & ~new_n648_;
  assign new_n653_ = ~new_n649_ & new_n652_;
  assign pv259_13_ = ~new_n651_ | ~new_n653_;
  assign new_n655_ = pv192_27_ & new_n338_;
  assign new_n656_ = pv128_27_ & new_n341_;
  assign new_n657_ = ~pv192_27_ & new_n343_;
  assign new_n658_ = pv160_27_ & new_n345_;
  assign new_n659_ = ~new_n347_ & ~new_n658_;
  assign new_n660_ = ~new_n655_ & ~new_n656_;
  assign new_n661_ = ~new_n657_ & new_n660_;
  assign pv259_31_ = ~new_n659_ | ~new_n661_;
  assign new_n663_ = pv192_8_ & new_n338_;
  assign new_n664_ = pv128_8_ & new_n341_;
  assign new_n665_ = ~pv192_8_ & new_n343_;
  assign new_n666_ = pv160_8_ & new_n345_;
  assign new_n667_ = ~new_n347_ & ~new_n666_;
  assign new_n668_ = ~new_n663_ & ~new_n664_;
  assign new_n669_ = ~new_n665_ & new_n668_;
  assign pv259_12_ = ~new_n667_ | ~new_n669_;
  assign new_n671_ = pv192_26_ & new_n338_;
  assign new_n672_ = pv128_26_ & new_n341_;
  assign new_n673_ = ~pv192_26_ & new_n343_;
  assign new_n674_ = pv160_26_ & new_n345_;
  assign new_n675_ = ~new_n347_ & ~new_n674_;
  assign new_n676_ = ~new_n671_ & ~new_n672_;
  assign new_n677_ = ~new_n673_ & new_n676_;
  assign pv259_30_ = ~new_n675_ | ~new_n677_;
  assign new_n679_ = pv32_9_ & new_n267_;
  assign new_n680_ = pv64_9_ & new_n269_;
  assign new_n681_ = pv96_9_ & new_n271_;
  assign new_n682_ = ~pv96_9_ & new_n273_;
  assign new_n683_ = ~new_n681_ & ~new_n682_;
  assign new_n684_ = ~new_n679_ & ~new_n680_;
  assign pv227_9_ = ~new_n683_ | ~new_n684_;
  assign new_n686_ = pv192_11_ & new_n338_;
  assign new_n687_ = pv128_11_ & new_n341_;
  assign new_n688_ = ~pv192_11_ & new_n343_;
  assign new_n689_ = pv160_11_ & new_n345_;
  assign new_n690_ = ~new_n347_ & ~new_n689_;
  assign new_n691_ = ~new_n686_ & ~new_n687_;
  assign new_n692_ = ~new_n688_ & new_n691_;
  assign pv259_15_ = ~new_n690_ | ~new_n692_;
  assign new_n694_ = pv192_16_ & new_n338_;
  assign new_n695_ = pv128_16_ & new_n341_;
  assign new_n696_ = ~pv192_16_ & new_n343_;
  assign new_n697_ = pv160_16_ & new_n345_;
  assign new_n698_ = ~new_n347_ & ~new_n697_;
  assign new_n699_ = ~new_n694_ & ~new_n695_;
  assign new_n700_ = ~new_n696_ & new_n699_;
  assign pv259_20_ = ~new_n698_ | ~new_n700_;
  assign new_n702_ = pv32_19_ & new_n267_;
  assign new_n703_ = pv64_19_ & new_n269_;
  assign new_n704_ = pv96_19_ & new_n271_;
  assign new_n705_ = ~pv96_19_ & new_n273_;
  assign new_n706_ = ~new_n704_ & ~new_n705_;
  assign new_n707_ = ~new_n702_ & ~new_n703_;
  assign pv227_19_ = ~new_n706_ | ~new_n707_;
  assign new_n709_ = pv192_10_ & new_n338_;
  assign new_n710_ = pv128_10_ & new_n341_;
  assign new_n711_ = ~pv192_10_ & new_n343_;
  assign new_n712_ = pv160_10_ & new_n345_;
  assign new_n713_ = ~new_n347_ & ~new_n712_;
  assign new_n714_ = ~new_n709_ & ~new_n710_;
  assign new_n715_ = ~new_n711_ & new_n714_;
  assign pv259_14_ = ~new_n713_ | ~new_n715_;
  assign new_n717_ = pv192_17_ & new_n338_;
  assign new_n718_ = pv128_17_ & new_n341_;
  assign new_n719_ = ~pv192_17_ & new_n343_;
  assign new_n720_ = pv160_17_ & new_n345_;
  assign new_n721_ = ~new_n347_ & ~new_n720_;
  assign new_n722_ = ~new_n717_ & ~new_n718_;
  assign new_n723_ = ~new_n719_ & new_n722_;
  assign pv259_21_ = ~new_n721_ | ~new_n723_;
  assign new_n725_ = pv192_0_ & new_n338_;
  assign new_n726_ = pv128_0_ & new_n341_;
  assign new_n727_ = ~pv192_0_ & new_n343_;
  assign new_n728_ = pv160_0_ & new_n345_;
  assign new_n729_ = ~new_n347_ & ~new_n728_;
  assign new_n730_ = ~new_n725_ & ~new_n726_;
  assign new_n731_ = ~new_n727_ & new_n730_;
  assign pv259_4_ = ~new_n729_ | ~new_n731_;
  assign new_n733_ = pv96_31_ & new_n338_;
  assign new_n734_ = pv32_31_ & new_n341_;
  assign new_n735_ = ~pv96_31_ & new_n343_;
  assign new_n736_ = pv64_31_ & new_n345_;
  assign new_n737_ = ~new_n347_ & ~new_n736_;
  assign new_n738_ = ~new_n733_ & ~new_n734_;
  assign new_n739_ = ~new_n735_ & new_n738_;
  assign pv259_3_ = ~new_n737_ | ~new_n739_;
  assign new_n741_ = pv192_2_ & new_n338_;
  assign new_n742_ = pv128_2_ & new_n341_;
  assign new_n743_ = ~pv192_2_ & new_n343_;
  assign new_n744_ = pv160_2_ & new_n345_;
  assign new_n745_ = ~new_n347_ & ~new_n744_;
  assign new_n746_ = ~new_n741_ & ~new_n742_;
  assign new_n747_ = ~new_n743_ & new_n746_;
  assign pv259_6_ = ~new_n745_ | ~new_n747_;
  assign new_n749_ = pv192_1_ & new_n338_;
  assign new_n750_ = pv128_1_ & new_n341_;
  assign new_n751_ = ~pv192_1_ & new_n343_;
  assign new_n752_ = pv160_1_ & new_n345_;
  assign new_n753_ = ~new_n347_ & ~new_n752_;
  assign new_n754_ = ~new_n749_ & ~new_n750_;
  assign new_n755_ = ~new_n751_ & new_n754_;
  assign pv259_5_ = ~new_n753_ | ~new_n755_;
  assign new_n757_ = pv192_4_ & new_n338_;
  assign new_n758_ = pv128_4_ & new_n341_;
  assign new_n759_ = ~pv192_4_ & new_n343_;
  assign new_n760_ = pv160_4_ & new_n345_;
  assign new_n761_ = ~new_n347_ & ~new_n760_;
  assign new_n762_ = ~new_n757_ & ~new_n758_;
  assign new_n763_ = ~new_n759_ & new_n762_;
  assign pv259_8_ = ~new_n761_ | ~new_n763_;
  assign new_n765_ = pv192_3_ & new_n338_;
  assign new_n766_ = pv128_3_ & new_n341_;
  assign new_n767_ = ~pv192_3_ & new_n343_;
  assign new_n768_ = pv160_3_ & new_n345_;
  assign new_n769_ = ~new_n347_ & ~new_n768_;
  assign new_n770_ = ~new_n765_ & ~new_n766_;
  assign new_n771_ = ~new_n767_ & new_n770_;
  assign pv259_7_ = ~new_n769_ | ~new_n771_;
  assign new_n773_ = pv192_5_ & new_n338_;
  assign new_n774_ = pv128_5_ & new_n341_;
  assign new_n775_ = ~pv192_5_ & new_n343_;
  assign new_n776_ = pv160_5_ & new_n345_;
  assign new_n777_ = ~new_n347_ & ~new_n776_;
  assign new_n778_ = ~new_n773_ & ~new_n774_;
  assign new_n779_ = ~new_n775_ & new_n778_;
  assign pv259_9_ = ~new_n777_ | ~new_n779_;
endmodule

