// Benchmark "testing" written by ABC on Thu Oct  8 22:16:41 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A140  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A140;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[442]_ , \new_[443]_ ,
    \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[453]_ , \new_[454]_ ,
    \new_[457]_ , \new_[460]_ , \new_[461]_ , \new_[462]_ , \new_[463]_ ,
    \new_[467]_ , \new_[468]_ , \new_[471]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[480]_ , \new_[481]_ , \new_[484]_ , \new_[487]_ ,
    \new_[488]_ , \new_[489]_ , \new_[490]_ , \new_[491]_ , \new_[495]_ ,
    \new_[496]_ , \new_[500]_ , \new_[501]_ , \new_[502]_ , \new_[506]_ ,
    \new_[507]_ , \new_[510]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[520]_ , \new_[521]_ , \new_[524]_ , \new_[527]_ ,
    \new_[528]_ , \new_[529]_ , \new_[533]_ , \new_[534]_ , \new_[537]_ ,
    \new_[540]_ , \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ ,
    \new_[545]_ , \new_[549]_ , \new_[550]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[560]_ , \new_[561]_ , \new_[564]_ , \new_[567]_ ,
    \new_[568]_ , \new_[569]_ , \new_[570]_ , \new_[574]_ , \new_[575]_ ,
    \new_[578]_ , \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[587]_ ,
    \new_[588]_ , \new_[591]_ , \new_[594]_ , \new_[595]_ , \new_[596]_ ,
    \new_[597]_ , \new_[598]_ , \new_[602]_ , \new_[603]_ , \new_[606]_ ,
    \new_[609]_ , \new_[610]_ , \new_[611]_ , \new_[615]_ , \new_[616]_ ,
    \new_[619]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[629]_ , \new_[630]_ , \new_[633]_ , \new_[636]_ , \new_[637]_ ,
    \new_[638]_ , \new_[642]_ , \new_[643]_ , \new_[646]_ , \new_[649]_ ,
    \new_[650]_ , \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ ,
    \new_[655]_ , \new_[659]_ , \new_[660]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[670]_ , \new_[671]_ , \new_[674]_ , \new_[677]_ ,
    \new_[678]_ , \new_[679]_ , \new_[680]_ , \new_[684]_ , \new_[685]_ ,
    \new_[688]_ , \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[697]_ ,
    \new_[698]_ , \new_[701]_ , \new_[704]_ , \new_[705]_ , \new_[706]_ ,
    \new_[707]_ , \new_[708]_ , \new_[712]_ , \new_[713]_ , \new_[716]_ ,
    \new_[719]_ , \new_[720]_ , \new_[721]_ , \new_[725]_ , \new_[726]_ ,
    \new_[729]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[739]_ , \new_[740]_ , \new_[743]_ , \new_[746]_ , \new_[747]_ ,
    \new_[748]_ , \new_[752]_ , \new_[753]_ , \new_[756]_ , \new_[759]_ ,
    \new_[760]_ , \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ ,
    \new_[768]_ , \new_[769]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[779]_ , \new_[780]_ , \new_[783]_ , \new_[786]_ , \new_[787]_ ,
    \new_[788]_ , \new_[789]_ , \new_[793]_ , \new_[794]_ , \new_[797]_ ,
    \new_[800]_ , \new_[801]_ , \new_[802]_ , \new_[806]_ , \new_[807]_ ,
    \new_[810]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ , \new_[816]_ ,
    \new_[817]_ , \new_[821]_ , \new_[822]_ , \new_[825]_ , \new_[828]_ ,
    \new_[829]_ , \new_[830]_ , \new_[834]_ , \new_[835]_ , \new_[838]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[848]_ ,
    \new_[849]_ , \new_[852]_ , \new_[855]_ , \new_[856]_ , \new_[857]_ ,
    \new_[861]_ , \new_[862]_ , \new_[865]_ , \new_[868]_ , \new_[869]_ ,
    \new_[870]_ , \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ ,
    \new_[875]_ , \new_[879]_ , \new_[880]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[890]_ , \new_[891]_ , \new_[894]_ , \new_[897]_ ,
    \new_[898]_ , \new_[899]_ , \new_[900]_ , \new_[904]_ , \new_[905]_ ,
    \new_[908]_ , \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[917]_ ,
    \new_[918]_ , \new_[921]_ , \new_[924]_ , \new_[925]_ , \new_[926]_ ,
    \new_[927]_ , \new_[928]_ , \new_[932]_ , \new_[933]_ , \new_[937]_ ,
    \new_[938]_ , \new_[939]_ , \new_[943]_ , \new_[944]_ , \new_[947]_ ,
    \new_[950]_ , \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[957]_ ,
    \new_[958]_ , \new_[961]_ , \new_[964]_ , \new_[965]_ , \new_[966]_ ,
    \new_[970]_ , \new_[971]_ , \new_[974]_ , \new_[977]_ , \new_[978]_ ,
    \new_[979]_ , \new_[980]_ , \new_[981]_ , \new_[982]_ , \new_[986]_ ,
    \new_[987]_ , \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[997]_ ,
    \new_[998]_ , \new_[1001]_ , \new_[1004]_ , \new_[1005]_ ,
    \new_[1006]_ , \new_[1007]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1015]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1024]_ , \new_[1025]_ , \new_[1028]_ , \new_[1031]_ ,
    \new_[1032]_ , \new_[1033]_ , \new_[1034]_ , \new_[1035]_ ,
    \new_[1039]_ , \new_[1040]_ , \new_[1043]_ , \new_[1046]_ ,
    \new_[1047]_ , \new_[1048]_ , \new_[1052]_ , \new_[1053]_ ,
    \new_[1056]_ , \new_[1059]_ , \new_[1060]_ , \new_[1061]_ ,
    \new_[1062]_ , \new_[1066]_ , \new_[1067]_ , \new_[1070]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1079]_ ,
    \new_[1080]_ , \new_[1083]_ , \new_[1086]_ , \new_[1087]_ ,
    \new_[1088]_ , \new_[1089]_ , \new_[1090]_ , \new_[1091]_ ,
    \new_[1092]_ , \new_[1096]_ , \new_[1097]_ , \new_[1101]_ ,
    \new_[1102]_ , \new_[1103]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1111]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1121]_ , \new_[1122]_ , \new_[1125]_ ,
    \new_[1128]_ , \new_[1129]_ , \new_[1130]_ , \new_[1134]_ ,
    \new_[1135]_ , \new_[1138]_ , \new_[1141]_ , \new_[1142]_ ,
    \new_[1143]_ , \new_[1144]_ , \new_[1145]_ , \new_[1149]_ ,
    \new_[1150]_ , \new_[1153]_ , \new_[1156]_ , \new_[1157]_ ,
    \new_[1158]_ , \new_[1162]_ , \new_[1163]_ , \new_[1166]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1176]_ , \new_[1177]_ , \new_[1180]_ , \new_[1183]_ ,
    \new_[1184]_ , \new_[1185]_ , \new_[1189]_ , \new_[1190]_ ,
    \new_[1193]_ , \new_[1196]_ , \new_[1197]_ , \new_[1198]_ ,
    \new_[1199]_ , \new_[1200]_ , \new_[1201]_ , \new_[1205]_ ,
    \new_[1206]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1216]_ , \new_[1217]_ , \new_[1220]_ , \new_[1223]_ ,
    \new_[1224]_ , \new_[1225]_ , \new_[1226]_ , \new_[1230]_ ,
    \new_[1231]_ , \new_[1234]_ , \new_[1237]_ , \new_[1238]_ ,
    \new_[1239]_ , \new_[1243]_ , \new_[1244]_ , \new_[1247]_ ,
    \new_[1250]_ , \new_[1251]_ , \new_[1252]_ , \new_[1253]_ ,
    \new_[1254]_ , \new_[1258]_ , \new_[1259]_ , \new_[1262]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1271]_ ,
    \new_[1272]_ , \new_[1275]_ , \new_[1278]_ , \new_[1279]_ ,
    \new_[1280]_ , \new_[1281]_ , \new_[1285]_ , \new_[1286]_ ,
    \new_[1289]_ , \new_[1292]_ , \new_[1293]_ , \new_[1294]_ ,
    \new_[1298]_ , \new_[1299]_ , \new_[1302]_ , \new_[1305]_ ,
    \new_[1306]_ , \new_[1307]_ , \new_[1308]_ , \new_[1309]_ ,
    \new_[1310]_ , \new_[1311]_ , \new_[1312]_ , \new_[1315]_ ,
    \new_[1318]_ , \new_[1321]_ , \new_[1324]_ , \new_[1327]_ ,
    \new_[1330]_ , \new_[1333]_ , \new_[1336]_ , \new_[1339]_ ,
    \new_[1343]_ , \new_[1344]_ , \new_[1347]_ , \new_[1351]_ ,
    \new_[1352]_ , \new_[1355]_ , \new_[1358]_ , \new_[1359]_ ,
    \new_[1362]_ , \new_[1365]_ , \new_[1366]_ , \new_[1369]_ ,
    \new_[1372]_ , \new_[1373]_ , \new_[1376]_ , \new_[1379]_ ,
    \new_[1380]_ , \new_[1383]_ , \new_[1386]_ , \new_[1387]_ ,
    \new_[1390]_ , \new_[1393]_ , \new_[1394]_ , \new_[1397]_ ,
    \new_[1400]_ , \new_[1401]_ , \new_[1404]_ , \new_[1407]_ ,
    \new_[1408]_ , \new_[1411]_ , \new_[1414]_ , \new_[1415]_ ,
    \new_[1418]_ , \new_[1421]_ , \new_[1422]_ , \new_[1425]_ ,
    \new_[1428]_ , \new_[1429]_ , \new_[1432]_ , \new_[1435]_ ,
    \new_[1436]_ , \new_[1439]_ , \new_[1442]_ , \new_[1443]_ ,
    \new_[1446]_ , \new_[1449]_ , \new_[1450]_ , \new_[1453]_ ,
    \new_[1456]_ , \new_[1457]_ , \new_[1460]_ , \new_[1463]_ ,
    \new_[1464]_ , \new_[1467]_ , \new_[1470]_ , \new_[1471]_ ,
    \new_[1474]_ , \new_[1477]_ , \new_[1478]_ , \new_[1481]_ ,
    \new_[1484]_ , \new_[1485]_ , \new_[1488]_ , \new_[1491]_ ,
    \new_[1492]_ , \new_[1495]_ , \new_[1498]_ , \new_[1499]_ ,
    \new_[1502]_ , \new_[1505]_ , \new_[1506]_ , \new_[1509]_ ,
    \new_[1512]_ , \new_[1513]_ , \new_[1516]_ , \new_[1519]_ ,
    \new_[1520]_ , \new_[1523]_ , \new_[1526]_ , \new_[1527]_ ,
    \new_[1530]_ , \new_[1533]_ , \new_[1534]_ , \new_[1537]_ ,
    \new_[1540]_ , \new_[1541]_ , \new_[1544]_ , \new_[1547]_ ,
    \new_[1548]_ , \new_[1551]_ , \new_[1554]_ , \new_[1555]_ ,
    \new_[1558]_ , \new_[1561]_ , \new_[1562]_ , \new_[1565]_ ,
    \new_[1568]_ , \new_[1569]_ , \new_[1572]_ , \new_[1575]_ ,
    \new_[1576]_ , \new_[1579]_ , \new_[1582]_ , \new_[1583]_ ,
    \new_[1586]_ , \new_[1589]_ , \new_[1590]_ , \new_[1593]_ ,
    \new_[1596]_ , \new_[1597]_ , \new_[1600]_ , \new_[1603]_ ,
    \new_[1604]_ , \new_[1607]_ , \new_[1610]_ , \new_[1611]_ ,
    \new_[1614]_ , \new_[1617]_ , \new_[1618]_ , \new_[1621]_ ,
    \new_[1624]_ , \new_[1625]_ , \new_[1628]_ , \new_[1631]_ ,
    \new_[1632]_ , \new_[1635]_ , \new_[1638]_ , \new_[1639]_ ,
    \new_[1642]_ , \new_[1645]_ , \new_[1646]_ , \new_[1649]_ ,
    \new_[1652]_ , \new_[1653]_ , \new_[1656]_ , \new_[1659]_ ,
    \new_[1660]_ , \new_[1663]_ , \new_[1666]_ , \new_[1667]_ ,
    \new_[1670]_ , \new_[1673]_ , \new_[1674]_ , \new_[1677]_ ,
    \new_[1680]_ , \new_[1681]_ , \new_[1684]_ , \new_[1687]_ ,
    \new_[1688]_ , \new_[1691]_ , \new_[1694]_ , \new_[1695]_ ,
    \new_[1698]_ , \new_[1701]_ , \new_[1702]_ , \new_[1705]_ ,
    \new_[1708]_ , \new_[1709]_ , \new_[1712]_ , \new_[1715]_ ,
    \new_[1716]_ , \new_[1719]_ , \new_[1722]_ , \new_[1723]_ ,
    \new_[1726]_ , \new_[1729]_ , \new_[1730]_ , \new_[1733]_ ,
    \new_[1736]_ , \new_[1737]_ , \new_[1740]_ , \new_[1743]_ ,
    \new_[1744]_ , \new_[1747]_ , \new_[1750]_ , \new_[1751]_ ,
    \new_[1754]_ , \new_[1757]_ , \new_[1758]_ , \new_[1761]_ ,
    \new_[1764]_ , \new_[1765]_ , \new_[1768]_ , \new_[1771]_ ,
    \new_[1772]_ , \new_[1775]_ , \new_[1778]_ , \new_[1779]_ ,
    \new_[1782]_ , \new_[1785]_ , \new_[1786]_ , \new_[1789]_ ,
    \new_[1792]_ , \new_[1793]_ , \new_[1796]_ , \new_[1799]_ ,
    \new_[1800]_ , \new_[1803]_ , \new_[1806]_ , \new_[1807]_ ,
    \new_[1810]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1819]_ , \new_[1822]_ , \new_[1823]_ , \new_[1826]_ ,
    \new_[1830]_ , \new_[1831]_ , \new_[1832]_ , \new_[1835]_ ,
    \new_[1838]_ , \new_[1839]_ , \new_[1842]_ , \new_[1846]_ ,
    \new_[1847]_ , \new_[1848]_ , \new_[1851]_ , \new_[1854]_ ,
    \new_[1855]_ , \new_[1858]_ , \new_[1862]_ , \new_[1863]_ ,
    \new_[1864]_ , \new_[1867]_ , \new_[1870]_ , \new_[1871]_ ,
    \new_[1874]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1883]_ , \new_[1886]_ , \new_[1887]_ , \new_[1890]_ ,
    \new_[1894]_ , \new_[1895]_ , \new_[1896]_ , \new_[1899]_ ,
    \new_[1902]_ , \new_[1903]_ , \new_[1906]_ , \new_[1910]_ ,
    \new_[1911]_ , \new_[1912]_ , \new_[1915]_ , \new_[1918]_ ,
    \new_[1919]_ , \new_[1922]_ , \new_[1926]_ , \new_[1927]_ ,
    \new_[1928]_ , \new_[1931]_ , \new_[1934]_ , \new_[1935]_ ,
    \new_[1938]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1947]_ , \new_[1950]_ , \new_[1951]_ , \new_[1954]_ ,
    \new_[1958]_ , \new_[1959]_ , \new_[1960]_ , \new_[1963]_ ,
    \new_[1966]_ , \new_[1967]_ , \new_[1970]_ , \new_[1974]_ ,
    \new_[1975]_ , \new_[1976]_ , \new_[1979]_ , \new_[1982]_ ,
    \new_[1983]_ , \new_[1986]_ , \new_[1990]_ , \new_[1991]_ ,
    \new_[1992]_ , \new_[1995]_ , \new_[1998]_ , \new_[1999]_ ,
    \new_[2002]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2011]_ , \new_[2014]_ , \new_[2015]_ , \new_[2018]_ ,
    \new_[2022]_ , \new_[2023]_ , \new_[2024]_ , \new_[2027]_ ,
    \new_[2030]_ , \new_[2031]_ , \new_[2034]_ , \new_[2038]_ ,
    \new_[2039]_ , \new_[2040]_ , \new_[2043]_ , \new_[2046]_ ,
    \new_[2047]_ , \new_[2050]_ , \new_[2054]_ , \new_[2055]_ ,
    \new_[2056]_ , \new_[2059]_ , \new_[2062]_ , \new_[2063]_ ,
    \new_[2066]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2075]_ , \new_[2078]_ , \new_[2079]_ , \new_[2082]_ ,
    \new_[2086]_ , \new_[2087]_ , \new_[2088]_ , \new_[2091]_ ,
    \new_[2094]_ , \new_[2095]_ , \new_[2098]_ , \new_[2102]_ ,
    \new_[2103]_ , \new_[2104]_ , \new_[2107]_ , \new_[2110]_ ,
    \new_[2111]_ , \new_[2114]_ , \new_[2118]_ , \new_[2119]_ ,
    \new_[2120]_ , \new_[2123]_ , \new_[2126]_ , \new_[2127]_ ,
    \new_[2130]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2139]_ , \new_[2142]_ , \new_[2143]_ , \new_[2146]_ ,
    \new_[2150]_ , \new_[2151]_ , \new_[2152]_ , \new_[2155]_ ,
    \new_[2158]_ , \new_[2159]_ , \new_[2162]_ , \new_[2166]_ ,
    \new_[2167]_ , \new_[2168]_ , \new_[2171]_ , \new_[2174]_ ,
    \new_[2175]_ , \new_[2178]_ , \new_[2182]_ , \new_[2183]_ ,
    \new_[2184]_ , \new_[2187]_ , \new_[2190]_ , \new_[2191]_ ,
    \new_[2194]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2203]_ , \new_[2206]_ , \new_[2207]_ , \new_[2210]_ ,
    \new_[2214]_ , \new_[2215]_ , \new_[2216]_ , \new_[2219]_ ,
    \new_[2222]_ , \new_[2223]_ , \new_[2226]_ , \new_[2230]_ ,
    \new_[2231]_ , \new_[2232]_ , \new_[2235]_ , \new_[2238]_ ,
    \new_[2239]_ , \new_[2242]_ , \new_[2246]_ , \new_[2247]_ ,
    \new_[2248]_ , \new_[2251]_ , \new_[2254]_ , \new_[2255]_ ,
    \new_[2258]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2267]_ , \new_[2270]_ , \new_[2271]_ , \new_[2274]_ ,
    \new_[2278]_ , \new_[2279]_ , \new_[2280]_ , \new_[2283]_ ,
    \new_[2286]_ , \new_[2287]_ , \new_[2290]_ , \new_[2294]_ ,
    \new_[2295]_ , \new_[2296]_ , \new_[2299]_ , \new_[2302]_ ,
    \new_[2303]_ , \new_[2306]_ , \new_[2310]_ , \new_[2311]_ ,
    \new_[2312]_ , \new_[2315]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2324]_ , \new_[2328]_ , \new_[2329]_ ,
    \new_[2330]_ , \new_[2333]_ , \new_[2337]_ , \new_[2338]_ ,
    \new_[2339]_ , \new_[2342]_ , \new_[2346]_ , \new_[2347]_ ,
    \new_[2348]_ , \new_[2351]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2360]_ , \new_[2364]_ , \new_[2365]_ ,
    \new_[2366]_ , \new_[2369]_ , \new_[2373]_ , \new_[2374]_ ,
    \new_[2375]_ , \new_[2378]_ , \new_[2382]_ , \new_[2383]_ ,
    \new_[2384]_ , \new_[2387]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2396]_ , \new_[2400]_ , \new_[2401]_ ,
    \new_[2402]_ , \new_[2405]_ , \new_[2409]_ , \new_[2410]_ ,
    \new_[2411]_ , \new_[2414]_ , \new_[2418]_ , \new_[2419]_ ,
    \new_[2420]_ , \new_[2423]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2432]_ , \new_[2436]_ , \new_[2437]_ ,
    \new_[2438]_ , \new_[2441]_ , \new_[2445]_ , \new_[2446]_ ,
    \new_[2447]_ , \new_[2450]_ , \new_[2454]_ , \new_[2455]_ ,
    \new_[2456]_ , \new_[2459]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2468]_ , \new_[2472]_ , \new_[2473]_ ,
    \new_[2474]_ , \new_[2477]_ , \new_[2481]_ , \new_[2482]_ ,
    \new_[2483]_ , \new_[2486]_ , \new_[2490]_ , \new_[2491]_ ,
    \new_[2492]_ , \new_[2495]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2504]_ , \new_[2508]_ , \new_[2509]_ ,
    \new_[2510]_ , \new_[2513]_ , \new_[2517]_ , \new_[2518]_ ,
    \new_[2519]_ , \new_[2522]_ , \new_[2526]_ , \new_[2527]_ ,
    \new_[2528]_ , \new_[2531]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2540]_ , \new_[2544]_ , \new_[2545]_ ,
    \new_[2546]_ , \new_[2549]_ , \new_[2553]_ , \new_[2554]_ ,
    \new_[2555]_ , \new_[2558]_ , \new_[2562]_ , \new_[2563]_ ,
    \new_[2564]_ , \new_[2567]_ , \new_[2571]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2576]_ , \new_[2580]_ , \new_[2581]_ ,
    \new_[2582]_ , \new_[2585]_ , \new_[2589]_ , \new_[2590]_ ,
    \new_[2591]_ , \new_[2594]_ , \new_[2598]_ , \new_[2599]_ ,
    \new_[2600]_ , \new_[2603]_ , \new_[2607]_ , \new_[2608]_ ,
    \new_[2609]_ , \new_[2612]_ , \new_[2616]_ , \new_[2617]_ ,
    \new_[2618]_ , \new_[2621]_ , \new_[2625]_ , \new_[2626]_ ,
    \new_[2627]_ , \new_[2630]_ , \new_[2634]_ , \new_[2635]_ ,
    \new_[2636]_ , \new_[2639]_ , \new_[2643]_ , \new_[2644]_ ,
    \new_[2645]_ , \new_[2648]_ , \new_[2652]_ , \new_[2653]_ ,
    \new_[2654]_ , \new_[2657]_ , \new_[2661]_ , \new_[2662]_ ,
    \new_[2663]_ , \new_[2666]_ , \new_[2670]_ , \new_[2671]_ ,
    \new_[2672]_ , \new_[2675]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2684]_ , \new_[2688]_ , \new_[2689]_ ,
    \new_[2690]_ , \new_[2693]_ , \new_[2697]_ , \new_[2698]_ ,
    \new_[2699]_ , \new_[2702]_ , \new_[2706]_ , \new_[2707]_ ,
    \new_[2708]_ , \new_[2711]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2720]_ , \new_[2724]_ , \new_[2725]_ ,
    \new_[2726]_ , \new_[2729]_ , \new_[2733]_ , \new_[2734]_ ,
    \new_[2735]_ , \new_[2738]_ , \new_[2742]_ , \new_[2743]_ ,
    \new_[2744]_ , \new_[2747]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2753]_ , \new_[2756]_ , \new_[2760]_ , \new_[2761]_ ,
    \new_[2762]_ , \new_[2765]_ , \new_[2769]_ , \new_[2770]_ ,
    \new_[2771]_ , \new_[2774]_ , \new_[2778]_ , \new_[2779]_ ,
    \new_[2780]_ , \new_[2783]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2792]_ , \new_[2796]_ , \new_[2797]_ ,
    \new_[2798]_ , \new_[2801]_ , \new_[2805]_ , \new_[2806]_ ,
    \new_[2807]_ , \new_[2810]_ , \new_[2814]_ , \new_[2815]_ ,
    \new_[2816]_ , \new_[2819]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2828]_ , \new_[2832]_ , \new_[2833]_ ,
    \new_[2834]_ , \new_[2837]_ , \new_[2841]_ , \new_[2842]_ ,
    \new_[2843]_ , \new_[2846]_ , \new_[2850]_ , \new_[2851]_ ,
    \new_[2852]_ , \new_[2855]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2861]_ , \new_[2864]_ , \new_[2868]_ , \new_[2869]_ ,
    \new_[2870]_ , \new_[2873]_ , \new_[2877]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2882]_ , \new_[2886]_ , \new_[2887]_ ,
    \new_[2888]_ , \new_[2891]_ , \new_[2895]_ , \new_[2896]_ ,
    \new_[2897]_ , \new_[2900]_ , \new_[2904]_ , \new_[2905]_ ,
    \new_[2906]_ , \new_[2909]_ , \new_[2913]_ , \new_[2914]_ ,
    \new_[2915]_ , \new_[2918]_ , \new_[2922]_ , \new_[2923]_ ,
    \new_[2924]_ , \new_[2927]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2936]_ , \new_[2940]_ , \new_[2941]_ ,
    \new_[2942]_ , \new_[2945]_ , \new_[2949]_ , \new_[2950]_ ,
    \new_[2951]_ , \new_[2954]_ , \new_[2958]_ , \new_[2959]_ ,
    \new_[2960]_ , \new_[2963]_ , \new_[2967]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2972]_ , \new_[2976]_ , \new_[2977]_ ,
    \new_[2978]_ , \new_[2981]_ , \new_[2985]_ , \new_[2986]_ ,
    \new_[2987]_ , \new_[2990]_ , \new_[2994]_ , \new_[2995]_ ,
    \new_[2996]_ , \new_[2999]_ , \new_[3003]_ , \new_[3004]_ ,
    \new_[3005]_ , \new_[3008]_ , \new_[3012]_ , \new_[3013]_ ,
    \new_[3014]_ , \new_[3017]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3023]_ , \new_[3026]_ , \new_[3030]_ , \new_[3031]_ ,
    \new_[3032]_ , \new_[3035]_ , \new_[3039]_ , \new_[3040]_ ,
    \new_[3041]_ , \new_[3044]_ , \new_[3048]_ , \new_[3049]_ ,
    \new_[3050]_ , \new_[3053]_ , \new_[3057]_ , \new_[3058]_ ,
    \new_[3059]_ , \new_[3062]_ , \new_[3066]_ , \new_[3067]_ ,
    \new_[3068]_ , \new_[3071]_ , \new_[3075]_ , \new_[3076]_ ,
    \new_[3077]_ , \new_[3080]_ , \new_[3084]_ , \new_[3085]_ ,
    \new_[3086]_ , \new_[3089]_ , \new_[3093]_ , \new_[3094]_ ,
    \new_[3095]_ , \new_[3098]_ , \new_[3102]_ , \new_[3103]_ ,
    \new_[3104]_ , \new_[3107]_ , \new_[3111]_ , \new_[3112]_ ,
    \new_[3113]_ , \new_[3116]_ , \new_[3120]_ , \new_[3121]_ ,
    \new_[3122]_ , \new_[3125]_ , \new_[3129]_ , \new_[3130]_ ,
    \new_[3131]_ , \new_[3134]_ , \new_[3138]_ , \new_[3139]_ ,
    \new_[3140]_ , \new_[3143]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3152]_ , \new_[3156]_ , \new_[3157]_ ,
    \new_[3158]_ , \new_[3161]_ , \new_[3165]_ , \new_[3166]_ ,
    \new_[3167]_ , \new_[3170]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3179]_ , \new_[3183]_ , \new_[3184]_ ,
    \new_[3185]_ , \new_[3188]_ , \new_[3192]_ , \new_[3193]_ ,
    \new_[3194]_ , \new_[3197]_ , \new_[3201]_ , \new_[3202]_ ,
    \new_[3203]_ , \new_[3206]_ , \new_[3210]_ , \new_[3211]_ ,
    \new_[3212]_ , \new_[3215]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3221]_ , \new_[3224]_ , \new_[3228]_ , \new_[3229]_ ,
    \new_[3230]_ , \new_[3233]_ , \new_[3237]_ , \new_[3238]_ ,
    \new_[3239]_ , \new_[3242]_ , \new_[3246]_ , \new_[3247]_ ,
    \new_[3248]_ , \new_[3251]_ , \new_[3255]_ , \new_[3256]_ ,
    \new_[3257]_ , \new_[3260]_ , \new_[3264]_ , \new_[3265]_ ,
    \new_[3266]_ , \new_[3269]_ , \new_[3273]_ , \new_[3274]_ ,
    \new_[3275]_ , \new_[3278]_ , \new_[3282]_ , \new_[3283]_ ,
    \new_[3284]_ , \new_[3287]_ , \new_[3291]_ , \new_[3292]_ ,
    \new_[3293]_ , \new_[3296]_ , \new_[3300]_ , \new_[3301]_ ,
    \new_[3302]_ , \new_[3305]_ , \new_[3309]_ , \new_[3310]_ ,
    \new_[3311]_ , \new_[3314]_ , \new_[3318]_ , \new_[3319]_ ,
    \new_[3320]_ , \new_[3323]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3332]_ , \new_[3336]_ , \new_[3337]_ ,
    \new_[3338]_ , \new_[3341]_ , \new_[3345]_ , \new_[3346]_ ,
    \new_[3347]_ , \new_[3350]_ , \new_[3354]_ , \new_[3355]_ ,
    \new_[3356]_ , \new_[3359]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3368]_ , \new_[3372]_ , \new_[3373]_ ,
    \new_[3374]_ , \new_[3377]_ , \new_[3381]_ , \new_[3382]_ ,
    \new_[3383]_ , \new_[3386]_ , \new_[3390]_ , \new_[3391]_ ,
    \new_[3392]_ , \new_[3395]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3404]_ , \new_[3408]_ , \new_[3409]_ ,
    \new_[3410]_ , \new_[3413]_ , \new_[3417]_ , \new_[3418]_ ,
    \new_[3419]_ , \new_[3422]_ , \new_[3426]_ , \new_[3427]_ ,
    \new_[3428]_ , \new_[3431]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3440]_ , \new_[3444]_ , \new_[3445]_ ,
    \new_[3446]_ , \new_[3449]_ , \new_[3453]_ , \new_[3454]_ ,
    \new_[3455]_ , \new_[3458]_ , \new_[3462]_ , \new_[3463]_ ,
    \new_[3464]_ , \new_[3467]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3476]_ , \new_[3480]_ , \new_[3481]_ ,
    \new_[3482]_ , \new_[3485]_ , \new_[3489]_ , \new_[3490]_ ,
    \new_[3491]_ , \new_[3494]_ , \new_[3498]_ , \new_[3499]_ ,
    \new_[3500]_ , \new_[3503]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3512]_ , \new_[3516]_ , \new_[3517]_ ,
    \new_[3518]_ , \new_[3521]_ , \new_[3525]_ , \new_[3526]_ ,
    \new_[3527]_ , \new_[3530]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3536]_ , \new_[3539]_ , \new_[3543]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3548]_ , \new_[3552]_ , \new_[3553]_ ,
    \new_[3554]_ , \new_[3557]_ , \new_[3561]_ , \new_[3562]_ ,
    \new_[3563]_ , \new_[3566]_ , \new_[3570]_ , \new_[3571]_ ,
    \new_[3572]_ , \new_[3575]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3584]_ , \new_[3588]_ , \new_[3589]_ ,
    \new_[3590]_ , \new_[3593]_ , \new_[3597]_ , \new_[3598]_ ,
    \new_[3599]_ , \new_[3602]_ , \new_[3606]_ , \new_[3607]_ ,
    \new_[3608]_ , \new_[3611]_ , \new_[3615]_ , \new_[3616]_ ,
    \new_[3617]_ , \new_[3620]_ , \new_[3624]_ , \new_[3625]_ ,
    \new_[3626]_ , \new_[3629]_ , \new_[3633]_ , \new_[3634]_ ,
    \new_[3635]_ , \new_[3638]_ , \new_[3642]_ , \new_[3643]_ ,
    \new_[3644]_ , \new_[3647]_ , \new_[3651]_ , \new_[3652]_ ,
    \new_[3653]_ , \new_[3656]_ , \new_[3660]_ , \new_[3661]_ ,
    \new_[3662]_ , \new_[3665]_ , \new_[3669]_ , \new_[3670]_ ,
    \new_[3671]_ , \new_[3674]_ , \new_[3678]_ , \new_[3679]_ ,
    \new_[3680]_ , \new_[3683]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3692]_ , \new_[3696]_ , \new_[3697]_ ,
    \new_[3698]_ , \new_[3701]_ , \new_[3705]_ , \new_[3706]_ ,
    \new_[3707]_ , \new_[3710]_ , \new_[3714]_ , \new_[3715]_ ,
    \new_[3716]_ , \new_[3719]_ , \new_[3723]_ , \new_[3724]_ ,
    \new_[3725]_ , \new_[3728]_ , \new_[3732]_ , \new_[3733]_ ,
    \new_[3734]_ , \new_[3737]_ , \new_[3741]_ , \new_[3742]_ ,
    \new_[3743]_ , \new_[3746]_ , \new_[3750]_ , \new_[3751]_ ,
    \new_[3752]_ , \new_[3755]_ , \new_[3759]_ , \new_[3760]_ ,
    \new_[3761]_ , \new_[3764]_ , \new_[3768]_ , \new_[3769]_ ,
    \new_[3770]_ , \new_[3773]_ , \new_[3777]_ , \new_[3778]_ ,
    \new_[3779]_ , \new_[3782]_ , \new_[3786]_ , \new_[3787]_ ,
    \new_[3788]_ , \new_[3791]_ , \new_[3795]_ , \new_[3796]_ ,
    \new_[3797]_ , \new_[3800]_ , \new_[3804]_ , \new_[3805]_ ,
    \new_[3806]_ , \new_[3809]_ , \new_[3813]_ , \new_[3814]_ ,
    \new_[3815]_ , \new_[3818]_ , \new_[3822]_ , \new_[3823]_ ,
    \new_[3824]_ , \new_[3827]_ , \new_[3831]_ , \new_[3832]_ ,
    \new_[3833]_ , \new_[3836]_ , \new_[3840]_ , \new_[3841]_ ,
    \new_[3842]_ , \new_[3845]_ , \new_[3849]_ , \new_[3850]_ ,
    \new_[3851]_ , \new_[3854]_ , \new_[3858]_ , \new_[3859]_ ,
    \new_[3860]_ , \new_[3863]_ , \new_[3867]_ , \new_[3868]_ ,
    \new_[3869]_ , \new_[3872]_ , \new_[3876]_ , \new_[3877]_ ,
    \new_[3878]_ , \new_[3881]_ , \new_[3885]_ , \new_[3886]_ ,
    \new_[3887]_ , \new_[3890]_ , \new_[3894]_ , \new_[3895]_ ,
    \new_[3896]_ , \new_[3899]_ , \new_[3903]_ , \new_[3904]_ ,
    \new_[3905]_ , \new_[3908]_ , \new_[3912]_ , \new_[3913]_ ,
    \new_[3914]_ , \new_[3917]_ , \new_[3921]_ , \new_[3922]_ ,
    \new_[3923]_ , \new_[3926]_ , \new_[3930]_ , \new_[3931]_ ,
    \new_[3932]_ , \new_[3935]_ , \new_[3939]_ , \new_[3940]_ ,
    \new_[3941]_ , \new_[3944]_ , \new_[3948]_ , \new_[3949]_ ,
    \new_[3950]_ , \new_[3953]_ , \new_[3957]_ , \new_[3958]_ ,
    \new_[3959]_ , \new_[3962]_ , \new_[3966]_ , \new_[3967]_ ,
    \new_[3968]_ , \new_[3971]_ , \new_[3975]_ , \new_[3976]_ ,
    \new_[3977]_ , \new_[3980]_ , \new_[3984]_ , \new_[3985]_ ,
    \new_[3986]_ , \new_[3989]_ , \new_[3993]_ , \new_[3994]_ ,
    \new_[3995]_ , \new_[3998]_ , \new_[4002]_ , \new_[4003]_ ,
    \new_[4004]_ , \new_[4007]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4013]_ , \new_[4016]_ , \new_[4020]_ , \new_[4021]_ ,
    \new_[4022]_ , \new_[4025]_ , \new_[4029]_ , \new_[4030]_ ,
    \new_[4031]_ , \new_[4034]_ , \new_[4038]_ , \new_[4039]_ ,
    \new_[4040]_ , \new_[4043]_ , \new_[4047]_ , \new_[4048]_ ,
    \new_[4049]_ , \new_[4052]_ , \new_[4056]_ , \new_[4057]_ ,
    \new_[4058]_ , \new_[4061]_ , \new_[4065]_ , \new_[4066]_ ,
    \new_[4067]_ , \new_[4070]_ , \new_[4074]_ , \new_[4075]_ ,
    \new_[4076]_ , \new_[4079]_ , \new_[4083]_ , \new_[4084]_ ,
    \new_[4085]_ , \new_[4088]_ , \new_[4092]_ , \new_[4093]_ ,
    \new_[4094]_ , \new_[4097]_ , \new_[4101]_ , \new_[4102]_ ,
    \new_[4103]_ , \new_[4106]_ , \new_[4110]_ , \new_[4111]_ ,
    \new_[4112]_ , \new_[4115]_ , \new_[4119]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4124]_ , \new_[4128]_ , \new_[4129]_ ,
    \new_[4130]_ , \new_[4133]_ , \new_[4137]_ , \new_[4138]_ ,
    \new_[4139]_ , \new_[4142]_ , \new_[4146]_ , \new_[4147]_ ,
    \new_[4148]_ , \new_[4151]_ , \new_[4155]_ , \new_[4156]_ ,
    \new_[4157]_ , \new_[4160]_ , \new_[4164]_ , \new_[4165]_ ,
    \new_[4166]_ , \new_[4169]_ , \new_[4173]_ , \new_[4174]_ ,
    \new_[4175]_ , \new_[4178]_ , \new_[4182]_ , \new_[4183]_ ,
    \new_[4184]_ , \new_[4187]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4193]_ , \new_[4196]_ , \new_[4200]_ , \new_[4201]_ ,
    \new_[4202]_ , \new_[4205]_ , \new_[4209]_ , \new_[4210]_ ,
    \new_[4211]_ , \new_[4214]_ , \new_[4218]_ , \new_[4219]_ ,
    \new_[4220]_ , \new_[4223]_ , \new_[4227]_ , \new_[4228]_ ,
    \new_[4229]_ , \new_[4232]_ , \new_[4236]_ , \new_[4237]_ ,
    \new_[4238]_ , \new_[4241]_ , \new_[4245]_ , \new_[4246]_ ,
    \new_[4247]_ , \new_[4250]_ , \new_[4254]_ , \new_[4255]_ ,
    \new_[4256]_ , \new_[4259]_ , \new_[4263]_ , \new_[4264]_ ,
    \new_[4265]_ , \new_[4268]_ , \new_[4272]_ , \new_[4273]_ ,
    \new_[4274]_ , \new_[4277]_ , \new_[4281]_ , \new_[4282]_ ,
    \new_[4283]_ , \new_[4286]_ , \new_[4290]_ , \new_[4291]_ ,
    \new_[4292]_ , \new_[4295]_ , \new_[4299]_ , \new_[4300]_ ,
    \new_[4301]_ , \new_[4304]_ , \new_[4308]_ , \new_[4309]_ ,
    \new_[4310]_ , \new_[4313]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4319]_ , \new_[4322]_ , \new_[4326]_ , \new_[4327]_ ,
    \new_[4328]_ , \new_[4331]_ , \new_[4335]_ , \new_[4336]_ ,
    \new_[4337]_ , \new_[4340]_ , \new_[4344]_ , \new_[4345]_ ,
    \new_[4346]_ , \new_[4349]_ , \new_[4353]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4358]_ , \new_[4362]_ , \new_[4363]_ ,
    \new_[4364]_ , \new_[4367]_ , \new_[4371]_ , \new_[4372]_ ,
    \new_[4373]_ , \new_[4376]_ , \new_[4380]_ , \new_[4381]_ ,
    \new_[4382]_ , \new_[4385]_ , \new_[4389]_ , \new_[4390]_ ,
    \new_[4391]_ , \new_[4394]_ , \new_[4398]_ , \new_[4399]_ ,
    \new_[4400]_ , \new_[4403]_ , \new_[4407]_ , \new_[4408]_ ,
    \new_[4409]_ , \new_[4412]_ , \new_[4416]_ , \new_[4417]_ ,
    \new_[4418]_ , \new_[4421]_ , \new_[4425]_ , \new_[4426]_ ,
    \new_[4427]_ , \new_[4430]_ , \new_[4434]_ , \new_[4435]_ ,
    \new_[4436]_ , \new_[4439]_ , \new_[4443]_ , \new_[4444]_ ,
    \new_[4445]_ , \new_[4448]_ , \new_[4452]_ , \new_[4453]_ ,
    \new_[4454]_ , \new_[4457]_ , \new_[4461]_ , \new_[4462]_ ,
    \new_[4463]_ , \new_[4466]_ , \new_[4470]_ , \new_[4471]_ ,
    \new_[4472]_ , \new_[4475]_ , \new_[4479]_ , \new_[4480]_ ,
    \new_[4481]_ , \new_[4484]_ , \new_[4488]_ , \new_[4489]_ ,
    \new_[4490]_ , \new_[4493]_ , \new_[4497]_ , \new_[4498]_ ,
    \new_[4499]_ , \new_[4502]_ , \new_[4506]_ , \new_[4507]_ ,
    \new_[4508]_ , \new_[4511]_ , \new_[4515]_ , \new_[4516]_ ,
    \new_[4517]_ , \new_[4520]_ , \new_[4524]_ , \new_[4525]_ ,
    \new_[4526]_ , \new_[4529]_ , \new_[4533]_ , \new_[4534]_ ,
    \new_[4535]_ , \new_[4538]_ , \new_[4542]_ , \new_[4543]_ ,
    \new_[4544]_ , \new_[4547]_ , \new_[4551]_ , \new_[4552]_ ,
    \new_[4553]_ , \new_[4556]_ , \new_[4560]_ , \new_[4561]_ ,
    \new_[4562]_ , \new_[4565]_ , \new_[4569]_ , \new_[4570]_ ,
    \new_[4571]_ , \new_[4574]_ , \new_[4578]_ , \new_[4579]_ ,
    \new_[4580]_ , \new_[4583]_ , \new_[4587]_ , \new_[4588]_ ,
    \new_[4589]_ , \new_[4592]_ , \new_[4596]_ , \new_[4597]_ ,
    \new_[4598]_ , \new_[4601]_ , \new_[4605]_ , \new_[4606]_ ,
    \new_[4607]_ , \new_[4610]_ , \new_[4614]_ , \new_[4615]_ ,
    \new_[4616]_ , \new_[4619]_ , \new_[4623]_ , \new_[4624]_ ,
    \new_[4625]_ , \new_[4628]_ , \new_[4632]_ , \new_[4633]_ ,
    \new_[4634]_ , \new_[4637]_ , \new_[4641]_ , \new_[4642]_ ,
    \new_[4643]_ , \new_[4646]_ , \new_[4650]_ , \new_[4651]_ ,
    \new_[4652]_ , \new_[4655]_ , \new_[4659]_ , \new_[4660]_ ,
    \new_[4661]_ , \new_[4664]_ , \new_[4668]_ , \new_[4669]_ ,
    \new_[4670]_ , \new_[4673]_ , \new_[4677]_ , \new_[4678]_ ,
    \new_[4679]_ , \new_[4682]_ , \new_[4686]_ , \new_[4687]_ ,
    \new_[4688]_ , \new_[4691]_ , \new_[4695]_ , \new_[4696]_ ,
    \new_[4697]_ , \new_[4700]_ , \new_[4704]_ , \new_[4705]_ ,
    \new_[4706]_ , \new_[4709]_ , \new_[4713]_ , \new_[4714]_ ,
    \new_[4715]_ , \new_[4718]_ , \new_[4722]_ , \new_[4723]_ ,
    \new_[4724]_ , \new_[4727]_ , \new_[4731]_ , \new_[4732]_ ,
    \new_[4733]_ , \new_[4736]_ , \new_[4740]_ , \new_[4741]_ ,
    \new_[4742]_ , \new_[4745]_ , \new_[4749]_ , \new_[4750]_ ,
    \new_[4751]_ , \new_[4754]_ , \new_[4758]_ , \new_[4759]_ ,
    \new_[4760]_ , \new_[4763]_ , \new_[4767]_ , \new_[4768]_ ,
    \new_[4769]_ , \new_[4773]_ , \new_[4774]_ , \new_[4778]_ ,
    \new_[4779]_ , \new_[4780]_ , \new_[4783]_ , \new_[4787]_ ,
    \new_[4788]_ , \new_[4789]_ , \new_[4793]_ , \new_[4794]_ ,
    \new_[4798]_ , \new_[4799]_ , \new_[4800]_ , \new_[4803]_ ,
    \new_[4807]_ , \new_[4808]_ , \new_[4809]_ , \new_[4813]_ ,
    \new_[4814]_ , \new_[4818]_ , \new_[4819]_ , \new_[4820]_ ,
    \new_[4823]_ , \new_[4827]_ , \new_[4828]_ , \new_[4829]_ ,
    \new_[4833]_ , \new_[4834]_ , \new_[4838]_ , \new_[4839]_ ,
    \new_[4840]_ , \new_[4843]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4849]_ , \new_[4853]_ , \new_[4854]_ , \new_[4858]_ ,
    \new_[4859]_ , \new_[4860]_ , \new_[4863]_ , \new_[4867]_ ,
    \new_[4868]_ , \new_[4869]_ , \new_[4873]_ , \new_[4874]_ ,
    \new_[4878]_ , \new_[4879]_ , \new_[4880]_ , \new_[4883]_ ,
    \new_[4887]_ , \new_[4888]_ , \new_[4889]_ , \new_[4893]_ ,
    \new_[4894]_ , \new_[4898]_ , \new_[4899]_ , \new_[4900]_ ,
    \new_[4903]_ , \new_[4907]_ , \new_[4908]_ , \new_[4909]_ ,
    \new_[4913]_ , \new_[4914]_ , \new_[4918]_ , \new_[4919]_ ,
    \new_[4920]_ , \new_[4923]_ , \new_[4927]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4933]_ , \new_[4934]_ , \new_[4938]_ ,
    \new_[4939]_ , \new_[4940]_ , \new_[4943]_ , \new_[4947]_ ,
    \new_[4948]_ , \new_[4949]_ , \new_[4953]_ , \new_[4954]_ ,
    \new_[4958]_ , \new_[4959]_ , \new_[4960]_ , \new_[4963]_ ,
    \new_[4967]_ , \new_[4968]_ , \new_[4969]_ , \new_[4973]_ ,
    \new_[4974]_ , \new_[4978]_ , \new_[4979]_ , \new_[4980]_ ,
    \new_[4983]_ , \new_[4987]_ , \new_[4988]_ , \new_[4989]_ ,
    \new_[4993]_ , \new_[4994]_ , \new_[4998]_ , \new_[4999]_ ,
    \new_[5000]_ , \new_[5003]_ , \new_[5007]_ , \new_[5008]_ ,
    \new_[5009]_ , \new_[5013]_ , \new_[5014]_ , \new_[5018]_ ,
    \new_[5019]_ , \new_[5020]_ , \new_[5023]_ , \new_[5027]_ ,
    \new_[5028]_ , \new_[5029]_ , \new_[5033]_ , \new_[5034]_ ,
    \new_[5038]_ , \new_[5039]_ , \new_[5040]_ , \new_[5043]_ ,
    \new_[5047]_ , \new_[5048]_ , \new_[5049]_ , \new_[5053]_ ,
    \new_[5054]_ , \new_[5058]_ , \new_[5059]_ , \new_[5060]_ ,
    \new_[5063]_ , \new_[5067]_ , \new_[5068]_ , \new_[5069]_ ,
    \new_[5073]_ , \new_[5074]_ , \new_[5078]_ , \new_[5079]_ ,
    \new_[5080]_ , \new_[5083]_ , \new_[5087]_ , \new_[5088]_ ,
    \new_[5089]_ , \new_[5093]_ , \new_[5094]_ , \new_[5098]_ ,
    \new_[5099]_ , \new_[5100]_ , \new_[5103]_ , \new_[5107]_ ,
    \new_[5108]_ , \new_[5109]_ , \new_[5113]_ , \new_[5114]_ ,
    \new_[5118]_ , \new_[5119]_ , \new_[5120]_ , \new_[5123]_ ,
    \new_[5127]_ , \new_[5128]_ , \new_[5129]_ , \new_[5133]_ ,
    \new_[5134]_ , \new_[5138]_ , \new_[5139]_ , \new_[5140]_ ,
    \new_[5143]_ , \new_[5147]_ , \new_[5148]_ , \new_[5149]_ ,
    \new_[5153]_ , \new_[5154]_ , \new_[5158]_ , \new_[5159]_ ,
    \new_[5160]_ , \new_[5163]_ , \new_[5167]_ , \new_[5168]_ ,
    \new_[5169]_ , \new_[5173]_ , \new_[5174]_ , \new_[5178]_ ,
    \new_[5179]_ , \new_[5180]_ , \new_[5183]_ , \new_[5187]_ ,
    \new_[5188]_ , \new_[5189]_ , \new_[5193]_ , \new_[5194]_ ,
    \new_[5198]_ , \new_[5199]_ , \new_[5200]_ , \new_[5203]_ ,
    \new_[5207]_ , \new_[5208]_ , \new_[5209]_ , \new_[5213]_ ,
    \new_[5214]_ , \new_[5218]_ , \new_[5219]_ , \new_[5220]_ ,
    \new_[5223]_ , \new_[5227]_ , \new_[5228]_ , \new_[5229]_ ,
    \new_[5233]_ , \new_[5234]_ , \new_[5238]_ , \new_[5239]_ ,
    \new_[5240]_ , \new_[5243]_ , \new_[5247]_ , \new_[5248]_ ,
    \new_[5249]_ , \new_[5253]_ , \new_[5254]_ , \new_[5258]_ ,
    \new_[5259]_ , \new_[5260]_ , \new_[5263]_ , \new_[5267]_ ,
    \new_[5268]_ , \new_[5269]_ , \new_[5273]_ , \new_[5274]_ ,
    \new_[5278]_ , \new_[5279]_ , \new_[5280]_ , \new_[5283]_ ,
    \new_[5287]_ , \new_[5288]_ , \new_[5289]_ , \new_[5293]_ ,
    \new_[5294]_ , \new_[5298]_ , \new_[5299]_ , \new_[5300]_ ,
    \new_[5303]_ , \new_[5307]_ , \new_[5308]_ , \new_[5309]_ ,
    \new_[5313]_ , \new_[5314]_ , \new_[5318]_ , \new_[5319]_ ,
    \new_[5320]_ , \new_[5323]_ , \new_[5327]_ , \new_[5328]_ ,
    \new_[5329]_ , \new_[5333]_ , \new_[5334]_ , \new_[5338]_ ,
    \new_[5339]_ , \new_[5340]_ , \new_[5343]_ , \new_[5347]_ ,
    \new_[5348]_ , \new_[5349]_ , \new_[5353]_ , \new_[5354]_ ,
    \new_[5358]_ , \new_[5359]_ , \new_[5360]_ , \new_[5363]_ ,
    \new_[5367]_ , \new_[5368]_ , \new_[5369]_ , \new_[5373]_ ,
    \new_[5374]_ , \new_[5378]_ , \new_[5379]_ , \new_[5380]_ ,
    \new_[5383]_ , \new_[5387]_ , \new_[5388]_ , \new_[5389]_ ,
    \new_[5393]_ , \new_[5394]_ , \new_[5398]_ , \new_[5399]_ ,
    \new_[5400]_ , \new_[5403]_ , \new_[5407]_ , \new_[5408]_ ,
    \new_[5409]_ , \new_[5413]_ , \new_[5414]_ , \new_[5418]_ ,
    \new_[5419]_ , \new_[5420]_ , \new_[5423]_ , \new_[5427]_ ,
    \new_[5428]_ , \new_[5429]_ , \new_[5433]_ , \new_[5434]_ ,
    \new_[5438]_ , \new_[5439]_ , \new_[5440]_ , \new_[5443]_ ,
    \new_[5447]_ , \new_[5448]_ , \new_[5449]_ , \new_[5453]_ ,
    \new_[5454]_ , \new_[5458]_ , \new_[5459]_ , \new_[5460]_ ,
    \new_[5463]_ , \new_[5467]_ , \new_[5468]_ , \new_[5469]_ ,
    \new_[5473]_ , \new_[5474]_ , \new_[5478]_ , \new_[5479]_ ,
    \new_[5480]_ , \new_[5483]_ , \new_[5487]_ , \new_[5488]_ ,
    \new_[5489]_ , \new_[5493]_ , \new_[5494]_ , \new_[5498]_ ,
    \new_[5499]_ , \new_[5500]_ , \new_[5503]_ , \new_[5507]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5513]_ , \new_[5514]_ ,
    \new_[5518]_ , \new_[5519]_ , \new_[5520]_ , \new_[5523]_ ,
    \new_[5527]_ , \new_[5528]_ , \new_[5529]_ , \new_[5533]_ ,
    \new_[5534]_ , \new_[5538]_ , \new_[5539]_ , \new_[5540]_ ,
    \new_[5543]_ , \new_[5547]_ , \new_[5548]_ , \new_[5549]_ ,
    \new_[5553]_ , \new_[5554]_ , \new_[5558]_ , \new_[5559]_ ,
    \new_[5560]_ , \new_[5563]_ , \new_[5567]_ , \new_[5568]_ ,
    \new_[5569]_ , \new_[5573]_ , \new_[5574]_ , \new_[5578]_ ,
    \new_[5579]_ , \new_[5580]_ , \new_[5583]_ , \new_[5587]_ ,
    \new_[5588]_ , \new_[5589]_ , \new_[5593]_ , \new_[5594]_ ,
    \new_[5598]_ , \new_[5599]_ , \new_[5600]_ , \new_[5603]_ ,
    \new_[5607]_ , \new_[5608]_ , \new_[5609]_ , \new_[5613]_ ,
    \new_[5614]_ , \new_[5618]_ , \new_[5619]_ , \new_[5620]_ ,
    \new_[5623]_ , \new_[5627]_ , \new_[5628]_ , \new_[5629]_ ,
    \new_[5633]_ , \new_[5634]_ , \new_[5638]_ , \new_[5639]_ ,
    \new_[5640]_ , \new_[5643]_ , \new_[5647]_ , \new_[5648]_ ,
    \new_[5649]_ , \new_[5653]_ , \new_[5654]_ , \new_[5658]_ ,
    \new_[5659]_ , \new_[5660]_ , \new_[5663]_ , \new_[5667]_ ,
    \new_[5668]_ , \new_[5669]_ , \new_[5673]_ , \new_[5674]_ ,
    \new_[5678]_ , \new_[5679]_ , \new_[5680]_ , \new_[5683]_ ,
    \new_[5687]_ , \new_[5688]_ , \new_[5689]_ , \new_[5693]_ ,
    \new_[5694]_ , \new_[5698]_ , \new_[5699]_ , \new_[5700]_ ,
    \new_[5703]_ , \new_[5707]_ , \new_[5708]_ , \new_[5709]_ ,
    \new_[5713]_ , \new_[5714]_ , \new_[5718]_ , \new_[5719]_ ,
    \new_[5720]_ , \new_[5723]_ , \new_[5727]_ , \new_[5728]_ ,
    \new_[5729]_ , \new_[5733]_ , \new_[5734]_ , \new_[5738]_ ,
    \new_[5739]_ , \new_[5740]_ , \new_[5743]_ , \new_[5747]_ ,
    \new_[5748]_ , \new_[5749]_ , \new_[5753]_ , \new_[5754]_ ,
    \new_[5758]_ , \new_[5759]_ , \new_[5760]_ , \new_[5763]_ ,
    \new_[5767]_ , \new_[5768]_ , \new_[5769]_ , \new_[5773]_ ,
    \new_[5774]_ , \new_[5778]_ , \new_[5779]_ , \new_[5780]_ ,
    \new_[5783]_ , \new_[5787]_ , \new_[5788]_ , \new_[5789]_ ,
    \new_[5793]_ , \new_[5794]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5800]_ , \new_[5803]_ , \new_[5807]_ , \new_[5808]_ ,
    \new_[5809]_ , \new_[5813]_ , \new_[5814]_ , \new_[5818]_ ,
    \new_[5819]_ , \new_[5820]_ , \new_[5823]_ , \new_[5827]_ ,
    \new_[5828]_ , \new_[5829]_ , \new_[5833]_ , \new_[5834]_ ,
    \new_[5838]_ , \new_[5839]_ , \new_[5840]_ , \new_[5843]_ ,
    \new_[5847]_ , \new_[5848]_ , \new_[5849]_ , \new_[5853]_ ,
    \new_[5854]_ , \new_[5858]_ , \new_[5859]_ , \new_[5860]_ ,
    \new_[5863]_ , \new_[5867]_ , \new_[5868]_ , \new_[5869]_ ,
    \new_[5873]_ , \new_[5874]_ , \new_[5878]_ , \new_[5879]_ ,
    \new_[5880]_ , \new_[5883]_ , \new_[5887]_ , \new_[5888]_ ,
    \new_[5889]_ , \new_[5893]_ , \new_[5894]_ , \new_[5898]_ ,
    \new_[5899]_ , \new_[5900]_ , \new_[5903]_ , \new_[5907]_ ,
    \new_[5908]_ , \new_[5909]_ , \new_[5913]_ , \new_[5914]_ ,
    \new_[5918]_ , \new_[5919]_ , \new_[5920]_ , \new_[5923]_ ,
    \new_[5927]_ , \new_[5928]_ , \new_[5929]_ , \new_[5933]_ ,
    \new_[5934]_ , \new_[5938]_ , \new_[5939]_ , \new_[5940]_ ,
    \new_[5943]_ , \new_[5947]_ , \new_[5948]_ , \new_[5949]_ ,
    \new_[5953]_ , \new_[5954]_ , \new_[5958]_ , \new_[5959]_ ,
    \new_[5960]_ , \new_[5963]_ , \new_[5967]_ , \new_[5968]_ ,
    \new_[5969]_ , \new_[5973]_ , \new_[5974]_ , \new_[5978]_ ,
    \new_[5979]_ , \new_[5980]_ , \new_[5983]_ , \new_[5987]_ ,
    \new_[5988]_ , \new_[5989]_ , \new_[5993]_ , \new_[5994]_ ,
    \new_[5998]_ , \new_[5999]_ , \new_[6000]_ , \new_[6003]_ ,
    \new_[6007]_ , \new_[6008]_ , \new_[6009]_ , \new_[6013]_ ,
    \new_[6014]_ , \new_[6018]_ , \new_[6019]_ , \new_[6020]_ ,
    \new_[6023]_ , \new_[6027]_ , \new_[6028]_ , \new_[6029]_ ,
    \new_[6033]_ , \new_[6034]_ , \new_[6038]_ , \new_[6039]_ ,
    \new_[6040]_ , \new_[6043]_ , \new_[6047]_ , \new_[6048]_ ,
    \new_[6049]_ , \new_[6053]_ , \new_[6054]_ , \new_[6058]_ ,
    \new_[6059]_ , \new_[6060]_ , \new_[6063]_ , \new_[6067]_ ,
    \new_[6068]_ , \new_[6069]_ , \new_[6073]_ , \new_[6074]_ ,
    \new_[6078]_ , \new_[6079]_ , \new_[6080]_ , \new_[6083]_ ,
    \new_[6087]_ , \new_[6088]_ , \new_[6089]_ , \new_[6093]_ ,
    \new_[6094]_ , \new_[6098]_ , \new_[6099]_ , \new_[6100]_ ,
    \new_[6103]_ , \new_[6107]_ , \new_[6108]_ , \new_[6109]_ ,
    \new_[6113]_ , \new_[6114]_ , \new_[6118]_ , \new_[6119]_ ,
    \new_[6120]_ , \new_[6123]_ , \new_[6127]_ , \new_[6128]_ ,
    \new_[6129]_ , \new_[6133]_ , \new_[6134]_ , \new_[6138]_ ,
    \new_[6139]_ , \new_[6140]_ , \new_[6143]_ , \new_[6147]_ ,
    \new_[6148]_ , \new_[6149]_ , \new_[6153]_ , \new_[6154]_ ,
    \new_[6158]_ , \new_[6159]_ , \new_[6160]_ , \new_[6163]_ ,
    \new_[6167]_ , \new_[6168]_ , \new_[6169]_ , \new_[6173]_ ,
    \new_[6174]_ , \new_[6178]_ , \new_[6179]_ , \new_[6180]_ ,
    \new_[6183]_ , \new_[6187]_ , \new_[6188]_ , \new_[6189]_ ,
    \new_[6193]_ , \new_[6194]_ , \new_[6198]_ , \new_[6199]_ ,
    \new_[6200]_ , \new_[6203]_ , \new_[6207]_ , \new_[6208]_ ,
    \new_[6209]_ , \new_[6213]_ , \new_[6214]_ , \new_[6218]_ ,
    \new_[6219]_ , \new_[6220]_ , \new_[6223]_ , \new_[6227]_ ,
    \new_[6228]_ , \new_[6229]_ , \new_[6233]_ , \new_[6234]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6240]_ , \new_[6243]_ ,
    \new_[6247]_ , \new_[6248]_ , \new_[6249]_ , \new_[6253]_ ,
    \new_[6254]_ , \new_[6258]_ , \new_[6259]_ , \new_[6260]_ ,
    \new_[6263]_ , \new_[6267]_ , \new_[6268]_ , \new_[6269]_ ,
    \new_[6273]_ , \new_[6274]_ , \new_[6278]_ , \new_[6279]_ ,
    \new_[6280]_ , \new_[6283]_ , \new_[6287]_ , \new_[6288]_ ,
    \new_[6289]_ , \new_[6293]_ , \new_[6294]_ , \new_[6298]_ ,
    \new_[6299]_ , \new_[6300]_ , \new_[6303]_ , \new_[6307]_ ,
    \new_[6308]_ , \new_[6309]_ , \new_[6313]_ , \new_[6314]_ ,
    \new_[6318]_ , \new_[6319]_ , \new_[6320]_ , \new_[6323]_ ,
    \new_[6327]_ , \new_[6328]_ , \new_[6329]_ , \new_[6333]_ ,
    \new_[6334]_ , \new_[6338]_ , \new_[6339]_ , \new_[6340]_ ,
    \new_[6343]_ , \new_[6347]_ , \new_[6348]_ , \new_[6349]_ ,
    \new_[6353]_ , \new_[6354]_ , \new_[6358]_ , \new_[6359]_ ,
    \new_[6360]_ , \new_[6363]_ , \new_[6367]_ , \new_[6368]_ ,
    \new_[6369]_ , \new_[6373]_ , \new_[6374]_ , \new_[6378]_ ,
    \new_[6379]_ , \new_[6380]_ , \new_[6383]_ , \new_[6387]_ ,
    \new_[6388]_ , \new_[6389]_ , \new_[6393]_ , \new_[6394]_ ,
    \new_[6398]_ , \new_[6399]_ , \new_[6400]_ , \new_[6403]_ ,
    \new_[6407]_ , \new_[6408]_ , \new_[6409]_ , \new_[6413]_ ,
    \new_[6414]_ , \new_[6418]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6423]_ , \new_[6427]_ , \new_[6428]_ , \new_[6429]_ ,
    \new_[6433]_ , \new_[6434]_ , \new_[6438]_ , \new_[6439]_ ,
    \new_[6440]_ , \new_[6443]_ , \new_[6447]_ , \new_[6448]_ ,
    \new_[6449]_ , \new_[6453]_ , \new_[6454]_ , \new_[6458]_ ,
    \new_[6459]_ , \new_[6460]_ , \new_[6463]_ , \new_[6467]_ ,
    \new_[6468]_ , \new_[6469]_ , \new_[6473]_ , \new_[6474]_ ,
    \new_[6478]_ , \new_[6479]_ , \new_[6480]_ , \new_[6483]_ ,
    \new_[6487]_ , \new_[6488]_ , \new_[6489]_ , \new_[6493]_ ,
    \new_[6494]_ , \new_[6498]_ , \new_[6499]_ , \new_[6500]_ ,
    \new_[6503]_ , \new_[6507]_ , \new_[6508]_ , \new_[6509]_ ,
    \new_[6513]_ , \new_[6514]_ , \new_[6518]_ , \new_[6519]_ ,
    \new_[6520]_ , \new_[6523]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6529]_ , \new_[6533]_ , \new_[6534]_ , \new_[6538]_ ,
    \new_[6539]_ , \new_[6540]_ , \new_[6543]_ , \new_[6547]_ ,
    \new_[6548]_ , \new_[6549]_ , \new_[6553]_ , \new_[6554]_ ,
    \new_[6558]_ , \new_[6559]_ , \new_[6560]_ , \new_[6563]_ ,
    \new_[6567]_ , \new_[6568]_ , \new_[6569]_ , \new_[6573]_ ,
    \new_[6574]_ , \new_[6578]_ , \new_[6579]_ , \new_[6580]_ ,
    \new_[6583]_ , \new_[6587]_ , \new_[6588]_ , \new_[6589]_ ,
    \new_[6593]_ , \new_[6594]_ , \new_[6598]_ , \new_[6599]_ ,
    \new_[6600]_ , \new_[6603]_ , \new_[6607]_ , \new_[6608]_ ,
    \new_[6609]_ , \new_[6613]_ , \new_[6614]_ , \new_[6618]_ ,
    \new_[6619]_ , \new_[6620]_ , \new_[6623]_ , \new_[6627]_ ,
    \new_[6628]_ , \new_[6629]_ , \new_[6633]_ , \new_[6634]_ ,
    \new_[6638]_ , \new_[6639]_ , \new_[6640]_ , \new_[6643]_ ,
    \new_[6647]_ , \new_[6648]_ , \new_[6649]_ , \new_[6653]_ ,
    \new_[6654]_ , \new_[6658]_ , \new_[6659]_ , \new_[6660]_ ,
    \new_[6663]_ , \new_[6667]_ , \new_[6668]_ , \new_[6669]_ ,
    \new_[6673]_ , \new_[6674]_ , \new_[6678]_ , \new_[6679]_ ,
    \new_[6680]_ , \new_[6683]_ , \new_[6687]_ , \new_[6688]_ ,
    \new_[6689]_ , \new_[6693]_ , \new_[6694]_ , \new_[6698]_ ,
    \new_[6699]_ , \new_[6700]_ , \new_[6703]_ , \new_[6707]_ ,
    \new_[6708]_ , \new_[6709]_ , \new_[6713]_ , \new_[6714]_ ,
    \new_[6718]_ , \new_[6719]_ , \new_[6720]_ , \new_[6723]_ ,
    \new_[6727]_ , \new_[6728]_ , \new_[6729]_ , \new_[6733]_ ,
    \new_[6734]_ , \new_[6738]_ , \new_[6739]_ , \new_[6740]_ ,
    \new_[6743]_ , \new_[6747]_ , \new_[6748]_ , \new_[6749]_ ,
    \new_[6753]_ , \new_[6754]_ , \new_[6758]_ , \new_[6759]_ ,
    \new_[6760]_ , \new_[6763]_ , \new_[6767]_ , \new_[6768]_ ,
    \new_[6769]_ , \new_[6773]_ , \new_[6774]_ , \new_[6778]_ ,
    \new_[6779]_ , \new_[6780]_ , \new_[6783]_ , \new_[6787]_ ,
    \new_[6788]_ , \new_[6789]_ , \new_[6793]_ , \new_[6794]_ ,
    \new_[6798]_ , \new_[6799]_ , \new_[6800]_ , \new_[6803]_ ,
    \new_[6807]_ , \new_[6808]_ , \new_[6809]_ , \new_[6813]_ ,
    \new_[6814]_ , \new_[6818]_ , \new_[6819]_ , \new_[6820]_ ,
    \new_[6823]_ , \new_[6827]_ , \new_[6828]_ , \new_[6829]_ ,
    \new_[6833]_ , \new_[6834]_ , \new_[6838]_ , \new_[6839]_ ,
    \new_[6840]_ , \new_[6843]_ , \new_[6847]_ , \new_[6848]_ ,
    \new_[6849]_ , \new_[6853]_ , \new_[6854]_ , \new_[6858]_ ,
    \new_[6859]_ , \new_[6860]_ , \new_[6863]_ , \new_[6867]_ ,
    \new_[6868]_ , \new_[6869]_ , \new_[6873]_ , \new_[6874]_ ,
    \new_[6878]_ , \new_[6879]_ , \new_[6880]_ , \new_[6883]_ ,
    \new_[6887]_ , \new_[6888]_ , \new_[6889]_ , \new_[6893]_ ,
    \new_[6894]_ , \new_[6898]_ , \new_[6899]_ , \new_[6900]_ ,
    \new_[6903]_ , \new_[6907]_ , \new_[6908]_ , \new_[6909]_ ,
    \new_[6913]_ , \new_[6914]_ , \new_[6918]_ , \new_[6919]_ ,
    \new_[6920]_ , \new_[6923]_ , \new_[6927]_ , \new_[6928]_ ,
    \new_[6929]_ , \new_[6933]_ , \new_[6934]_ , \new_[6938]_ ,
    \new_[6939]_ , \new_[6940]_ , \new_[6943]_ , \new_[6947]_ ,
    \new_[6948]_ , \new_[6949]_ , \new_[6953]_ , \new_[6954]_ ,
    \new_[6958]_ , \new_[6959]_ , \new_[6960]_ , \new_[6963]_ ,
    \new_[6967]_ , \new_[6968]_ , \new_[6969]_ , \new_[6973]_ ,
    \new_[6974]_ , \new_[6978]_ , \new_[6979]_ , \new_[6980]_ ,
    \new_[6983]_ , \new_[6987]_ , \new_[6988]_ , \new_[6989]_ ,
    \new_[6993]_ , \new_[6994]_ , \new_[6998]_ , \new_[6999]_ ,
    \new_[7000]_ , \new_[7003]_ , \new_[7007]_ , \new_[7008]_ ,
    \new_[7009]_ , \new_[7013]_ , \new_[7014]_ , \new_[7018]_ ,
    \new_[7019]_ , \new_[7020]_ , \new_[7023]_ , \new_[7027]_ ,
    \new_[7028]_ , \new_[7029]_ , \new_[7033]_ , \new_[7034]_ ,
    \new_[7038]_ , \new_[7039]_ , \new_[7040]_ , \new_[7043]_ ,
    \new_[7047]_ , \new_[7048]_ , \new_[7049]_ , \new_[7053]_ ,
    \new_[7054]_ , \new_[7058]_ , \new_[7059]_ , \new_[7060]_ ,
    \new_[7063]_ , \new_[7067]_ , \new_[7068]_ , \new_[7069]_ ,
    \new_[7073]_ , \new_[7074]_ , \new_[7078]_ , \new_[7079]_ ,
    \new_[7080]_ , \new_[7083]_ , \new_[7087]_ , \new_[7088]_ ,
    \new_[7089]_ , \new_[7093]_ , \new_[7094]_ , \new_[7098]_ ,
    \new_[7099]_ , \new_[7100]_ , \new_[7103]_ , \new_[7107]_ ,
    \new_[7108]_ , \new_[7109]_ , \new_[7113]_ , \new_[7114]_ ,
    \new_[7118]_ , \new_[7119]_ , \new_[7120]_ , \new_[7123]_ ,
    \new_[7127]_ , \new_[7128]_ , \new_[7129]_ , \new_[7133]_ ,
    \new_[7134]_ , \new_[7138]_ , \new_[7139]_ , \new_[7140]_ ,
    \new_[7143]_ , \new_[7147]_ , \new_[7148]_ , \new_[7149]_ ,
    \new_[7153]_ , \new_[7154]_ , \new_[7158]_ , \new_[7159]_ ,
    \new_[7160]_ , \new_[7163]_ , \new_[7167]_ , \new_[7168]_ ,
    \new_[7169]_ , \new_[7173]_ , \new_[7174]_ , \new_[7178]_ ,
    \new_[7179]_ , \new_[7180]_ , \new_[7183]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7189]_ , \new_[7193]_ , \new_[7194]_ ,
    \new_[7198]_ , \new_[7199]_ , \new_[7200]_ , \new_[7203]_ ,
    \new_[7207]_ , \new_[7208]_ , \new_[7209]_ , \new_[7213]_ ,
    \new_[7214]_ , \new_[7218]_ , \new_[7219]_ , \new_[7220]_ ,
    \new_[7223]_ , \new_[7227]_ , \new_[7228]_ , \new_[7229]_ ,
    \new_[7233]_ , \new_[7234]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7243]_ , \new_[7247]_ , \new_[7248]_ ,
    \new_[7249]_ , \new_[7253]_ , \new_[7254]_ , \new_[7258]_ ,
    \new_[7259]_ , \new_[7260]_ , \new_[7263]_ , \new_[7267]_ ,
    \new_[7268]_ , \new_[7269]_ , \new_[7273]_ , \new_[7274]_ ,
    \new_[7278]_ , \new_[7279]_ , \new_[7280]_ , \new_[7283]_ ,
    \new_[7287]_ , \new_[7288]_ , \new_[7289]_ , \new_[7293]_ ,
    \new_[7294]_ , \new_[7298]_ , \new_[7299]_ , \new_[7300]_ ,
    \new_[7303]_ , \new_[7307]_ , \new_[7308]_ , \new_[7309]_ ,
    \new_[7313]_ , \new_[7314]_ , \new_[7318]_ , \new_[7319]_ ,
    \new_[7320]_ , \new_[7323]_ , \new_[7327]_ , \new_[7328]_ ,
    \new_[7329]_ , \new_[7333]_ , \new_[7334]_ , \new_[7338]_ ,
    \new_[7339]_ , \new_[7340]_ , \new_[7343]_ , \new_[7347]_ ,
    \new_[7348]_ , \new_[7349]_ , \new_[7353]_ , \new_[7354]_ ,
    \new_[7358]_ , \new_[7359]_ , \new_[7360]_ , \new_[7363]_ ,
    \new_[7367]_ , \new_[7368]_ , \new_[7369]_ , \new_[7373]_ ,
    \new_[7374]_ , \new_[7378]_ , \new_[7379]_ , \new_[7380]_ ,
    \new_[7383]_ , \new_[7387]_ , \new_[7388]_ , \new_[7389]_ ,
    \new_[7393]_ , \new_[7394]_ , \new_[7398]_ , \new_[7399]_ ,
    \new_[7400]_ , \new_[7403]_ , \new_[7407]_ , \new_[7408]_ ,
    \new_[7409]_ , \new_[7413]_ , \new_[7414]_ , \new_[7418]_ ,
    \new_[7419]_ , \new_[7420]_ , \new_[7423]_ , \new_[7427]_ ,
    \new_[7428]_ , \new_[7429]_ , \new_[7433]_ , \new_[7434]_ ,
    \new_[7438]_ , \new_[7439]_ , \new_[7440]_ , \new_[7443]_ ,
    \new_[7447]_ , \new_[7448]_ , \new_[7449]_ , \new_[7453]_ ,
    \new_[7454]_ , \new_[7458]_ , \new_[7459]_ , \new_[7460]_ ,
    \new_[7463]_ , \new_[7467]_ , \new_[7468]_ , \new_[7469]_ ,
    \new_[7473]_ , \new_[7474]_ , \new_[7478]_ , \new_[7479]_ ,
    \new_[7480]_ , \new_[7483]_ , \new_[7487]_ , \new_[7488]_ ,
    \new_[7489]_ , \new_[7493]_ , \new_[7494]_ , \new_[7498]_ ,
    \new_[7499]_ , \new_[7500]_ , \new_[7503]_ , \new_[7507]_ ,
    \new_[7508]_ , \new_[7509]_ , \new_[7513]_ , \new_[7514]_ ,
    \new_[7518]_ , \new_[7519]_ , \new_[7520]_ , \new_[7523]_ ,
    \new_[7527]_ , \new_[7528]_ , \new_[7529]_ , \new_[7533]_ ,
    \new_[7534]_ , \new_[7538]_ , \new_[7539]_ , \new_[7540]_ ,
    \new_[7543]_ , \new_[7547]_ , \new_[7548]_ , \new_[7549]_ ,
    \new_[7553]_ , \new_[7554]_ , \new_[7558]_ , \new_[7559]_ ,
    \new_[7560]_ , \new_[7563]_ , \new_[7567]_ , \new_[7568]_ ,
    \new_[7569]_ , \new_[7573]_ , \new_[7574]_ , \new_[7578]_ ,
    \new_[7579]_ , \new_[7580]_ , \new_[7583]_ , \new_[7587]_ ,
    \new_[7588]_ , \new_[7589]_ , \new_[7593]_ , \new_[7594]_ ,
    \new_[7598]_ , \new_[7599]_ , \new_[7600]_ , \new_[7603]_ ,
    \new_[7607]_ , \new_[7608]_ , \new_[7609]_ , \new_[7613]_ ,
    \new_[7614]_ , \new_[7618]_ , \new_[7619]_ , \new_[7620]_ ,
    \new_[7623]_ , \new_[7627]_ , \new_[7628]_ , \new_[7629]_ ,
    \new_[7633]_ , \new_[7634]_ , \new_[7638]_ , \new_[7639]_ ,
    \new_[7640]_ , \new_[7643]_ , \new_[7647]_ , \new_[7648]_ ,
    \new_[7649]_ , \new_[7653]_ , \new_[7654]_ , \new_[7658]_ ,
    \new_[7659]_ , \new_[7660]_ , \new_[7663]_ , \new_[7667]_ ,
    \new_[7668]_ , \new_[7669]_ , \new_[7673]_ , \new_[7674]_ ,
    \new_[7678]_ , \new_[7679]_ , \new_[7680]_ , \new_[7683]_ ,
    \new_[7687]_ , \new_[7688]_ , \new_[7689]_ , \new_[7693]_ ,
    \new_[7694]_ , \new_[7698]_ , \new_[7699]_ , \new_[7700]_ ,
    \new_[7703]_ , \new_[7707]_ , \new_[7708]_ , \new_[7709]_ ,
    \new_[7713]_ , \new_[7714]_ , \new_[7718]_ , \new_[7719]_ ,
    \new_[7720]_ , \new_[7723]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7733]_ , \new_[7734]_ , \new_[7738]_ ,
    \new_[7739]_ , \new_[7740]_ , \new_[7743]_ , \new_[7747]_ ,
    \new_[7748]_ , \new_[7749]_ , \new_[7753]_ , \new_[7754]_ ,
    \new_[7758]_ , \new_[7759]_ , \new_[7760]_ , \new_[7763]_ ,
    \new_[7767]_ , \new_[7768]_ , \new_[7769]_ , \new_[7773]_ ,
    \new_[7774]_ , \new_[7778]_ , \new_[7779]_ , \new_[7780]_ ,
    \new_[7783]_ , \new_[7787]_ , \new_[7788]_ , \new_[7789]_ ,
    \new_[7793]_ , \new_[7794]_ , \new_[7798]_ , \new_[7799]_ ,
    \new_[7800]_ , \new_[7803]_ , \new_[7807]_ , \new_[7808]_ ,
    \new_[7809]_ , \new_[7813]_ , \new_[7814]_ , \new_[7818]_ ,
    \new_[7819]_ , \new_[7820]_ , \new_[7823]_ , \new_[7827]_ ,
    \new_[7828]_ , \new_[7829]_ , \new_[7833]_ , \new_[7834]_ ,
    \new_[7838]_ , \new_[7839]_ , \new_[7840]_ , \new_[7843]_ ,
    \new_[7847]_ , \new_[7848]_ , \new_[7849]_ , \new_[7853]_ ,
    \new_[7854]_ , \new_[7858]_ , \new_[7859]_ , \new_[7860]_ ,
    \new_[7863]_ , \new_[7867]_ , \new_[7868]_ , \new_[7869]_ ,
    \new_[7873]_ , \new_[7874]_ , \new_[7878]_ , \new_[7879]_ ,
    \new_[7880]_ , \new_[7883]_ , \new_[7887]_ , \new_[7888]_ ,
    \new_[7889]_ , \new_[7893]_ , \new_[7894]_ , \new_[7898]_ ,
    \new_[7899]_ , \new_[7900]_ , \new_[7903]_ , \new_[7907]_ ,
    \new_[7908]_ , \new_[7909]_ , \new_[7913]_ , \new_[7914]_ ,
    \new_[7918]_ , \new_[7919]_ , \new_[7920]_ , \new_[7923]_ ,
    \new_[7927]_ , \new_[7928]_ , \new_[7929]_ , \new_[7933]_ ,
    \new_[7934]_ , \new_[7938]_ , \new_[7939]_ , \new_[7940]_ ,
    \new_[7943]_ , \new_[7947]_ , \new_[7948]_ , \new_[7949]_ ,
    \new_[7953]_ , \new_[7954]_ , \new_[7958]_ , \new_[7959]_ ,
    \new_[7960]_ , \new_[7964]_ , \new_[7965]_ , \new_[7969]_ ,
    \new_[7970]_ , \new_[7971]_ , \new_[7975]_ , \new_[7976]_ ,
    \new_[7980]_ , \new_[7981]_ , \new_[7982]_ , \new_[7986]_ ,
    \new_[7987]_ , \new_[7991]_ , \new_[7992]_ , \new_[7993]_ ,
    \new_[7997]_ , \new_[7998]_ , \new_[8002]_ , \new_[8003]_ ,
    \new_[8004]_ , \new_[8008]_ , \new_[8009]_ , \new_[8013]_ ,
    \new_[8014]_ , \new_[8015]_ , \new_[8019]_ , \new_[8020]_ ,
    \new_[8024]_ , \new_[8025]_ , \new_[8026]_ , \new_[8030]_ ,
    \new_[8031]_ , \new_[8035]_ , \new_[8036]_ , \new_[8037]_ ,
    \new_[8041]_ , \new_[8042]_ , \new_[8046]_ , \new_[8047]_ ,
    \new_[8048]_ , \new_[8052]_ , \new_[8053]_ , \new_[8057]_ ,
    \new_[8058]_ , \new_[8059]_ , \new_[8063]_ , \new_[8064]_ ,
    \new_[8068]_ , \new_[8069]_ , \new_[8070]_ , \new_[8074]_ ,
    \new_[8075]_ , \new_[8079]_ , \new_[8080]_ , \new_[8081]_ ,
    \new_[8085]_ , \new_[8086]_ , \new_[8090]_ , \new_[8091]_ ,
    \new_[8092]_ , \new_[8096]_ , \new_[8097]_ , \new_[8101]_ ,
    \new_[8102]_ , \new_[8103]_ , \new_[8107]_ , \new_[8108]_ ,
    \new_[8112]_ , \new_[8113]_ , \new_[8114]_ , \new_[8118]_ ,
    \new_[8119]_ , \new_[8123]_ , \new_[8124]_ , \new_[8125]_ ,
    \new_[8129]_ , \new_[8130]_ , \new_[8134]_ , \new_[8135]_ ,
    \new_[8136]_ , \new_[8140]_ , \new_[8141]_ , \new_[8145]_ ,
    \new_[8146]_ , \new_[8147]_ , \new_[8151]_ , \new_[8152]_ ,
    \new_[8156]_ , \new_[8157]_ , \new_[8158]_ , \new_[8162]_ ,
    \new_[8163]_ , \new_[8167]_ , \new_[8168]_ , \new_[8169]_ ,
    \new_[8173]_ , \new_[8174]_ , \new_[8178]_ , \new_[8179]_ ,
    \new_[8180]_ , \new_[8184]_ , \new_[8185]_ , \new_[8189]_ ,
    \new_[8190]_ , \new_[8191]_ , \new_[8195]_ , \new_[8196]_ ,
    \new_[8200]_ , \new_[8201]_ , \new_[8202]_ , \new_[8206]_ ,
    \new_[8207]_ , \new_[8211]_ , \new_[8212]_ , \new_[8213]_ ,
    \new_[8217]_ , \new_[8218]_ , \new_[8222]_ , \new_[8223]_ ,
    \new_[8224]_ , \new_[8228]_ , \new_[8229]_ , \new_[8233]_ ,
    \new_[8234]_ , \new_[8235]_ , \new_[8239]_ , \new_[8240]_ ,
    \new_[8244]_ , \new_[8245]_ , \new_[8246]_ , \new_[8250]_ ,
    \new_[8251]_ , \new_[8255]_ , \new_[8256]_ , \new_[8257]_ ,
    \new_[8261]_ , \new_[8262]_ , \new_[8266]_ , \new_[8267]_ ,
    \new_[8268]_ , \new_[8272]_ , \new_[8273]_ , \new_[8277]_ ,
    \new_[8278]_ , \new_[8279]_ , \new_[8283]_ , \new_[8284]_ ,
    \new_[8288]_ , \new_[8289]_ , \new_[8290]_ , \new_[8294]_ ,
    \new_[8295]_ , \new_[8299]_ , \new_[8300]_ , \new_[8301]_ ,
    \new_[8305]_ , \new_[8306]_ , \new_[8310]_ , \new_[8311]_ ,
    \new_[8312]_ , \new_[8316]_ , \new_[8317]_ , \new_[8321]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8327]_ , \new_[8328]_ ,
    \new_[8332]_ , \new_[8333]_ , \new_[8334]_ , \new_[8338]_ ,
    \new_[8339]_ , \new_[8343]_ , \new_[8344]_ , \new_[8345]_ ,
    \new_[8349]_ , \new_[8350]_ , \new_[8354]_ , \new_[8355]_ ,
    \new_[8356]_ , \new_[8360]_ , \new_[8361]_ , \new_[8365]_ ,
    \new_[8366]_ , \new_[8367]_ , \new_[8371]_ , \new_[8372]_ ,
    \new_[8376]_ , \new_[8377]_ , \new_[8378]_ , \new_[8382]_ ,
    \new_[8383]_ , \new_[8387]_ , \new_[8388]_ , \new_[8389]_ ,
    \new_[8393]_ , \new_[8394]_ , \new_[8398]_ , \new_[8399]_ ,
    \new_[8400]_ , \new_[8404]_ , \new_[8405]_ , \new_[8409]_ ,
    \new_[8410]_ , \new_[8411]_ , \new_[8415]_ , \new_[8416]_ ,
    \new_[8420]_ , \new_[8421]_ , \new_[8422]_ , \new_[8426]_ ,
    \new_[8427]_ , \new_[8431]_ , \new_[8432]_ , \new_[8433]_ ,
    \new_[8437]_ , \new_[8438]_ , \new_[8442]_ , \new_[8443]_ ,
    \new_[8444]_ , \new_[8448]_ , \new_[8449]_ , \new_[8453]_ ,
    \new_[8454]_ , \new_[8455]_ , \new_[8459]_ , \new_[8460]_ ,
    \new_[8464]_ , \new_[8465]_ , \new_[8466]_ , \new_[8470]_ ,
    \new_[8471]_ , \new_[8475]_ , \new_[8476]_ , \new_[8477]_ ,
    \new_[8481]_ , \new_[8482]_ , \new_[8486]_ , \new_[8487]_ ,
    \new_[8488]_ , \new_[8492]_ , \new_[8493]_ , \new_[8497]_ ,
    \new_[8498]_ , \new_[8499]_ , \new_[8503]_ , \new_[8504]_ ,
    \new_[8508]_ , \new_[8509]_ , \new_[8510]_ , \new_[8514]_ ,
    \new_[8515]_ , \new_[8519]_ , \new_[8520]_ , \new_[8521]_ ,
    \new_[8525]_ , \new_[8526]_ , \new_[8530]_ , \new_[8531]_ ,
    \new_[8532]_ , \new_[8536]_ , \new_[8537]_ , \new_[8541]_ ,
    \new_[8542]_ , \new_[8543]_ , \new_[8547]_ , \new_[8548]_ ,
    \new_[8552]_ , \new_[8553]_ , \new_[8554]_ , \new_[8558]_ ,
    \new_[8559]_ , \new_[8563]_ , \new_[8564]_ , \new_[8565]_ ,
    \new_[8569]_ , \new_[8570]_ , \new_[8574]_ , \new_[8575]_ ,
    \new_[8576]_ , \new_[8580]_ , \new_[8581]_ , \new_[8585]_ ,
    \new_[8586]_ , \new_[8587]_ , \new_[8591]_ , \new_[8592]_ ,
    \new_[8596]_ , \new_[8597]_ , \new_[8598]_ , \new_[8602]_ ,
    \new_[8603]_ , \new_[8607]_ , \new_[8608]_ , \new_[8609]_ ,
    \new_[8613]_ , \new_[8614]_ , \new_[8618]_ , \new_[8619]_ ,
    \new_[8620]_ , \new_[8624]_ , \new_[8625]_ , \new_[8629]_ ,
    \new_[8630]_ , \new_[8631]_ , \new_[8635]_ , \new_[8636]_ ,
    \new_[8640]_ , \new_[8641]_ , \new_[8642]_ , \new_[8646]_ ,
    \new_[8647]_ , \new_[8651]_ , \new_[8652]_ , \new_[8653]_ ,
    \new_[8657]_ , \new_[8658]_ , \new_[8662]_ , \new_[8663]_ ,
    \new_[8664]_ , \new_[8668]_ , \new_[8669]_ , \new_[8673]_ ,
    \new_[8674]_ , \new_[8675]_ , \new_[8679]_ , \new_[8680]_ ,
    \new_[8684]_ , \new_[8685]_ , \new_[8686]_ , \new_[8690]_ ,
    \new_[8691]_ , \new_[8695]_ , \new_[8696]_ , \new_[8697]_ ,
    \new_[8701]_ , \new_[8702]_ , \new_[8706]_ , \new_[8707]_ ,
    \new_[8708]_ , \new_[8712]_ , \new_[8713]_ , \new_[8717]_ ,
    \new_[8718]_ , \new_[8719]_ , \new_[8723]_ , \new_[8724]_ ,
    \new_[8728]_ , \new_[8729]_ , \new_[8730]_ , \new_[8734]_ ,
    \new_[8735]_ , \new_[8739]_ , \new_[8740]_ , \new_[8741]_ ,
    \new_[8745]_ , \new_[8746]_ , \new_[8750]_ , \new_[8751]_ ,
    \new_[8752]_ , \new_[8756]_ , \new_[8757]_ , \new_[8761]_ ,
    \new_[8762]_ , \new_[8763]_ , \new_[8767]_ , \new_[8768]_ ,
    \new_[8772]_ , \new_[8773]_ , \new_[8774]_ , \new_[8778]_ ,
    \new_[8779]_ , \new_[8783]_ , \new_[8784]_ , \new_[8785]_ ,
    \new_[8789]_ , \new_[8790]_ , \new_[8794]_ , \new_[8795]_ ,
    \new_[8796]_ , \new_[8800]_ , \new_[8801]_ , \new_[8805]_ ,
    \new_[8806]_ , \new_[8807]_ , \new_[8811]_ , \new_[8812]_ ,
    \new_[8816]_ , \new_[8817]_ , \new_[8818]_ , \new_[8822]_ ,
    \new_[8823]_ , \new_[8827]_ , \new_[8828]_ , \new_[8829]_ ,
    \new_[8833]_ , \new_[8834]_ , \new_[8838]_ , \new_[8839]_ ,
    \new_[8840]_ , \new_[8844]_ , \new_[8845]_ , \new_[8849]_ ,
    \new_[8850]_ , \new_[8851]_ , \new_[8855]_ , \new_[8856]_ ,
    \new_[8860]_ , \new_[8861]_ , \new_[8862]_ , \new_[8866]_ ,
    \new_[8867]_ , \new_[8871]_ , \new_[8872]_ , \new_[8873]_ ,
    \new_[8877]_ , \new_[8878]_ , \new_[8882]_ , \new_[8883]_ ,
    \new_[8884]_ , \new_[8888]_ , \new_[8889]_ , \new_[8893]_ ,
    \new_[8894]_ , \new_[8895]_ , \new_[8899]_ , \new_[8900]_ ,
    \new_[8904]_ , \new_[8905]_ , \new_[8906]_ , \new_[8910]_ ,
    \new_[8911]_ , \new_[8915]_ , \new_[8916]_ , \new_[8917]_ ,
    \new_[8921]_ , \new_[8922]_ , \new_[8926]_ , \new_[8927]_ ,
    \new_[8928]_ , \new_[8932]_ , \new_[8933]_ , \new_[8937]_ ,
    \new_[8938]_ , \new_[8939]_ , \new_[8943]_ , \new_[8944]_ ,
    \new_[8948]_ , \new_[8949]_ , \new_[8950]_ , \new_[8954]_ ,
    \new_[8955]_ , \new_[8959]_ , \new_[8960]_ , \new_[8961]_ ,
    \new_[8965]_ , \new_[8966]_ , \new_[8970]_ , \new_[8971]_ ,
    \new_[8972]_ , \new_[8976]_ , \new_[8977]_ , \new_[8981]_ ,
    \new_[8982]_ , \new_[8983]_ , \new_[8987]_ , \new_[8988]_ ,
    \new_[8992]_ , \new_[8993]_ , \new_[8994]_ , \new_[8998]_ ,
    \new_[8999]_ , \new_[9003]_ , \new_[9004]_ , \new_[9005]_ ,
    \new_[9009]_ , \new_[9010]_ , \new_[9014]_ , \new_[9015]_ ,
    \new_[9016]_ , \new_[9020]_ , \new_[9021]_ , \new_[9025]_ ,
    \new_[9026]_ , \new_[9027]_ , \new_[9031]_ , \new_[9032]_ ,
    \new_[9036]_ , \new_[9037]_ , \new_[9038]_ , \new_[9042]_ ,
    \new_[9043]_ , \new_[9047]_ , \new_[9048]_ , \new_[9049]_ ,
    \new_[9053]_ , \new_[9054]_ , \new_[9058]_ , \new_[9059]_ ,
    \new_[9060]_ , \new_[9064]_ , \new_[9065]_ , \new_[9069]_ ,
    \new_[9070]_ , \new_[9071]_ , \new_[9075]_ , \new_[9076]_ ,
    \new_[9080]_ , \new_[9081]_ , \new_[9082]_ , \new_[9086]_ ,
    \new_[9087]_ , \new_[9091]_ , \new_[9092]_ , \new_[9093]_ ,
    \new_[9097]_ , \new_[9098]_ , \new_[9102]_ , \new_[9103]_ ,
    \new_[9104]_ , \new_[9108]_ , \new_[9109]_ , \new_[9113]_ ,
    \new_[9114]_ , \new_[9115]_ , \new_[9119]_ , \new_[9120]_ ,
    \new_[9124]_ , \new_[9125]_ , \new_[9126]_ , \new_[9130]_ ,
    \new_[9131]_ , \new_[9135]_ , \new_[9136]_ , \new_[9137]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9146]_ , \new_[9147]_ ,
    \new_[9148]_ , \new_[9152]_ , \new_[9153]_ , \new_[9157]_ ,
    \new_[9158]_ , \new_[9159]_ , \new_[9163]_ , \new_[9164]_ ,
    \new_[9168]_ , \new_[9169]_ , \new_[9170]_ , \new_[9174]_ ,
    \new_[9175]_ , \new_[9179]_ , \new_[9180]_ , \new_[9181]_ ,
    \new_[9185]_ , \new_[9186]_ , \new_[9190]_ , \new_[9191]_ ,
    \new_[9192]_ , \new_[9196]_ , \new_[9197]_ , \new_[9201]_ ,
    \new_[9202]_ , \new_[9203]_ , \new_[9207]_ , \new_[9208]_ ,
    \new_[9212]_ , \new_[9213]_ , \new_[9214]_ , \new_[9218]_ ,
    \new_[9219]_ , \new_[9223]_ , \new_[9224]_ , \new_[9225]_ ,
    \new_[9229]_ , \new_[9230]_ , \new_[9234]_ , \new_[9235]_ ,
    \new_[9236]_ , \new_[9240]_ , \new_[9241]_ , \new_[9245]_ ,
    \new_[9246]_ , \new_[9247]_ , \new_[9251]_ , \new_[9252]_ ,
    \new_[9256]_ , \new_[9257]_ , \new_[9258]_ , \new_[9262]_ ,
    \new_[9263]_ , \new_[9267]_ , \new_[9268]_ , \new_[9269]_ ,
    \new_[9273]_ , \new_[9274]_ , \new_[9278]_ , \new_[9279]_ ,
    \new_[9280]_ , \new_[9284]_ , \new_[9285]_ , \new_[9289]_ ,
    \new_[9290]_ , \new_[9291]_ , \new_[9295]_ , \new_[9296]_ ,
    \new_[9300]_ , \new_[9301]_ , \new_[9302]_ , \new_[9306]_ ,
    \new_[9307]_ , \new_[9311]_ , \new_[9312]_ , \new_[9313]_ ,
    \new_[9317]_ , \new_[9318]_ , \new_[9322]_ , \new_[9323]_ ,
    \new_[9324]_ , \new_[9328]_ , \new_[9329]_ , \new_[9333]_ ,
    \new_[9334]_ , \new_[9335]_ , \new_[9339]_ , \new_[9340]_ ,
    \new_[9344]_ , \new_[9345]_ , \new_[9346]_ , \new_[9350]_ ,
    \new_[9351]_ , \new_[9355]_ , \new_[9356]_ , \new_[9357]_ ,
    \new_[9361]_ , \new_[9362]_ , \new_[9366]_ , \new_[9367]_ ,
    \new_[9368]_ , \new_[9372]_ , \new_[9373]_ , \new_[9377]_ ,
    \new_[9378]_ , \new_[9379]_ , \new_[9383]_ , \new_[9384]_ ,
    \new_[9387]_ , \new_[9390]_ , \new_[9391]_ , \new_[9392]_ ,
    \new_[9396]_ , \new_[9397]_ , \new_[9401]_ , \new_[9402]_ ,
    \new_[9403]_ , \new_[9407]_ , \new_[9408]_ , \new_[9411]_ ,
    \new_[9414]_ , \new_[9415]_ , \new_[9416]_ , \new_[9420]_ ,
    \new_[9421]_ , \new_[9425]_ , \new_[9426]_ , \new_[9427]_ ,
    \new_[9431]_ , \new_[9432]_ , \new_[9435]_ , \new_[9438]_ ,
    \new_[9439]_ , \new_[9440]_ , \new_[9444]_ , \new_[9445]_ ,
    \new_[9449]_ , \new_[9450]_ , \new_[9451]_ , \new_[9455]_ ,
    \new_[9456]_ , \new_[9459]_ , \new_[9462]_ , \new_[9463]_ ,
    \new_[9464]_ , \new_[9468]_ , \new_[9469]_ , \new_[9473]_ ,
    \new_[9474]_ , \new_[9475]_ , \new_[9479]_ , \new_[9480]_ ,
    \new_[9483]_ , \new_[9486]_ , \new_[9487]_ , \new_[9488]_ ,
    \new_[9492]_ , \new_[9493]_ , \new_[9497]_ , \new_[9498]_ ,
    \new_[9499]_ , \new_[9503]_ , \new_[9504]_ , \new_[9507]_ ,
    \new_[9510]_ , \new_[9511]_ , \new_[9512]_ , \new_[9516]_ ,
    \new_[9517]_ , \new_[9521]_ , \new_[9522]_ , \new_[9523]_ ,
    \new_[9527]_ , \new_[9528]_ , \new_[9531]_ , \new_[9534]_ ,
    \new_[9535]_ , \new_[9536]_ , \new_[9540]_ , \new_[9541]_ ,
    \new_[9545]_ , \new_[9546]_ , \new_[9547]_ , \new_[9551]_ ,
    \new_[9552]_ , \new_[9555]_ , \new_[9558]_ , \new_[9559]_ ,
    \new_[9560]_ ;
  assign A140 = \new_[1312]_  | \new_[875]_ ;
  assign \new_[1]_  = \new_[9560]_  & \new_[9547]_ ;
  assign \new_[2]_  = \new_[9536]_  & \new_[9523]_ ;
  assign \new_[3]_  = \new_[9512]_  & \new_[9499]_ ;
  assign \new_[4]_  = \new_[9488]_  & \new_[9475]_ ;
  assign \new_[5]_  = \new_[9464]_  & \new_[9451]_ ;
  assign \new_[6]_  = \new_[9440]_  & \new_[9427]_ ;
  assign \new_[7]_  = \new_[9416]_  & \new_[9403]_ ;
  assign \new_[8]_  = \new_[9392]_  & \new_[9379]_ ;
  assign \new_[9]_  = \new_[9368]_  & \new_[9357]_ ;
  assign \new_[10]_  = \new_[9346]_  & \new_[9335]_ ;
  assign \new_[11]_  = \new_[9324]_  & \new_[9313]_ ;
  assign \new_[12]_  = \new_[9302]_  & \new_[9291]_ ;
  assign \new_[13]_  = \new_[9280]_  & \new_[9269]_ ;
  assign \new_[14]_  = \new_[9258]_  & \new_[9247]_ ;
  assign \new_[15]_  = \new_[9236]_  & \new_[9225]_ ;
  assign \new_[16]_  = \new_[9214]_  & \new_[9203]_ ;
  assign \new_[17]_  = \new_[9192]_  & \new_[9181]_ ;
  assign \new_[18]_  = \new_[9170]_  & \new_[9159]_ ;
  assign \new_[19]_  = \new_[9148]_  & \new_[9137]_ ;
  assign \new_[20]_  = \new_[9126]_  & \new_[9115]_ ;
  assign \new_[21]_  = \new_[9104]_  & \new_[9093]_ ;
  assign \new_[22]_  = \new_[9082]_  & \new_[9071]_ ;
  assign \new_[23]_  = \new_[9060]_  & \new_[9049]_ ;
  assign \new_[24]_  = \new_[9038]_  & \new_[9027]_ ;
  assign \new_[25]_  = \new_[9016]_  & \new_[9005]_ ;
  assign \new_[26]_  = \new_[8994]_  & \new_[8983]_ ;
  assign \new_[27]_  = \new_[8972]_  & \new_[8961]_ ;
  assign \new_[28]_  = \new_[8950]_  & \new_[8939]_ ;
  assign \new_[29]_  = \new_[8928]_  & \new_[8917]_ ;
  assign \new_[30]_  = \new_[8906]_  & \new_[8895]_ ;
  assign \new_[31]_  = \new_[8884]_  & \new_[8873]_ ;
  assign \new_[32]_  = \new_[8862]_  & \new_[8851]_ ;
  assign \new_[33]_  = \new_[8840]_  & \new_[8829]_ ;
  assign \new_[34]_  = \new_[8818]_  & \new_[8807]_ ;
  assign \new_[35]_  = \new_[8796]_  & \new_[8785]_ ;
  assign \new_[36]_  = \new_[8774]_  & \new_[8763]_ ;
  assign \new_[37]_  = \new_[8752]_  & \new_[8741]_ ;
  assign \new_[38]_  = \new_[8730]_  & \new_[8719]_ ;
  assign \new_[39]_  = \new_[8708]_  & \new_[8697]_ ;
  assign \new_[40]_  = \new_[8686]_  & \new_[8675]_ ;
  assign \new_[41]_  = \new_[8664]_  & \new_[8653]_ ;
  assign \new_[42]_  = \new_[8642]_  & \new_[8631]_ ;
  assign \new_[43]_  = \new_[8620]_  & \new_[8609]_ ;
  assign \new_[44]_  = \new_[8598]_  & \new_[8587]_ ;
  assign \new_[45]_  = \new_[8576]_  & \new_[8565]_ ;
  assign \new_[46]_  = \new_[8554]_  & \new_[8543]_ ;
  assign \new_[47]_  = \new_[8532]_  & \new_[8521]_ ;
  assign \new_[48]_  = \new_[8510]_  & \new_[8499]_ ;
  assign \new_[49]_  = \new_[8488]_  & \new_[8477]_ ;
  assign \new_[50]_  = \new_[8466]_  & \new_[8455]_ ;
  assign \new_[51]_  = \new_[8444]_  & \new_[8433]_ ;
  assign \new_[52]_  = \new_[8422]_  & \new_[8411]_ ;
  assign \new_[53]_  = \new_[8400]_  & \new_[8389]_ ;
  assign \new_[54]_  = \new_[8378]_  & \new_[8367]_ ;
  assign \new_[55]_  = \new_[8356]_  & \new_[8345]_ ;
  assign \new_[56]_  = \new_[8334]_  & \new_[8323]_ ;
  assign \new_[57]_  = \new_[8312]_  & \new_[8301]_ ;
  assign \new_[58]_  = \new_[8290]_  & \new_[8279]_ ;
  assign \new_[59]_  = \new_[8268]_  & \new_[8257]_ ;
  assign \new_[60]_  = \new_[8246]_  & \new_[8235]_ ;
  assign \new_[61]_  = \new_[8224]_  & \new_[8213]_ ;
  assign \new_[62]_  = \new_[8202]_  & \new_[8191]_ ;
  assign \new_[63]_  = \new_[8180]_  & \new_[8169]_ ;
  assign \new_[64]_  = \new_[8158]_  & \new_[8147]_ ;
  assign \new_[65]_  = \new_[8136]_  & \new_[8125]_ ;
  assign \new_[66]_  = \new_[8114]_  & \new_[8103]_ ;
  assign \new_[67]_  = \new_[8092]_  & \new_[8081]_ ;
  assign \new_[68]_  = \new_[8070]_  & \new_[8059]_ ;
  assign \new_[69]_  = \new_[8048]_  & \new_[8037]_ ;
  assign \new_[70]_  = \new_[8026]_  & \new_[8015]_ ;
  assign \new_[71]_  = \new_[8004]_  & \new_[7993]_ ;
  assign \new_[72]_  = \new_[7982]_  & \new_[7971]_ ;
  assign \new_[73]_  = \new_[7960]_  & \new_[7949]_ ;
  assign \new_[74]_  = \new_[7940]_  & \new_[7929]_ ;
  assign \new_[75]_  = \new_[7920]_  & \new_[7909]_ ;
  assign \new_[76]_  = \new_[7900]_  & \new_[7889]_ ;
  assign \new_[77]_  = \new_[7880]_  & \new_[7869]_ ;
  assign \new_[78]_  = \new_[7860]_  & \new_[7849]_ ;
  assign \new_[79]_  = \new_[7840]_  & \new_[7829]_ ;
  assign \new_[80]_  = \new_[7820]_  & \new_[7809]_ ;
  assign \new_[81]_  = \new_[7800]_  & \new_[7789]_ ;
  assign \new_[82]_  = \new_[7780]_  & \new_[7769]_ ;
  assign \new_[83]_  = \new_[7760]_  & \new_[7749]_ ;
  assign \new_[84]_  = \new_[7740]_  & \new_[7729]_ ;
  assign \new_[85]_  = \new_[7720]_  & \new_[7709]_ ;
  assign \new_[86]_  = \new_[7700]_  & \new_[7689]_ ;
  assign \new_[87]_  = \new_[7680]_  & \new_[7669]_ ;
  assign \new_[88]_  = \new_[7660]_  & \new_[7649]_ ;
  assign \new_[89]_  = \new_[7640]_  & \new_[7629]_ ;
  assign \new_[90]_  = \new_[7620]_  & \new_[7609]_ ;
  assign \new_[91]_  = \new_[7600]_  & \new_[7589]_ ;
  assign \new_[92]_  = \new_[7580]_  & \new_[7569]_ ;
  assign \new_[93]_  = \new_[7560]_  & \new_[7549]_ ;
  assign \new_[94]_  = \new_[7540]_  & \new_[7529]_ ;
  assign \new_[95]_  = \new_[7520]_  & \new_[7509]_ ;
  assign \new_[96]_  = \new_[7500]_  & \new_[7489]_ ;
  assign \new_[97]_  = \new_[7480]_  & \new_[7469]_ ;
  assign \new_[98]_  = \new_[7460]_  & \new_[7449]_ ;
  assign \new_[99]_  = \new_[7440]_  & \new_[7429]_ ;
  assign \new_[100]_  = \new_[7420]_  & \new_[7409]_ ;
  assign \new_[101]_  = \new_[7400]_  & \new_[7389]_ ;
  assign \new_[102]_  = \new_[7380]_  & \new_[7369]_ ;
  assign \new_[103]_  = \new_[7360]_  & \new_[7349]_ ;
  assign \new_[104]_  = \new_[7340]_  & \new_[7329]_ ;
  assign \new_[105]_  = \new_[7320]_  & \new_[7309]_ ;
  assign \new_[106]_  = \new_[7300]_  & \new_[7289]_ ;
  assign \new_[107]_  = \new_[7280]_  & \new_[7269]_ ;
  assign \new_[108]_  = \new_[7260]_  & \new_[7249]_ ;
  assign \new_[109]_  = \new_[7240]_  & \new_[7229]_ ;
  assign \new_[110]_  = \new_[7220]_  & \new_[7209]_ ;
  assign \new_[111]_  = \new_[7200]_  & \new_[7189]_ ;
  assign \new_[112]_  = \new_[7180]_  & \new_[7169]_ ;
  assign \new_[113]_  = \new_[7160]_  & \new_[7149]_ ;
  assign \new_[114]_  = \new_[7140]_  & \new_[7129]_ ;
  assign \new_[115]_  = \new_[7120]_  & \new_[7109]_ ;
  assign \new_[116]_  = \new_[7100]_  & \new_[7089]_ ;
  assign \new_[117]_  = \new_[7080]_  & \new_[7069]_ ;
  assign \new_[118]_  = \new_[7060]_  & \new_[7049]_ ;
  assign \new_[119]_  = \new_[7040]_  & \new_[7029]_ ;
  assign \new_[120]_  = \new_[7020]_  & \new_[7009]_ ;
  assign \new_[121]_  = \new_[7000]_  & \new_[6989]_ ;
  assign \new_[122]_  = \new_[6980]_  & \new_[6969]_ ;
  assign \new_[123]_  = \new_[6960]_  & \new_[6949]_ ;
  assign \new_[124]_  = \new_[6940]_  & \new_[6929]_ ;
  assign \new_[125]_  = \new_[6920]_  & \new_[6909]_ ;
  assign \new_[126]_  = \new_[6900]_  & \new_[6889]_ ;
  assign \new_[127]_  = \new_[6880]_  & \new_[6869]_ ;
  assign \new_[128]_  = \new_[6860]_  & \new_[6849]_ ;
  assign \new_[129]_  = \new_[6840]_  & \new_[6829]_ ;
  assign \new_[130]_  = \new_[6820]_  & \new_[6809]_ ;
  assign \new_[131]_  = \new_[6800]_  & \new_[6789]_ ;
  assign \new_[132]_  = \new_[6780]_  & \new_[6769]_ ;
  assign \new_[133]_  = \new_[6760]_  & \new_[6749]_ ;
  assign \new_[134]_  = \new_[6740]_  & \new_[6729]_ ;
  assign \new_[135]_  = \new_[6720]_  & \new_[6709]_ ;
  assign \new_[136]_  = \new_[6700]_  & \new_[6689]_ ;
  assign \new_[137]_  = \new_[6680]_  & \new_[6669]_ ;
  assign \new_[138]_  = \new_[6660]_  & \new_[6649]_ ;
  assign \new_[139]_  = \new_[6640]_  & \new_[6629]_ ;
  assign \new_[140]_  = \new_[6620]_  & \new_[6609]_ ;
  assign \new_[141]_  = \new_[6600]_  & \new_[6589]_ ;
  assign \new_[142]_  = \new_[6580]_  & \new_[6569]_ ;
  assign \new_[143]_  = \new_[6560]_  & \new_[6549]_ ;
  assign \new_[144]_  = \new_[6540]_  & \new_[6529]_ ;
  assign \new_[145]_  = \new_[6520]_  & \new_[6509]_ ;
  assign \new_[146]_  = \new_[6500]_  & \new_[6489]_ ;
  assign \new_[147]_  = \new_[6480]_  & \new_[6469]_ ;
  assign \new_[148]_  = \new_[6460]_  & \new_[6449]_ ;
  assign \new_[149]_  = \new_[6440]_  & \new_[6429]_ ;
  assign \new_[150]_  = \new_[6420]_  & \new_[6409]_ ;
  assign \new_[151]_  = \new_[6400]_  & \new_[6389]_ ;
  assign \new_[152]_  = \new_[6380]_  & \new_[6369]_ ;
  assign \new_[153]_  = \new_[6360]_  & \new_[6349]_ ;
  assign \new_[154]_  = \new_[6340]_  & \new_[6329]_ ;
  assign \new_[155]_  = \new_[6320]_  & \new_[6309]_ ;
  assign \new_[156]_  = \new_[6300]_  & \new_[6289]_ ;
  assign \new_[157]_  = \new_[6280]_  & \new_[6269]_ ;
  assign \new_[158]_  = \new_[6260]_  & \new_[6249]_ ;
  assign \new_[159]_  = \new_[6240]_  & \new_[6229]_ ;
  assign \new_[160]_  = \new_[6220]_  & \new_[6209]_ ;
  assign \new_[161]_  = \new_[6200]_  & \new_[6189]_ ;
  assign \new_[162]_  = \new_[6180]_  & \new_[6169]_ ;
  assign \new_[163]_  = \new_[6160]_  & \new_[6149]_ ;
  assign \new_[164]_  = \new_[6140]_  & \new_[6129]_ ;
  assign \new_[165]_  = \new_[6120]_  & \new_[6109]_ ;
  assign \new_[166]_  = \new_[6100]_  & \new_[6089]_ ;
  assign \new_[167]_  = \new_[6080]_  & \new_[6069]_ ;
  assign \new_[168]_  = \new_[6060]_  & \new_[6049]_ ;
  assign \new_[169]_  = \new_[6040]_  & \new_[6029]_ ;
  assign \new_[170]_  = \new_[6020]_  & \new_[6009]_ ;
  assign \new_[171]_  = \new_[6000]_  & \new_[5989]_ ;
  assign \new_[172]_  = \new_[5980]_  & \new_[5969]_ ;
  assign \new_[173]_  = \new_[5960]_  & \new_[5949]_ ;
  assign \new_[174]_  = \new_[5940]_  & \new_[5929]_ ;
  assign \new_[175]_  = \new_[5920]_  & \new_[5909]_ ;
  assign \new_[176]_  = \new_[5900]_  & \new_[5889]_ ;
  assign \new_[177]_  = \new_[5880]_  & \new_[5869]_ ;
  assign \new_[178]_  = \new_[5860]_  & \new_[5849]_ ;
  assign \new_[179]_  = \new_[5840]_  & \new_[5829]_ ;
  assign \new_[180]_  = \new_[5820]_  & \new_[5809]_ ;
  assign \new_[181]_  = \new_[5800]_  & \new_[5789]_ ;
  assign \new_[182]_  = \new_[5780]_  & \new_[5769]_ ;
  assign \new_[183]_  = \new_[5760]_  & \new_[5749]_ ;
  assign \new_[184]_  = \new_[5740]_  & \new_[5729]_ ;
  assign \new_[185]_  = \new_[5720]_  & \new_[5709]_ ;
  assign \new_[186]_  = \new_[5700]_  & \new_[5689]_ ;
  assign \new_[187]_  = \new_[5680]_  & \new_[5669]_ ;
  assign \new_[188]_  = \new_[5660]_  & \new_[5649]_ ;
  assign \new_[189]_  = \new_[5640]_  & \new_[5629]_ ;
  assign \new_[190]_  = \new_[5620]_  & \new_[5609]_ ;
  assign \new_[191]_  = \new_[5600]_  & \new_[5589]_ ;
  assign \new_[192]_  = \new_[5580]_  & \new_[5569]_ ;
  assign \new_[193]_  = \new_[5560]_  & \new_[5549]_ ;
  assign \new_[194]_  = \new_[5540]_  & \new_[5529]_ ;
  assign \new_[195]_  = \new_[5520]_  & \new_[5509]_ ;
  assign \new_[196]_  = \new_[5500]_  & \new_[5489]_ ;
  assign \new_[197]_  = \new_[5480]_  & \new_[5469]_ ;
  assign \new_[198]_  = \new_[5460]_  & \new_[5449]_ ;
  assign \new_[199]_  = \new_[5440]_  & \new_[5429]_ ;
  assign \new_[200]_  = \new_[5420]_  & \new_[5409]_ ;
  assign \new_[201]_  = \new_[5400]_  & \new_[5389]_ ;
  assign \new_[202]_  = \new_[5380]_  & \new_[5369]_ ;
  assign \new_[203]_  = \new_[5360]_  & \new_[5349]_ ;
  assign \new_[204]_  = \new_[5340]_  & \new_[5329]_ ;
  assign \new_[205]_  = \new_[5320]_  & \new_[5309]_ ;
  assign \new_[206]_  = \new_[5300]_  & \new_[5289]_ ;
  assign \new_[207]_  = \new_[5280]_  & \new_[5269]_ ;
  assign \new_[208]_  = \new_[5260]_  & \new_[5249]_ ;
  assign \new_[209]_  = \new_[5240]_  & \new_[5229]_ ;
  assign \new_[210]_  = \new_[5220]_  & \new_[5209]_ ;
  assign \new_[211]_  = \new_[5200]_  & \new_[5189]_ ;
  assign \new_[212]_  = \new_[5180]_  & \new_[5169]_ ;
  assign \new_[213]_  = \new_[5160]_  & \new_[5149]_ ;
  assign \new_[214]_  = \new_[5140]_  & \new_[5129]_ ;
  assign \new_[215]_  = \new_[5120]_  & \new_[5109]_ ;
  assign \new_[216]_  = \new_[5100]_  & \new_[5089]_ ;
  assign \new_[217]_  = \new_[5080]_  & \new_[5069]_ ;
  assign \new_[218]_  = \new_[5060]_  & \new_[5049]_ ;
  assign \new_[219]_  = \new_[5040]_  & \new_[5029]_ ;
  assign \new_[220]_  = \new_[5020]_  & \new_[5009]_ ;
  assign \new_[221]_  = \new_[5000]_  & \new_[4989]_ ;
  assign \new_[222]_  = \new_[4980]_  & \new_[4969]_ ;
  assign \new_[223]_  = \new_[4960]_  & \new_[4949]_ ;
  assign \new_[224]_  = \new_[4940]_  & \new_[4929]_ ;
  assign \new_[225]_  = \new_[4920]_  & \new_[4909]_ ;
  assign \new_[226]_  = \new_[4900]_  & \new_[4889]_ ;
  assign \new_[227]_  = \new_[4880]_  & \new_[4869]_ ;
  assign \new_[228]_  = \new_[4860]_  & \new_[4849]_ ;
  assign \new_[229]_  = \new_[4840]_  & \new_[4829]_ ;
  assign \new_[230]_  = \new_[4820]_  & \new_[4809]_ ;
  assign \new_[231]_  = \new_[4800]_  & \new_[4789]_ ;
  assign \new_[232]_  = \new_[4780]_  & \new_[4769]_ ;
  assign \new_[233]_  = \new_[4760]_  & \new_[4751]_ ;
  assign \new_[234]_  = \new_[4742]_  & \new_[4733]_ ;
  assign \new_[235]_  = \new_[4724]_  & \new_[4715]_ ;
  assign \new_[236]_  = \new_[4706]_  & \new_[4697]_ ;
  assign \new_[237]_  = \new_[4688]_  & \new_[4679]_ ;
  assign \new_[238]_  = \new_[4670]_  & \new_[4661]_ ;
  assign \new_[239]_  = \new_[4652]_  & \new_[4643]_ ;
  assign \new_[240]_  = \new_[4634]_  & \new_[4625]_ ;
  assign \new_[241]_  = \new_[4616]_  & \new_[4607]_ ;
  assign \new_[242]_  = \new_[4598]_  & \new_[4589]_ ;
  assign \new_[243]_  = \new_[4580]_  & \new_[4571]_ ;
  assign \new_[244]_  = \new_[4562]_  & \new_[4553]_ ;
  assign \new_[245]_  = \new_[4544]_  & \new_[4535]_ ;
  assign \new_[246]_  = \new_[4526]_  & \new_[4517]_ ;
  assign \new_[247]_  = \new_[4508]_  & \new_[4499]_ ;
  assign \new_[248]_  = \new_[4490]_  & \new_[4481]_ ;
  assign \new_[249]_  = \new_[4472]_  & \new_[4463]_ ;
  assign \new_[250]_  = \new_[4454]_  & \new_[4445]_ ;
  assign \new_[251]_  = \new_[4436]_  & \new_[4427]_ ;
  assign \new_[252]_  = \new_[4418]_  & \new_[4409]_ ;
  assign \new_[253]_  = \new_[4400]_  & \new_[4391]_ ;
  assign \new_[254]_  = \new_[4382]_  & \new_[4373]_ ;
  assign \new_[255]_  = \new_[4364]_  & \new_[4355]_ ;
  assign \new_[256]_  = \new_[4346]_  & \new_[4337]_ ;
  assign \new_[257]_  = \new_[4328]_  & \new_[4319]_ ;
  assign \new_[258]_  = \new_[4310]_  & \new_[4301]_ ;
  assign \new_[259]_  = \new_[4292]_  & \new_[4283]_ ;
  assign \new_[260]_  = \new_[4274]_  & \new_[4265]_ ;
  assign \new_[261]_  = \new_[4256]_  & \new_[4247]_ ;
  assign \new_[262]_  = \new_[4238]_  & \new_[4229]_ ;
  assign \new_[263]_  = \new_[4220]_  & \new_[4211]_ ;
  assign \new_[264]_  = \new_[4202]_  & \new_[4193]_ ;
  assign \new_[265]_  = \new_[4184]_  & \new_[4175]_ ;
  assign \new_[266]_  = \new_[4166]_  & \new_[4157]_ ;
  assign \new_[267]_  = \new_[4148]_  & \new_[4139]_ ;
  assign \new_[268]_  = \new_[4130]_  & \new_[4121]_ ;
  assign \new_[269]_  = \new_[4112]_  & \new_[4103]_ ;
  assign \new_[270]_  = \new_[4094]_  & \new_[4085]_ ;
  assign \new_[271]_  = \new_[4076]_  & \new_[4067]_ ;
  assign \new_[272]_  = \new_[4058]_  & \new_[4049]_ ;
  assign \new_[273]_  = \new_[4040]_  & \new_[4031]_ ;
  assign \new_[274]_  = \new_[4022]_  & \new_[4013]_ ;
  assign \new_[275]_  = \new_[4004]_  & \new_[3995]_ ;
  assign \new_[276]_  = \new_[3986]_  & \new_[3977]_ ;
  assign \new_[277]_  = \new_[3968]_  & \new_[3959]_ ;
  assign \new_[278]_  = \new_[3950]_  & \new_[3941]_ ;
  assign \new_[279]_  = \new_[3932]_  & \new_[3923]_ ;
  assign \new_[280]_  = \new_[3914]_  & \new_[3905]_ ;
  assign \new_[281]_  = \new_[3896]_  & \new_[3887]_ ;
  assign \new_[282]_  = \new_[3878]_  & \new_[3869]_ ;
  assign \new_[283]_  = \new_[3860]_  & \new_[3851]_ ;
  assign \new_[284]_  = \new_[3842]_  & \new_[3833]_ ;
  assign \new_[285]_  = \new_[3824]_  & \new_[3815]_ ;
  assign \new_[286]_  = \new_[3806]_  & \new_[3797]_ ;
  assign \new_[287]_  = \new_[3788]_  & \new_[3779]_ ;
  assign \new_[288]_  = \new_[3770]_  & \new_[3761]_ ;
  assign \new_[289]_  = \new_[3752]_  & \new_[3743]_ ;
  assign \new_[290]_  = \new_[3734]_  & \new_[3725]_ ;
  assign \new_[291]_  = \new_[3716]_  & \new_[3707]_ ;
  assign \new_[292]_  = \new_[3698]_  & \new_[3689]_ ;
  assign \new_[293]_  = \new_[3680]_  & \new_[3671]_ ;
  assign \new_[294]_  = \new_[3662]_  & \new_[3653]_ ;
  assign \new_[295]_  = \new_[3644]_  & \new_[3635]_ ;
  assign \new_[296]_  = \new_[3626]_  & \new_[3617]_ ;
  assign \new_[297]_  = \new_[3608]_  & \new_[3599]_ ;
  assign \new_[298]_  = \new_[3590]_  & \new_[3581]_ ;
  assign \new_[299]_  = \new_[3572]_  & \new_[3563]_ ;
  assign \new_[300]_  = \new_[3554]_  & \new_[3545]_ ;
  assign \new_[301]_  = \new_[3536]_  & \new_[3527]_ ;
  assign \new_[302]_  = \new_[3518]_  & \new_[3509]_ ;
  assign \new_[303]_  = \new_[3500]_  & \new_[3491]_ ;
  assign \new_[304]_  = \new_[3482]_  & \new_[3473]_ ;
  assign \new_[305]_  = \new_[3464]_  & \new_[3455]_ ;
  assign \new_[306]_  = \new_[3446]_  & \new_[3437]_ ;
  assign \new_[307]_  = \new_[3428]_  & \new_[3419]_ ;
  assign \new_[308]_  = \new_[3410]_  & \new_[3401]_ ;
  assign \new_[309]_  = \new_[3392]_  & \new_[3383]_ ;
  assign \new_[310]_  = \new_[3374]_  & \new_[3365]_ ;
  assign \new_[311]_  = \new_[3356]_  & \new_[3347]_ ;
  assign \new_[312]_  = \new_[3338]_  & \new_[3329]_ ;
  assign \new_[313]_  = \new_[3320]_  & \new_[3311]_ ;
  assign \new_[314]_  = \new_[3302]_  & \new_[3293]_ ;
  assign \new_[315]_  = \new_[3284]_  & \new_[3275]_ ;
  assign \new_[316]_  = \new_[3266]_  & \new_[3257]_ ;
  assign \new_[317]_  = \new_[3248]_  & \new_[3239]_ ;
  assign \new_[318]_  = \new_[3230]_  & \new_[3221]_ ;
  assign \new_[319]_  = \new_[3212]_  & \new_[3203]_ ;
  assign \new_[320]_  = \new_[3194]_  & \new_[3185]_ ;
  assign \new_[321]_  = \new_[3176]_  & \new_[3167]_ ;
  assign \new_[322]_  = \new_[3158]_  & \new_[3149]_ ;
  assign \new_[323]_  = \new_[3140]_  & \new_[3131]_ ;
  assign \new_[324]_  = \new_[3122]_  & \new_[3113]_ ;
  assign \new_[325]_  = \new_[3104]_  & \new_[3095]_ ;
  assign \new_[326]_  = \new_[3086]_  & \new_[3077]_ ;
  assign \new_[327]_  = \new_[3068]_  & \new_[3059]_ ;
  assign \new_[328]_  = \new_[3050]_  & \new_[3041]_ ;
  assign \new_[329]_  = \new_[3032]_  & \new_[3023]_ ;
  assign \new_[330]_  = \new_[3014]_  & \new_[3005]_ ;
  assign \new_[331]_  = \new_[2996]_  & \new_[2987]_ ;
  assign \new_[332]_  = \new_[2978]_  & \new_[2969]_ ;
  assign \new_[333]_  = \new_[2960]_  & \new_[2951]_ ;
  assign \new_[334]_  = \new_[2942]_  & \new_[2933]_ ;
  assign \new_[335]_  = \new_[2924]_  & \new_[2915]_ ;
  assign \new_[336]_  = \new_[2906]_  & \new_[2897]_ ;
  assign \new_[337]_  = \new_[2888]_  & \new_[2879]_ ;
  assign \new_[338]_  = \new_[2870]_  & \new_[2861]_ ;
  assign \new_[339]_  = \new_[2852]_  & \new_[2843]_ ;
  assign \new_[340]_  = \new_[2834]_  & \new_[2825]_ ;
  assign \new_[341]_  = \new_[2816]_  & \new_[2807]_ ;
  assign \new_[342]_  = \new_[2798]_  & \new_[2789]_ ;
  assign \new_[343]_  = \new_[2780]_  & \new_[2771]_ ;
  assign \new_[344]_  = \new_[2762]_  & \new_[2753]_ ;
  assign \new_[345]_  = \new_[2744]_  & \new_[2735]_ ;
  assign \new_[346]_  = \new_[2726]_  & \new_[2717]_ ;
  assign \new_[347]_  = \new_[2708]_  & \new_[2699]_ ;
  assign \new_[348]_  = \new_[2690]_  & \new_[2681]_ ;
  assign \new_[349]_  = \new_[2672]_  & \new_[2663]_ ;
  assign \new_[350]_  = \new_[2654]_  & \new_[2645]_ ;
  assign \new_[351]_  = \new_[2636]_  & \new_[2627]_ ;
  assign \new_[352]_  = \new_[2618]_  & \new_[2609]_ ;
  assign \new_[353]_  = \new_[2600]_  & \new_[2591]_ ;
  assign \new_[354]_  = \new_[2582]_  & \new_[2573]_ ;
  assign \new_[355]_  = \new_[2564]_  & \new_[2555]_ ;
  assign \new_[356]_  = \new_[2546]_  & \new_[2537]_ ;
  assign \new_[357]_  = \new_[2528]_  & \new_[2519]_ ;
  assign \new_[358]_  = \new_[2510]_  & \new_[2501]_ ;
  assign \new_[359]_  = \new_[2492]_  & \new_[2483]_ ;
  assign \new_[360]_  = \new_[2474]_  & \new_[2465]_ ;
  assign \new_[361]_  = \new_[2456]_  & \new_[2447]_ ;
  assign \new_[362]_  = \new_[2438]_  & \new_[2429]_ ;
  assign \new_[363]_  = \new_[2420]_  & \new_[2411]_ ;
  assign \new_[364]_  = \new_[2402]_  & \new_[2393]_ ;
  assign \new_[365]_  = \new_[2384]_  & \new_[2375]_ ;
  assign \new_[366]_  = \new_[2366]_  & \new_[2357]_ ;
  assign \new_[367]_  = \new_[2348]_  & \new_[2339]_ ;
  assign \new_[368]_  = \new_[2330]_  & \new_[2321]_ ;
  assign \new_[369]_  = \new_[2312]_  & \new_[2303]_ ;
  assign \new_[370]_  = \new_[2296]_  & \new_[2287]_ ;
  assign \new_[371]_  = \new_[2280]_  & \new_[2271]_ ;
  assign \new_[372]_  = \new_[2264]_  & \new_[2255]_ ;
  assign \new_[373]_  = \new_[2248]_  & \new_[2239]_ ;
  assign \new_[374]_  = \new_[2232]_  & \new_[2223]_ ;
  assign \new_[375]_  = \new_[2216]_  & \new_[2207]_ ;
  assign \new_[376]_  = \new_[2200]_  & \new_[2191]_ ;
  assign \new_[377]_  = \new_[2184]_  & \new_[2175]_ ;
  assign \new_[378]_  = \new_[2168]_  & \new_[2159]_ ;
  assign \new_[379]_  = \new_[2152]_  & \new_[2143]_ ;
  assign \new_[380]_  = \new_[2136]_  & \new_[2127]_ ;
  assign \new_[381]_  = \new_[2120]_  & \new_[2111]_ ;
  assign \new_[382]_  = \new_[2104]_  & \new_[2095]_ ;
  assign \new_[383]_  = \new_[2088]_  & \new_[2079]_ ;
  assign \new_[384]_  = \new_[2072]_  & \new_[2063]_ ;
  assign \new_[385]_  = \new_[2056]_  & \new_[2047]_ ;
  assign \new_[386]_  = \new_[2040]_  & \new_[2031]_ ;
  assign \new_[387]_  = \new_[2024]_  & \new_[2015]_ ;
  assign \new_[388]_  = \new_[2008]_  & \new_[1999]_ ;
  assign \new_[389]_  = \new_[1992]_  & \new_[1983]_ ;
  assign \new_[390]_  = \new_[1976]_  & \new_[1967]_ ;
  assign \new_[391]_  = \new_[1960]_  & \new_[1951]_ ;
  assign \new_[392]_  = \new_[1944]_  & \new_[1935]_ ;
  assign \new_[393]_  = \new_[1928]_  & \new_[1919]_ ;
  assign \new_[394]_  = \new_[1912]_  & \new_[1903]_ ;
  assign \new_[395]_  = \new_[1896]_  & \new_[1887]_ ;
  assign \new_[396]_  = \new_[1880]_  & \new_[1871]_ ;
  assign \new_[397]_  = \new_[1864]_  & \new_[1855]_ ;
  assign \new_[398]_  = \new_[1848]_  & \new_[1839]_ ;
  assign \new_[399]_  = \new_[1832]_  & \new_[1823]_ ;
  assign \new_[400]_  = \new_[1816]_  & \new_[1807]_ ;
  assign \new_[401]_  = \new_[1800]_  & \new_[1793]_ ;
  assign \new_[402]_  = \new_[1786]_  & \new_[1779]_ ;
  assign \new_[403]_  = \new_[1772]_  & \new_[1765]_ ;
  assign \new_[404]_  = \new_[1758]_  & \new_[1751]_ ;
  assign \new_[405]_  = \new_[1744]_  & \new_[1737]_ ;
  assign \new_[406]_  = \new_[1730]_  & \new_[1723]_ ;
  assign \new_[407]_  = \new_[1716]_  & \new_[1709]_ ;
  assign \new_[408]_  = \new_[1702]_  & \new_[1695]_ ;
  assign \new_[409]_  = \new_[1688]_  & \new_[1681]_ ;
  assign \new_[410]_  = \new_[1674]_  & \new_[1667]_ ;
  assign \new_[411]_  = \new_[1660]_  & \new_[1653]_ ;
  assign \new_[412]_  = \new_[1646]_  & \new_[1639]_ ;
  assign \new_[413]_  = \new_[1632]_  & \new_[1625]_ ;
  assign \new_[414]_  = \new_[1618]_  & \new_[1611]_ ;
  assign \new_[415]_  = \new_[1604]_  & \new_[1597]_ ;
  assign \new_[416]_  = \new_[1590]_  & \new_[1583]_ ;
  assign \new_[417]_  = \new_[1576]_  & \new_[1569]_ ;
  assign \new_[418]_  = \new_[1562]_  & \new_[1555]_ ;
  assign \new_[419]_  = \new_[1548]_  & \new_[1541]_ ;
  assign \new_[420]_  = \new_[1534]_  & \new_[1527]_ ;
  assign \new_[421]_  = \new_[1520]_  & \new_[1513]_ ;
  assign \new_[422]_  = \new_[1506]_  & \new_[1499]_ ;
  assign \new_[423]_  = \new_[1492]_  & \new_[1485]_ ;
  assign \new_[424]_  = \new_[1478]_  & \new_[1471]_ ;
  assign \new_[425]_  = \new_[1464]_  & \new_[1457]_ ;
  assign \new_[426]_  = \new_[1450]_  & \new_[1443]_ ;
  assign \new_[427]_  = \new_[1436]_  & \new_[1429]_ ;
  assign \new_[428]_  = \new_[1422]_  & \new_[1415]_ ;
  assign \new_[429]_  = \new_[1408]_  & \new_[1401]_ ;
  assign \new_[430]_  = \new_[1394]_  & \new_[1387]_ ;
  assign \new_[431]_  = \new_[1380]_  & \new_[1373]_ ;
  assign \new_[432]_  = \new_[1366]_  & \new_[1359]_ ;
  assign \new_[433]_  = \new_[1352]_  & \new_[1347]_ ;
  assign \new_[434]_  = \new_[1344]_  & \new_[1339]_ ;
  assign \new_[435]_  = \new_[1336]_  & \new_[1333]_ ;
  assign \new_[436]_  = \new_[1330]_  & \new_[1327]_ ;
  assign \new_[437]_  = \new_[1324]_  & \new_[1321]_ ;
  assign \new_[438]_  = \new_[1318]_  & \new_[1315]_ ;
  assign \new_[442]_  = \new_[436]_  | \new_[437]_ ;
  assign \new_[443]_  = \new_[438]_  | \new_[442]_ ;
  assign \new_[447]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[448]_  = \new_[435]_  | \new_[447]_ ;
  assign \new_[449]_  = \new_[448]_  | \new_[443]_ ;
  assign \new_[453]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[454]_  = \new_[432]_  | \new_[453]_ ;
  assign \new_[457]_  = \new_[428]_  | \new_[429]_ ;
  assign \new_[460]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[461]_  = \new_[460]_  | \new_[457]_ ;
  assign \new_[462]_  = \new_[461]_  | \new_[454]_ ;
  assign \new_[463]_  = \new_[462]_  | \new_[449]_ ;
  assign \new_[467]_  = \new_[423]_  | \new_[424]_ ;
  assign \new_[468]_  = \new_[425]_  | \new_[467]_ ;
  assign \new_[471]_  = \new_[421]_  | \new_[422]_ ;
  assign \new_[474]_  = \new_[419]_  | \new_[420]_ ;
  assign \new_[475]_  = \new_[474]_  | \new_[471]_ ;
  assign \new_[476]_  = \new_[475]_  | \new_[468]_ ;
  assign \new_[480]_  = \new_[416]_  | \new_[417]_ ;
  assign \new_[481]_  = \new_[418]_  | \new_[480]_ ;
  assign \new_[484]_  = \new_[414]_  | \new_[415]_ ;
  assign \new_[487]_  = \new_[412]_  | \new_[413]_ ;
  assign \new_[488]_  = \new_[487]_  | \new_[484]_ ;
  assign \new_[489]_  = \new_[488]_  | \new_[481]_ ;
  assign \new_[490]_  = \new_[489]_  | \new_[476]_ ;
  assign \new_[491]_  = \new_[490]_  | \new_[463]_ ;
  assign \new_[495]_  = \new_[409]_  | \new_[410]_ ;
  assign \new_[496]_  = \new_[411]_  | \new_[495]_ ;
  assign \new_[500]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[501]_  = \new_[408]_  | \new_[500]_ ;
  assign \new_[502]_  = \new_[501]_  | \new_[496]_ ;
  assign \new_[506]_  = \new_[403]_  | \new_[404]_ ;
  assign \new_[507]_  = \new_[405]_  | \new_[506]_ ;
  assign \new_[510]_  = \new_[401]_  | \new_[402]_ ;
  assign \new_[513]_  = \new_[399]_  | \new_[400]_ ;
  assign \new_[514]_  = \new_[513]_  | \new_[510]_ ;
  assign \new_[515]_  = \new_[514]_  | \new_[507]_ ;
  assign \new_[516]_  = \new_[515]_  | \new_[502]_ ;
  assign \new_[520]_  = \new_[396]_  | \new_[397]_ ;
  assign \new_[521]_  = \new_[398]_  | \new_[520]_ ;
  assign \new_[524]_  = \new_[394]_  | \new_[395]_ ;
  assign \new_[527]_  = \new_[392]_  | \new_[393]_ ;
  assign \new_[528]_  = \new_[527]_  | \new_[524]_ ;
  assign \new_[529]_  = \new_[528]_  | \new_[521]_ ;
  assign \new_[533]_  = \new_[389]_  | \new_[390]_ ;
  assign \new_[534]_  = \new_[391]_  | \new_[533]_ ;
  assign \new_[537]_  = \new_[387]_  | \new_[388]_ ;
  assign \new_[540]_  = \new_[385]_  | \new_[386]_ ;
  assign \new_[541]_  = \new_[540]_  | \new_[537]_ ;
  assign \new_[542]_  = \new_[541]_  | \new_[534]_ ;
  assign \new_[543]_  = \new_[542]_  | \new_[529]_ ;
  assign \new_[544]_  = \new_[543]_  | \new_[516]_ ;
  assign \new_[545]_  = \new_[544]_  | \new_[491]_ ;
  assign \new_[549]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[550]_  = \new_[384]_  | \new_[549]_ ;
  assign \new_[554]_  = \new_[379]_  | \new_[380]_ ;
  assign \new_[555]_  = \new_[381]_  | \new_[554]_ ;
  assign \new_[556]_  = \new_[555]_  | \new_[550]_ ;
  assign \new_[560]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[561]_  = \new_[378]_  | \new_[560]_ ;
  assign \new_[564]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[567]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[568]_  = \new_[567]_  | \new_[564]_ ;
  assign \new_[569]_  = \new_[568]_  | \new_[561]_ ;
  assign \new_[570]_  = \new_[569]_  | \new_[556]_ ;
  assign \new_[574]_  = \new_[369]_  | \new_[370]_ ;
  assign \new_[575]_  = \new_[371]_  | \new_[574]_ ;
  assign \new_[578]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[581]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[582]_  = \new_[581]_  | \new_[578]_ ;
  assign \new_[583]_  = \new_[582]_  | \new_[575]_ ;
  assign \new_[587]_  = \new_[362]_  | \new_[363]_ ;
  assign \new_[588]_  = \new_[364]_  | \new_[587]_ ;
  assign \new_[591]_  = \new_[360]_  | \new_[361]_ ;
  assign \new_[594]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[595]_  = \new_[594]_  | \new_[591]_ ;
  assign \new_[596]_  = \new_[595]_  | \new_[588]_ ;
  assign \new_[597]_  = \new_[596]_  | \new_[583]_ ;
  assign \new_[598]_  = \new_[597]_  | \new_[570]_ ;
  assign \new_[602]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[603]_  = \new_[357]_  | \new_[602]_ ;
  assign \new_[606]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[609]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[610]_  = \new_[609]_  | \new_[606]_ ;
  assign \new_[611]_  = \new_[610]_  | \new_[603]_ ;
  assign \new_[615]_  = \new_[348]_  | \new_[349]_ ;
  assign \new_[616]_  = \new_[350]_  | \new_[615]_ ;
  assign \new_[619]_  = \new_[346]_  | \new_[347]_ ;
  assign \new_[622]_  = \new_[344]_  | \new_[345]_ ;
  assign \new_[623]_  = \new_[622]_  | \new_[619]_ ;
  assign \new_[624]_  = \new_[623]_  | \new_[616]_ ;
  assign \new_[625]_  = \new_[624]_  | \new_[611]_ ;
  assign \new_[629]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[630]_  = \new_[343]_  | \new_[629]_ ;
  assign \new_[633]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[636]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[637]_  = \new_[636]_  | \new_[633]_ ;
  assign \new_[638]_  = \new_[637]_  | \new_[630]_ ;
  assign \new_[642]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[643]_  = \new_[336]_  | \new_[642]_ ;
  assign \new_[646]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[649]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[650]_  = \new_[649]_  | \new_[646]_ ;
  assign \new_[651]_  = \new_[650]_  | \new_[643]_ ;
  assign \new_[652]_  = \new_[651]_  | \new_[638]_ ;
  assign \new_[653]_  = \new_[652]_  | \new_[625]_ ;
  assign \new_[654]_  = \new_[653]_  | \new_[598]_ ;
  assign \new_[655]_  = \new_[654]_  | \new_[545]_ ;
  assign \new_[659]_  = \new_[327]_  | \new_[328]_ ;
  assign \new_[660]_  = \new_[329]_  | \new_[659]_ ;
  assign \new_[664]_  = \new_[324]_  | \new_[325]_ ;
  assign \new_[665]_  = \new_[326]_  | \new_[664]_ ;
  assign \new_[666]_  = \new_[665]_  | \new_[660]_ ;
  assign \new_[670]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[671]_  = \new_[323]_  | \new_[670]_ ;
  assign \new_[674]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[677]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[678]_  = \new_[677]_  | \new_[674]_ ;
  assign \new_[679]_  = \new_[678]_  | \new_[671]_ ;
  assign \new_[680]_  = \new_[679]_  | \new_[666]_ ;
  assign \new_[684]_  = \new_[314]_  | \new_[315]_ ;
  assign \new_[685]_  = \new_[316]_  | \new_[684]_ ;
  assign \new_[688]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[691]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[692]_  = \new_[691]_  | \new_[688]_ ;
  assign \new_[693]_  = \new_[692]_  | \new_[685]_ ;
  assign \new_[697]_  = \new_[307]_  | \new_[308]_ ;
  assign \new_[698]_  = \new_[309]_  | \new_[697]_ ;
  assign \new_[701]_  = \new_[305]_  | \new_[306]_ ;
  assign \new_[704]_  = \new_[303]_  | \new_[304]_ ;
  assign \new_[705]_  = \new_[704]_  | \new_[701]_ ;
  assign \new_[706]_  = \new_[705]_  | \new_[698]_ ;
  assign \new_[707]_  = \new_[706]_  | \new_[693]_ ;
  assign \new_[708]_  = \new_[707]_  | \new_[680]_ ;
  assign \new_[712]_  = \new_[300]_  | \new_[301]_ ;
  assign \new_[713]_  = \new_[302]_  | \new_[712]_ ;
  assign \new_[716]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[719]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[720]_  = \new_[719]_  | \new_[716]_ ;
  assign \new_[721]_  = \new_[720]_  | \new_[713]_ ;
  assign \new_[725]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[726]_  = \new_[295]_  | \new_[725]_ ;
  assign \new_[729]_  = \new_[291]_  | \new_[292]_ ;
  assign \new_[732]_  = \new_[289]_  | \new_[290]_ ;
  assign \new_[733]_  = \new_[732]_  | \new_[729]_ ;
  assign \new_[734]_  = \new_[733]_  | \new_[726]_ ;
  assign \new_[735]_  = \new_[734]_  | \new_[721]_ ;
  assign \new_[739]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[740]_  = \new_[288]_  | \new_[739]_ ;
  assign \new_[743]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[746]_  = \new_[282]_  | \new_[283]_ ;
  assign \new_[747]_  = \new_[746]_  | \new_[743]_ ;
  assign \new_[748]_  = \new_[747]_  | \new_[740]_ ;
  assign \new_[752]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[753]_  = \new_[281]_  | \new_[752]_ ;
  assign \new_[756]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[759]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[760]_  = \new_[759]_  | \new_[756]_ ;
  assign \new_[761]_  = \new_[760]_  | \new_[753]_ ;
  assign \new_[762]_  = \new_[761]_  | \new_[748]_ ;
  assign \new_[763]_  = \new_[762]_  | \new_[735]_ ;
  assign \new_[764]_  = \new_[763]_  | \new_[708]_ ;
  assign \new_[768]_  = \new_[272]_  | \new_[273]_ ;
  assign \new_[769]_  = \new_[274]_  | \new_[768]_ ;
  assign \new_[773]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[774]_  = \new_[271]_  | \new_[773]_ ;
  assign \new_[775]_  = \new_[774]_  | \new_[769]_ ;
  assign \new_[779]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[780]_  = \new_[268]_  | \new_[779]_ ;
  assign \new_[783]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[786]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[787]_  = \new_[786]_  | \new_[783]_ ;
  assign \new_[788]_  = \new_[787]_  | \new_[780]_ ;
  assign \new_[789]_  = \new_[788]_  | \new_[775]_ ;
  assign \new_[793]_  = \new_[259]_  | \new_[260]_ ;
  assign \new_[794]_  = \new_[261]_  | \new_[793]_ ;
  assign \new_[797]_  = \new_[257]_  | \new_[258]_ ;
  assign \new_[800]_  = \new_[255]_  | \new_[256]_ ;
  assign \new_[801]_  = \new_[800]_  | \new_[797]_ ;
  assign \new_[802]_  = \new_[801]_  | \new_[794]_ ;
  assign \new_[806]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[807]_  = \new_[254]_  | \new_[806]_ ;
  assign \new_[810]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[813]_  = \new_[248]_  | \new_[249]_ ;
  assign \new_[814]_  = \new_[813]_  | \new_[810]_ ;
  assign \new_[815]_  = \new_[814]_  | \new_[807]_ ;
  assign \new_[816]_  = \new_[815]_  | \new_[802]_ ;
  assign \new_[817]_  = \new_[816]_  | \new_[789]_ ;
  assign \new_[821]_  = \new_[245]_  | \new_[246]_ ;
  assign \new_[822]_  = \new_[247]_  | \new_[821]_ ;
  assign \new_[825]_  = \new_[243]_  | \new_[244]_ ;
  assign \new_[828]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[829]_  = \new_[828]_  | \new_[825]_ ;
  assign \new_[830]_  = \new_[829]_  | \new_[822]_ ;
  assign \new_[834]_  = \new_[238]_  | \new_[239]_ ;
  assign \new_[835]_  = \new_[240]_  | \new_[834]_ ;
  assign \new_[838]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[841]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[842]_  = \new_[841]_  | \new_[838]_ ;
  assign \new_[843]_  = \new_[842]_  | \new_[835]_ ;
  assign \new_[844]_  = \new_[843]_  | \new_[830]_ ;
  assign \new_[848]_  = \new_[231]_  | \new_[232]_ ;
  assign \new_[849]_  = \new_[233]_  | \new_[848]_ ;
  assign \new_[852]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[855]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[856]_  = \new_[855]_  | \new_[852]_ ;
  assign \new_[857]_  = \new_[856]_  | \new_[849]_ ;
  assign \new_[861]_  = \new_[224]_  | \new_[225]_ ;
  assign \new_[862]_  = \new_[226]_  | \new_[861]_ ;
  assign \new_[865]_  = \new_[222]_  | \new_[223]_ ;
  assign \new_[868]_  = \new_[220]_  | \new_[221]_ ;
  assign \new_[869]_  = \new_[868]_  | \new_[865]_ ;
  assign \new_[870]_  = \new_[869]_  | \new_[862]_ ;
  assign \new_[871]_  = \new_[870]_  | \new_[857]_ ;
  assign \new_[872]_  = \new_[871]_  | \new_[844]_ ;
  assign \new_[873]_  = \new_[872]_  | \new_[817]_ ;
  assign \new_[874]_  = \new_[873]_  | \new_[764]_ ;
  assign \new_[875]_  = \new_[874]_  | \new_[655]_ ;
  assign \new_[879]_  = \new_[217]_  | \new_[218]_ ;
  assign \new_[880]_  = \new_[219]_  | \new_[879]_ ;
  assign \new_[884]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[885]_  = \new_[216]_  | \new_[884]_ ;
  assign \new_[886]_  = \new_[885]_  | \new_[880]_ ;
  assign \new_[890]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[891]_  = \new_[213]_  | \new_[890]_ ;
  assign \new_[894]_  = \new_[209]_  | \new_[210]_ ;
  assign \new_[897]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[898]_  = \new_[897]_  | \new_[894]_ ;
  assign \new_[899]_  = \new_[898]_  | \new_[891]_ ;
  assign \new_[900]_  = \new_[899]_  | \new_[886]_ ;
  assign \new_[904]_  = \new_[204]_  | \new_[205]_ ;
  assign \new_[905]_  = \new_[206]_  | \new_[904]_ ;
  assign \new_[908]_  = \new_[202]_  | \new_[203]_ ;
  assign \new_[911]_  = \new_[200]_  | \new_[201]_ ;
  assign \new_[912]_  = \new_[911]_  | \new_[908]_ ;
  assign \new_[913]_  = \new_[912]_  | \new_[905]_ ;
  assign \new_[917]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[918]_  = \new_[199]_  | \new_[917]_ ;
  assign \new_[921]_  = \new_[195]_  | \new_[196]_ ;
  assign \new_[924]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[925]_  = \new_[924]_  | \new_[921]_ ;
  assign \new_[926]_  = \new_[925]_  | \new_[918]_ ;
  assign \new_[927]_  = \new_[926]_  | \new_[913]_ ;
  assign \new_[928]_  = \new_[927]_  | \new_[900]_ ;
  assign \new_[932]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[933]_  = \new_[192]_  | \new_[932]_ ;
  assign \new_[937]_  = \new_[187]_  | \new_[188]_ ;
  assign \new_[938]_  = \new_[189]_  | \new_[937]_ ;
  assign \new_[939]_  = \new_[938]_  | \new_[933]_ ;
  assign \new_[943]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[944]_  = \new_[186]_  | \new_[943]_ ;
  assign \new_[947]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[950]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[951]_  = \new_[950]_  | \new_[947]_ ;
  assign \new_[952]_  = \new_[951]_  | \new_[944]_ ;
  assign \new_[953]_  = \new_[952]_  | \new_[939]_ ;
  assign \new_[957]_  = \new_[177]_  | \new_[178]_ ;
  assign \new_[958]_  = \new_[179]_  | \new_[957]_ ;
  assign \new_[961]_  = \new_[175]_  | \new_[176]_ ;
  assign \new_[964]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[965]_  = \new_[964]_  | \new_[961]_ ;
  assign \new_[966]_  = \new_[965]_  | \new_[958]_ ;
  assign \new_[970]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[971]_  = \new_[172]_  | \new_[970]_ ;
  assign \new_[974]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[977]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[978]_  = \new_[977]_  | \new_[974]_ ;
  assign \new_[979]_  = \new_[978]_  | \new_[971]_ ;
  assign \new_[980]_  = \new_[979]_  | \new_[966]_ ;
  assign \new_[981]_  = \new_[980]_  | \new_[953]_ ;
  assign \new_[982]_  = \new_[981]_  | \new_[928]_ ;
  assign \new_[986]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[987]_  = \new_[165]_  | \new_[986]_ ;
  assign \new_[991]_  = \new_[160]_  | \new_[161]_ ;
  assign \new_[992]_  = \new_[162]_  | \new_[991]_ ;
  assign \new_[993]_  = \new_[992]_  | \new_[987]_ ;
  assign \new_[997]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[998]_  = \new_[159]_  | \new_[997]_ ;
  assign \new_[1001]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[1004]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[1005]_  = \new_[1004]_  | \new_[1001]_ ;
  assign \new_[1006]_  = \new_[1005]_  | \new_[998]_ ;
  assign \new_[1007]_  = \new_[1006]_  | \new_[993]_ ;
  assign \new_[1011]_  = \new_[150]_  | \new_[151]_ ;
  assign \new_[1012]_  = \new_[152]_  | \new_[1011]_ ;
  assign \new_[1015]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[1018]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[1019]_  = \new_[1018]_  | \new_[1015]_ ;
  assign \new_[1020]_  = \new_[1019]_  | \new_[1012]_ ;
  assign \new_[1024]_  = \new_[143]_  | \new_[144]_ ;
  assign \new_[1025]_  = \new_[145]_  | \new_[1024]_ ;
  assign \new_[1028]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[1031]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[1032]_  = \new_[1031]_  | \new_[1028]_ ;
  assign \new_[1033]_  = \new_[1032]_  | \new_[1025]_ ;
  assign \new_[1034]_  = \new_[1033]_  | \new_[1020]_ ;
  assign \new_[1035]_  = \new_[1034]_  | \new_[1007]_ ;
  assign \new_[1039]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[1040]_  = \new_[138]_  | \new_[1039]_ ;
  assign \new_[1043]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[1046]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[1047]_  = \new_[1046]_  | \new_[1043]_ ;
  assign \new_[1048]_  = \new_[1047]_  | \new_[1040]_ ;
  assign \new_[1052]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[1053]_  = \new_[131]_  | \new_[1052]_ ;
  assign \new_[1056]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[1059]_  = \new_[125]_  | \new_[126]_ ;
  assign \new_[1060]_  = \new_[1059]_  | \new_[1056]_ ;
  assign \new_[1061]_  = \new_[1060]_  | \new_[1053]_ ;
  assign \new_[1062]_  = \new_[1061]_  | \new_[1048]_ ;
  assign \new_[1066]_  = \new_[122]_  | \new_[123]_ ;
  assign \new_[1067]_  = \new_[124]_  | \new_[1066]_ ;
  assign \new_[1070]_  = \new_[120]_  | \new_[121]_ ;
  assign \new_[1073]_  = \new_[118]_  | \new_[119]_ ;
  assign \new_[1074]_  = \new_[1073]_  | \new_[1070]_ ;
  assign \new_[1075]_  = \new_[1074]_  | \new_[1067]_ ;
  assign \new_[1079]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[1080]_  = \new_[117]_  | \new_[1079]_ ;
  assign \new_[1083]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[1086]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[1087]_  = \new_[1086]_  | \new_[1083]_ ;
  assign \new_[1088]_  = \new_[1087]_  | \new_[1080]_ ;
  assign \new_[1089]_  = \new_[1088]_  | \new_[1075]_ ;
  assign \new_[1090]_  = \new_[1089]_  | \new_[1062]_ ;
  assign \new_[1091]_  = \new_[1090]_  | \new_[1035]_ ;
  assign \new_[1092]_  = \new_[1091]_  | \new_[982]_ ;
  assign \new_[1096]_  = \new_[108]_  | \new_[109]_ ;
  assign \new_[1097]_  = \new_[110]_  | \new_[1096]_ ;
  assign \new_[1101]_  = \new_[105]_  | \new_[106]_ ;
  assign \new_[1102]_  = \new_[107]_  | \new_[1101]_ ;
  assign \new_[1103]_  = \new_[1102]_  | \new_[1097]_ ;
  assign \new_[1107]_  = \new_[102]_  | \new_[103]_ ;
  assign \new_[1108]_  = \new_[104]_  | \new_[1107]_ ;
  assign \new_[1111]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[1114]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[1115]_  = \new_[1114]_  | \new_[1111]_ ;
  assign \new_[1116]_  = \new_[1115]_  | \new_[1108]_ ;
  assign \new_[1117]_  = \new_[1116]_  | \new_[1103]_ ;
  assign \new_[1121]_  = \new_[95]_  | \new_[96]_ ;
  assign \new_[1122]_  = \new_[97]_  | \new_[1121]_ ;
  assign \new_[1125]_  = \new_[93]_  | \new_[94]_ ;
  assign \new_[1128]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[1129]_  = \new_[1128]_  | \new_[1125]_ ;
  assign \new_[1130]_  = \new_[1129]_  | \new_[1122]_ ;
  assign \new_[1134]_  = \new_[88]_  | \new_[89]_ ;
  assign \new_[1135]_  = \new_[90]_  | \new_[1134]_ ;
  assign \new_[1138]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[1141]_  = \new_[84]_  | \new_[85]_ ;
  assign \new_[1142]_  = \new_[1141]_  | \new_[1138]_ ;
  assign \new_[1143]_  = \new_[1142]_  | \new_[1135]_ ;
  assign \new_[1144]_  = \new_[1143]_  | \new_[1130]_ ;
  assign \new_[1145]_  = \new_[1144]_  | \new_[1117]_ ;
  assign \new_[1149]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[1150]_  = \new_[83]_  | \new_[1149]_ ;
  assign \new_[1153]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[1156]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[1157]_  = \new_[1156]_  | \new_[1153]_ ;
  assign \new_[1158]_  = \new_[1157]_  | \new_[1150]_ ;
  assign \new_[1162]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[1163]_  = \new_[76]_  | \new_[1162]_ ;
  assign \new_[1166]_  = \new_[72]_  | \new_[73]_ ;
  assign \new_[1169]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[1170]_  = \new_[1169]_  | \new_[1166]_ ;
  assign \new_[1171]_  = \new_[1170]_  | \new_[1163]_ ;
  assign \new_[1172]_  = \new_[1171]_  | \new_[1158]_ ;
  assign \new_[1176]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[1177]_  = \new_[69]_  | \new_[1176]_ ;
  assign \new_[1180]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[1183]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[1184]_  = \new_[1183]_  | \new_[1180]_ ;
  assign \new_[1185]_  = \new_[1184]_  | \new_[1177]_ ;
  assign \new_[1189]_  = \new_[60]_  | \new_[61]_ ;
  assign \new_[1190]_  = \new_[62]_  | \new_[1189]_ ;
  assign \new_[1193]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[1196]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[1197]_  = \new_[1196]_  | \new_[1193]_ ;
  assign \new_[1198]_  = \new_[1197]_  | \new_[1190]_ ;
  assign \new_[1199]_  = \new_[1198]_  | \new_[1185]_ ;
  assign \new_[1200]_  = \new_[1199]_  | \new_[1172]_ ;
  assign \new_[1201]_  = \new_[1200]_  | \new_[1145]_ ;
  assign \new_[1205]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[1206]_  = \new_[55]_  | \new_[1205]_ ;
  assign \new_[1210]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[1211]_  = \new_[52]_  | \new_[1210]_ ;
  assign \new_[1212]_  = \new_[1211]_  | \new_[1206]_ ;
  assign \new_[1216]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[1217]_  = \new_[49]_  | \new_[1216]_ ;
  assign \new_[1220]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[1223]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[1224]_  = \new_[1223]_  | \new_[1220]_ ;
  assign \new_[1225]_  = \new_[1224]_  | \new_[1217]_ ;
  assign \new_[1226]_  = \new_[1225]_  | \new_[1212]_ ;
  assign \new_[1230]_  = \new_[40]_  | \new_[41]_ ;
  assign \new_[1231]_  = \new_[42]_  | \new_[1230]_ ;
  assign \new_[1234]_  = \new_[38]_  | \new_[39]_ ;
  assign \new_[1237]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[1238]_  = \new_[1237]_  | \new_[1234]_ ;
  assign \new_[1239]_  = \new_[1238]_  | \new_[1231]_ ;
  assign \new_[1243]_  = \new_[33]_  | \new_[34]_ ;
  assign \new_[1244]_  = \new_[35]_  | \new_[1243]_ ;
  assign \new_[1247]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[1250]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[1251]_  = \new_[1250]_  | \new_[1247]_ ;
  assign \new_[1252]_  = \new_[1251]_  | \new_[1244]_ ;
  assign \new_[1253]_  = \new_[1252]_  | \new_[1239]_ ;
  assign \new_[1254]_  = \new_[1253]_  | \new_[1226]_ ;
  assign \new_[1258]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[1259]_  = \new_[28]_  | \new_[1258]_ ;
  assign \new_[1262]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[1265]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[1266]_  = \new_[1265]_  | \new_[1262]_ ;
  assign \new_[1267]_  = \new_[1266]_  | \new_[1259]_ ;
  assign \new_[1271]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[1272]_  = \new_[21]_  | \new_[1271]_ ;
  assign \new_[1275]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[1278]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[1279]_  = \new_[1278]_  | \new_[1275]_ ;
  assign \new_[1280]_  = \new_[1279]_  | \new_[1272]_ ;
  assign \new_[1281]_  = \new_[1280]_  | \new_[1267]_ ;
  assign \new_[1285]_  = \new_[12]_  | \new_[13]_ ;
  assign \new_[1286]_  = \new_[14]_  | \new_[1285]_ ;
  assign \new_[1289]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[1292]_  = \new_[8]_  | \new_[9]_ ;
  assign \new_[1293]_  = \new_[1292]_  | \new_[1289]_ ;
  assign \new_[1294]_  = \new_[1293]_  | \new_[1286]_ ;
  assign \new_[1298]_  = \new_[5]_  | \new_[6]_ ;
  assign \new_[1299]_  = \new_[7]_  | \new_[1298]_ ;
  assign \new_[1302]_  = \new_[3]_  | \new_[4]_ ;
  assign \new_[1305]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[1306]_  = \new_[1305]_  | \new_[1302]_ ;
  assign \new_[1307]_  = \new_[1306]_  | \new_[1299]_ ;
  assign \new_[1308]_  = \new_[1307]_  | \new_[1294]_ ;
  assign \new_[1309]_  = \new_[1308]_  | \new_[1281]_ ;
  assign \new_[1310]_  = \new_[1309]_  | \new_[1254]_ ;
  assign \new_[1311]_  = \new_[1310]_  | \new_[1201]_ ;
  assign \new_[1312]_  = \new_[1311]_  | \new_[1092]_ ;
  assign \new_[1315]_  = A266 & ~A265;
  assign \new_[1318]_  = A268 & A267;
  assign \new_[1321]_  = A266 & ~A265;
  assign \new_[1324]_  = A269 & A267;
  assign \new_[1327]_  = ~A266 & A265;
  assign \new_[1330]_  = A268 & A267;
  assign \new_[1333]_  = ~A266 & A265;
  assign \new_[1336]_  = A269 & A267;
  assign \new_[1339]_  = A266 & ~A265;
  assign \new_[1343]_  = ~A269 & ~A268;
  assign \new_[1344]_  = ~A267 & \new_[1343]_ ;
  assign \new_[1347]_  = ~A266 & A265;
  assign \new_[1351]_  = ~A269 & ~A268;
  assign \new_[1352]_  = ~A267 & \new_[1351]_ ;
  assign \new_[1355]_  = A200 & ~A199;
  assign \new_[1358]_  = A202 & A201;
  assign \new_[1359]_  = \new_[1358]_  & \new_[1355]_ ;
  assign \new_[1362]_  = A233 & ~A232;
  assign \new_[1365]_  = A235 & A234;
  assign \new_[1366]_  = \new_[1365]_  & \new_[1362]_ ;
  assign \new_[1369]_  = A200 & ~A199;
  assign \new_[1372]_  = A202 & A201;
  assign \new_[1373]_  = \new_[1372]_  & \new_[1369]_ ;
  assign \new_[1376]_  = A233 & ~A232;
  assign \new_[1379]_  = A236 & A234;
  assign \new_[1380]_  = \new_[1379]_  & \new_[1376]_ ;
  assign \new_[1383]_  = A200 & ~A199;
  assign \new_[1386]_  = A202 & A201;
  assign \new_[1387]_  = \new_[1386]_  & \new_[1383]_ ;
  assign \new_[1390]_  = ~A233 & A232;
  assign \new_[1393]_  = A235 & A234;
  assign \new_[1394]_  = \new_[1393]_  & \new_[1390]_ ;
  assign \new_[1397]_  = A200 & ~A199;
  assign \new_[1400]_  = A202 & A201;
  assign \new_[1401]_  = \new_[1400]_  & \new_[1397]_ ;
  assign \new_[1404]_  = ~A233 & A232;
  assign \new_[1407]_  = A236 & A234;
  assign \new_[1408]_  = \new_[1407]_  & \new_[1404]_ ;
  assign \new_[1411]_  = A200 & ~A199;
  assign \new_[1414]_  = A203 & A201;
  assign \new_[1415]_  = \new_[1414]_  & \new_[1411]_ ;
  assign \new_[1418]_  = A233 & ~A232;
  assign \new_[1421]_  = A235 & A234;
  assign \new_[1422]_  = \new_[1421]_  & \new_[1418]_ ;
  assign \new_[1425]_  = A200 & ~A199;
  assign \new_[1428]_  = A203 & A201;
  assign \new_[1429]_  = \new_[1428]_  & \new_[1425]_ ;
  assign \new_[1432]_  = A233 & ~A232;
  assign \new_[1435]_  = A236 & A234;
  assign \new_[1436]_  = \new_[1435]_  & \new_[1432]_ ;
  assign \new_[1439]_  = A200 & ~A199;
  assign \new_[1442]_  = A203 & A201;
  assign \new_[1443]_  = \new_[1442]_  & \new_[1439]_ ;
  assign \new_[1446]_  = ~A233 & A232;
  assign \new_[1449]_  = A235 & A234;
  assign \new_[1450]_  = \new_[1449]_  & \new_[1446]_ ;
  assign \new_[1453]_  = A200 & ~A199;
  assign \new_[1456]_  = A203 & A201;
  assign \new_[1457]_  = \new_[1456]_  & \new_[1453]_ ;
  assign \new_[1460]_  = ~A233 & A232;
  assign \new_[1463]_  = A236 & A234;
  assign \new_[1464]_  = \new_[1463]_  & \new_[1460]_ ;
  assign \new_[1467]_  = ~A200 & A199;
  assign \new_[1470]_  = A202 & A201;
  assign \new_[1471]_  = \new_[1470]_  & \new_[1467]_ ;
  assign \new_[1474]_  = A233 & ~A232;
  assign \new_[1477]_  = A235 & A234;
  assign \new_[1478]_  = \new_[1477]_  & \new_[1474]_ ;
  assign \new_[1481]_  = ~A200 & A199;
  assign \new_[1484]_  = A202 & A201;
  assign \new_[1485]_  = \new_[1484]_  & \new_[1481]_ ;
  assign \new_[1488]_  = A233 & ~A232;
  assign \new_[1491]_  = A236 & A234;
  assign \new_[1492]_  = \new_[1491]_  & \new_[1488]_ ;
  assign \new_[1495]_  = ~A200 & A199;
  assign \new_[1498]_  = A202 & A201;
  assign \new_[1499]_  = \new_[1498]_  & \new_[1495]_ ;
  assign \new_[1502]_  = ~A233 & A232;
  assign \new_[1505]_  = A235 & A234;
  assign \new_[1506]_  = \new_[1505]_  & \new_[1502]_ ;
  assign \new_[1509]_  = ~A200 & A199;
  assign \new_[1512]_  = A202 & A201;
  assign \new_[1513]_  = \new_[1512]_  & \new_[1509]_ ;
  assign \new_[1516]_  = ~A233 & A232;
  assign \new_[1519]_  = A236 & A234;
  assign \new_[1520]_  = \new_[1519]_  & \new_[1516]_ ;
  assign \new_[1523]_  = ~A200 & A199;
  assign \new_[1526]_  = A203 & A201;
  assign \new_[1527]_  = \new_[1526]_  & \new_[1523]_ ;
  assign \new_[1530]_  = A233 & ~A232;
  assign \new_[1533]_  = A235 & A234;
  assign \new_[1534]_  = \new_[1533]_  & \new_[1530]_ ;
  assign \new_[1537]_  = ~A200 & A199;
  assign \new_[1540]_  = A203 & A201;
  assign \new_[1541]_  = \new_[1540]_  & \new_[1537]_ ;
  assign \new_[1544]_  = A233 & ~A232;
  assign \new_[1547]_  = A236 & A234;
  assign \new_[1548]_  = \new_[1547]_  & \new_[1544]_ ;
  assign \new_[1551]_  = ~A200 & A199;
  assign \new_[1554]_  = A203 & A201;
  assign \new_[1555]_  = \new_[1554]_  & \new_[1551]_ ;
  assign \new_[1558]_  = ~A233 & A232;
  assign \new_[1561]_  = A235 & A234;
  assign \new_[1562]_  = \new_[1561]_  & \new_[1558]_ ;
  assign \new_[1565]_  = ~A200 & A199;
  assign \new_[1568]_  = A203 & A201;
  assign \new_[1569]_  = \new_[1568]_  & \new_[1565]_ ;
  assign \new_[1572]_  = ~A233 & A232;
  assign \new_[1575]_  = A236 & A234;
  assign \new_[1576]_  = \new_[1575]_  & \new_[1572]_ ;
  assign \new_[1579]_  = A168 & ~A170;
  assign \new_[1582]_  = ~A166 & A167;
  assign \new_[1583]_  = \new_[1582]_  & \new_[1579]_ ;
  assign \new_[1586]_  = A233 & ~A232;
  assign \new_[1589]_  = A235 & A234;
  assign \new_[1590]_  = \new_[1589]_  & \new_[1586]_ ;
  assign \new_[1593]_  = A168 & ~A170;
  assign \new_[1596]_  = ~A166 & A167;
  assign \new_[1597]_  = \new_[1596]_  & \new_[1593]_ ;
  assign \new_[1600]_  = A233 & ~A232;
  assign \new_[1603]_  = A236 & A234;
  assign \new_[1604]_  = \new_[1603]_  & \new_[1600]_ ;
  assign \new_[1607]_  = A168 & ~A170;
  assign \new_[1610]_  = ~A166 & A167;
  assign \new_[1611]_  = \new_[1610]_  & \new_[1607]_ ;
  assign \new_[1614]_  = ~A233 & A232;
  assign \new_[1617]_  = A235 & A234;
  assign \new_[1618]_  = \new_[1617]_  & \new_[1614]_ ;
  assign \new_[1621]_  = A168 & ~A170;
  assign \new_[1624]_  = ~A166 & A167;
  assign \new_[1625]_  = \new_[1624]_  & \new_[1621]_ ;
  assign \new_[1628]_  = ~A233 & A232;
  assign \new_[1631]_  = A236 & A234;
  assign \new_[1632]_  = \new_[1631]_  & \new_[1628]_ ;
  assign \new_[1635]_  = A168 & ~A170;
  assign \new_[1638]_  = A166 & ~A167;
  assign \new_[1639]_  = \new_[1638]_  & \new_[1635]_ ;
  assign \new_[1642]_  = A233 & ~A232;
  assign \new_[1645]_  = A235 & A234;
  assign \new_[1646]_  = \new_[1645]_  & \new_[1642]_ ;
  assign \new_[1649]_  = A168 & ~A170;
  assign \new_[1652]_  = A166 & ~A167;
  assign \new_[1653]_  = \new_[1652]_  & \new_[1649]_ ;
  assign \new_[1656]_  = A233 & ~A232;
  assign \new_[1659]_  = A236 & A234;
  assign \new_[1660]_  = \new_[1659]_  & \new_[1656]_ ;
  assign \new_[1663]_  = A168 & ~A170;
  assign \new_[1666]_  = A166 & ~A167;
  assign \new_[1667]_  = \new_[1666]_  & \new_[1663]_ ;
  assign \new_[1670]_  = ~A233 & A232;
  assign \new_[1673]_  = A235 & A234;
  assign \new_[1674]_  = \new_[1673]_  & \new_[1670]_ ;
  assign \new_[1677]_  = A168 & ~A170;
  assign \new_[1680]_  = A166 & ~A167;
  assign \new_[1681]_  = \new_[1680]_  & \new_[1677]_ ;
  assign \new_[1684]_  = ~A233 & A232;
  assign \new_[1687]_  = A236 & A234;
  assign \new_[1688]_  = \new_[1687]_  & \new_[1684]_ ;
  assign \new_[1691]_  = A168 & A169;
  assign \new_[1694]_  = ~A166 & A167;
  assign \new_[1695]_  = \new_[1694]_  & \new_[1691]_ ;
  assign \new_[1698]_  = A233 & ~A232;
  assign \new_[1701]_  = A235 & A234;
  assign \new_[1702]_  = \new_[1701]_  & \new_[1698]_ ;
  assign \new_[1705]_  = A168 & A169;
  assign \new_[1708]_  = ~A166 & A167;
  assign \new_[1709]_  = \new_[1708]_  & \new_[1705]_ ;
  assign \new_[1712]_  = A233 & ~A232;
  assign \new_[1715]_  = A236 & A234;
  assign \new_[1716]_  = \new_[1715]_  & \new_[1712]_ ;
  assign \new_[1719]_  = A168 & A169;
  assign \new_[1722]_  = ~A166 & A167;
  assign \new_[1723]_  = \new_[1722]_  & \new_[1719]_ ;
  assign \new_[1726]_  = ~A233 & A232;
  assign \new_[1729]_  = A235 & A234;
  assign \new_[1730]_  = \new_[1729]_  & \new_[1726]_ ;
  assign \new_[1733]_  = A168 & A169;
  assign \new_[1736]_  = ~A166 & A167;
  assign \new_[1737]_  = \new_[1736]_  & \new_[1733]_ ;
  assign \new_[1740]_  = ~A233 & A232;
  assign \new_[1743]_  = A236 & A234;
  assign \new_[1744]_  = \new_[1743]_  & \new_[1740]_ ;
  assign \new_[1747]_  = A168 & A169;
  assign \new_[1750]_  = A166 & ~A167;
  assign \new_[1751]_  = \new_[1750]_  & \new_[1747]_ ;
  assign \new_[1754]_  = A233 & ~A232;
  assign \new_[1757]_  = A235 & A234;
  assign \new_[1758]_  = \new_[1757]_  & \new_[1754]_ ;
  assign \new_[1761]_  = A168 & A169;
  assign \new_[1764]_  = A166 & ~A167;
  assign \new_[1765]_  = \new_[1764]_  & \new_[1761]_ ;
  assign \new_[1768]_  = A233 & ~A232;
  assign \new_[1771]_  = A236 & A234;
  assign \new_[1772]_  = \new_[1771]_  & \new_[1768]_ ;
  assign \new_[1775]_  = A168 & A169;
  assign \new_[1778]_  = A166 & ~A167;
  assign \new_[1779]_  = \new_[1778]_  & \new_[1775]_ ;
  assign \new_[1782]_  = ~A233 & A232;
  assign \new_[1785]_  = A235 & A234;
  assign \new_[1786]_  = \new_[1785]_  & \new_[1782]_ ;
  assign \new_[1789]_  = A168 & A169;
  assign \new_[1792]_  = A166 & ~A167;
  assign \new_[1793]_  = \new_[1792]_  & \new_[1789]_ ;
  assign \new_[1796]_  = ~A233 & A232;
  assign \new_[1799]_  = A236 & A234;
  assign \new_[1800]_  = \new_[1799]_  & \new_[1796]_ ;
  assign \new_[1803]_  = A200 & ~A199;
  assign \new_[1806]_  = A202 & A201;
  assign \new_[1807]_  = \new_[1806]_  & \new_[1803]_ ;
  assign \new_[1810]_  = A233 & ~A232;
  assign \new_[1814]_  = ~A236 & ~A235;
  assign \new_[1815]_  = ~A234 & \new_[1814]_ ;
  assign \new_[1816]_  = \new_[1815]_  & \new_[1810]_ ;
  assign \new_[1819]_  = A200 & ~A199;
  assign \new_[1822]_  = A202 & A201;
  assign \new_[1823]_  = \new_[1822]_  & \new_[1819]_ ;
  assign \new_[1826]_  = ~A233 & A232;
  assign \new_[1830]_  = ~A236 & ~A235;
  assign \new_[1831]_  = ~A234 & \new_[1830]_ ;
  assign \new_[1832]_  = \new_[1831]_  & \new_[1826]_ ;
  assign \new_[1835]_  = A200 & ~A199;
  assign \new_[1838]_  = A203 & A201;
  assign \new_[1839]_  = \new_[1838]_  & \new_[1835]_ ;
  assign \new_[1842]_  = A233 & ~A232;
  assign \new_[1846]_  = ~A236 & ~A235;
  assign \new_[1847]_  = ~A234 & \new_[1846]_ ;
  assign \new_[1848]_  = \new_[1847]_  & \new_[1842]_ ;
  assign \new_[1851]_  = A200 & ~A199;
  assign \new_[1854]_  = A203 & A201;
  assign \new_[1855]_  = \new_[1854]_  & \new_[1851]_ ;
  assign \new_[1858]_  = ~A233 & A232;
  assign \new_[1862]_  = ~A236 & ~A235;
  assign \new_[1863]_  = ~A234 & \new_[1862]_ ;
  assign \new_[1864]_  = \new_[1863]_  & \new_[1858]_ ;
  assign \new_[1867]_  = A200 & ~A199;
  assign \new_[1870]_  = ~A202 & ~A201;
  assign \new_[1871]_  = \new_[1870]_  & \new_[1867]_ ;
  assign \new_[1874]_  = ~A232 & ~A203;
  assign \new_[1878]_  = A235 & A234;
  assign \new_[1879]_  = A233 & \new_[1878]_ ;
  assign \new_[1880]_  = \new_[1879]_  & \new_[1874]_ ;
  assign \new_[1883]_  = A200 & ~A199;
  assign \new_[1886]_  = ~A202 & ~A201;
  assign \new_[1887]_  = \new_[1886]_  & \new_[1883]_ ;
  assign \new_[1890]_  = ~A232 & ~A203;
  assign \new_[1894]_  = A236 & A234;
  assign \new_[1895]_  = A233 & \new_[1894]_ ;
  assign \new_[1896]_  = \new_[1895]_  & \new_[1890]_ ;
  assign \new_[1899]_  = A200 & ~A199;
  assign \new_[1902]_  = ~A202 & ~A201;
  assign \new_[1903]_  = \new_[1902]_  & \new_[1899]_ ;
  assign \new_[1906]_  = A232 & ~A203;
  assign \new_[1910]_  = A235 & A234;
  assign \new_[1911]_  = ~A233 & \new_[1910]_ ;
  assign \new_[1912]_  = \new_[1911]_  & \new_[1906]_ ;
  assign \new_[1915]_  = A200 & ~A199;
  assign \new_[1918]_  = ~A202 & ~A201;
  assign \new_[1919]_  = \new_[1918]_  & \new_[1915]_ ;
  assign \new_[1922]_  = A232 & ~A203;
  assign \new_[1926]_  = A236 & A234;
  assign \new_[1927]_  = ~A233 & \new_[1926]_ ;
  assign \new_[1928]_  = \new_[1927]_  & \new_[1922]_ ;
  assign \new_[1931]_  = ~A200 & A199;
  assign \new_[1934]_  = A202 & A201;
  assign \new_[1935]_  = \new_[1934]_  & \new_[1931]_ ;
  assign \new_[1938]_  = A233 & ~A232;
  assign \new_[1942]_  = ~A236 & ~A235;
  assign \new_[1943]_  = ~A234 & \new_[1942]_ ;
  assign \new_[1944]_  = \new_[1943]_  & \new_[1938]_ ;
  assign \new_[1947]_  = ~A200 & A199;
  assign \new_[1950]_  = A202 & A201;
  assign \new_[1951]_  = \new_[1950]_  & \new_[1947]_ ;
  assign \new_[1954]_  = ~A233 & A232;
  assign \new_[1958]_  = ~A236 & ~A235;
  assign \new_[1959]_  = ~A234 & \new_[1958]_ ;
  assign \new_[1960]_  = \new_[1959]_  & \new_[1954]_ ;
  assign \new_[1963]_  = ~A200 & A199;
  assign \new_[1966]_  = A203 & A201;
  assign \new_[1967]_  = \new_[1966]_  & \new_[1963]_ ;
  assign \new_[1970]_  = A233 & ~A232;
  assign \new_[1974]_  = ~A236 & ~A235;
  assign \new_[1975]_  = ~A234 & \new_[1974]_ ;
  assign \new_[1976]_  = \new_[1975]_  & \new_[1970]_ ;
  assign \new_[1979]_  = ~A200 & A199;
  assign \new_[1982]_  = A203 & A201;
  assign \new_[1983]_  = \new_[1982]_  & \new_[1979]_ ;
  assign \new_[1986]_  = ~A233 & A232;
  assign \new_[1990]_  = ~A236 & ~A235;
  assign \new_[1991]_  = ~A234 & \new_[1990]_ ;
  assign \new_[1992]_  = \new_[1991]_  & \new_[1986]_ ;
  assign \new_[1995]_  = ~A200 & A199;
  assign \new_[1998]_  = ~A202 & ~A201;
  assign \new_[1999]_  = \new_[1998]_  & \new_[1995]_ ;
  assign \new_[2002]_  = ~A232 & ~A203;
  assign \new_[2006]_  = A235 & A234;
  assign \new_[2007]_  = A233 & \new_[2006]_ ;
  assign \new_[2008]_  = \new_[2007]_  & \new_[2002]_ ;
  assign \new_[2011]_  = ~A200 & A199;
  assign \new_[2014]_  = ~A202 & ~A201;
  assign \new_[2015]_  = \new_[2014]_  & \new_[2011]_ ;
  assign \new_[2018]_  = ~A232 & ~A203;
  assign \new_[2022]_  = A236 & A234;
  assign \new_[2023]_  = A233 & \new_[2022]_ ;
  assign \new_[2024]_  = \new_[2023]_  & \new_[2018]_ ;
  assign \new_[2027]_  = ~A200 & A199;
  assign \new_[2030]_  = ~A202 & ~A201;
  assign \new_[2031]_  = \new_[2030]_  & \new_[2027]_ ;
  assign \new_[2034]_  = A232 & ~A203;
  assign \new_[2038]_  = A235 & A234;
  assign \new_[2039]_  = ~A233 & \new_[2038]_ ;
  assign \new_[2040]_  = \new_[2039]_  & \new_[2034]_ ;
  assign \new_[2043]_  = ~A200 & A199;
  assign \new_[2046]_  = ~A202 & ~A201;
  assign \new_[2047]_  = \new_[2046]_  & \new_[2043]_ ;
  assign \new_[2050]_  = A232 & ~A203;
  assign \new_[2054]_  = A236 & A234;
  assign \new_[2055]_  = ~A233 & \new_[2054]_ ;
  assign \new_[2056]_  = \new_[2055]_  & \new_[2050]_ ;
  assign \new_[2059]_  = A168 & ~A170;
  assign \new_[2062]_  = ~A166 & A167;
  assign \new_[2063]_  = \new_[2062]_  & \new_[2059]_ ;
  assign \new_[2066]_  = A233 & ~A232;
  assign \new_[2070]_  = ~A236 & ~A235;
  assign \new_[2071]_  = ~A234 & \new_[2070]_ ;
  assign \new_[2072]_  = \new_[2071]_  & \new_[2066]_ ;
  assign \new_[2075]_  = A168 & ~A170;
  assign \new_[2078]_  = ~A166 & A167;
  assign \new_[2079]_  = \new_[2078]_  & \new_[2075]_ ;
  assign \new_[2082]_  = ~A233 & A232;
  assign \new_[2086]_  = ~A236 & ~A235;
  assign \new_[2087]_  = ~A234 & \new_[2086]_ ;
  assign \new_[2088]_  = \new_[2087]_  & \new_[2082]_ ;
  assign \new_[2091]_  = A168 & ~A170;
  assign \new_[2094]_  = A166 & ~A167;
  assign \new_[2095]_  = \new_[2094]_  & \new_[2091]_ ;
  assign \new_[2098]_  = A233 & ~A232;
  assign \new_[2102]_  = ~A236 & ~A235;
  assign \new_[2103]_  = ~A234 & \new_[2102]_ ;
  assign \new_[2104]_  = \new_[2103]_  & \new_[2098]_ ;
  assign \new_[2107]_  = A168 & ~A170;
  assign \new_[2110]_  = A166 & ~A167;
  assign \new_[2111]_  = \new_[2110]_  & \new_[2107]_ ;
  assign \new_[2114]_  = ~A233 & A232;
  assign \new_[2118]_  = ~A236 & ~A235;
  assign \new_[2119]_  = ~A234 & \new_[2118]_ ;
  assign \new_[2120]_  = \new_[2119]_  & \new_[2114]_ ;
  assign \new_[2123]_  = A168 & A169;
  assign \new_[2126]_  = ~A166 & A167;
  assign \new_[2127]_  = \new_[2126]_  & \new_[2123]_ ;
  assign \new_[2130]_  = A233 & ~A232;
  assign \new_[2134]_  = ~A236 & ~A235;
  assign \new_[2135]_  = ~A234 & \new_[2134]_ ;
  assign \new_[2136]_  = \new_[2135]_  & \new_[2130]_ ;
  assign \new_[2139]_  = A168 & A169;
  assign \new_[2142]_  = ~A166 & A167;
  assign \new_[2143]_  = \new_[2142]_  & \new_[2139]_ ;
  assign \new_[2146]_  = ~A233 & A232;
  assign \new_[2150]_  = ~A236 & ~A235;
  assign \new_[2151]_  = ~A234 & \new_[2150]_ ;
  assign \new_[2152]_  = \new_[2151]_  & \new_[2146]_ ;
  assign \new_[2155]_  = A168 & A169;
  assign \new_[2158]_  = A166 & ~A167;
  assign \new_[2159]_  = \new_[2158]_  & \new_[2155]_ ;
  assign \new_[2162]_  = A233 & ~A232;
  assign \new_[2166]_  = ~A236 & ~A235;
  assign \new_[2167]_  = ~A234 & \new_[2166]_ ;
  assign \new_[2168]_  = \new_[2167]_  & \new_[2162]_ ;
  assign \new_[2171]_  = A168 & A169;
  assign \new_[2174]_  = A166 & ~A167;
  assign \new_[2175]_  = \new_[2174]_  & \new_[2171]_ ;
  assign \new_[2178]_  = ~A233 & A232;
  assign \new_[2182]_  = ~A236 & ~A235;
  assign \new_[2183]_  = ~A234 & \new_[2182]_ ;
  assign \new_[2184]_  = \new_[2183]_  & \new_[2178]_ ;
  assign \new_[2187]_  = ~A169 & A170;
  assign \new_[2190]_  = A167 & ~A168;
  assign \new_[2191]_  = \new_[2190]_  & \new_[2187]_ ;
  assign \new_[2194]_  = ~A232 & ~A166;
  assign \new_[2198]_  = A235 & A234;
  assign \new_[2199]_  = A233 & \new_[2198]_ ;
  assign \new_[2200]_  = \new_[2199]_  & \new_[2194]_ ;
  assign \new_[2203]_  = ~A169 & A170;
  assign \new_[2206]_  = A167 & ~A168;
  assign \new_[2207]_  = \new_[2206]_  & \new_[2203]_ ;
  assign \new_[2210]_  = ~A232 & ~A166;
  assign \new_[2214]_  = A236 & A234;
  assign \new_[2215]_  = A233 & \new_[2214]_ ;
  assign \new_[2216]_  = \new_[2215]_  & \new_[2210]_ ;
  assign \new_[2219]_  = ~A169 & A170;
  assign \new_[2222]_  = A167 & ~A168;
  assign \new_[2223]_  = \new_[2222]_  & \new_[2219]_ ;
  assign \new_[2226]_  = A232 & ~A166;
  assign \new_[2230]_  = A235 & A234;
  assign \new_[2231]_  = ~A233 & \new_[2230]_ ;
  assign \new_[2232]_  = \new_[2231]_  & \new_[2226]_ ;
  assign \new_[2235]_  = ~A169 & A170;
  assign \new_[2238]_  = A167 & ~A168;
  assign \new_[2239]_  = \new_[2238]_  & \new_[2235]_ ;
  assign \new_[2242]_  = A232 & ~A166;
  assign \new_[2246]_  = A236 & A234;
  assign \new_[2247]_  = ~A233 & \new_[2246]_ ;
  assign \new_[2248]_  = \new_[2247]_  & \new_[2242]_ ;
  assign \new_[2251]_  = ~A169 & A170;
  assign \new_[2254]_  = ~A167 & ~A168;
  assign \new_[2255]_  = \new_[2254]_  & \new_[2251]_ ;
  assign \new_[2258]_  = ~A232 & A166;
  assign \new_[2262]_  = A235 & A234;
  assign \new_[2263]_  = A233 & \new_[2262]_ ;
  assign \new_[2264]_  = \new_[2263]_  & \new_[2258]_ ;
  assign \new_[2267]_  = ~A169 & A170;
  assign \new_[2270]_  = ~A167 & ~A168;
  assign \new_[2271]_  = \new_[2270]_  & \new_[2267]_ ;
  assign \new_[2274]_  = ~A232 & A166;
  assign \new_[2278]_  = A236 & A234;
  assign \new_[2279]_  = A233 & \new_[2278]_ ;
  assign \new_[2280]_  = \new_[2279]_  & \new_[2274]_ ;
  assign \new_[2283]_  = ~A169 & A170;
  assign \new_[2286]_  = ~A167 & ~A168;
  assign \new_[2287]_  = \new_[2286]_  & \new_[2283]_ ;
  assign \new_[2290]_  = A232 & A166;
  assign \new_[2294]_  = A235 & A234;
  assign \new_[2295]_  = ~A233 & \new_[2294]_ ;
  assign \new_[2296]_  = \new_[2295]_  & \new_[2290]_ ;
  assign \new_[2299]_  = ~A169 & A170;
  assign \new_[2302]_  = ~A167 & ~A168;
  assign \new_[2303]_  = \new_[2302]_  & \new_[2299]_ ;
  assign \new_[2306]_  = A232 & A166;
  assign \new_[2310]_  = A236 & A234;
  assign \new_[2311]_  = ~A233 & \new_[2310]_ ;
  assign \new_[2312]_  = \new_[2311]_  & \new_[2306]_ ;
  assign \new_[2315]_  = A200 & ~A199;
  assign \new_[2319]_  = ~A203 & ~A202;
  assign \new_[2320]_  = ~A201 & \new_[2319]_ ;
  assign \new_[2321]_  = \new_[2320]_  & \new_[2315]_ ;
  assign \new_[2324]_  = A233 & ~A232;
  assign \new_[2328]_  = ~A236 & ~A235;
  assign \new_[2329]_  = ~A234 & \new_[2328]_ ;
  assign \new_[2330]_  = \new_[2329]_  & \new_[2324]_ ;
  assign \new_[2333]_  = A200 & ~A199;
  assign \new_[2337]_  = ~A203 & ~A202;
  assign \new_[2338]_  = ~A201 & \new_[2337]_ ;
  assign \new_[2339]_  = \new_[2338]_  & \new_[2333]_ ;
  assign \new_[2342]_  = ~A233 & A232;
  assign \new_[2346]_  = ~A236 & ~A235;
  assign \new_[2347]_  = ~A234 & \new_[2346]_ ;
  assign \new_[2348]_  = \new_[2347]_  & \new_[2342]_ ;
  assign \new_[2351]_  = ~A200 & A199;
  assign \new_[2355]_  = ~A203 & ~A202;
  assign \new_[2356]_  = ~A201 & \new_[2355]_ ;
  assign \new_[2357]_  = \new_[2356]_  & \new_[2351]_ ;
  assign \new_[2360]_  = A233 & ~A232;
  assign \new_[2364]_  = ~A236 & ~A235;
  assign \new_[2365]_  = ~A234 & \new_[2364]_ ;
  assign \new_[2366]_  = \new_[2365]_  & \new_[2360]_ ;
  assign \new_[2369]_  = ~A200 & A199;
  assign \new_[2373]_  = ~A203 & ~A202;
  assign \new_[2374]_  = ~A201 & \new_[2373]_ ;
  assign \new_[2375]_  = \new_[2374]_  & \new_[2369]_ ;
  assign \new_[2378]_  = ~A233 & A232;
  assign \new_[2382]_  = ~A236 & ~A235;
  assign \new_[2383]_  = ~A234 & \new_[2382]_ ;
  assign \new_[2384]_  = \new_[2383]_  & \new_[2378]_ ;
  assign \new_[2387]_  = A166 & A167;
  assign \new_[2391]_  = A201 & A200;
  assign \new_[2392]_  = ~A199 & \new_[2391]_ ;
  assign \new_[2393]_  = \new_[2392]_  & \new_[2387]_ ;
  assign \new_[2396]_  = A298 & A202;
  assign \new_[2400]_  = A301 & A300;
  assign \new_[2401]_  = ~A299 & \new_[2400]_ ;
  assign \new_[2402]_  = \new_[2401]_  & \new_[2396]_ ;
  assign \new_[2405]_  = A166 & A167;
  assign \new_[2409]_  = A201 & A200;
  assign \new_[2410]_  = ~A199 & \new_[2409]_ ;
  assign \new_[2411]_  = \new_[2410]_  & \new_[2405]_ ;
  assign \new_[2414]_  = A298 & A202;
  assign \new_[2418]_  = A302 & A300;
  assign \new_[2419]_  = ~A299 & \new_[2418]_ ;
  assign \new_[2420]_  = \new_[2419]_  & \new_[2414]_ ;
  assign \new_[2423]_  = A166 & A167;
  assign \new_[2427]_  = A201 & A200;
  assign \new_[2428]_  = ~A199 & \new_[2427]_ ;
  assign \new_[2429]_  = \new_[2428]_  & \new_[2423]_ ;
  assign \new_[2432]_  = ~A298 & A202;
  assign \new_[2436]_  = A301 & A300;
  assign \new_[2437]_  = A299 & \new_[2436]_ ;
  assign \new_[2438]_  = \new_[2437]_  & \new_[2432]_ ;
  assign \new_[2441]_  = A166 & A167;
  assign \new_[2445]_  = A201 & A200;
  assign \new_[2446]_  = ~A199 & \new_[2445]_ ;
  assign \new_[2447]_  = \new_[2446]_  & \new_[2441]_ ;
  assign \new_[2450]_  = ~A298 & A202;
  assign \new_[2454]_  = A302 & A300;
  assign \new_[2455]_  = A299 & \new_[2454]_ ;
  assign \new_[2456]_  = \new_[2455]_  & \new_[2450]_ ;
  assign \new_[2459]_  = A166 & A167;
  assign \new_[2463]_  = A201 & A200;
  assign \new_[2464]_  = ~A199 & \new_[2463]_ ;
  assign \new_[2465]_  = \new_[2464]_  & \new_[2459]_ ;
  assign \new_[2468]_  = A298 & A203;
  assign \new_[2472]_  = A301 & A300;
  assign \new_[2473]_  = ~A299 & \new_[2472]_ ;
  assign \new_[2474]_  = \new_[2473]_  & \new_[2468]_ ;
  assign \new_[2477]_  = A166 & A167;
  assign \new_[2481]_  = A201 & A200;
  assign \new_[2482]_  = ~A199 & \new_[2481]_ ;
  assign \new_[2483]_  = \new_[2482]_  & \new_[2477]_ ;
  assign \new_[2486]_  = A298 & A203;
  assign \new_[2490]_  = A302 & A300;
  assign \new_[2491]_  = ~A299 & \new_[2490]_ ;
  assign \new_[2492]_  = \new_[2491]_  & \new_[2486]_ ;
  assign \new_[2495]_  = A166 & A167;
  assign \new_[2499]_  = A201 & A200;
  assign \new_[2500]_  = ~A199 & \new_[2499]_ ;
  assign \new_[2501]_  = \new_[2500]_  & \new_[2495]_ ;
  assign \new_[2504]_  = ~A298 & A203;
  assign \new_[2508]_  = A301 & A300;
  assign \new_[2509]_  = A299 & \new_[2508]_ ;
  assign \new_[2510]_  = \new_[2509]_  & \new_[2504]_ ;
  assign \new_[2513]_  = A166 & A167;
  assign \new_[2517]_  = A201 & A200;
  assign \new_[2518]_  = ~A199 & \new_[2517]_ ;
  assign \new_[2519]_  = \new_[2518]_  & \new_[2513]_ ;
  assign \new_[2522]_  = ~A298 & A203;
  assign \new_[2526]_  = A302 & A300;
  assign \new_[2527]_  = A299 & \new_[2526]_ ;
  assign \new_[2528]_  = \new_[2527]_  & \new_[2522]_ ;
  assign \new_[2531]_  = A166 & A167;
  assign \new_[2535]_  = A201 & ~A200;
  assign \new_[2536]_  = A199 & \new_[2535]_ ;
  assign \new_[2537]_  = \new_[2536]_  & \new_[2531]_ ;
  assign \new_[2540]_  = A298 & A202;
  assign \new_[2544]_  = A301 & A300;
  assign \new_[2545]_  = ~A299 & \new_[2544]_ ;
  assign \new_[2546]_  = \new_[2545]_  & \new_[2540]_ ;
  assign \new_[2549]_  = A166 & A167;
  assign \new_[2553]_  = A201 & ~A200;
  assign \new_[2554]_  = A199 & \new_[2553]_ ;
  assign \new_[2555]_  = \new_[2554]_  & \new_[2549]_ ;
  assign \new_[2558]_  = A298 & A202;
  assign \new_[2562]_  = A302 & A300;
  assign \new_[2563]_  = ~A299 & \new_[2562]_ ;
  assign \new_[2564]_  = \new_[2563]_  & \new_[2558]_ ;
  assign \new_[2567]_  = A166 & A167;
  assign \new_[2571]_  = A201 & ~A200;
  assign \new_[2572]_  = A199 & \new_[2571]_ ;
  assign \new_[2573]_  = \new_[2572]_  & \new_[2567]_ ;
  assign \new_[2576]_  = ~A298 & A202;
  assign \new_[2580]_  = A301 & A300;
  assign \new_[2581]_  = A299 & \new_[2580]_ ;
  assign \new_[2582]_  = \new_[2581]_  & \new_[2576]_ ;
  assign \new_[2585]_  = A166 & A167;
  assign \new_[2589]_  = A201 & ~A200;
  assign \new_[2590]_  = A199 & \new_[2589]_ ;
  assign \new_[2591]_  = \new_[2590]_  & \new_[2585]_ ;
  assign \new_[2594]_  = ~A298 & A202;
  assign \new_[2598]_  = A302 & A300;
  assign \new_[2599]_  = A299 & \new_[2598]_ ;
  assign \new_[2600]_  = \new_[2599]_  & \new_[2594]_ ;
  assign \new_[2603]_  = A166 & A167;
  assign \new_[2607]_  = A201 & ~A200;
  assign \new_[2608]_  = A199 & \new_[2607]_ ;
  assign \new_[2609]_  = \new_[2608]_  & \new_[2603]_ ;
  assign \new_[2612]_  = A298 & A203;
  assign \new_[2616]_  = A301 & A300;
  assign \new_[2617]_  = ~A299 & \new_[2616]_ ;
  assign \new_[2618]_  = \new_[2617]_  & \new_[2612]_ ;
  assign \new_[2621]_  = A166 & A167;
  assign \new_[2625]_  = A201 & ~A200;
  assign \new_[2626]_  = A199 & \new_[2625]_ ;
  assign \new_[2627]_  = \new_[2626]_  & \new_[2621]_ ;
  assign \new_[2630]_  = A298 & A203;
  assign \new_[2634]_  = A302 & A300;
  assign \new_[2635]_  = ~A299 & \new_[2634]_ ;
  assign \new_[2636]_  = \new_[2635]_  & \new_[2630]_ ;
  assign \new_[2639]_  = A166 & A167;
  assign \new_[2643]_  = A201 & ~A200;
  assign \new_[2644]_  = A199 & \new_[2643]_ ;
  assign \new_[2645]_  = \new_[2644]_  & \new_[2639]_ ;
  assign \new_[2648]_  = ~A298 & A203;
  assign \new_[2652]_  = A301 & A300;
  assign \new_[2653]_  = A299 & \new_[2652]_ ;
  assign \new_[2654]_  = \new_[2653]_  & \new_[2648]_ ;
  assign \new_[2657]_  = A166 & A167;
  assign \new_[2661]_  = A201 & ~A200;
  assign \new_[2662]_  = A199 & \new_[2661]_ ;
  assign \new_[2663]_  = \new_[2662]_  & \new_[2657]_ ;
  assign \new_[2666]_  = ~A298 & A203;
  assign \new_[2670]_  = A302 & A300;
  assign \new_[2671]_  = A299 & \new_[2670]_ ;
  assign \new_[2672]_  = \new_[2671]_  & \new_[2666]_ ;
  assign \new_[2675]_  = ~A166 & ~A167;
  assign \new_[2679]_  = A201 & A200;
  assign \new_[2680]_  = ~A199 & \new_[2679]_ ;
  assign \new_[2681]_  = \new_[2680]_  & \new_[2675]_ ;
  assign \new_[2684]_  = A298 & A202;
  assign \new_[2688]_  = A301 & A300;
  assign \new_[2689]_  = ~A299 & \new_[2688]_ ;
  assign \new_[2690]_  = \new_[2689]_  & \new_[2684]_ ;
  assign \new_[2693]_  = ~A166 & ~A167;
  assign \new_[2697]_  = A201 & A200;
  assign \new_[2698]_  = ~A199 & \new_[2697]_ ;
  assign \new_[2699]_  = \new_[2698]_  & \new_[2693]_ ;
  assign \new_[2702]_  = A298 & A202;
  assign \new_[2706]_  = A302 & A300;
  assign \new_[2707]_  = ~A299 & \new_[2706]_ ;
  assign \new_[2708]_  = \new_[2707]_  & \new_[2702]_ ;
  assign \new_[2711]_  = ~A166 & ~A167;
  assign \new_[2715]_  = A201 & A200;
  assign \new_[2716]_  = ~A199 & \new_[2715]_ ;
  assign \new_[2717]_  = \new_[2716]_  & \new_[2711]_ ;
  assign \new_[2720]_  = ~A298 & A202;
  assign \new_[2724]_  = A301 & A300;
  assign \new_[2725]_  = A299 & \new_[2724]_ ;
  assign \new_[2726]_  = \new_[2725]_  & \new_[2720]_ ;
  assign \new_[2729]_  = ~A166 & ~A167;
  assign \new_[2733]_  = A201 & A200;
  assign \new_[2734]_  = ~A199 & \new_[2733]_ ;
  assign \new_[2735]_  = \new_[2734]_  & \new_[2729]_ ;
  assign \new_[2738]_  = ~A298 & A202;
  assign \new_[2742]_  = A302 & A300;
  assign \new_[2743]_  = A299 & \new_[2742]_ ;
  assign \new_[2744]_  = \new_[2743]_  & \new_[2738]_ ;
  assign \new_[2747]_  = ~A166 & ~A167;
  assign \new_[2751]_  = A201 & A200;
  assign \new_[2752]_  = ~A199 & \new_[2751]_ ;
  assign \new_[2753]_  = \new_[2752]_  & \new_[2747]_ ;
  assign \new_[2756]_  = A298 & A203;
  assign \new_[2760]_  = A301 & A300;
  assign \new_[2761]_  = ~A299 & \new_[2760]_ ;
  assign \new_[2762]_  = \new_[2761]_  & \new_[2756]_ ;
  assign \new_[2765]_  = ~A166 & ~A167;
  assign \new_[2769]_  = A201 & A200;
  assign \new_[2770]_  = ~A199 & \new_[2769]_ ;
  assign \new_[2771]_  = \new_[2770]_  & \new_[2765]_ ;
  assign \new_[2774]_  = A298 & A203;
  assign \new_[2778]_  = A302 & A300;
  assign \new_[2779]_  = ~A299 & \new_[2778]_ ;
  assign \new_[2780]_  = \new_[2779]_  & \new_[2774]_ ;
  assign \new_[2783]_  = ~A166 & ~A167;
  assign \new_[2787]_  = A201 & A200;
  assign \new_[2788]_  = ~A199 & \new_[2787]_ ;
  assign \new_[2789]_  = \new_[2788]_  & \new_[2783]_ ;
  assign \new_[2792]_  = ~A298 & A203;
  assign \new_[2796]_  = A301 & A300;
  assign \new_[2797]_  = A299 & \new_[2796]_ ;
  assign \new_[2798]_  = \new_[2797]_  & \new_[2792]_ ;
  assign \new_[2801]_  = ~A166 & ~A167;
  assign \new_[2805]_  = A201 & A200;
  assign \new_[2806]_  = ~A199 & \new_[2805]_ ;
  assign \new_[2807]_  = \new_[2806]_  & \new_[2801]_ ;
  assign \new_[2810]_  = ~A298 & A203;
  assign \new_[2814]_  = A302 & A300;
  assign \new_[2815]_  = A299 & \new_[2814]_ ;
  assign \new_[2816]_  = \new_[2815]_  & \new_[2810]_ ;
  assign \new_[2819]_  = ~A166 & ~A167;
  assign \new_[2823]_  = A201 & ~A200;
  assign \new_[2824]_  = A199 & \new_[2823]_ ;
  assign \new_[2825]_  = \new_[2824]_  & \new_[2819]_ ;
  assign \new_[2828]_  = A298 & A202;
  assign \new_[2832]_  = A301 & A300;
  assign \new_[2833]_  = ~A299 & \new_[2832]_ ;
  assign \new_[2834]_  = \new_[2833]_  & \new_[2828]_ ;
  assign \new_[2837]_  = ~A166 & ~A167;
  assign \new_[2841]_  = A201 & ~A200;
  assign \new_[2842]_  = A199 & \new_[2841]_ ;
  assign \new_[2843]_  = \new_[2842]_  & \new_[2837]_ ;
  assign \new_[2846]_  = A298 & A202;
  assign \new_[2850]_  = A302 & A300;
  assign \new_[2851]_  = ~A299 & \new_[2850]_ ;
  assign \new_[2852]_  = \new_[2851]_  & \new_[2846]_ ;
  assign \new_[2855]_  = ~A166 & ~A167;
  assign \new_[2859]_  = A201 & ~A200;
  assign \new_[2860]_  = A199 & \new_[2859]_ ;
  assign \new_[2861]_  = \new_[2860]_  & \new_[2855]_ ;
  assign \new_[2864]_  = ~A298 & A202;
  assign \new_[2868]_  = A301 & A300;
  assign \new_[2869]_  = A299 & \new_[2868]_ ;
  assign \new_[2870]_  = \new_[2869]_  & \new_[2864]_ ;
  assign \new_[2873]_  = ~A166 & ~A167;
  assign \new_[2877]_  = A201 & ~A200;
  assign \new_[2878]_  = A199 & \new_[2877]_ ;
  assign \new_[2879]_  = \new_[2878]_  & \new_[2873]_ ;
  assign \new_[2882]_  = ~A298 & A202;
  assign \new_[2886]_  = A302 & A300;
  assign \new_[2887]_  = A299 & \new_[2886]_ ;
  assign \new_[2888]_  = \new_[2887]_  & \new_[2882]_ ;
  assign \new_[2891]_  = ~A166 & ~A167;
  assign \new_[2895]_  = A201 & ~A200;
  assign \new_[2896]_  = A199 & \new_[2895]_ ;
  assign \new_[2897]_  = \new_[2896]_  & \new_[2891]_ ;
  assign \new_[2900]_  = A298 & A203;
  assign \new_[2904]_  = A301 & A300;
  assign \new_[2905]_  = ~A299 & \new_[2904]_ ;
  assign \new_[2906]_  = \new_[2905]_  & \new_[2900]_ ;
  assign \new_[2909]_  = ~A166 & ~A167;
  assign \new_[2913]_  = A201 & ~A200;
  assign \new_[2914]_  = A199 & \new_[2913]_ ;
  assign \new_[2915]_  = \new_[2914]_  & \new_[2909]_ ;
  assign \new_[2918]_  = A298 & A203;
  assign \new_[2922]_  = A302 & A300;
  assign \new_[2923]_  = ~A299 & \new_[2922]_ ;
  assign \new_[2924]_  = \new_[2923]_  & \new_[2918]_ ;
  assign \new_[2927]_  = ~A166 & ~A167;
  assign \new_[2931]_  = A201 & ~A200;
  assign \new_[2932]_  = A199 & \new_[2931]_ ;
  assign \new_[2933]_  = \new_[2932]_  & \new_[2927]_ ;
  assign \new_[2936]_  = ~A298 & A203;
  assign \new_[2940]_  = A301 & A300;
  assign \new_[2941]_  = A299 & \new_[2940]_ ;
  assign \new_[2942]_  = \new_[2941]_  & \new_[2936]_ ;
  assign \new_[2945]_  = ~A166 & ~A167;
  assign \new_[2949]_  = A201 & ~A200;
  assign \new_[2950]_  = A199 & \new_[2949]_ ;
  assign \new_[2951]_  = \new_[2950]_  & \new_[2945]_ ;
  assign \new_[2954]_  = ~A298 & A203;
  assign \new_[2958]_  = A302 & A300;
  assign \new_[2959]_  = A299 & \new_[2958]_ ;
  assign \new_[2960]_  = \new_[2959]_  & \new_[2954]_ ;
  assign \new_[2963]_  = A168 & ~A170;
  assign \new_[2967]_  = ~A201 & ~A166;
  assign \new_[2968]_  = A167 & \new_[2967]_ ;
  assign \new_[2969]_  = \new_[2968]_  & \new_[2963]_ ;
  assign \new_[2972]_  = A298 & A202;
  assign \new_[2976]_  = A301 & A300;
  assign \new_[2977]_  = ~A299 & \new_[2976]_ ;
  assign \new_[2978]_  = \new_[2977]_  & \new_[2972]_ ;
  assign \new_[2981]_  = A168 & ~A170;
  assign \new_[2985]_  = ~A201 & ~A166;
  assign \new_[2986]_  = A167 & \new_[2985]_ ;
  assign \new_[2987]_  = \new_[2986]_  & \new_[2981]_ ;
  assign \new_[2990]_  = A298 & A202;
  assign \new_[2994]_  = A302 & A300;
  assign \new_[2995]_  = ~A299 & \new_[2994]_ ;
  assign \new_[2996]_  = \new_[2995]_  & \new_[2990]_ ;
  assign \new_[2999]_  = A168 & ~A170;
  assign \new_[3003]_  = ~A201 & ~A166;
  assign \new_[3004]_  = A167 & \new_[3003]_ ;
  assign \new_[3005]_  = \new_[3004]_  & \new_[2999]_ ;
  assign \new_[3008]_  = ~A298 & A202;
  assign \new_[3012]_  = A301 & A300;
  assign \new_[3013]_  = A299 & \new_[3012]_ ;
  assign \new_[3014]_  = \new_[3013]_  & \new_[3008]_ ;
  assign \new_[3017]_  = A168 & ~A170;
  assign \new_[3021]_  = ~A201 & ~A166;
  assign \new_[3022]_  = A167 & \new_[3021]_ ;
  assign \new_[3023]_  = \new_[3022]_  & \new_[3017]_ ;
  assign \new_[3026]_  = ~A298 & A202;
  assign \new_[3030]_  = A302 & A300;
  assign \new_[3031]_  = A299 & \new_[3030]_ ;
  assign \new_[3032]_  = \new_[3031]_  & \new_[3026]_ ;
  assign \new_[3035]_  = A168 & ~A170;
  assign \new_[3039]_  = ~A201 & ~A166;
  assign \new_[3040]_  = A167 & \new_[3039]_ ;
  assign \new_[3041]_  = \new_[3040]_  & \new_[3035]_ ;
  assign \new_[3044]_  = A298 & A203;
  assign \new_[3048]_  = A301 & A300;
  assign \new_[3049]_  = ~A299 & \new_[3048]_ ;
  assign \new_[3050]_  = \new_[3049]_  & \new_[3044]_ ;
  assign \new_[3053]_  = A168 & ~A170;
  assign \new_[3057]_  = ~A201 & ~A166;
  assign \new_[3058]_  = A167 & \new_[3057]_ ;
  assign \new_[3059]_  = \new_[3058]_  & \new_[3053]_ ;
  assign \new_[3062]_  = A298 & A203;
  assign \new_[3066]_  = A302 & A300;
  assign \new_[3067]_  = ~A299 & \new_[3066]_ ;
  assign \new_[3068]_  = \new_[3067]_  & \new_[3062]_ ;
  assign \new_[3071]_  = A168 & ~A170;
  assign \new_[3075]_  = ~A201 & ~A166;
  assign \new_[3076]_  = A167 & \new_[3075]_ ;
  assign \new_[3077]_  = \new_[3076]_  & \new_[3071]_ ;
  assign \new_[3080]_  = ~A298 & A203;
  assign \new_[3084]_  = A301 & A300;
  assign \new_[3085]_  = A299 & \new_[3084]_ ;
  assign \new_[3086]_  = \new_[3085]_  & \new_[3080]_ ;
  assign \new_[3089]_  = A168 & ~A170;
  assign \new_[3093]_  = ~A201 & ~A166;
  assign \new_[3094]_  = A167 & \new_[3093]_ ;
  assign \new_[3095]_  = \new_[3094]_  & \new_[3089]_ ;
  assign \new_[3098]_  = ~A298 & A203;
  assign \new_[3102]_  = A302 & A300;
  assign \new_[3103]_  = A299 & \new_[3102]_ ;
  assign \new_[3104]_  = \new_[3103]_  & \new_[3098]_ ;
  assign \new_[3107]_  = A168 & ~A170;
  assign \new_[3111]_  = A199 & ~A166;
  assign \new_[3112]_  = A167 & \new_[3111]_ ;
  assign \new_[3113]_  = \new_[3112]_  & \new_[3107]_ ;
  assign \new_[3116]_  = A298 & A200;
  assign \new_[3120]_  = A301 & A300;
  assign \new_[3121]_  = ~A299 & \new_[3120]_ ;
  assign \new_[3122]_  = \new_[3121]_  & \new_[3116]_ ;
  assign \new_[3125]_  = A168 & ~A170;
  assign \new_[3129]_  = A199 & ~A166;
  assign \new_[3130]_  = A167 & \new_[3129]_ ;
  assign \new_[3131]_  = \new_[3130]_  & \new_[3125]_ ;
  assign \new_[3134]_  = A298 & A200;
  assign \new_[3138]_  = A302 & A300;
  assign \new_[3139]_  = ~A299 & \new_[3138]_ ;
  assign \new_[3140]_  = \new_[3139]_  & \new_[3134]_ ;
  assign \new_[3143]_  = A168 & ~A170;
  assign \new_[3147]_  = A199 & ~A166;
  assign \new_[3148]_  = A167 & \new_[3147]_ ;
  assign \new_[3149]_  = \new_[3148]_  & \new_[3143]_ ;
  assign \new_[3152]_  = ~A298 & A200;
  assign \new_[3156]_  = A301 & A300;
  assign \new_[3157]_  = A299 & \new_[3156]_ ;
  assign \new_[3158]_  = \new_[3157]_  & \new_[3152]_ ;
  assign \new_[3161]_  = A168 & ~A170;
  assign \new_[3165]_  = A199 & ~A166;
  assign \new_[3166]_  = A167 & \new_[3165]_ ;
  assign \new_[3167]_  = \new_[3166]_  & \new_[3161]_ ;
  assign \new_[3170]_  = ~A298 & A200;
  assign \new_[3174]_  = A302 & A300;
  assign \new_[3175]_  = A299 & \new_[3174]_ ;
  assign \new_[3176]_  = \new_[3175]_  & \new_[3170]_ ;
  assign \new_[3179]_  = A168 & ~A170;
  assign \new_[3183]_  = ~A199 & ~A166;
  assign \new_[3184]_  = A167 & \new_[3183]_ ;
  assign \new_[3185]_  = \new_[3184]_  & \new_[3179]_ ;
  assign \new_[3188]_  = A298 & ~A200;
  assign \new_[3192]_  = A301 & A300;
  assign \new_[3193]_  = ~A299 & \new_[3192]_ ;
  assign \new_[3194]_  = \new_[3193]_  & \new_[3188]_ ;
  assign \new_[3197]_  = A168 & ~A170;
  assign \new_[3201]_  = ~A199 & ~A166;
  assign \new_[3202]_  = A167 & \new_[3201]_ ;
  assign \new_[3203]_  = \new_[3202]_  & \new_[3197]_ ;
  assign \new_[3206]_  = A298 & ~A200;
  assign \new_[3210]_  = A302 & A300;
  assign \new_[3211]_  = ~A299 & \new_[3210]_ ;
  assign \new_[3212]_  = \new_[3211]_  & \new_[3206]_ ;
  assign \new_[3215]_  = A168 & ~A170;
  assign \new_[3219]_  = ~A199 & ~A166;
  assign \new_[3220]_  = A167 & \new_[3219]_ ;
  assign \new_[3221]_  = \new_[3220]_  & \new_[3215]_ ;
  assign \new_[3224]_  = ~A298 & ~A200;
  assign \new_[3228]_  = A301 & A300;
  assign \new_[3229]_  = A299 & \new_[3228]_ ;
  assign \new_[3230]_  = \new_[3229]_  & \new_[3224]_ ;
  assign \new_[3233]_  = A168 & ~A170;
  assign \new_[3237]_  = ~A199 & ~A166;
  assign \new_[3238]_  = A167 & \new_[3237]_ ;
  assign \new_[3239]_  = \new_[3238]_  & \new_[3233]_ ;
  assign \new_[3242]_  = ~A298 & ~A200;
  assign \new_[3246]_  = A302 & A300;
  assign \new_[3247]_  = A299 & \new_[3246]_ ;
  assign \new_[3248]_  = \new_[3247]_  & \new_[3242]_ ;
  assign \new_[3251]_  = A168 & ~A170;
  assign \new_[3255]_  = ~A201 & A166;
  assign \new_[3256]_  = ~A167 & \new_[3255]_ ;
  assign \new_[3257]_  = \new_[3256]_  & \new_[3251]_ ;
  assign \new_[3260]_  = A298 & A202;
  assign \new_[3264]_  = A301 & A300;
  assign \new_[3265]_  = ~A299 & \new_[3264]_ ;
  assign \new_[3266]_  = \new_[3265]_  & \new_[3260]_ ;
  assign \new_[3269]_  = A168 & ~A170;
  assign \new_[3273]_  = ~A201 & A166;
  assign \new_[3274]_  = ~A167 & \new_[3273]_ ;
  assign \new_[3275]_  = \new_[3274]_  & \new_[3269]_ ;
  assign \new_[3278]_  = A298 & A202;
  assign \new_[3282]_  = A302 & A300;
  assign \new_[3283]_  = ~A299 & \new_[3282]_ ;
  assign \new_[3284]_  = \new_[3283]_  & \new_[3278]_ ;
  assign \new_[3287]_  = A168 & ~A170;
  assign \new_[3291]_  = ~A201 & A166;
  assign \new_[3292]_  = ~A167 & \new_[3291]_ ;
  assign \new_[3293]_  = \new_[3292]_  & \new_[3287]_ ;
  assign \new_[3296]_  = ~A298 & A202;
  assign \new_[3300]_  = A301 & A300;
  assign \new_[3301]_  = A299 & \new_[3300]_ ;
  assign \new_[3302]_  = \new_[3301]_  & \new_[3296]_ ;
  assign \new_[3305]_  = A168 & ~A170;
  assign \new_[3309]_  = ~A201 & A166;
  assign \new_[3310]_  = ~A167 & \new_[3309]_ ;
  assign \new_[3311]_  = \new_[3310]_  & \new_[3305]_ ;
  assign \new_[3314]_  = ~A298 & A202;
  assign \new_[3318]_  = A302 & A300;
  assign \new_[3319]_  = A299 & \new_[3318]_ ;
  assign \new_[3320]_  = \new_[3319]_  & \new_[3314]_ ;
  assign \new_[3323]_  = A168 & ~A170;
  assign \new_[3327]_  = ~A201 & A166;
  assign \new_[3328]_  = ~A167 & \new_[3327]_ ;
  assign \new_[3329]_  = \new_[3328]_  & \new_[3323]_ ;
  assign \new_[3332]_  = A298 & A203;
  assign \new_[3336]_  = A301 & A300;
  assign \new_[3337]_  = ~A299 & \new_[3336]_ ;
  assign \new_[3338]_  = \new_[3337]_  & \new_[3332]_ ;
  assign \new_[3341]_  = A168 & ~A170;
  assign \new_[3345]_  = ~A201 & A166;
  assign \new_[3346]_  = ~A167 & \new_[3345]_ ;
  assign \new_[3347]_  = \new_[3346]_  & \new_[3341]_ ;
  assign \new_[3350]_  = A298 & A203;
  assign \new_[3354]_  = A302 & A300;
  assign \new_[3355]_  = ~A299 & \new_[3354]_ ;
  assign \new_[3356]_  = \new_[3355]_  & \new_[3350]_ ;
  assign \new_[3359]_  = A168 & ~A170;
  assign \new_[3363]_  = ~A201 & A166;
  assign \new_[3364]_  = ~A167 & \new_[3363]_ ;
  assign \new_[3365]_  = \new_[3364]_  & \new_[3359]_ ;
  assign \new_[3368]_  = ~A298 & A203;
  assign \new_[3372]_  = A301 & A300;
  assign \new_[3373]_  = A299 & \new_[3372]_ ;
  assign \new_[3374]_  = \new_[3373]_  & \new_[3368]_ ;
  assign \new_[3377]_  = A168 & ~A170;
  assign \new_[3381]_  = ~A201 & A166;
  assign \new_[3382]_  = ~A167 & \new_[3381]_ ;
  assign \new_[3383]_  = \new_[3382]_  & \new_[3377]_ ;
  assign \new_[3386]_  = ~A298 & A203;
  assign \new_[3390]_  = A302 & A300;
  assign \new_[3391]_  = A299 & \new_[3390]_ ;
  assign \new_[3392]_  = \new_[3391]_  & \new_[3386]_ ;
  assign \new_[3395]_  = A168 & ~A170;
  assign \new_[3399]_  = A199 & A166;
  assign \new_[3400]_  = ~A167 & \new_[3399]_ ;
  assign \new_[3401]_  = \new_[3400]_  & \new_[3395]_ ;
  assign \new_[3404]_  = A298 & A200;
  assign \new_[3408]_  = A301 & A300;
  assign \new_[3409]_  = ~A299 & \new_[3408]_ ;
  assign \new_[3410]_  = \new_[3409]_  & \new_[3404]_ ;
  assign \new_[3413]_  = A168 & ~A170;
  assign \new_[3417]_  = A199 & A166;
  assign \new_[3418]_  = ~A167 & \new_[3417]_ ;
  assign \new_[3419]_  = \new_[3418]_  & \new_[3413]_ ;
  assign \new_[3422]_  = A298 & A200;
  assign \new_[3426]_  = A302 & A300;
  assign \new_[3427]_  = ~A299 & \new_[3426]_ ;
  assign \new_[3428]_  = \new_[3427]_  & \new_[3422]_ ;
  assign \new_[3431]_  = A168 & ~A170;
  assign \new_[3435]_  = A199 & A166;
  assign \new_[3436]_  = ~A167 & \new_[3435]_ ;
  assign \new_[3437]_  = \new_[3436]_  & \new_[3431]_ ;
  assign \new_[3440]_  = ~A298 & A200;
  assign \new_[3444]_  = A301 & A300;
  assign \new_[3445]_  = A299 & \new_[3444]_ ;
  assign \new_[3446]_  = \new_[3445]_  & \new_[3440]_ ;
  assign \new_[3449]_  = A168 & ~A170;
  assign \new_[3453]_  = A199 & A166;
  assign \new_[3454]_  = ~A167 & \new_[3453]_ ;
  assign \new_[3455]_  = \new_[3454]_  & \new_[3449]_ ;
  assign \new_[3458]_  = ~A298 & A200;
  assign \new_[3462]_  = A302 & A300;
  assign \new_[3463]_  = A299 & \new_[3462]_ ;
  assign \new_[3464]_  = \new_[3463]_  & \new_[3458]_ ;
  assign \new_[3467]_  = A168 & ~A170;
  assign \new_[3471]_  = ~A199 & A166;
  assign \new_[3472]_  = ~A167 & \new_[3471]_ ;
  assign \new_[3473]_  = \new_[3472]_  & \new_[3467]_ ;
  assign \new_[3476]_  = A298 & ~A200;
  assign \new_[3480]_  = A301 & A300;
  assign \new_[3481]_  = ~A299 & \new_[3480]_ ;
  assign \new_[3482]_  = \new_[3481]_  & \new_[3476]_ ;
  assign \new_[3485]_  = A168 & ~A170;
  assign \new_[3489]_  = ~A199 & A166;
  assign \new_[3490]_  = ~A167 & \new_[3489]_ ;
  assign \new_[3491]_  = \new_[3490]_  & \new_[3485]_ ;
  assign \new_[3494]_  = A298 & ~A200;
  assign \new_[3498]_  = A302 & A300;
  assign \new_[3499]_  = ~A299 & \new_[3498]_ ;
  assign \new_[3500]_  = \new_[3499]_  & \new_[3494]_ ;
  assign \new_[3503]_  = A168 & ~A170;
  assign \new_[3507]_  = ~A199 & A166;
  assign \new_[3508]_  = ~A167 & \new_[3507]_ ;
  assign \new_[3509]_  = \new_[3508]_  & \new_[3503]_ ;
  assign \new_[3512]_  = ~A298 & ~A200;
  assign \new_[3516]_  = A301 & A300;
  assign \new_[3517]_  = A299 & \new_[3516]_ ;
  assign \new_[3518]_  = \new_[3517]_  & \new_[3512]_ ;
  assign \new_[3521]_  = A168 & ~A170;
  assign \new_[3525]_  = ~A199 & A166;
  assign \new_[3526]_  = ~A167 & \new_[3525]_ ;
  assign \new_[3527]_  = \new_[3526]_  & \new_[3521]_ ;
  assign \new_[3530]_  = ~A298 & ~A200;
  assign \new_[3534]_  = A302 & A300;
  assign \new_[3535]_  = A299 & \new_[3534]_ ;
  assign \new_[3536]_  = \new_[3535]_  & \new_[3530]_ ;
  assign \new_[3539]_  = ~A168 & ~A170;
  assign \new_[3543]_  = A201 & A200;
  assign \new_[3544]_  = ~A199 & \new_[3543]_ ;
  assign \new_[3545]_  = \new_[3544]_  & \new_[3539]_ ;
  assign \new_[3548]_  = A298 & A202;
  assign \new_[3552]_  = A301 & A300;
  assign \new_[3553]_  = ~A299 & \new_[3552]_ ;
  assign \new_[3554]_  = \new_[3553]_  & \new_[3548]_ ;
  assign \new_[3557]_  = ~A168 & ~A170;
  assign \new_[3561]_  = A201 & A200;
  assign \new_[3562]_  = ~A199 & \new_[3561]_ ;
  assign \new_[3563]_  = \new_[3562]_  & \new_[3557]_ ;
  assign \new_[3566]_  = A298 & A202;
  assign \new_[3570]_  = A302 & A300;
  assign \new_[3571]_  = ~A299 & \new_[3570]_ ;
  assign \new_[3572]_  = \new_[3571]_  & \new_[3566]_ ;
  assign \new_[3575]_  = ~A168 & ~A170;
  assign \new_[3579]_  = A201 & A200;
  assign \new_[3580]_  = ~A199 & \new_[3579]_ ;
  assign \new_[3581]_  = \new_[3580]_  & \new_[3575]_ ;
  assign \new_[3584]_  = ~A298 & A202;
  assign \new_[3588]_  = A301 & A300;
  assign \new_[3589]_  = A299 & \new_[3588]_ ;
  assign \new_[3590]_  = \new_[3589]_  & \new_[3584]_ ;
  assign \new_[3593]_  = ~A168 & ~A170;
  assign \new_[3597]_  = A201 & A200;
  assign \new_[3598]_  = ~A199 & \new_[3597]_ ;
  assign \new_[3599]_  = \new_[3598]_  & \new_[3593]_ ;
  assign \new_[3602]_  = ~A298 & A202;
  assign \new_[3606]_  = A302 & A300;
  assign \new_[3607]_  = A299 & \new_[3606]_ ;
  assign \new_[3608]_  = \new_[3607]_  & \new_[3602]_ ;
  assign \new_[3611]_  = ~A168 & ~A170;
  assign \new_[3615]_  = A201 & A200;
  assign \new_[3616]_  = ~A199 & \new_[3615]_ ;
  assign \new_[3617]_  = \new_[3616]_  & \new_[3611]_ ;
  assign \new_[3620]_  = A298 & A203;
  assign \new_[3624]_  = A301 & A300;
  assign \new_[3625]_  = ~A299 & \new_[3624]_ ;
  assign \new_[3626]_  = \new_[3625]_  & \new_[3620]_ ;
  assign \new_[3629]_  = ~A168 & ~A170;
  assign \new_[3633]_  = A201 & A200;
  assign \new_[3634]_  = ~A199 & \new_[3633]_ ;
  assign \new_[3635]_  = \new_[3634]_  & \new_[3629]_ ;
  assign \new_[3638]_  = A298 & A203;
  assign \new_[3642]_  = A302 & A300;
  assign \new_[3643]_  = ~A299 & \new_[3642]_ ;
  assign \new_[3644]_  = \new_[3643]_  & \new_[3638]_ ;
  assign \new_[3647]_  = ~A168 & ~A170;
  assign \new_[3651]_  = A201 & A200;
  assign \new_[3652]_  = ~A199 & \new_[3651]_ ;
  assign \new_[3653]_  = \new_[3652]_  & \new_[3647]_ ;
  assign \new_[3656]_  = ~A298 & A203;
  assign \new_[3660]_  = A301 & A300;
  assign \new_[3661]_  = A299 & \new_[3660]_ ;
  assign \new_[3662]_  = \new_[3661]_  & \new_[3656]_ ;
  assign \new_[3665]_  = ~A168 & ~A170;
  assign \new_[3669]_  = A201 & A200;
  assign \new_[3670]_  = ~A199 & \new_[3669]_ ;
  assign \new_[3671]_  = \new_[3670]_  & \new_[3665]_ ;
  assign \new_[3674]_  = ~A298 & A203;
  assign \new_[3678]_  = A302 & A300;
  assign \new_[3679]_  = A299 & \new_[3678]_ ;
  assign \new_[3680]_  = \new_[3679]_  & \new_[3674]_ ;
  assign \new_[3683]_  = ~A168 & ~A170;
  assign \new_[3687]_  = A201 & ~A200;
  assign \new_[3688]_  = A199 & \new_[3687]_ ;
  assign \new_[3689]_  = \new_[3688]_  & \new_[3683]_ ;
  assign \new_[3692]_  = A298 & A202;
  assign \new_[3696]_  = A301 & A300;
  assign \new_[3697]_  = ~A299 & \new_[3696]_ ;
  assign \new_[3698]_  = \new_[3697]_  & \new_[3692]_ ;
  assign \new_[3701]_  = ~A168 & ~A170;
  assign \new_[3705]_  = A201 & ~A200;
  assign \new_[3706]_  = A199 & \new_[3705]_ ;
  assign \new_[3707]_  = \new_[3706]_  & \new_[3701]_ ;
  assign \new_[3710]_  = A298 & A202;
  assign \new_[3714]_  = A302 & A300;
  assign \new_[3715]_  = ~A299 & \new_[3714]_ ;
  assign \new_[3716]_  = \new_[3715]_  & \new_[3710]_ ;
  assign \new_[3719]_  = ~A168 & ~A170;
  assign \new_[3723]_  = A201 & ~A200;
  assign \new_[3724]_  = A199 & \new_[3723]_ ;
  assign \new_[3725]_  = \new_[3724]_  & \new_[3719]_ ;
  assign \new_[3728]_  = ~A298 & A202;
  assign \new_[3732]_  = A301 & A300;
  assign \new_[3733]_  = A299 & \new_[3732]_ ;
  assign \new_[3734]_  = \new_[3733]_  & \new_[3728]_ ;
  assign \new_[3737]_  = ~A168 & ~A170;
  assign \new_[3741]_  = A201 & ~A200;
  assign \new_[3742]_  = A199 & \new_[3741]_ ;
  assign \new_[3743]_  = \new_[3742]_  & \new_[3737]_ ;
  assign \new_[3746]_  = ~A298 & A202;
  assign \new_[3750]_  = A302 & A300;
  assign \new_[3751]_  = A299 & \new_[3750]_ ;
  assign \new_[3752]_  = \new_[3751]_  & \new_[3746]_ ;
  assign \new_[3755]_  = ~A168 & ~A170;
  assign \new_[3759]_  = A201 & ~A200;
  assign \new_[3760]_  = A199 & \new_[3759]_ ;
  assign \new_[3761]_  = \new_[3760]_  & \new_[3755]_ ;
  assign \new_[3764]_  = A298 & A203;
  assign \new_[3768]_  = A301 & A300;
  assign \new_[3769]_  = ~A299 & \new_[3768]_ ;
  assign \new_[3770]_  = \new_[3769]_  & \new_[3764]_ ;
  assign \new_[3773]_  = ~A168 & ~A170;
  assign \new_[3777]_  = A201 & ~A200;
  assign \new_[3778]_  = A199 & \new_[3777]_ ;
  assign \new_[3779]_  = \new_[3778]_  & \new_[3773]_ ;
  assign \new_[3782]_  = A298 & A203;
  assign \new_[3786]_  = A302 & A300;
  assign \new_[3787]_  = ~A299 & \new_[3786]_ ;
  assign \new_[3788]_  = \new_[3787]_  & \new_[3782]_ ;
  assign \new_[3791]_  = ~A168 & ~A170;
  assign \new_[3795]_  = A201 & ~A200;
  assign \new_[3796]_  = A199 & \new_[3795]_ ;
  assign \new_[3797]_  = \new_[3796]_  & \new_[3791]_ ;
  assign \new_[3800]_  = ~A298 & A203;
  assign \new_[3804]_  = A301 & A300;
  assign \new_[3805]_  = A299 & \new_[3804]_ ;
  assign \new_[3806]_  = \new_[3805]_  & \new_[3800]_ ;
  assign \new_[3809]_  = ~A168 & ~A170;
  assign \new_[3813]_  = A201 & ~A200;
  assign \new_[3814]_  = A199 & \new_[3813]_ ;
  assign \new_[3815]_  = \new_[3814]_  & \new_[3809]_ ;
  assign \new_[3818]_  = ~A298 & A203;
  assign \new_[3822]_  = A302 & A300;
  assign \new_[3823]_  = A299 & \new_[3822]_ ;
  assign \new_[3824]_  = \new_[3823]_  & \new_[3818]_ ;
  assign \new_[3827]_  = A168 & A169;
  assign \new_[3831]_  = ~A201 & ~A166;
  assign \new_[3832]_  = A167 & \new_[3831]_ ;
  assign \new_[3833]_  = \new_[3832]_  & \new_[3827]_ ;
  assign \new_[3836]_  = A298 & A202;
  assign \new_[3840]_  = A301 & A300;
  assign \new_[3841]_  = ~A299 & \new_[3840]_ ;
  assign \new_[3842]_  = \new_[3841]_  & \new_[3836]_ ;
  assign \new_[3845]_  = A168 & A169;
  assign \new_[3849]_  = ~A201 & ~A166;
  assign \new_[3850]_  = A167 & \new_[3849]_ ;
  assign \new_[3851]_  = \new_[3850]_  & \new_[3845]_ ;
  assign \new_[3854]_  = A298 & A202;
  assign \new_[3858]_  = A302 & A300;
  assign \new_[3859]_  = ~A299 & \new_[3858]_ ;
  assign \new_[3860]_  = \new_[3859]_  & \new_[3854]_ ;
  assign \new_[3863]_  = A168 & A169;
  assign \new_[3867]_  = ~A201 & ~A166;
  assign \new_[3868]_  = A167 & \new_[3867]_ ;
  assign \new_[3869]_  = \new_[3868]_  & \new_[3863]_ ;
  assign \new_[3872]_  = ~A298 & A202;
  assign \new_[3876]_  = A301 & A300;
  assign \new_[3877]_  = A299 & \new_[3876]_ ;
  assign \new_[3878]_  = \new_[3877]_  & \new_[3872]_ ;
  assign \new_[3881]_  = A168 & A169;
  assign \new_[3885]_  = ~A201 & ~A166;
  assign \new_[3886]_  = A167 & \new_[3885]_ ;
  assign \new_[3887]_  = \new_[3886]_  & \new_[3881]_ ;
  assign \new_[3890]_  = ~A298 & A202;
  assign \new_[3894]_  = A302 & A300;
  assign \new_[3895]_  = A299 & \new_[3894]_ ;
  assign \new_[3896]_  = \new_[3895]_  & \new_[3890]_ ;
  assign \new_[3899]_  = A168 & A169;
  assign \new_[3903]_  = ~A201 & ~A166;
  assign \new_[3904]_  = A167 & \new_[3903]_ ;
  assign \new_[3905]_  = \new_[3904]_  & \new_[3899]_ ;
  assign \new_[3908]_  = A298 & A203;
  assign \new_[3912]_  = A301 & A300;
  assign \new_[3913]_  = ~A299 & \new_[3912]_ ;
  assign \new_[3914]_  = \new_[3913]_  & \new_[3908]_ ;
  assign \new_[3917]_  = A168 & A169;
  assign \new_[3921]_  = ~A201 & ~A166;
  assign \new_[3922]_  = A167 & \new_[3921]_ ;
  assign \new_[3923]_  = \new_[3922]_  & \new_[3917]_ ;
  assign \new_[3926]_  = A298 & A203;
  assign \new_[3930]_  = A302 & A300;
  assign \new_[3931]_  = ~A299 & \new_[3930]_ ;
  assign \new_[3932]_  = \new_[3931]_  & \new_[3926]_ ;
  assign \new_[3935]_  = A168 & A169;
  assign \new_[3939]_  = ~A201 & ~A166;
  assign \new_[3940]_  = A167 & \new_[3939]_ ;
  assign \new_[3941]_  = \new_[3940]_  & \new_[3935]_ ;
  assign \new_[3944]_  = ~A298 & A203;
  assign \new_[3948]_  = A301 & A300;
  assign \new_[3949]_  = A299 & \new_[3948]_ ;
  assign \new_[3950]_  = \new_[3949]_  & \new_[3944]_ ;
  assign \new_[3953]_  = A168 & A169;
  assign \new_[3957]_  = ~A201 & ~A166;
  assign \new_[3958]_  = A167 & \new_[3957]_ ;
  assign \new_[3959]_  = \new_[3958]_  & \new_[3953]_ ;
  assign \new_[3962]_  = ~A298 & A203;
  assign \new_[3966]_  = A302 & A300;
  assign \new_[3967]_  = A299 & \new_[3966]_ ;
  assign \new_[3968]_  = \new_[3967]_  & \new_[3962]_ ;
  assign \new_[3971]_  = A168 & A169;
  assign \new_[3975]_  = A199 & ~A166;
  assign \new_[3976]_  = A167 & \new_[3975]_ ;
  assign \new_[3977]_  = \new_[3976]_  & \new_[3971]_ ;
  assign \new_[3980]_  = A298 & A200;
  assign \new_[3984]_  = A301 & A300;
  assign \new_[3985]_  = ~A299 & \new_[3984]_ ;
  assign \new_[3986]_  = \new_[3985]_  & \new_[3980]_ ;
  assign \new_[3989]_  = A168 & A169;
  assign \new_[3993]_  = A199 & ~A166;
  assign \new_[3994]_  = A167 & \new_[3993]_ ;
  assign \new_[3995]_  = \new_[3994]_  & \new_[3989]_ ;
  assign \new_[3998]_  = A298 & A200;
  assign \new_[4002]_  = A302 & A300;
  assign \new_[4003]_  = ~A299 & \new_[4002]_ ;
  assign \new_[4004]_  = \new_[4003]_  & \new_[3998]_ ;
  assign \new_[4007]_  = A168 & A169;
  assign \new_[4011]_  = A199 & ~A166;
  assign \new_[4012]_  = A167 & \new_[4011]_ ;
  assign \new_[4013]_  = \new_[4012]_  & \new_[4007]_ ;
  assign \new_[4016]_  = ~A298 & A200;
  assign \new_[4020]_  = A301 & A300;
  assign \new_[4021]_  = A299 & \new_[4020]_ ;
  assign \new_[4022]_  = \new_[4021]_  & \new_[4016]_ ;
  assign \new_[4025]_  = A168 & A169;
  assign \new_[4029]_  = A199 & ~A166;
  assign \new_[4030]_  = A167 & \new_[4029]_ ;
  assign \new_[4031]_  = \new_[4030]_  & \new_[4025]_ ;
  assign \new_[4034]_  = ~A298 & A200;
  assign \new_[4038]_  = A302 & A300;
  assign \new_[4039]_  = A299 & \new_[4038]_ ;
  assign \new_[4040]_  = \new_[4039]_  & \new_[4034]_ ;
  assign \new_[4043]_  = A168 & A169;
  assign \new_[4047]_  = ~A199 & ~A166;
  assign \new_[4048]_  = A167 & \new_[4047]_ ;
  assign \new_[4049]_  = \new_[4048]_  & \new_[4043]_ ;
  assign \new_[4052]_  = A298 & ~A200;
  assign \new_[4056]_  = A301 & A300;
  assign \new_[4057]_  = ~A299 & \new_[4056]_ ;
  assign \new_[4058]_  = \new_[4057]_  & \new_[4052]_ ;
  assign \new_[4061]_  = A168 & A169;
  assign \new_[4065]_  = ~A199 & ~A166;
  assign \new_[4066]_  = A167 & \new_[4065]_ ;
  assign \new_[4067]_  = \new_[4066]_  & \new_[4061]_ ;
  assign \new_[4070]_  = A298 & ~A200;
  assign \new_[4074]_  = A302 & A300;
  assign \new_[4075]_  = ~A299 & \new_[4074]_ ;
  assign \new_[4076]_  = \new_[4075]_  & \new_[4070]_ ;
  assign \new_[4079]_  = A168 & A169;
  assign \new_[4083]_  = ~A199 & ~A166;
  assign \new_[4084]_  = A167 & \new_[4083]_ ;
  assign \new_[4085]_  = \new_[4084]_  & \new_[4079]_ ;
  assign \new_[4088]_  = ~A298 & ~A200;
  assign \new_[4092]_  = A301 & A300;
  assign \new_[4093]_  = A299 & \new_[4092]_ ;
  assign \new_[4094]_  = \new_[4093]_  & \new_[4088]_ ;
  assign \new_[4097]_  = A168 & A169;
  assign \new_[4101]_  = ~A199 & ~A166;
  assign \new_[4102]_  = A167 & \new_[4101]_ ;
  assign \new_[4103]_  = \new_[4102]_  & \new_[4097]_ ;
  assign \new_[4106]_  = ~A298 & ~A200;
  assign \new_[4110]_  = A302 & A300;
  assign \new_[4111]_  = A299 & \new_[4110]_ ;
  assign \new_[4112]_  = \new_[4111]_  & \new_[4106]_ ;
  assign \new_[4115]_  = A168 & A169;
  assign \new_[4119]_  = ~A201 & A166;
  assign \new_[4120]_  = ~A167 & \new_[4119]_ ;
  assign \new_[4121]_  = \new_[4120]_  & \new_[4115]_ ;
  assign \new_[4124]_  = A298 & A202;
  assign \new_[4128]_  = A301 & A300;
  assign \new_[4129]_  = ~A299 & \new_[4128]_ ;
  assign \new_[4130]_  = \new_[4129]_  & \new_[4124]_ ;
  assign \new_[4133]_  = A168 & A169;
  assign \new_[4137]_  = ~A201 & A166;
  assign \new_[4138]_  = ~A167 & \new_[4137]_ ;
  assign \new_[4139]_  = \new_[4138]_  & \new_[4133]_ ;
  assign \new_[4142]_  = A298 & A202;
  assign \new_[4146]_  = A302 & A300;
  assign \new_[4147]_  = ~A299 & \new_[4146]_ ;
  assign \new_[4148]_  = \new_[4147]_  & \new_[4142]_ ;
  assign \new_[4151]_  = A168 & A169;
  assign \new_[4155]_  = ~A201 & A166;
  assign \new_[4156]_  = ~A167 & \new_[4155]_ ;
  assign \new_[4157]_  = \new_[4156]_  & \new_[4151]_ ;
  assign \new_[4160]_  = ~A298 & A202;
  assign \new_[4164]_  = A301 & A300;
  assign \new_[4165]_  = A299 & \new_[4164]_ ;
  assign \new_[4166]_  = \new_[4165]_  & \new_[4160]_ ;
  assign \new_[4169]_  = A168 & A169;
  assign \new_[4173]_  = ~A201 & A166;
  assign \new_[4174]_  = ~A167 & \new_[4173]_ ;
  assign \new_[4175]_  = \new_[4174]_  & \new_[4169]_ ;
  assign \new_[4178]_  = ~A298 & A202;
  assign \new_[4182]_  = A302 & A300;
  assign \new_[4183]_  = A299 & \new_[4182]_ ;
  assign \new_[4184]_  = \new_[4183]_  & \new_[4178]_ ;
  assign \new_[4187]_  = A168 & A169;
  assign \new_[4191]_  = ~A201 & A166;
  assign \new_[4192]_  = ~A167 & \new_[4191]_ ;
  assign \new_[4193]_  = \new_[4192]_  & \new_[4187]_ ;
  assign \new_[4196]_  = A298 & A203;
  assign \new_[4200]_  = A301 & A300;
  assign \new_[4201]_  = ~A299 & \new_[4200]_ ;
  assign \new_[4202]_  = \new_[4201]_  & \new_[4196]_ ;
  assign \new_[4205]_  = A168 & A169;
  assign \new_[4209]_  = ~A201 & A166;
  assign \new_[4210]_  = ~A167 & \new_[4209]_ ;
  assign \new_[4211]_  = \new_[4210]_  & \new_[4205]_ ;
  assign \new_[4214]_  = A298 & A203;
  assign \new_[4218]_  = A302 & A300;
  assign \new_[4219]_  = ~A299 & \new_[4218]_ ;
  assign \new_[4220]_  = \new_[4219]_  & \new_[4214]_ ;
  assign \new_[4223]_  = A168 & A169;
  assign \new_[4227]_  = ~A201 & A166;
  assign \new_[4228]_  = ~A167 & \new_[4227]_ ;
  assign \new_[4229]_  = \new_[4228]_  & \new_[4223]_ ;
  assign \new_[4232]_  = ~A298 & A203;
  assign \new_[4236]_  = A301 & A300;
  assign \new_[4237]_  = A299 & \new_[4236]_ ;
  assign \new_[4238]_  = \new_[4237]_  & \new_[4232]_ ;
  assign \new_[4241]_  = A168 & A169;
  assign \new_[4245]_  = ~A201 & A166;
  assign \new_[4246]_  = ~A167 & \new_[4245]_ ;
  assign \new_[4247]_  = \new_[4246]_  & \new_[4241]_ ;
  assign \new_[4250]_  = ~A298 & A203;
  assign \new_[4254]_  = A302 & A300;
  assign \new_[4255]_  = A299 & \new_[4254]_ ;
  assign \new_[4256]_  = \new_[4255]_  & \new_[4250]_ ;
  assign \new_[4259]_  = A168 & A169;
  assign \new_[4263]_  = A199 & A166;
  assign \new_[4264]_  = ~A167 & \new_[4263]_ ;
  assign \new_[4265]_  = \new_[4264]_  & \new_[4259]_ ;
  assign \new_[4268]_  = A298 & A200;
  assign \new_[4272]_  = A301 & A300;
  assign \new_[4273]_  = ~A299 & \new_[4272]_ ;
  assign \new_[4274]_  = \new_[4273]_  & \new_[4268]_ ;
  assign \new_[4277]_  = A168 & A169;
  assign \new_[4281]_  = A199 & A166;
  assign \new_[4282]_  = ~A167 & \new_[4281]_ ;
  assign \new_[4283]_  = \new_[4282]_  & \new_[4277]_ ;
  assign \new_[4286]_  = A298 & A200;
  assign \new_[4290]_  = A302 & A300;
  assign \new_[4291]_  = ~A299 & \new_[4290]_ ;
  assign \new_[4292]_  = \new_[4291]_  & \new_[4286]_ ;
  assign \new_[4295]_  = A168 & A169;
  assign \new_[4299]_  = A199 & A166;
  assign \new_[4300]_  = ~A167 & \new_[4299]_ ;
  assign \new_[4301]_  = \new_[4300]_  & \new_[4295]_ ;
  assign \new_[4304]_  = ~A298 & A200;
  assign \new_[4308]_  = A301 & A300;
  assign \new_[4309]_  = A299 & \new_[4308]_ ;
  assign \new_[4310]_  = \new_[4309]_  & \new_[4304]_ ;
  assign \new_[4313]_  = A168 & A169;
  assign \new_[4317]_  = A199 & A166;
  assign \new_[4318]_  = ~A167 & \new_[4317]_ ;
  assign \new_[4319]_  = \new_[4318]_  & \new_[4313]_ ;
  assign \new_[4322]_  = ~A298 & A200;
  assign \new_[4326]_  = A302 & A300;
  assign \new_[4327]_  = A299 & \new_[4326]_ ;
  assign \new_[4328]_  = \new_[4327]_  & \new_[4322]_ ;
  assign \new_[4331]_  = A168 & A169;
  assign \new_[4335]_  = ~A199 & A166;
  assign \new_[4336]_  = ~A167 & \new_[4335]_ ;
  assign \new_[4337]_  = \new_[4336]_  & \new_[4331]_ ;
  assign \new_[4340]_  = A298 & ~A200;
  assign \new_[4344]_  = A301 & A300;
  assign \new_[4345]_  = ~A299 & \new_[4344]_ ;
  assign \new_[4346]_  = \new_[4345]_  & \new_[4340]_ ;
  assign \new_[4349]_  = A168 & A169;
  assign \new_[4353]_  = ~A199 & A166;
  assign \new_[4354]_  = ~A167 & \new_[4353]_ ;
  assign \new_[4355]_  = \new_[4354]_  & \new_[4349]_ ;
  assign \new_[4358]_  = A298 & ~A200;
  assign \new_[4362]_  = A302 & A300;
  assign \new_[4363]_  = ~A299 & \new_[4362]_ ;
  assign \new_[4364]_  = \new_[4363]_  & \new_[4358]_ ;
  assign \new_[4367]_  = A168 & A169;
  assign \new_[4371]_  = ~A199 & A166;
  assign \new_[4372]_  = ~A167 & \new_[4371]_ ;
  assign \new_[4373]_  = \new_[4372]_  & \new_[4367]_ ;
  assign \new_[4376]_  = ~A298 & ~A200;
  assign \new_[4380]_  = A301 & A300;
  assign \new_[4381]_  = A299 & \new_[4380]_ ;
  assign \new_[4382]_  = \new_[4381]_  & \new_[4376]_ ;
  assign \new_[4385]_  = A168 & A169;
  assign \new_[4389]_  = ~A199 & A166;
  assign \new_[4390]_  = ~A167 & \new_[4389]_ ;
  assign \new_[4391]_  = \new_[4390]_  & \new_[4385]_ ;
  assign \new_[4394]_  = ~A298 & ~A200;
  assign \new_[4398]_  = A302 & A300;
  assign \new_[4399]_  = A299 & \new_[4398]_ ;
  assign \new_[4400]_  = \new_[4399]_  & \new_[4394]_ ;
  assign \new_[4403]_  = ~A168 & A169;
  assign \new_[4407]_  = A201 & A200;
  assign \new_[4408]_  = ~A199 & \new_[4407]_ ;
  assign \new_[4409]_  = \new_[4408]_  & \new_[4403]_ ;
  assign \new_[4412]_  = A298 & A202;
  assign \new_[4416]_  = A301 & A300;
  assign \new_[4417]_  = ~A299 & \new_[4416]_ ;
  assign \new_[4418]_  = \new_[4417]_  & \new_[4412]_ ;
  assign \new_[4421]_  = ~A168 & A169;
  assign \new_[4425]_  = A201 & A200;
  assign \new_[4426]_  = ~A199 & \new_[4425]_ ;
  assign \new_[4427]_  = \new_[4426]_  & \new_[4421]_ ;
  assign \new_[4430]_  = A298 & A202;
  assign \new_[4434]_  = A302 & A300;
  assign \new_[4435]_  = ~A299 & \new_[4434]_ ;
  assign \new_[4436]_  = \new_[4435]_  & \new_[4430]_ ;
  assign \new_[4439]_  = ~A168 & A169;
  assign \new_[4443]_  = A201 & A200;
  assign \new_[4444]_  = ~A199 & \new_[4443]_ ;
  assign \new_[4445]_  = \new_[4444]_  & \new_[4439]_ ;
  assign \new_[4448]_  = ~A298 & A202;
  assign \new_[4452]_  = A301 & A300;
  assign \new_[4453]_  = A299 & \new_[4452]_ ;
  assign \new_[4454]_  = \new_[4453]_  & \new_[4448]_ ;
  assign \new_[4457]_  = ~A168 & A169;
  assign \new_[4461]_  = A201 & A200;
  assign \new_[4462]_  = ~A199 & \new_[4461]_ ;
  assign \new_[4463]_  = \new_[4462]_  & \new_[4457]_ ;
  assign \new_[4466]_  = ~A298 & A202;
  assign \new_[4470]_  = A302 & A300;
  assign \new_[4471]_  = A299 & \new_[4470]_ ;
  assign \new_[4472]_  = \new_[4471]_  & \new_[4466]_ ;
  assign \new_[4475]_  = ~A168 & A169;
  assign \new_[4479]_  = A201 & A200;
  assign \new_[4480]_  = ~A199 & \new_[4479]_ ;
  assign \new_[4481]_  = \new_[4480]_  & \new_[4475]_ ;
  assign \new_[4484]_  = A298 & A203;
  assign \new_[4488]_  = A301 & A300;
  assign \new_[4489]_  = ~A299 & \new_[4488]_ ;
  assign \new_[4490]_  = \new_[4489]_  & \new_[4484]_ ;
  assign \new_[4493]_  = ~A168 & A169;
  assign \new_[4497]_  = A201 & A200;
  assign \new_[4498]_  = ~A199 & \new_[4497]_ ;
  assign \new_[4499]_  = \new_[4498]_  & \new_[4493]_ ;
  assign \new_[4502]_  = A298 & A203;
  assign \new_[4506]_  = A302 & A300;
  assign \new_[4507]_  = ~A299 & \new_[4506]_ ;
  assign \new_[4508]_  = \new_[4507]_  & \new_[4502]_ ;
  assign \new_[4511]_  = ~A168 & A169;
  assign \new_[4515]_  = A201 & A200;
  assign \new_[4516]_  = ~A199 & \new_[4515]_ ;
  assign \new_[4517]_  = \new_[4516]_  & \new_[4511]_ ;
  assign \new_[4520]_  = ~A298 & A203;
  assign \new_[4524]_  = A301 & A300;
  assign \new_[4525]_  = A299 & \new_[4524]_ ;
  assign \new_[4526]_  = \new_[4525]_  & \new_[4520]_ ;
  assign \new_[4529]_  = ~A168 & A169;
  assign \new_[4533]_  = A201 & A200;
  assign \new_[4534]_  = ~A199 & \new_[4533]_ ;
  assign \new_[4535]_  = \new_[4534]_  & \new_[4529]_ ;
  assign \new_[4538]_  = ~A298 & A203;
  assign \new_[4542]_  = A302 & A300;
  assign \new_[4543]_  = A299 & \new_[4542]_ ;
  assign \new_[4544]_  = \new_[4543]_  & \new_[4538]_ ;
  assign \new_[4547]_  = ~A168 & A169;
  assign \new_[4551]_  = A201 & ~A200;
  assign \new_[4552]_  = A199 & \new_[4551]_ ;
  assign \new_[4553]_  = \new_[4552]_  & \new_[4547]_ ;
  assign \new_[4556]_  = A298 & A202;
  assign \new_[4560]_  = A301 & A300;
  assign \new_[4561]_  = ~A299 & \new_[4560]_ ;
  assign \new_[4562]_  = \new_[4561]_  & \new_[4556]_ ;
  assign \new_[4565]_  = ~A168 & A169;
  assign \new_[4569]_  = A201 & ~A200;
  assign \new_[4570]_  = A199 & \new_[4569]_ ;
  assign \new_[4571]_  = \new_[4570]_  & \new_[4565]_ ;
  assign \new_[4574]_  = A298 & A202;
  assign \new_[4578]_  = A302 & A300;
  assign \new_[4579]_  = ~A299 & \new_[4578]_ ;
  assign \new_[4580]_  = \new_[4579]_  & \new_[4574]_ ;
  assign \new_[4583]_  = ~A168 & A169;
  assign \new_[4587]_  = A201 & ~A200;
  assign \new_[4588]_  = A199 & \new_[4587]_ ;
  assign \new_[4589]_  = \new_[4588]_  & \new_[4583]_ ;
  assign \new_[4592]_  = ~A298 & A202;
  assign \new_[4596]_  = A301 & A300;
  assign \new_[4597]_  = A299 & \new_[4596]_ ;
  assign \new_[4598]_  = \new_[4597]_  & \new_[4592]_ ;
  assign \new_[4601]_  = ~A168 & A169;
  assign \new_[4605]_  = A201 & ~A200;
  assign \new_[4606]_  = A199 & \new_[4605]_ ;
  assign \new_[4607]_  = \new_[4606]_  & \new_[4601]_ ;
  assign \new_[4610]_  = ~A298 & A202;
  assign \new_[4614]_  = A302 & A300;
  assign \new_[4615]_  = A299 & \new_[4614]_ ;
  assign \new_[4616]_  = \new_[4615]_  & \new_[4610]_ ;
  assign \new_[4619]_  = ~A168 & A169;
  assign \new_[4623]_  = A201 & ~A200;
  assign \new_[4624]_  = A199 & \new_[4623]_ ;
  assign \new_[4625]_  = \new_[4624]_  & \new_[4619]_ ;
  assign \new_[4628]_  = A298 & A203;
  assign \new_[4632]_  = A301 & A300;
  assign \new_[4633]_  = ~A299 & \new_[4632]_ ;
  assign \new_[4634]_  = \new_[4633]_  & \new_[4628]_ ;
  assign \new_[4637]_  = ~A168 & A169;
  assign \new_[4641]_  = A201 & ~A200;
  assign \new_[4642]_  = A199 & \new_[4641]_ ;
  assign \new_[4643]_  = \new_[4642]_  & \new_[4637]_ ;
  assign \new_[4646]_  = A298 & A203;
  assign \new_[4650]_  = A302 & A300;
  assign \new_[4651]_  = ~A299 & \new_[4650]_ ;
  assign \new_[4652]_  = \new_[4651]_  & \new_[4646]_ ;
  assign \new_[4655]_  = ~A168 & A169;
  assign \new_[4659]_  = A201 & ~A200;
  assign \new_[4660]_  = A199 & \new_[4659]_ ;
  assign \new_[4661]_  = \new_[4660]_  & \new_[4655]_ ;
  assign \new_[4664]_  = ~A298 & A203;
  assign \new_[4668]_  = A301 & A300;
  assign \new_[4669]_  = A299 & \new_[4668]_ ;
  assign \new_[4670]_  = \new_[4669]_  & \new_[4664]_ ;
  assign \new_[4673]_  = ~A168 & A169;
  assign \new_[4677]_  = A201 & ~A200;
  assign \new_[4678]_  = A199 & \new_[4677]_ ;
  assign \new_[4679]_  = \new_[4678]_  & \new_[4673]_ ;
  assign \new_[4682]_  = ~A298 & A203;
  assign \new_[4686]_  = A302 & A300;
  assign \new_[4687]_  = A299 & \new_[4686]_ ;
  assign \new_[4688]_  = \new_[4687]_  & \new_[4682]_ ;
  assign \new_[4691]_  = ~A169 & A170;
  assign \new_[4695]_  = ~A166 & A167;
  assign \new_[4696]_  = ~A168 & \new_[4695]_ ;
  assign \new_[4697]_  = \new_[4696]_  & \new_[4691]_ ;
  assign \new_[4700]_  = A233 & ~A232;
  assign \new_[4704]_  = ~A236 & ~A235;
  assign \new_[4705]_  = ~A234 & \new_[4704]_ ;
  assign \new_[4706]_  = \new_[4705]_  & \new_[4700]_ ;
  assign \new_[4709]_  = ~A169 & A170;
  assign \new_[4713]_  = ~A166 & A167;
  assign \new_[4714]_  = ~A168 & \new_[4713]_ ;
  assign \new_[4715]_  = \new_[4714]_  & \new_[4709]_ ;
  assign \new_[4718]_  = ~A233 & A232;
  assign \new_[4722]_  = ~A236 & ~A235;
  assign \new_[4723]_  = ~A234 & \new_[4722]_ ;
  assign \new_[4724]_  = \new_[4723]_  & \new_[4718]_ ;
  assign \new_[4727]_  = ~A169 & A170;
  assign \new_[4731]_  = A166 & ~A167;
  assign \new_[4732]_  = ~A168 & \new_[4731]_ ;
  assign \new_[4733]_  = \new_[4732]_  & \new_[4727]_ ;
  assign \new_[4736]_  = A233 & ~A232;
  assign \new_[4740]_  = ~A236 & ~A235;
  assign \new_[4741]_  = ~A234 & \new_[4740]_ ;
  assign \new_[4742]_  = \new_[4741]_  & \new_[4736]_ ;
  assign \new_[4745]_  = ~A169 & A170;
  assign \new_[4749]_  = A166 & ~A167;
  assign \new_[4750]_  = ~A168 & \new_[4749]_ ;
  assign \new_[4751]_  = \new_[4750]_  & \new_[4745]_ ;
  assign \new_[4754]_  = ~A233 & A232;
  assign \new_[4758]_  = ~A236 & ~A235;
  assign \new_[4759]_  = ~A234 & \new_[4758]_ ;
  assign \new_[4760]_  = \new_[4759]_  & \new_[4754]_ ;
  assign \new_[4763]_  = A166 & A167;
  assign \new_[4767]_  = A201 & A200;
  assign \new_[4768]_  = ~A199 & \new_[4767]_ ;
  assign \new_[4769]_  = \new_[4768]_  & \new_[4763]_ ;
  assign \new_[4773]_  = ~A299 & A298;
  assign \new_[4774]_  = A202 & \new_[4773]_ ;
  assign \new_[4778]_  = ~A302 & ~A301;
  assign \new_[4779]_  = ~A300 & \new_[4778]_ ;
  assign \new_[4780]_  = \new_[4779]_  & \new_[4774]_ ;
  assign \new_[4783]_  = A166 & A167;
  assign \new_[4787]_  = A201 & A200;
  assign \new_[4788]_  = ~A199 & \new_[4787]_ ;
  assign \new_[4789]_  = \new_[4788]_  & \new_[4783]_ ;
  assign \new_[4793]_  = A299 & ~A298;
  assign \new_[4794]_  = A202 & \new_[4793]_ ;
  assign \new_[4798]_  = ~A302 & ~A301;
  assign \new_[4799]_  = ~A300 & \new_[4798]_ ;
  assign \new_[4800]_  = \new_[4799]_  & \new_[4794]_ ;
  assign \new_[4803]_  = A166 & A167;
  assign \new_[4807]_  = A201 & A200;
  assign \new_[4808]_  = ~A199 & \new_[4807]_ ;
  assign \new_[4809]_  = \new_[4808]_  & \new_[4803]_ ;
  assign \new_[4813]_  = ~A299 & A298;
  assign \new_[4814]_  = A203 & \new_[4813]_ ;
  assign \new_[4818]_  = ~A302 & ~A301;
  assign \new_[4819]_  = ~A300 & \new_[4818]_ ;
  assign \new_[4820]_  = \new_[4819]_  & \new_[4814]_ ;
  assign \new_[4823]_  = A166 & A167;
  assign \new_[4827]_  = A201 & A200;
  assign \new_[4828]_  = ~A199 & \new_[4827]_ ;
  assign \new_[4829]_  = \new_[4828]_  & \new_[4823]_ ;
  assign \new_[4833]_  = A299 & ~A298;
  assign \new_[4834]_  = A203 & \new_[4833]_ ;
  assign \new_[4838]_  = ~A302 & ~A301;
  assign \new_[4839]_  = ~A300 & \new_[4838]_ ;
  assign \new_[4840]_  = \new_[4839]_  & \new_[4834]_ ;
  assign \new_[4843]_  = A166 & A167;
  assign \new_[4847]_  = ~A201 & A200;
  assign \new_[4848]_  = ~A199 & \new_[4847]_ ;
  assign \new_[4849]_  = \new_[4848]_  & \new_[4843]_ ;
  assign \new_[4853]_  = A298 & ~A203;
  assign \new_[4854]_  = ~A202 & \new_[4853]_ ;
  assign \new_[4858]_  = A301 & A300;
  assign \new_[4859]_  = ~A299 & \new_[4858]_ ;
  assign \new_[4860]_  = \new_[4859]_  & \new_[4854]_ ;
  assign \new_[4863]_  = A166 & A167;
  assign \new_[4867]_  = ~A201 & A200;
  assign \new_[4868]_  = ~A199 & \new_[4867]_ ;
  assign \new_[4869]_  = \new_[4868]_  & \new_[4863]_ ;
  assign \new_[4873]_  = A298 & ~A203;
  assign \new_[4874]_  = ~A202 & \new_[4873]_ ;
  assign \new_[4878]_  = A302 & A300;
  assign \new_[4879]_  = ~A299 & \new_[4878]_ ;
  assign \new_[4880]_  = \new_[4879]_  & \new_[4874]_ ;
  assign \new_[4883]_  = A166 & A167;
  assign \new_[4887]_  = ~A201 & A200;
  assign \new_[4888]_  = ~A199 & \new_[4887]_ ;
  assign \new_[4889]_  = \new_[4888]_  & \new_[4883]_ ;
  assign \new_[4893]_  = ~A298 & ~A203;
  assign \new_[4894]_  = ~A202 & \new_[4893]_ ;
  assign \new_[4898]_  = A301 & A300;
  assign \new_[4899]_  = A299 & \new_[4898]_ ;
  assign \new_[4900]_  = \new_[4899]_  & \new_[4894]_ ;
  assign \new_[4903]_  = A166 & A167;
  assign \new_[4907]_  = ~A201 & A200;
  assign \new_[4908]_  = ~A199 & \new_[4907]_ ;
  assign \new_[4909]_  = \new_[4908]_  & \new_[4903]_ ;
  assign \new_[4913]_  = ~A298 & ~A203;
  assign \new_[4914]_  = ~A202 & \new_[4913]_ ;
  assign \new_[4918]_  = A302 & A300;
  assign \new_[4919]_  = A299 & \new_[4918]_ ;
  assign \new_[4920]_  = \new_[4919]_  & \new_[4914]_ ;
  assign \new_[4923]_  = A166 & A167;
  assign \new_[4927]_  = A201 & ~A200;
  assign \new_[4928]_  = A199 & \new_[4927]_ ;
  assign \new_[4929]_  = \new_[4928]_  & \new_[4923]_ ;
  assign \new_[4933]_  = ~A299 & A298;
  assign \new_[4934]_  = A202 & \new_[4933]_ ;
  assign \new_[4938]_  = ~A302 & ~A301;
  assign \new_[4939]_  = ~A300 & \new_[4938]_ ;
  assign \new_[4940]_  = \new_[4939]_  & \new_[4934]_ ;
  assign \new_[4943]_  = A166 & A167;
  assign \new_[4947]_  = A201 & ~A200;
  assign \new_[4948]_  = A199 & \new_[4947]_ ;
  assign \new_[4949]_  = \new_[4948]_  & \new_[4943]_ ;
  assign \new_[4953]_  = A299 & ~A298;
  assign \new_[4954]_  = A202 & \new_[4953]_ ;
  assign \new_[4958]_  = ~A302 & ~A301;
  assign \new_[4959]_  = ~A300 & \new_[4958]_ ;
  assign \new_[4960]_  = \new_[4959]_  & \new_[4954]_ ;
  assign \new_[4963]_  = A166 & A167;
  assign \new_[4967]_  = A201 & ~A200;
  assign \new_[4968]_  = A199 & \new_[4967]_ ;
  assign \new_[4969]_  = \new_[4968]_  & \new_[4963]_ ;
  assign \new_[4973]_  = ~A299 & A298;
  assign \new_[4974]_  = A203 & \new_[4973]_ ;
  assign \new_[4978]_  = ~A302 & ~A301;
  assign \new_[4979]_  = ~A300 & \new_[4978]_ ;
  assign \new_[4980]_  = \new_[4979]_  & \new_[4974]_ ;
  assign \new_[4983]_  = A166 & A167;
  assign \new_[4987]_  = A201 & ~A200;
  assign \new_[4988]_  = A199 & \new_[4987]_ ;
  assign \new_[4989]_  = \new_[4988]_  & \new_[4983]_ ;
  assign \new_[4993]_  = A299 & ~A298;
  assign \new_[4994]_  = A203 & \new_[4993]_ ;
  assign \new_[4998]_  = ~A302 & ~A301;
  assign \new_[4999]_  = ~A300 & \new_[4998]_ ;
  assign \new_[5000]_  = \new_[4999]_  & \new_[4994]_ ;
  assign \new_[5003]_  = A166 & A167;
  assign \new_[5007]_  = ~A201 & ~A200;
  assign \new_[5008]_  = A199 & \new_[5007]_ ;
  assign \new_[5009]_  = \new_[5008]_  & \new_[5003]_ ;
  assign \new_[5013]_  = A298 & ~A203;
  assign \new_[5014]_  = ~A202 & \new_[5013]_ ;
  assign \new_[5018]_  = A301 & A300;
  assign \new_[5019]_  = ~A299 & \new_[5018]_ ;
  assign \new_[5020]_  = \new_[5019]_  & \new_[5014]_ ;
  assign \new_[5023]_  = A166 & A167;
  assign \new_[5027]_  = ~A201 & ~A200;
  assign \new_[5028]_  = A199 & \new_[5027]_ ;
  assign \new_[5029]_  = \new_[5028]_  & \new_[5023]_ ;
  assign \new_[5033]_  = A298 & ~A203;
  assign \new_[5034]_  = ~A202 & \new_[5033]_ ;
  assign \new_[5038]_  = A302 & A300;
  assign \new_[5039]_  = ~A299 & \new_[5038]_ ;
  assign \new_[5040]_  = \new_[5039]_  & \new_[5034]_ ;
  assign \new_[5043]_  = A166 & A167;
  assign \new_[5047]_  = ~A201 & ~A200;
  assign \new_[5048]_  = A199 & \new_[5047]_ ;
  assign \new_[5049]_  = \new_[5048]_  & \new_[5043]_ ;
  assign \new_[5053]_  = ~A298 & ~A203;
  assign \new_[5054]_  = ~A202 & \new_[5053]_ ;
  assign \new_[5058]_  = A301 & A300;
  assign \new_[5059]_  = A299 & \new_[5058]_ ;
  assign \new_[5060]_  = \new_[5059]_  & \new_[5054]_ ;
  assign \new_[5063]_  = A166 & A167;
  assign \new_[5067]_  = ~A201 & ~A200;
  assign \new_[5068]_  = A199 & \new_[5067]_ ;
  assign \new_[5069]_  = \new_[5068]_  & \new_[5063]_ ;
  assign \new_[5073]_  = ~A298 & ~A203;
  assign \new_[5074]_  = ~A202 & \new_[5073]_ ;
  assign \new_[5078]_  = A302 & A300;
  assign \new_[5079]_  = A299 & \new_[5078]_ ;
  assign \new_[5080]_  = \new_[5079]_  & \new_[5074]_ ;
  assign \new_[5083]_  = ~A166 & ~A167;
  assign \new_[5087]_  = A201 & A200;
  assign \new_[5088]_  = ~A199 & \new_[5087]_ ;
  assign \new_[5089]_  = \new_[5088]_  & \new_[5083]_ ;
  assign \new_[5093]_  = ~A299 & A298;
  assign \new_[5094]_  = A202 & \new_[5093]_ ;
  assign \new_[5098]_  = ~A302 & ~A301;
  assign \new_[5099]_  = ~A300 & \new_[5098]_ ;
  assign \new_[5100]_  = \new_[5099]_  & \new_[5094]_ ;
  assign \new_[5103]_  = ~A166 & ~A167;
  assign \new_[5107]_  = A201 & A200;
  assign \new_[5108]_  = ~A199 & \new_[5107]_ ;
  assign \new_[5109]_  = \new_[5108]_  & \new_[5103]_ ;
  assign \new_[5113]_  = A299 & ~A298;
  assign \new_[5114]_  = A202 & \new_[5113]_ ;
  assign \new_[5118]_  = ~A302 & ~A301;
  assign \new_[5119]_  = ~A300 & \new_[5118]_ ;
  assign \new_[5120]_  = \new_[5119]_  & \new_[5114]_ ;
  assign \new_[5123]_  = ~A166 & ~A167;
  assign \new_[5127]_  = A201 & A200;
  assign \new_[5128]_  = ~A199 & \new_[5127]_ ;
  assign \new_[5129]_  = \new_[5128]_  & \new_[5123]_ ;
  assign \new_[5133]_  = ~A299 & A298;
  assign \new_[5134]_  = A203 & \new_[5133]_ ;
  assign \new_[5138]_  = ~A302 & ~A301;
  assign \new_[5139]_  = ~A300 & \new_[5138]_ ;
  assign \new_[5140]_  = \new_[5139]_  & \new_[5134]_ ;
  assign \new_[5143]_  = ~A166 & ~A167;
  assign \new_[5147]_  = A201 & A200;
  assign \new_[5148]_  = ~A199 & \new_[5147]_ ;
  assign \new_[5149]_  = \new_[5148]_  & \new_[5143]_ ;
  assign \new_[5153]_  = A299 & ~A298;
  assign \new_[5154]_  = A203 & \new_[5153]_ ;
  assign \new_[5158]_  = ~A302 & ~A301;
  assign \new_[5159]_  = ~A300 & \new_[5158]_ ;
  assign \new_[5160]_  = \new_[5159]_  & \new_[5154]_ ;
  assign \new_[5163]_  = ~A166 & ~A167;
  assign \new_[5167]_  = ~A201 & A200;
  assign \new_[5168]_  = ~A199 & \new_[5167]_ ;
  assign \new_[5169]_  = \new_[5168]_  & \new_[5163]_ ;
  assign \new_[5173]_  = A298 & ~A203;
  assign \new_[5174]_  = ~A202 & \new_[5173]_ ;
  assign \new_[5178]_  = A301 & A300;
  assign \new_[5179]_  = ~A299 & \new_[5178]_ ;
  assign \new_[5180]_  = \new_[5179]_  & \new_[5174]_ ;
  assign \new_[5183]_  = ~A166 & ~A167;
  assign \new_[5187]_  = ~A201 & A200;
  assign \new_[5188]_  = ~A199 & \new_[5187]_ ;
  assign \new_[5189]_  = \new_[5188]_  & \new_[5183]_ ;
  assign \new_[5193]_  = A298 & ~A203;
  assign \new_[5194]_  = ~A202 & \new_[5193]_ ;
  assign \new_[5198]_  = A302 & A300;
  assign \new_[5199]_  = ~A299 & \new_[5198]_ ;
  assign \new_[5200]_  = \new_[5199]_  & \new_[5194]_ ;
  assign \new_[5203]_  = ~A166 & ~A167;
  assign \new_[5207]_  = ~A201 & A200;
  assign \new_[5208]_  = ~A199 & \new_[5207]_ ;
  assign \new_[5209]_  = \new_[5208]_  & \new_[5203]_ ;
  assign \new_[5213]_  = ~A298 & ~A203;
  assign \new_[5214]_  = ~A202 & \new_[5213]_ ;
  assign \new_[5218]_  = A301 & A300;
  assign \new_[5219]_  = A299 & \new_[5218]_ ;
  assign \new_[5220]_  = \new_[5219]_  & \new_[5214]_ ;
  assign \new_[5223]_  = ~A166 & ~A167;
  assign \new_[5227]_  = ~A201 & A200;
  assign \new_[5228]_  = ~A199 & \new_[5227]_ ;
  assign \new_[5229]_  = \new_[5228]_  & \new_[5223]_ ;
  assign \new_[5233]_  = ~A298 & ~A203;
  assign \new_[5234]_  = ~A202 & \new_[5233]_ ;
  assign \new_[5238]_  = A302 & A300;
  assign \new_[5239]_  = A299 & \new_[5238]_ ;
  assign \new_[5240]_  = \new_[5239]_  & \new_[5234]_ ;
  assign \new_[5243]_  = ~A166 & ~A167;
  assign \new_[5247]_  = A201 & ~A200;
  assign \new_[5248]_  = A199 & \new_[5247]_ ;
  assign \new_[5249]_  = \new_[5248]_  & \new_[5243]_ ;
  assign \new_[5253]_  = ~A299 & A298;
  assign \new_[5254]_  = A202 & \new_[5253]_ ;
  assign \new_[5258]_  = ~A302 & ~A301;
  assign \new_[5259]_  = ~A300 & \new_[5258]_ ;
  assign \new_[5260]_  = \new_[5259]_  & \new_[5254]_ ;
  assign \new_[5263]_  = ~A166 & ~A167;
  assign \new_[5267]_  = A201 & ~A200;
  assign \new_[5268]_  = A199 & \new_[5267]_ ;
  assign \new_[5269]_  = \new_[5268]_  & \new_[5263]_ ;
  assign \new_[5273]_  = A299 & ~A298;
  assign \new_[5274]_  = A202 & \new_[5273]_ ;
  assign \new_[5278]_  = ~A302 & ~A301;
  assign \new_[5279]_  = ~A300 & \new_[5278]_ ;
  assign \new_[5280]_  = \new_[5279]_  & \new_[5274]_ ;
  assign \new_[5283]_  = ~A166 & ~A167;
  assign \new_[5287]_  = A201 & ~A200;
  assign \new_[5288]_  = A199 & \new_[5287]_ ;
  assign \new_[5289]_  = \new_[5288]_  & \new_[5283]_ ;
  assign \new_[5293]_  = ~A299 & A298;
  assign \new_[5294]_  = A203 & \new_[5293]_ ;
  assign \new_[5298]_  = ~A302 & ~A301;
  assign \new_[5299]_  = ~A300 & \new_[5298]_ ;
  assign \new_[5300]_  = \new_[5299]_  & \new_[5294]_ ;
  assign \new_[5303]_  = ~A166 & ~A167;
  assign \new_[5307]_  = A201 & ~A200;
  assign \new_[5308]_  = A199 & \new_[5307]_ ;
  assign \new_[5309]_  = \new_[5308]_  & \new_[5303]_ ;
  assign \new_[5313]_  = A299 & ~A298;
  assign \new_[5314]_  = A203 & \new_[5313]_ ;
  assign \new_[5318]_  = ~A302 & ~A301;
  assign \new_[5319]_  = ~A300 & \new_[5318]_ ;
  assign \new_[5320]_  = \new_[5319]_  & \new_[5314]_ ;
  assign \new_[5323]_  = ~A166 & ~A167;
  assign \new_[5327]_  = ~A201 & ~A200;
  assign \new_[5328]_  = A199 & \new_[5327]_ ;
  assign \new_[5329]_  = \new_[5328]_  & \new_[5323]_ ;
  assign \new_[5333]_  = A298 & ~A203;
  assign \new_[5334]_  = ~A202 & \new_[5333]_ ;
  assign \new_[5338]_  = A301 & A300;
  assign \new_[5339]_  = ~A299 & \new_[5338]_ ;
  assign \new_[5340]_  = \new_[5339]_  & \new_[5334]_ ;
  assign \new_[5343]_  = ~A166 & ~A167;
  assign \new_[5347]_  = ~A201 & ~A200;
  assign \new_[5348]_  = A199 & \new_[5347]_ ;
  assign \new_[5349]_  = \new_[5348]_  & \new_[5343]_ ;
  assign \new_[5353]_  = A298 & ~A203;
  assign \new_[5354]_  = ~A202 & \new_[5353]_ ;
  assign \new_[5358]_  = A302 & A300;
  assign \new_[5359]_  = ~A299 & \new_[5358]_ ;
  assign \new_[5360]_  = \new_[5359]_  & \new_[5354]_ ;
  assign \new_[5363]_  = ~A166 & ~A167;
  assign \new_[5367]_  = ~A201 & ~A200;
  assign \new_[5368]_  = A199 & \new_[5367]_ ;
  assign \new_[5369]_  = \new_[5368]_  & \new_[5363]_ ;
  assign \new_[5373]_  = ~A298 & ~A203;
  assign \new_[5374]_  = ~A202 & \new_[5373]_ ;
  assign \new_[5378]_  = A301 & A300;
  assign \new_[5379]_  = A299 & \new_[5378]_ ;
  assign \new_[5380]_  = \new_[5379]_  & \new_[5374]_ ;
  assign \new_[5383]_  = ~A166 & ~A167;
  assign \new_[5387]_  = ~A201 & ~A200;
  assign \new_[5388]_  = A199 & \new_[5387]_ ;
  assign \new_[5389]_  = \new_[5388]_  & \new_[5383]_ ;
  assign \new_[5393]_  = ~A298 & ~A203;
  assign \new_[5394]_  = ~A202 & \new_[5393]_ ;
  assign \new_[5398]_  = A302 & A300;
  assign \new_[5399]_  = A299 & \new_[5398]_ ;
  assign \new_[5400]_  = \new_[5399]_  & \new_[5394]_ ;
  assign \new_[5403]_  = A168 & ~A170;
  assign \new_[5407]_  = A201 & ~A166;
  assign \new_[5408]_  = A167 & \new_[5407]_ ;
  assign \new_[5409]_  = \new_[5408]_  & \new_[5403]_ ;
  assign \new_[5413]_  = A298 & ~A203;
  assign \new_[5414]_  = ~A202 & \new_[5413]_ ;
  assign \new_[5418]_  = A301 & A300;
  assign \new_[5419]_  = ~A299 & \new_[5418]_ ;
  assign \new_[5420]_  = \new_[5419]_  & \new_[5414]_ ;
  assign \new_[5423]_  = A168 & ~A170;
  assign \new_[5427]_  = A201 & ~A166;
  assign \new_[5428]_  = A167 & \new_[5427]_ ;
  assign \new_[5429]_  = \new_[5428]_  & \new_[5423]_ ;
  assign \new_[5433]_  = A298 & ~A203;
  assign \new_[5434]_  = ~A202 & \new_[5433]_ ;
  assign \new_[5438]_  = A302 & A300;
  assign \new_[5439]_  = ~A299 & \new_[5438]_ ;
  assign \new_[5440]_  = \new_[5439]_  & \new_[5434]_ ;
  assign \new_[5443]_  = A168 & ~A170;
  assign \new_[5447]_  = A201 & ~A166;
  assign \new_[5448]_  = A167 & \new_[5447]_ ;
  assign \new_[5449]_  = \new_[5448]_  & \new_[5443]_ ;
  assign \new_[5453]_  = ~A298 & ~A203;
  assign \new_[5454]_  = ~A202 & \new_[5453]_ ;
  assign \new_[5458]_  = A301 & A300;
  assign \new_[5459]_  = A299 & \new_[5458]_ ;
  assign \new_[5460]_  = \new_[5459]_  & \new_[5454]_ ;
  assign \new_[5463]_  = A168 & ~A170;
  assign \new_[5467]_  = A201 & ~A166;
  assign \new_[5468]_  = A167 & \new_[5467]_ ;
  assign \new_[5469]_  = \new_[5468]_  & \new_[5463]_ ;
  assign \new_[5473]_  = ~A298 & ~A203;
  assign \new_[5474]_  = ~A202 & \new_[5473]_ ;
  assign \new_[5478]_  = A302 & A300;
  assign \new_[5479]_  = A299 & \new_[5478]_ ;
  assign \new_[5480]_  = \new_[5479]_  & \new_[5474]_ ;
  assign \new_[5483]_  = A168 & ~A170;
  assign \new_[5487]_  = ~A201 & ~A166;
  assign \new_[5488]_  = A167 & \new_[5487]_ ;
  assign \new_[5489]_  = \new_[5488]_  & \new_[5483]_ ;
  assign \new_[5493]_  = ~A299 & A298;
  assign \new_[5494]_  = A202 & \new_[5493]_ ;
  assign \new_[5498]_  = ~A302 & ~A301;
  assign \new_[5499]_  = ~A300 & \new_[5498]_ ;
  assign \new_[5500]_  = \new_[5499]_  & \new_[5494]_ ;
  assign \new_[5503]_  = A168 & ~A170;
  assign \new_[5507]_  = ~A201 & ~A166;
  assign \new_[5508]_  = A167 & \new_[5507]_ ;
  assign \new_[5509]_  = \new_[5508]_  & \new_[5503]_ ;
  assign \new_[5513]_  = A299 & ~A298;
  assign \new_[5514]_  = A202 & \new_[5513]_ ;
  assign \new_[5518]_  = ~A302 & ~A301;
  assign \new_[5519]_  = ~A300 & \new_[5518]_ ;
  assign \new_[5520]_  = \new_[5519]_  & \new_[5514]_ ;
  assign \new_[5523]_  = A168 & ~A170;
  assign \new_[5527]_  = ~A201 & ~A166;
  assign \new_[5528]_  = A167 & \new_[5527]_ ;
  assign \new_[5529]_  = \new_[5528]_  & \new_[5523]_ ;
  assign \new_[5533]_  = ~A299 & A298;
  assign \new_[5534]_  = A203 & \new_[5533]_ ;
  assign \new_[5538]_  = ~A302 & ~A301;
  assign \new_[5539]_  = ~A300 & \new_[5538]_ ;
  assign \new_[5540]_  = \new_[5539]_  & \new_[5534]_ ;
  assign \new_[5543]_  = A168 & ~A170;
  assign \new_[5547]_  = ~A201 & ~A166;
  assign \new_[5548]_  = A167 & \new_[5547]_ ;
  assign \new_[5549]_  = \new_[5548]_  & \new_[5543]_ ;
  assign \new_[5553]_  = A299 & ~A298;
  assign \new_[5554]_  = A203 & \new_[5553]_ ;
  assign \new_[5558]_  = ~A302 & ~A301;
  assign \new_[5559]_  = ~A300 & \new_[5558]_ ;
  assign \new_[5560]_  = \new_[5559]_  & \new_[5554]_ ;
  assign \new_[5563]_  = A168 & ~A170;
  assign \new_[5567]_  = A199 & ~A166;
  assign \new_[5568]_  = A167 & \new_[5567]_ ;
  assign \new_[5569]_  = \new_[5568]_  & \new_[5563]_ ;
  assign \new_[5573]_  = ~A299 & A298;
  assign \new_[5574]_  = A200 & \new_[5573]_ ;
  assign \new_[5578]_  = ~A302 & ~A301;
  assign \new_[5579]_  = ~A300 & \new_[5578]_ ;
  assign \new_[5580]_  = \new_[5579]_  & \new_[5574]_ ;
  assign \new_[5583]_  = A168 & ~A170;
  assign \new_[5587]_  = A199 & ~A166;
  assign \new_[5588]_  = A167 & \new_[5587]_ ;
  assign \new_[5589]_  = \new_[5588]_  & \new_[5583]_ ;
  assign \new_[5593]_  = A299 & ~A298;
  assign \new_[5594]_  = A200 & \new_[5593]_ ;
  assign \new_[5598]_  = ~A302 & ~A301;
  assign \new_[5599]_  = ~A300 & \new_[5598]_ ;
  assign \new_[5600]_  = \new_[5599]_  & \new_[5594]_ ;
  assign \new_[5603]_  = A168 & ~A170;
  assign \new_[5607]_  = ~A199 & ~A166;
  assign \new_[5608]_  = A167 & \new_[5607]_ ;
  assign \new_[5609]_  = \new_[5608]_  & \new_[5603]_ ;
  assign \new_[5613]_  = ~A299 & A298;
  assign \new_[5614]_  = ~A200 & \new_[5613]_ ;
  assign \new_[5618]_  = ~A302 & ~A301;
  assign \new_[5619]_  = ~A300 & \new_[5618]_ ;
  assign \new_[5620]_  = \new_[5619]_  & \new_[5614]_ ;
  assign \new_[5623]_  = A168 & ~A170;
  assign \new_[5627]_  = ~A199 & ~A166;
  assign \new_[5628]_  = A167 & \new_[5627]_ ;
  assign \new_[5629]_  = \new_[5628]_  & \new_[5623]_ ;
  assign \new_[5633]_  = A299 & ~A298;
  assign \new_[5634]_  = ~A200 & \new_[5633]_ ;
  assign \new_[5638]_  = ~A302 & ~A301;
  assign \new_[5639]_  = ~A300 & \new_[5638]_ ;
  assign \new_[5640]_  = \new_[5639]_  & \new_[5634]_ ;
  assign \new_[5643]_  = A168 & ~A170;
  assign \new_[5647]_  = A201 & A166;
  assign \new_[5648]_  = ~A167 & \new_[5647]_ ;
  assign \new_[5649]_  = \new_[5648]_  & \new_[5643]_ ;
  assign \new_[5653]_  = A298 & ~A203;
  assign \new_[5654]_  = ~A202 & \new_[5653]_ ;
  assign \new_[5658]_  = A301 & A300;
  assign \new_[5659]_  = ~A299 & \new_[5658]_ ;
  assign \new_[5660]_  = \new_[5659]_  & \new_[5654]_ ;
  assign \new_[5663]_  = A168 & ~A170;
  assign \new_[5667]_  = A201 & A166;
  assign \new_[5668]_  = ~A167 & \new_[5667]_ ;
  assign \new_[5669]_  = \new_[5668]_  & \new_[5663]_ ;
  assign \new_[5673]_  = A298 & ~A203;
  assign \new_[5674]_  = ~A202 & \new_[5673]_ ;
  assign \new_[5678]_  = A302 & A300;
  assign \new_[5679]_  = ~A299 & \new_[5678]_ ;
  assign \new_[5680]_  = \new_[5679]_  & \new_[5674]_ ;
  assign \new_[5683]_  = A168 & ~A170;
  assign \new_[5687]_  = A201 & A166;
  assign \new_[5688]_  = ~A167 & \new_[5687]_ ;
  assign \new_[5689]_  = \new_[5688]_  & \new_[5683]_ ;
  assign \new_[5693]_  = ~A298 & ~A203;
  assign \new_[5694]_  = ~A202 & \new_[5693]_ ;
  assign \new_[5698]_  = A301 & A300;
  assign \new_[5699]_  = A299 & \new_[5698]_ ;
  assign \new_[5700]_  = \new_[5699]_  & \new_[5694]_ ;
  assign \new_[5703]_  = A168 & ~A170;
  assign \new_[5707]_  = A201 & A166;
  assign \new_[5708]_  = ~A167 & \new_[5707]_ ;
  assign \new_[5709]_  = \new_[5708]_  & \new_[5703]_ ;
  assign \new_[5713]_  = ~A298 & ~A203;
  assign \new_[5714]_  = ~A202 & \new_[5713]_ ;
  assign \new_[5718]_  = A302 & A300;
  assign \new_[5719]_  = A299 & \new_[5718]_ ;
  assign \new_[5720]_  = \new_[5719]_  & \new_[5714]_ ;
  assign \new_[5723]_  = A168 & ~A170;
  assign \new_[5727]_  = ~A201 & A166;
  assign \new_[5728]_  = ~A167 & \new_[5727]_ ;
  assign \new_[5729]_  = \new_[5728]_  & \new_[5723]_ ;
  assign \new_[5733]_  = ~A299 & A298;
  assign \new_[5734]_  = A202 & \new_[5733]_ ;
  assign \new_[5738]_  = ~A302 & ~A301;
  assign \new_[5739]_  = ~A300 & \new_[5738]_ ;
  assign \new_[5740]_  = \new_[5739]_  & \new_[5734]_ ;
  assign \new_[5743]_  = A168 & ~A170;
  assign \new_[5747]_  = ~A201 & A166;
  assign \new_[5748]_  = ~A167 & \new_[5747]_ ;
  assign \new_[5749]_  = \new_[5748]_  & \new_[5743]_ ;
  assign \new_[5753]_  = A299 & ~A298;
  assign \new_[5754]_  = A202 & \new_[5753]_ ;
  assign \new_[5758]_  = ~A302 & ~A301;
  assign \new_[5759]_  = ~A300 & \new_[5758]_ ;
  assign \new_[5760]_  = \new_[5759]_  & \new_[5754]_ ;
  assign \new_[5763]_  = A168 & ~A170;
  assign \new_[5767]_  = ~A201 & A166;
  assign \new_[5768]_  = ~A167 & \new_[5767]_ ;
  assign \new_[5769]_  = \new_[5768]_  & \new_[5763]_ ;
  assign \new_[5773]_  = ~A299 & A298;
  assign \new_[5774]_  = A203 & \new_[5773]_ ;
  assign \new_[5778]_  = ~A302 & ~A301;
  assign \new_[5779]_  = ~A300 & \new_[5778]_ ;
  assign \new_[5780]_  = \new_[5779]_  & \new_[5774]_ ;
  assign \new_[5783]_  = A168 & ~A170;
  assign \new_[5787]_  = ~A201 & A166;
  assign \new_[5788]_  = ~A167 & \new_[5787]_ ;
  assign \new_[5789]_  = \new_[5788]_  & \new_[5783]_ ;
  assign \new_[5793]_  = A299 & ~A298;
  assign \new_[5794]_  = A203 & \new_[5793]_ ;
  assign \new_[5798]_  = ~A302 & ~A301;
  assign \new_[5799]_  = ~A300 & \new_[5798]_ ;
  assign \new_[5800]_  = \new_[5799]_  & \new_[5794]_ ;
  assign \new_[5803]_  = A168 & ~A170;
  assign \new_[5807]_  = A199 & A166;
  assign \new_[5808]_  = ~A167 & \new_[5807]_ ;
  assign \new_[5809]_  = \new_[5808]_  & \new_[5803]_ ;
  assign \new_[5813]_  = ~A299 & A298;
  assign \new_[5814]_  = A200 & \new_[5813]_ ;
  assign \new_[5818]_  = ~A302 & ~A301;
  assign \new_[5819]_  = ~A300 & \new_[5818]_ ;
  assign \new_[5820]_  = \new_[5819]_  & \new_[5814]_ ;
  assign \new_[5823]_  = A168 & ~A170;
  assign \new_[5827]_  = A199 & A166;
  assign \new_[5828]_  = ~A167 & \new_[5827]_ ;
  assign \new_[5829]_  = \new_[5828]_  & \new_[5823]_ ;
  assign \new_[5833]_  = A299 & ~A298;
  assign \new_[5834]_  = A200 & \new_[5833]_ ;
  assign \new_[5838]_  = ~A302 & ~A301;
  assign \new_[5839]_  = ~A300 & \new_[5838]_ ;
  assign \new_[5840]_  = \new_[5839]_  & \new_[5834]_ ;
  assign \new_[5843]_  = A168 & ~A170;
  assign \new_[5847]_  = ~A199 & A166;
  assign \new_[5848]_  = ~A167 & \new_[5847]_ ;
  assign \new_[5849]_  = \new_[5848]_  & \new_[5843]_ ;
  assign \new_[5853]_  = ~A299 & A298;
  assign \new_[5854]_  = ~A200 & \new_[5853]_ ;
  assign \new_[5858]_  = ~A302 & ~A301;
  assign \new_[5859]_  = ~A300 & \new_[5858]_ ;
  assign \new_[5860]_  = \new_[5859]_  & \new_[5854]_ ;
  assign \new_[5863]_  = A168 & ~A170;
  assign \new_[5867]_  = ~A199 & A166;
  assign \new_[5868]_  = ~A167 & \new_[5867]_ ;
  assign \new_[5869]_  = \new_[5868]_  & \new_[5863]_ ;
  assign \new_[5873]_  = A299 & ~A298;
  assign \new_[5874]_  = ~A200 & \new_[5873]_ ;
  assign \new_[5878]_  = ~A302 & ~A301;
  assign \new_[5879]_  = ~A300 & \new_[5878]_ ;
  assign \new_[5880]_  = \new_[5879]_  & \new_[5874]_ ;
  assign \new_[5883]_  = ~A168 & ~A170;
  assign \new_[5887]_  = A201 & A200;
  assign \new_[5888]_  = ~A199 & \new_[5887]_ ;
  assign \new_[5889]_  = \new_[5888]_  & \new_[5883]_ ;
  assign \new_[5893]_  = ~A299 & A298;
  assign \new_[5894]_  = A202 & \new_[5893]_ ;
  assign \new_[5898]_  = ~A302 & ~A301;
  assign \new_[5899]_  = ~A300 & \new_[5898]_ ;
  assign \new_[5900]_  = \new_[5899]_  & \new_[5894]_ ;
  assign \new_[5903]_  = ~A168 & ~A170;
  assign \new_[5907]_  = A201 & A200;
  assign \new_[5908]_  = ~A199 & \new_[5907]_ ;
  assign \new_[5909]_  = \new_[5908]_  & \new_[5903]_ ;
  assign \new_[5913]_  = A299 & ~A298;
  assign \new_[5914]_  = A202 & \new_[5913]_ ;
  assign \new_[5918]_  = ~A302 & ~A301;
  assign \new_[5919]_  = ~A300 & \new_[5918]_ ;
  assign \new_[5920]_  = \new_[5919]_  & \new_[5914]_ ;
  assign \new_[5923]_  = ~A168 & ~A170;
  assign \new_[5927]_  = A201 & A200;
  assign \new_[5928]_  = ~A199 & \new_[5927]_ ;
  assign \new_[5929]_  = \new_[5928]_  & \new_[5923]_ ;
  assign \new_[5933]_  = ~A299 & A298;
  assign \new_[5934]_  = A203 & \new_[5933]_ ;
  assign \new_[5938]_  = ~A302 & ~A301;
  assign \new_[5939]_  = ~A300 & \new_[5938]_ ;
  assign \new_[5940]_  = \new_[5939]_  & \new_[5934]_ ;
  assign \new_[5943]_  = ~A168 & ~A170;
  assign \new_[5947]_  = A201 & A200;
  assign \new_[5948]_  = ~A199 & \new_[5947]_ ;
  assign \new_[5949]_  = \new_[5948]_  & \new_[5943]_ ;
  assign \new_[5953]_  = A299 & ~A298;
  assign \new_[5954]_  = A203 & \new_[5953]_ ;
  assign \new_[5958]_  = ~A302 & ~A301;
  assign \new_[5959]_  = ~A300 & \new_[5958]_ ;
  assign \new_[5960]_  = \new_[5959]_  & \new_[5954]_ ;
  assign \new_[5963]_  = ~A168 & ~A170;
  assign \new_[5967]_  = ~A201 & A200;
  assign \new_[5968]_  = ~A199 & \new_[5967]_ ;
  assign \new_[5969]_  = \new_[5968]_  & \new_[5963]_ ;
  assign \new_[5973]_  = A298 & ~A203;
  assign \new_[5974]_  = ~A202 & \new_[5973]_ ;
  assign \new_[5978]_  = A301 & A300;
  assign \new_[5979]_  = ~A299 & \new_[5978]_ ;
  assign \new_[5980]_  = \new_[5979]_  & \new_[5974]_ ;
  assign \new_[5983]_  = ~A168 & ~A170;
  assign \new_[5987]_  = ~A201 & A200;
  assign \new_[5988]_  = ~A199 & \new_[5987]_ ;
  assign \new_[5989]_  = \new_[5988]_  & \new_[5983]_ ;
  assign \new_[5993]_  = A298 & ~A203;
  assign \new_[5994]_  = ~A202 & \new_[5993]_ ;
  assign \new_[5998]_  = A302 & A300;
  assign \new_[5999]_  = ~A299 & \new_[5998]_ ;
  assign \new_[6000]_  = \new_[5999]_  & \new_[5994]_ ;
  assign \new_[6003]_  = ~A168 & ~A170;
  assign \new_[6007]_  = ~A201 & A200;
  assign \new_[6008]_  = ~A199 & \new_[6007]_ ;
  assign \new_[6009]_  = \new_[6008]_  & \new_[6003]_ ;
  assign \new_[6013]_  = ~A298 & ~A203;
  assign \new_[6014]_  = ~A202 & \new_[6013]_ ;
  assign \new_[6018]_  = A301 & A300;
  assign \new_[6019]_  = A299 & \new_[6018]_ ;
  assign \new_[6020]_  = \new_[6019]_  & \new_[6014]_ ;
  assign \new_[6023]_  = ~A168 & ~A170;
  assign \new_[6027]_  = ~A201 & A200;
  assign \new_[6028]_  = ~A199 & \new_[6027]_ ;
  assign \new_[6029]_  = \new_[6028]_  & \new_[6023]_ ;
  assign \new_[6033]_  = ~A298 & ~A203;
  assign \new_[6034]_  = ~A202 & \new_[6033]_ ;
  assign \new_[6038]_  = A302 & A300;
  assign \new_[6039]_  = A299 & \new_[6038]_ ;
  assign \new_[6040]_  = \new_[6039]_  & \new_[6034]_ ;
  assign \new_[6043]_  = ~A168 & ~A170;
  assign \new_[6047]_  = A201 & ~A200;
  assign \new_[6048]_  = A199 & \new_[6047]_ ;
  assign \new_[6049]_  = \new_[6048]_  & \new_[6043]_ ;
  assign \new_[6053]_  = ~A299 & A298;
  assign \new_[6054]_  = A202 & \new_[6053]_ ;
  assign \new_[6058]_  = ~A302 & ~A301;
  assign \new_[6059]_  = ~A300 & \new_[6058]_ ;
  assign \new_[6060]_  = \new_[6059]_  & \new_[6054]_ ;
  assign \new_[6063]_  = ~A168 & ~A170;
  assign \new_[6067]_  = A201 & ~A200;
  assign \new_[6068]_  = A199 & \new_[6067]_ ;
  assign \new_[6069]_  = \new_[6068]_  & \new_[6063]_ ;
  assign \new_[6073]_  = A299 & ~A298;
  assign \new_[6074]_  = A202 & \new_[6073]_ ;
  assign \new_[6078]_  = ~A302 & ~A301;
  assign \new_[6079]_  = ~A300 & \new_[6078]_ ;
  assign \new_[6080]_  = \new_[6079]_  & \new_[6074]_ ;
  assign \new_[6083]_  = ~A168 & ~A170;
  assign \new_[6087]_  = A201 & ~A200;
  assign \new_[6088]_  = A199 & \new_[6087]_ ;
  assign \new_[6089]_  = \new_[6088]_  & \new_[6083]_ ;
  assign \new_[6093]_  = ~A299 & A298;
  assign \new_[6094]_  = A203 & \new_[6093]_ ;
  assign \new_[6098]_  = ~A302 & ~A301;
  assign \new_[6099]_  = ~A300 & \new_[6098]_ ;
  assign \new_[6100]_  = \new_[6099]_  & \new_[6094]_ ;
  assign \new_[6103]_  = ~A168 & ~A170;
  assign \new_[6107]_  = A201 & ~A200;
  assign \new_[6108]_  = A199 & \new_[6107]_ ;
  assign \new_[6109]_  = \new_[6108]_  & \new_[6103]_ ;
  assign \new_[6113]_  = A299 & ~A298;
  assign \new_[6114]_  = A203 & \new_[6113]_ ;
  assign \new_[6118]_  = ~A302 & ~A301;
  assign \new_[6119]_  = ~A300 & \new_[6118]_ ;
  assign \new_[6120]_  = \new_[6119]_  & \new_[6114]_ ;
  assign \new_[6123]_  = ~A168 & ~A170;
  assign \new_[6127]_  = ~A201 & ~A200;
  assign \new_[6128]_  = A199 & \new_[6127]_ ;
  assign \new_[6129]_  = \new_[6128]_  & \new_[6123]_ ;
  assign \new_[6133]_  = A298 & ~A203;
  assign \new_[6134]_  = ~A202 & \new_[6133]_ ;
  assign \new_[6138]_  = A301 & A300;
  assign \new_[6139]_  = ~A299 & \new_[6138]_ ;
  assign \new_[6140]_  = \new_[6139]_  & \new_[6134]_ ;
  assign \new_[6143]_  = ~A168 & ~A170;
  assign \new_[6147]_  = ~A201 & ~A200;
  assign \new_[6148]_  = A199 & \new_[6147]_ ;
  assign \new_[6149]_  = \new_[6148]_  & \new_[6143]_ ;
  assign \new_[6153]_  = A298 & ~A203;
  assign \new_[6154]_  = ~A202 & \new_[6153]_ ;
  assign \new_[6158]_  = A302 & A300;
  assign \new_[6159]_  = ~A299 & \new_[6158]_ ;
  assign \new_[6160]_  = \new_[6159]_  & \new_[6154]_ ;
  assign \new_[6163]_  = ~A168 & ~A170;
  assign \new_[6167]_  = ~A201 & ~A200;
  assign \new_[6168]_  = A199 & \new_[6167]_ ;
  assign \new_[6169]_  = \new_[6168]_  & \new_[6163]_ ;
  assign \new_[6173]_  = ~A298 & ~A203;
  assign \new_[6174]_  = ~A202 & \new_[6173]_ ;
  assign \new_[6178]_  = A301 & A300;
  assign \new_[6179]_  = A299 & \new_[6178]_ ;
  assign \new_[6180]_  = \new_[6179]_  & \new_[6174]_ ;
  assign \new_[6183]_  = ~A168 & ~A170;
  assign \new_[6187]_  = ~A201 & ~A200;
  assign \new_[6188]_  = A199 & \new_[6187]_ ;
  assign \new_[6189]_  = \new_[6188]_  & \new_[6183]_ ;
  assign \new_[6193]_  = ~A298 & ~A203;
  assign \new_[6194]_  = ~A202 & \new_[6193]_ ;
  assign \new_[6198]_  = A302 & A300;
  assign \new_[6199]_  = A299 & \new_[6198]_ ;
  assign \new_[6200]_  = \new_[6199]_  & \new_[6194]_ ;
  assign \new_[6203]_  = A168 & A169;
  assign \new_[6207]_  = A201 & ~A166;
  assign \new_[6208]_  = A167 & \new_[6207]_ ;
  assign \new_[6209]_  = \new_[6208]_  & \new_[6203]_ ;
  assign \new_[6213]_  = A298 & ~A203;
  assign \new_[6214]_  = ~A202 & \new_[6213]_ ;
  assign \new_[6218]_  = A301 & A300;
  assign \new_[6219]_  = ~A299 & \new_[6218]_ ;
  assign \new_[6220]_  = \new_[6219]_  & \new_[6214]_ ;
  assign \new_[6223]_  = A168 & A169;
  assign \new_[6227]_  = A201 & ~A166;
  assign \new_[6228]_  = A167 & \new_[6227]_ ;
  assign \new_[6229]_  = \new_[6228]_  & \new_[6223]_ ;
  assign \new_[6233]_  = A298 & ~A203;
  assign \new_[6234]_  = ~A202 & \new_[6233]_ ;
  assign \new_[6238]_  = A302 & A300;
  assign \new_[6239]_  = ~A299 & \new_[6238]_ ;
  assign \new_[6240]_  = \new_[6239]_  & \new_[6234]_ ;
  assign \new_[6243]_  = A168 & A169;
  assign \new_[6247]_  = A201 & ~A166;
  assign \new_[6248]_  = A167 & \new_[6247]_ ;
  assign \new_[6249]_  = \new_[6248]_  & \new_[6243]_ ;
  assign \new_[6253]_  = ~A298 & ~A203;
  assign \new_[6254]_  = ~A202 & \new_[6253]_ ;
  assign \new_[6258]_  = A301 & A300;
  assign \new_[6259]_  = A299 & \new_[6258]_ ;
  assign \new_[6260]_  = \new_[6259]_  & \new_[6254]_ ;
  assign \new_[6263]_  = A168 & A169;
  assign \new_[6267]_  = A201 & ~A166;
  assign \new_[6268]_  = A167 & \new_[6267]_ ;
  assign \new_[6269]_  = \new_[6268]_  & \new_[6263]_ ;
  assign \new_[6273]_  = ~A298 & ~A203;
  assign \new_[6274]_  = ~A202 & \new_[6273]_ ;
  assign \new_[6278]_  = A302 & A300;
  assign \new_[6279]_  = A299 & \new_[6278]_ ;
  assign \new_[6280]_  = \new_[6279]_  & \new_[6274]_ ;
  assign \new_[6283]_  = A168 & A169;
  assign \new_[6287]_  = ~A201 & ~A166;
  assign \new_[6288]_  = A167 & \new_[6287]_ ;
  assign \new_[6289]_  = \new_[6288]_  & \new_[6283]_ ;
  assign \new_[6293]_  = ~A299 & A298;
  assign \new_[6294]_  = A202 & \new_[6293]_ ;
  assign \new_[6298]_  = ~A302 & ~A301;
  assign \new_[6299]_  = ~A300 & \new_[6298]_ ;
  assign \new_[6300]_  = \new_[6299]_  & \new_[6294]_ ;
  assign \new_[6303]_  = A168 & A169;
  assign \new_[6307]_  = ~A201 & ~A166;
  assign \new_[6308]_  = A167 & \new_[6307]_ ;
  assign \new_[6309]_  = \new_[6308]_  & \new_[6303]_ ;
  assign \new_[6313]_  = A299 & ~A298;
  assign \new_[6314]_  = A202 & \new_[6313]_ ;
  assign \new_[6318]_  = ~A302 & ~A301;
  assign \new_[6319]_  = ~A300 & \new_[6318]_ ;
  assign \new_[6320]_  = \new_[6319]_  & \new_[6314]_ ;
  assign \new_[6323]_  = A168 & A169;
  assign \new_[6327]_  = ~A201 & ~A166;
  assign \new_[6328]_  = A167 & \new_[6327]_ ;
  assign \new_[6329]_  = \new_[6328]_  & \new_[6323]_ ;
  assign \new_[6333]_  = ~A299 & A298;
  assign \new_[6334]_  = A203 & \new_[6333]_ ;
  assign \new_[6338]_  = ~A302 & ~A301;
  assign \new_[6339]_  = ~A300 & \new_[6338]_ ;
  assign \new_[6340]_  = \new_[6339]_  & \new_[6334]_ ;
  assign \new_[6343]_  = A168 & A169;
  assign \new_[6347]_  = ~A201 & ~A166;
  assign \new_[6348]_  = A167 & \new_[6347]_ ;
  assign \new_[6349]_  = \new_[6348]_  & \new_[6343]_ ;
  assign \new_[6353]_  = A299 & ~A298;
  assign \new_[6354]_  = A203 & \new_[6353]_ ;
  assign \new_[6358]_  = ~A302 & ~A301;
  assign \new_[6359]_  = ~A300 & \new_[6358]_ ;
  assign \new_[6360]_  = \new_[6359]_  & \new_[6354]_ ;
  assign \new_[6363]_  = A168 & A169;
  assign \new_[6367]_  = A199 & ~A166;
  assign \new_[6368]_  = A167 & \new_[6367]_ ;
  assign \new_[6369]_  = \new_[6368]_  & \new_[6363]_ ;
  assign \new_[6373]_  = ~A299 & A298;
  assign \new_[6374]_  = A200 & \new_[6373]_ ;
  assign \new_[6378]_  = ~A302 & ~A301;
  assign \new_[6379]_  = ~A300 & \new_[6378]_ ;
  assign \new_[6380]_  = \new_[6379]_  & \new_[6374]_ ;
  assign \new_[6383]_  = A168 & A169;
  assign \new_[6387]_  = A199 & ~A166;
  assign \new_[6388]_  = A167 & \new_[6387]_ ;
  assign \new_[6389]_  = \new_[6388]_  & \new_[6383]_ ;
  assign \new_[6393]_  = A299 & ~A298;
  assign \new_[6394]_  = A200 & \new_[6393]_ ;
  assign \new_[6398]_  = ~A302 & ~A301;
  assign \new_[6399]_  = ~A300 & \new_[6398]_ ;
  assign \new_[6400]_  = \new_[6399]_  & \new_[6394]_ ;
  assign \new_[6403]_  = A168 & A169;
  assign \new_[6407]_  = ~A199 & ~A166;
  assign \new_[6408]_  = A167 & \new_[6407]_ ;
  assign \new_[6409]_  = \new_[6408]_  & \new_[6403]_ ;
  assign \new_[6413]_  = ~A299 & A298;
  assign \new_[6414]_  = ~A200 & \new_[6413]_ ;
  assign \new_[6418]_  = ~A302 & ~A301;
  assign \new_[6419]_  = ~A300 & \new_[6418]_ ;
  assign \new_[6420]_  = \new_[6419]_  & \new_[6414]_ ;
  assign \new_[6423]_  = A168 & A169;
  assign \new_[6427]_  = ~A199 & ~A166;
  assign \new_[6428]_  = A167 & \new_[6427]_ ;
  assign \new_[6429]_  = \new_[6428]_  & \new_[6423]_ ;
  assign \new_[6433]_  = A299 & ~A298;
  assign \new_[6434]_  = ~A200 & \new_[6433]_ ;
  assign \new_[6438]_  = ~A302 & ~A301;
  assign \new_[6439]_  = ~A300 & \new_[6438]_ ;
  assign \new_[6440]_  = \new_[6439]_  & \new_[6434]_ ;
  assign \new_[6443]_  = A168 & A169;
  assign \new_[6447]_  = A201 & A166;
  assign \new_[6448]_  = ~A167 & \new_[6447]_ ;
  assign \new_[6449]_  = \new_[6448]_  & \new_[6443]_ ;
  assign \new_[6453]_  = A298 & ~A203;
  assign \new_[6454]_  = ~A202 & \new_[6453]_ ;
  assign \new_[6458]_  = A301 & A300;
  assign \new_[6459]_  = ~A299 & \new_[6458]_ ;
  assign \new_[6460]_  = \new_[6459]_  & \new_[6454]_ ;
  assign \new_[6463]_  = A168 & A169;
  assign \new_[6467]_  = A201 & A166;
  assign \new_[6468]_  = ~A167 & \new_[6467]_ ;
  assign \new_[6469]_  = \new_[6468]_  & \new_[6463]_ ;
  assign \new_[6473]_  = A298 & ~A203;
  assign \new_[6474]_  = ~A202 & \new_[6473]_ ;
  assign \new_[6478]_  = A302 & A300;
  assign \new_[6479]_  = ~A299 & \new_[6478]_ ;
  assign \new_[6480]_  = \new_[6479]_  & \new_[6474]_ ;
  assign \new_[6483]_  = A168 & A169;
  assign \new_[6487]_  = A201 & A166;
  assign \new_[6488]_  = ~A167 & \new_[6487]_ ;
  assign \new_[6489]_  = \new_[6488]_  & \new_[6483]_ ;
  assign \new_[6493]_  = ~A298 & ~A203;
  assign \new_[6494]_  = ~A202 & \new_[6493]_ ;
  assign \new_[6498]_  = A301 & A300;
  assign \new_[6499]_  = A299 & \new_[6498]_ ;
  assign \new_[6500]_  = \new_[6499]_  & \new_[6494]_ ;
  assign \new_[6503]_  = A168 & A169;
  assign \new_[6507]_  = A201 & A166;
  assign \new_[6508]_  = ~A167 & \new_[6507]_ ;
  assign \new_[6509]_  = \new_[6508]_  & \new_[6503]_ ;
  assign \new_[6513]_  = ~A298 & ~A203;
  assign \new_[6514]_  = ~A202 & \new_[6513]_ ;
  assign \new_[6518]_  = A302 & A300;
  assign \new_[6519]_  = A299 & \new_[6518]_ ;
  assign \new_[6520]_  = \new_[6519]_  & \new_[6514]_ ;
  assign \new_[6523]_  = A168 & A169;
  assign \new_[6527]_  = ~A201 & A166;
  assign \new_[6528]_  = ~A167 & \new_[6527]_ ;
  assign \new_[6529]_  = \new_[6528]_  & \new_[6523]_ ;
  assign \new_[6533]_  = ~A299 & A298;
  assign \new_[6534]_  = A202 & \new_[6533]_ ;
  assign \new_[6538]_  = ~A302 & ~A301;
  assign \new_[6539]_  = ~A300 & \new_[6538]_ ;
  assign \new_[6540]_  = \new_[6539]_  & \new_[6534]_ ;
  assign \new_[6543]_  = A168 & A169;
  assign \new_[6547]_  = ~A201 & A166;
  assign \new_[6548]_  = ~A167 & \new_[6547]_ ;
  assign \new_[6549]_  = \new_[6548]_  & \new_[6543]_ ;
  assign \new_[6553]_  = A299 & ~A298;
  assign \new_[6554]_  = A202 & \new_[6553]_ ;
  assign \new_[6558]_  = ~A302 & ~A301;
  assign \new_[6559]_  = ~A300 & \new_[6558]_ ;
  assign \new_[6560]_  = \new_[6559]_  & \new_[6554]_ ;
  assign \new_[6563]_  = A168 & A169;
  assign \new_[6567]_  = ~A201 & A166;
  assign \new_[6568]_  = ~A167 & \new_[6567]_ ;
  assign \new_[6569]_  = \new_[6568]_  & \new_[6563]_ ;
  assign \new_[6573]_  = ~A299 & A298;
  assign \new_[6574]_  = A203 & \new_[6573]_ ;
  assign \new_[6578]_  = ~A302 & ~A301;
  assign \new_[6579]_  = ~A300 & \new_[6578]_ ;
  assign \new_[6580]_  = \new_[6579]_  & \new_[6574]_ ;
  assign \new_[6583]_  = A168 & A169;
  assign \new_[6587]_  = ~A201 & A166;
  assign \new_[6588]_  = ~A167 & \new_[6587]_ ;
  assign \new_[6589]_  = \new_[6588]_  & \new_[6583]_ ;
  assign \new_[6593]_  = A299 & ~A298;
  assign \new_[6594]_  = A203 & \new_[6593]_ ;
  assign \new_[6598]_  = ~A302 & ~A301;
  assign \new_[6599]_  = ~A300 & \new_[6598]_ ;
  assign \new_[6600]_  = \new_[6599]_  & \new_[6594]_ ;
  assign \new_[6603]_  = A168 & A169;
  assign \new_[6607]_  = A199 & A166;
  assign \new_[6608]_  = ~A167 & \new_[6607]_ ;
  assign \new_[6609]_  = \new_[6608]_  & \new_[6603]_ ;
  assign \new_[6613]_  = ~A299 & A298;
  assign \new_[6614]_  = A200 & \new_[6613]_ ;
  assign \new_[6618]_  = ~A302 & ~A301;
  assign \new_[6619]_  = ~A300 & \new_[6618]_ ;
  assign \new_[6620]_  = \new_[6619]_  & \new_[6614]_ ;
  assign \new_[6623]_  = A168 & A169;
  assign \new_[6627]_  = A199 & A166;
  assign \new_[6628]_  = ~A167 & \new_[6627]_ ;
  assign \new_[6629]_  = \new_[6628]_  & \new_[6623]_ ;
  assign \new_[6633]_  = A299 & ~A298;
  assign \new_[6634]_  = A200 & \new_[6633]_ ;
  assign \new_[6638]_  = ~A302 & ~A301;
  assign \new_[6639]_  = ~A300 & \new_[6638]_ ;
  assign \new_[6640]_  = \new_[6639]_  & \new_[6634]_ ;
  assign \new_[6643]_  = A168 & A169;
  assign \new_[6647]_  = ~A199 & A166;
  assign \new_[6648]_  = ~A167 & \new_[6647]_ ;
  assign \new_[6649]_  = \new_[6648]_  & \new_[6643]_ ;
  assign \new_[6653]_  = ~A299 & A298;
  assign \new_[6654]_  = ~A200 & \new_[6653]_ ;
  assign \new_[6658]_  = ~A302 & ~A301;
  assign \new_[6659]_  = ~A300 & \new_[6658]_ ;
  assign \new_[6660]_  = \new_[6659]_  & \new_[6654]_ ;
  assign \new_[6663]_  = A168 & A169;
  assign \new_[6667]_  = ~A199 & A166;
  assign \new_[6668]_  = ~A167 & \new_[6667]_ ;
  assign \new_[6669]_  = \new_[6668]_  & \new_[6663]_ ;
  assign \new_[6673]_  = A299 & ~A298;
  assign \new_[6674]_  = ~A200 & \new_[6673]_ ;
  assign \new_[6678]_  = ~A302 & ~A301;
  assign \new_[6679]_  = ~A300 & \new_[6678]_ ;
  assign \new_[6680]_  = \new_[6679]_  & \new_[6674]_ ;
  assign \new_[6683]_  = ~A168 & A169;
  assign \new_[6687]_  = A201 & A200;
  assign \new_[6688]_  = ~A199 & \new_[6687]_ ;
  assign \new_[6689]_  = \new_[6688]_  & \new_[6683]_ ;
  assign \new_[6693]_  = ~A299 & A298;
  assign \new_[6694]_  = A202 & \new_[6693]_ ;
  assign \new_[6698]_  = ~A302 & ~A301;
  assign \new_[6699]_  = ~A300 & \new_[6698]_ ;
  assign \new_[6700]_  = \new_[6699]_  & \new_[6694]_ ;
  assign \new_[6703]_  = ~A168 & A169;
  assign \new_[6707]_  = A201 & A200;
  assign \new_[6708]_  = ~A199 & \new_[6707]_ ;
  assign \new_[6709]_  = \new_[6708]_  & \new_[6703]_ ;
  assign \new_[6713]_  = A299 & ~A298;
  assign \new_[6714]_  = A202 & \new_[6713]_ ;
  assign \new_[6718]_  = ~A302 & ~A301;
  assign \new_[6719]_  = ~A300 & \new_[6718]_ ;
  assign \new_[6720]_  = \new_[6719]_  & \new_[6714]_ ;
  assign \new_[6723]_  = ~A168 & A169;
  assign \new_[6727]_  = A201 & A200;
  assign \new_[6728]_  = ~A199 & \new_[6727]_ ;
  assign \new_[6729]_  = \new_[6728]_  & \new_[6723]_ ;
  assign \new_[6733]_  = ~A299 & A298;
  assign \new_[6734]_  = A203 & \new_[6733]_ ;
  assign \new_[6738]_  = ~A302 & ~A301;
  assign \new_[6739]_  = ~A300 & \new_[6738]_ ;
  assign \new_[6740]_  = \new_[6739]_  & \new_[6734]_ ;
  assign \new_[6743]_  = ~A168 & A169;
  assign \new_[6747]_  = A201 & A200;
  assign \new_[6748]_  = ~A199 & \new_[6747]_ ;
  assign \new_[6749]_  = \new_[6748]_  & \new_[6743]_ ;
  assign \new_[6753]_  = A299 & ~A298;
  assign \new_[6754]_  = A203 & \new_[6753]_ ;
  assign \new_[6758]_  = ~A302 & ~A301;
  assign \new_[6759]_  = ~A300 & \new_[6758]_ ;
  assign \new_[6760]_  = \new_[6759]_  & \new_[6754]_ ;
  assign \new_[6763]_  = ~A168 & A169;
  assign \new_[6767]_  = ~A201 & A200;
  assign \new_[6768]_  = ~A199 & \new_[6767]_ ;
  assign \new_[6769]_  = \new_[6768]_  & \new_[6763]_ ;
  assign \new_[6773]_  = A298 & ~A203;
  assign \new_[6774]_  = ~A202 & \new_[6773]_ ;
  assign \new_[6778]_  = A301 & A300;
  assign \new_[6779]_  = ~A299 & \new_[6778]_ ;
  assign \new_[6780]_  = \new_[6779]_  & \new_[6774]_ ;
  assign \new_[6783]_  = ~A168 & A169;
  assign \new_[6787]_  = ~A201 & A200;
  assign \new_[6788]_  = ~A199 & \new_[6787]_ ;
  assign \new_[6789]_  = \new_[6788]_  & \new_[6783]_ ;
  assign \new_[6793]_  = A298 & ~A203;
  assign \new_[6794]_  = ~A202 & \new_[6793]_ ;
  assign \new_[6798]_  = A302 & A300;
  assign \new_[6799]_  = ~A299 & \new_[6798]_ ;
  assign \new_[6800]_  = \new_[6799]_  & \new_[6794]_ ;
  assign \new_[6803]_  = ~A168 & A169;
  assign \new_[6807]_  = ~A201 & A200;
  assign \new_[6808]_  = ~A199 & \new_[6807]_ ;
  assign \new_[6809]_  = \new_[6808]_  & \new_[6803]_ ;
  assign \new_[6813]_  = ~A298 & ~A203;
  assign \new_[6814]_  = ~A202 & \new_[6813]_ ;
  assign \new_[6818]_  = A301 & A300;
  assign \new_[6819]_  = A299 & \new_[6818]_ ;
  assign \new_[6820]_  = \new_[6819]_  & \new_[6814]_ ;
  assign \new_[6823]_  = ~A168 & A169;
  assign \new_[6827]_  = ~A201 & A200;
  assign \new_[6828]_  = ~A199 & \new_[6827]_ ;
  assign \new_[6829]_  = \new_[6828]_  & \new_[6823]_ ;
  assign \new_[6833]_  = ~A298 & ~A203;
  assign \new_[6834]_  = ~A202 & \new_[6833]_ ;
  assign \new_[6838]_  = A302 & A300;
  assign \new_[6839]_  = A299 & \new_[6838]_ ;
  assign \new_[6840]_  = \new_[6839]_  & \new_[6834]_ ;
  assign \new_[6843]_  = ~A168 & A169;
  assign \new_[6847]_  = A201 & ~A200;
  assign \new_[6848]_  = A199 & \new_[6847]_ ;
  assign \new_[6849]_  = \new_[6848]_  & \new_[6843]_ ;
  assign \new_[6853]_  = ~A299 & A298;
  assign \new_[6854]_  = A202 & \new_[6853]_ ;
  assign \new_[6858]_  = ~A302 & ~A301;
  assign \new_[6859]_  = ~A300 & \new_[6858]_ ;
  assign \new_[6860]_  = \new_[6859]_  & \new_[6854]_ ;
  assign \new_[6863]_  = ~A168 & A169;
  assign \new_[6867]_  = A201 & ~A200;
  assign \new_[6868]_  = A199 & \new_[6867]_ ;
  assign \new_[6869]_  = \new_[6868]_  & \new_[6863]_ ;
  assign \new_[6873]_  = A299 & ~A298;
  assign \new_[6874]_  = A202 & \new_[6873]_ ;
  assign \new_[6878]_  = ~A302 & ~A301;
  assign \new_[6879]_  = ~A300 & \new_[6878]_ ;
  assign \new_[6880]_  = \new_[6879]_  & \new_[6874]_ ;
  assign \new_[6883]_  = ~A168 & A169;
  assign \new_[6887]_  = A201 & ~A200;
  assign \new_[6888]_  = A199 & \new_[6887]_ ;
  assign \new_[6889]_  = \new_[6888]_  & \new_[6883]_ ;
  assign \new_[6893]_  = ~A299 & A298;
  assign \new_[6894]_  = A203 & \new_[6893]_ ;
  assign \new_[6898]_  = ~A302 & ~A301;
  assign \new_[6899]_  = ~A300 & \new_[6898]_ ;
  assign \new_[6900]_  = \new_[6899]_  & \new_[6894]_ ;
  assign \new_[6903]_  = ~A168 & A169;
  assign \new_[6907]_  = A201 & ~A200;
  assign \new_[6908]_  = A199 & \new_[6907]_ ;
  assign \new_[6909]_  = \new_[6908]_  & \new_[6903]_ ;
  assign \new_[6913]_  = A299 & ~A298;
  assign \new_[6914]_  = A203 & \new_[6913]_ ;
  assign \new_[6918]_  = ~A302 & ~A301;
  assign \new_[6919]_  = ~A300 & \new_[6918]_ ;
  assign \new_[6920]_  = \new_[6919]_  & \new_[6914]_ ;
  assign \new_[6923]_  = ~A168 & A169;
  assign \new_[6927]_  = ~A201 & ~A200;
  assign \new_[6928]_  = A199 & \new_[6927]_ ;
  assign \new_[6929]_  = \new_[6928]_  & \new_[6923]_ ;
  assign \new_[6933]_  = A298 & ~A203;
  assign \new_[6934]_  = ~A202 & \new_[6933]_ ;
  assign \new_[6938]_  = A301 & A300;
  assign \new_[6939]_  = ~A299 & \new_[6938]_ ;
  assign \new_[6940]_  = \new_[6939]_  & \new_[6934]_ ;
  assign \new_[6943]_  = ~A168 & A169;
  assign \new_[6947]_  = ~A201 & ~A200;
  assign \new_[6948]_  = A199 & \new_[6947]_ ;
  assign \new_[6949]_  = \new_[6948]_  & \new_[6943]_ ;
  assign \new_[6953]_  = A298 & ~A203;
  assign \new_[6954]_  = ~A202 & \new_[6953]_ ;
  assign \new_[6958]_  = A302 & A300;
  assign \new_[6959]_  = ~A299 & \new_[6958]_ ;
  assign \new_[6960]_  = \new_[6959]_  & \new_[6954]_ ;
  assign \new_[6963]_  = ~A168 & A169;
  assign \new_[6967]_  = ~A201 & ~A200;
  assign \new_[6968]_  = A199 & \new_[6967]_ ;
  assign \new_[6969]_  = \new_[6968]_  & \new_[6963]_ ;
  assign \new_[6973]_  = ~A298 & ~A203;
  assign \new_[6974]_  = ~A202 & \new_[6973]_ ;
  assign \new_[6978]_  = A301 & A300;
  assign \new_[6979]_  = A299 & \new_[6978]_ ;
  assign \new_[6980]_  = \new_[6979]_  & \new_[6974]_ ;
  assign \new_[6983]_  = ~A168 & A169;
  assign \new_[6987]_  = ~A201 & ~A200;
  assign \new_[6988]_  = A199 & \new_[6987]_ ;
  assign \new_[6989]_  = \new_[6988]_  & \new_[6983]_ ;
  assign \new_[6993]_  = ~A298 & ~A203;
  assign \new_[6994]_  = ~A202 & \new_[6993]_ ;
  assign \new_[6998]_  = A302 & A300;
  assign \new_[6999]_  = A299 & \new_[6998]_ ;
  assign \new_[7000]_  = \new_[6999]_  & \new_[6994]_ ;
  assign \new_[7003]_  = ~A169 & A170;
  assign \new_[7007]_  = A200 & ~A199;
  assign \new_[7008]_  = A168 & \new_[7007]_ ;
  assign \new_[7009]_  = \new_[7008]_  & \new_[7003]_ ;
  assign \new_[7013]_  = A298 & A202;
  assign \new_[7014]_  = A201 & \new_[7013]_ ;
  assign \new_[7018]_  = A301 & A300;
  assign \new_[7019]_  = ~A299 & \new_[7018]_ ;
  assign \new_[7020]_  = \new_[7019]_  & \new_[7014]_ ;
  assign \new_[7023]_  = ~A169 & A170;
  assign \new_[7027]_  = A200 & ~A199;
  assign \new_[7028]_  = A168 & \new_[7027]_ ;
  assign \new_[7029]_  = \new_[7028]_  & \new_[7023]_ ;
  assign \new_[7033]_  = A298 & A202;
  assign \new_[7034]_  = A201 & \new_[7033]_ ;
  assign \new_[7038]_  = A302 & A300;
  assign \new_[7039]_  = ~A299 & \new_[7038]_ ;
  assign \new_[7040]_  = \new_[7039]_  & \new_[7034]_ ;
  assign \new_[7043]_  = ~A169 & A170;
  assign \new_[7047]_  = A200 & ~A199;
  assign \new_[7048]_  = A168 & \new_[7047]_ ;
  assign \new_[7049]_  = \new_[7048]_  & \new_[7043]_ ;
  assign \new_[7053]_  = ~A298 & A202;
  assign \new_[7054]_  = A201 & \new_[7053]_ ;
  assign \new_[7058]_  = A301 & A300;
  assign \new_[7059]_  = A299 & \new_[7058]_ ;
  assign \new_[7060]_  = \new_[7059]_  & \new_[7054]_ ;
  assign \new_[7063]_  = ~A169 & A170;
  assign \new_[7067]_  = A200 & ~A199;
  assign \new_[7068]_  = A168 & \new_[7067]_ ;
  assign \new_[7069]_  = \new_[7068]_  & \new_[7063]_ ;
  assign \new_[7073]_  = ~A298 & A202;
  assign \new_[7074]_  = A201 & \new_[7073]_ ;
  assign \new_[7078]_  = A302 & A300;
  assign \new_[7079]_  = A299 & \new_[7078]_ ;
  assign \new_[7080]_  = \new_[7079]_  & \new_[7074]_ ;
  assign \new_[7083]_  = ~A169 & A170;
  assign \new_[7087]_  = A200 & ~A199;
  assign \new_[7088]_  = A168 & \new_[7087]_ ;
  assign \new_[7089]_  = \new_[7088]_  & \new_[7083]_ ;
  assign \new_[7093]_  = A298 & A203;
  assign \new_[7094]_  = A201 & \new_[7093]_ ;
  assign \new_[7098]_  = A301 & A300;
  assign \new_[7099]_  = ~A299 & \new_[7098]_ ;
  assign \new_[7100]_  = \new_[7099]_  & \new_[7094]_ ;
  assign \new_[7103]_  = ~A169 & A170;
  assign \new_[7107]_  = A200 & ~A199;
  assign \new_[7108]_  = A168 & \new_[7107]_ ;
  assign \new_[7109]_  = \new_[7108]_  & \new_[7103]_ ;
  assign \new_[7113]_  = A298 & A203;
  assign \new_[7114]_  = A201 & \new_[7113]_ ;
  assign \new_[7118]_  = A302 & A300;
  assign \new_[7119]_  = ~A299 & \new_[7118]_ ;
  assign \new_[7120]_  = \new_[7119]_  & \new_[7114]_ ;
  assign \new_[7123]_  = ~A169 & A170;
  assign \new_[7127]_  = A200 & ~A199;
  assign \new_[7128]_  = A168 & \new_[7127]_ ;
  assign \new_[7129]_  = \new_[7128]_  & \new_[7123]_ ;
  assign \new_[7133]_  = ~A298 & A203;
  assign \new_[7134]_  = A201 & \new_[7133]_ ;
  assign \new_[7138]_  = A301 & A300;
  assign \new_[7139]_  = A299 & \new_[7138]_ ;
  assign \new_[7140]_  = \new_[7139]_  & \new_[7134]_ ;
  assign \new_[7143]_  = ~A169 & A170;
  assign \new_[7147]_  = A200 & ~A199;
  assign \new_[7148]_  = A168 & \new_[7147]_ ;
  assign \new_[7149]_  = \new_[7148]_  & \new_[7143]_ ;
  assign \new_[7153]_  = ~A298 & A203;
  assign \new_[7154]_  = A201 & \new_[7153]_ ;
  assign \new_[7158]_  = A302 & A300;
  assign \new_[7159]_  = A299 & \new_[7158]_ ;
  assign \new_[7160]_  = \new_[7159]_  & \new_[7154]_ ;
  assign \new_[7163]_  = ~A169 & A170;
  assign \new_[7167]_  = ~A200 & A199;
  assign \new_[7168]_  = A168 & \new_[7167]_ ;
  assign \new_[7169]_  = \new_[7168]_  & \new_[7163]_ ;
  assign \new_[7173]_  = A298 & A202;
  assign \new_[7174]_  = A201 & \new_[7173]_ ;
  assign \new_[7178]_  = A301 & A300;
  assign \new_[7179]_  = ~A299 & \new_[7178]_ ;
  assign \new_[7180]_  = \new_[7179]_  & \new_[7174]_ ;
  assign \new_[7183]_  = ~A169 & A170;
  assign \new_[7187]_  = ~A200 & A199;
  assign \new_[7188]_  = A168 & \new_[7187]_ ;
  assign \new_[7189]_  = \new_[7188]_  & \new_[7183]_ ;
  assign \new_[7193]_  = A298 & A202;
  assign \new_[7194]_  = A201 & \new_[7193]_ ;
  assign \new_[7198]_  = A302 & A300;
  assign \new_[7199]_  = ~A299 & \new_[7198]_ ;
  assign \new_[7200]_  = \new_[7199]_  & \new_[7194]_ ;
  assign \new_[7203]_  = ~A169 & A170;
  assign \new_[7207]_  = ~A200 & A199;
  assign \new_[7208]_  = A168 & \new_[7207]_ ;
  assign \new_[7209]_  = \new_[7208]_  & \new_[7203]_ ;
  assign \new_[7213]_  = ~A298 & A202;
  assign \new_[7214]_  = A201 & \new_[7213]_ ;
  assign \new_[7218]_  = A301 & A300;
  assign \new_[7219]_  = A299 & \new_[7218]_ ;
  assign \new_[7220]_  = \new_[7219]_  & \new_[7214]_ ;
  assign \new_[7223]_  = ~A169 & A170;
  assign \new_[7227]_  = ~A200 & A199;
  assign \new_[7228]_  = A168 & \new_[7227]_ ;
  assign \new_[7229]_  = \new_[7228]_  & \new_[7223]_ ;
  assign \new_[7233]_  = ~A298 & A202;
  assign \new_[7234]_  = A201 & \new_[7233]_ ;
  assign \new_[7238]_  = A302 & A300;
  assign \new_[7239]_  = A299 & \new_[7238]_ ;
  assign \new_[7240]_  = \new_[7239]_  & \new_[7234]_ ;
  assign \new_[7243]_  = ~A169 & A170;
  assign \new_[7247]_  = ~A200 & A199;
  assign \new_[7248]_  = A168 & \new_[7247]_ ;
  assign \new_[7249]_  = \new_[7248]_  & \new_[7243]_ ;
  assign \new_[7253]_  = A298 & A203;
  assign \new_[7254]_  = A201 & \new_[7253]_ ;
  assign \new_[7258]_  = A301 & A300;
  assign \new_[7259]_  = ~A299 & \new_[7258]_ ;
  assign \new_[7260]_  = \new_[7259]_  & \new_[7254]_ ;
  assign \new_[7263]_  = ~A169 & A170;
  assign \new_[7267]_  = ~A200 & A199;
  assign \new_[7268]_  = A168 & \new_[7267]_ ;
  assign \new_[7269]_  = \new_[7268]_  & \new_[7263]_ ;
  assign \new_[7273]_  = A298 & A203;
  assign \new_[7274]_  = A201 & \new_[7273]_ ;
  assign \new_[7278]_  = A302 & A300;
  assign \new_[7279]_  = ~A299 & \new_[7278]_ ;
  assign \new_[7280]_  = \new_[7279]_  & \new_[7274]_ ;
  assign \new_[7283]_  = ~A169 & A170;
  assign \new_[7287]_  = ~A200 & A199;
  assign \new_[7288]_  = A168 & \new_[7287]_ ;
  assign \new_[7289]_  = \new_[7288]_  & \new_[7283]_ ;
  assign \new_[7293]_  = ~A298 & A203;
  assign \new_[7294]_  = A201 & \new_[7293]_ ;
  assign \new_[7298]_  = A301 & A300;
  assign \new_[7299]_  = A299 & \new_[7298]_ ;
  assign \new_[7300]_  = \new_[7299]_  & \new_[7294]_ ;
  assign \new_[7303]_  = ~A169 & A170;
  assign \new_[7307]_  = ~A200 & A199;
  assign \new_[7308]_  = A168 & \new_[7307]_ ;
  assign \new_[7309]_  = \new_[7308]_  & \new_[7303]_ ;
  assign \new_[7313]_  = ~A298 & A203;
  assign \new_[7314]_  = A201 & \new_[7313]_ ;
  assign \new_[7318]_  = A302 & A300;
  assign \new_[7319]_  = A299 & \new_[7318]_ ;
  assign \new_[7320]_  = \new_[7319]_  & \new_[7314]_ ;
  assign \new_[7323]_  = ~A169 & A170;
  assign \new_[7327]_  = ~A166 & A167;
  assign \new_[7328]_  = ~A168 & \new_[7327]_ ;
  assign \new_[7329]_  = \new_[7328]_  & \new_[7323]_ ;
  assign \new_[7333]_  = A298 & A202;
  assign \new_[7334]_  = ~A201 & \new_[7333]_ ;
  assign \new_[7338]_  = A301 & A300;
  assign \new_[7339]_  = ~A299 & \new_[7338]_ ;
  assign \new_[7340]_  = \new_[7339]_  & \new_[7334]_ ;
  assign \new_[7343]_  = ~A169 & A170;
  assign \new_[7347]_  = ~A166 & A167;
  assign \new_[7348]_  = ~A168 & \new_[7347]_ ;
  assign \new_[7349]_  = \new_[7348]_  & \new_[7343]_ ;
  assign \new_[7353]_  = A298 & A202;
  assign \new_[7354]_  = ~A201 & \new_[7353]_ ;
  assign \new_[7358]_  = A302 & A300;
  assign \new_[7359]_  = ~A299 & \new_[7358]_ ;
  assign \new_[7360]_  = \new_[7359]_  & \new_[7354]_ ;
  assign \new_[7363]_  = ~A169 & A170;
  assign \new_[7367]_  = ~A166 & A167;
  assign \new_[7368]_  = ~A168 & \new_[7367]_ ;
  assign \new_[7369]_  = \new_[7368]_  & \new_[7363]_ ;
  assign \new_[7373]_  = ~A298 & A202;
  assign \new_[7374]_  = ~A201 & \new_[7373]_ ;
  assign \new_[7378]_  = A301 & A300;
  assign \new_[7379]_  = A299 & \new_[7378]_ ;
  assign \new_[7380]_  = \new_[7379]_  & \new_[7374]_ ;
  assign \new_[7383]_  = ~A169 & A170;
  assign \new_[7387]_  = ~A166 & A167;
  assign \new_[7388]_  = ~A168 & \new_[7387]_ ;
  assign \new_[7389]_  = \new_[7388]_  & \new_[7383]_ ;
  assign \new_[7393]_  = ~A298 & A202;
  assign \new_[7394]_  = ~A201 & \new_[7393]_ ;
  assign \new_[7398]_  = A302 & A300;
  assign \new_[7399]_  = A299 & \new_[7398]_ ;
  assign \new_[7400]_  = \new_[7399]_  & \new_[7394]_ ;
  assign \new_[7403]_  = ~A169 & A170;
  assign \new_[7407]_  = ~A166 & A167;
  assign \new_[7408]_  = ~A168 & \new_[7407]_ ;
  assign \new_[7409]_  = \new_[7408]_  & \new_[7403]_ ;
  assign \new_[7413]_  = A298 & A203;
  assign \new_[7414]_  = ~A201 & \new_[7413]_ ;
  assign \new_[7418]_  = A301 & A300;
  assign \new_[7419]_  = ~A299 & \new_[7418]_ ;
  assign \new_[7420]_  = \new_[7419]_  & \new_[7414]_ ;
  assign \new_[7423]_  = ~A169 & A170;
  assign \new_[7427]_  = ~A166 & A167;
  assign \new_[7428]_  = ~A168 & \new_[7427]_ ;
  assign \new_[7429]_  = \new_[7428]_  & \new_[7423]_ ;
  assign \new_[7433]_  = A298 & A203;
  assign \new_[7434]_  = ~A201 & \new_[7433]_ ;
  assign \new_[7438]_  = A302 & A300;
  assign \new_[7439]_  = ~A299 & \new_[7438]_ ;
  assign \new_[7440]_  = \new_[7439]_  & \new_[7434]_ ;
  assign \new_[7443]_  = ~A169 & A170;
  assign \new_[7447]_  = ~A166 & A167;
  assign \new_[7448]_  = ~A168 & \new_[7447]_ ;
  assign \new_[7449]_  = \new_[7448]_  & \new_[7443]_ ;
  assign \new_[7453]_  = ~A298 & A203;
  assign \new_[7454]_  = ~A201 & \new_[7453]_ ;
  assign \new_[7458]_  = A301 & A300;
  assign \new_[7459]_  = A299 & \new_[7458]_ ;
  assign \new_[7460]_  = \new_[7459]_  & \new_[7454]_ ;
  assign \new_[7463]_  = ~A169 & A170;
  assign \new_[7467]_  = ~A166 & A167;
  assign \new_[7468]_  = ~A168 & \new_[7467]_ ;
  assign \new_[7469]_  = \new_[7468]_  & \new_[7463]_ ;
  assign \new_[7473]_  = ~A298 & A203;
  assign \new_[7474]_  = ~A201 & \new_[7473]_ ;
  assign \new_[7478]_  = A302 & A300;
  assign \new_[7479]_  = A299 & \new_[7478]_ ;
  assign \new_[7480]_  = \new_[7479]_  & \new_[7474]_ ;
  assign \new_[7483]_  = ~A169 & A170;
  assign \new_[7487]_  = ~A166 & A167;
  assign \new_[7488]_  = ~A168 & \new_[7487]_ ;
  assign \new_[7489]_  = \new_[7488]_  & \new_[7483]_ ;
  assign \new_[7493]_  = A298 & A200;
  assign \new_[7494]_  = A199 & \new_[7493]_ ;
  assign \new_[7498]_  = A301 & A300;
  assign \new_[7499]_  = ~A299 & \new_[7498]_ ;
  assign \new_[7500]_  = \new_[7499]_  & \new_[7494]_ ;
  assign \new_[7503]_  = ~A169 & A170;
  assign \new_[7507]_  = ~A166 & A167;
  assign \new_[7508]_  = ~A168 & \new_[7507]_ ;
  assign \new_[7509]_  = \new_[7508]_  & \new_[7503]_ ;
  assign \new_[7513]_  = A298 & A200;
  assign \new_[7514]_  = A199 & \new_[7513]_ ;
  assign \new_[7518]_  = A302 & A300;
  assign \new_[7519]_  = ~A299 & \new_[7518]_ ;
  assign \new_[7520]_  = \new_[7519]_  & \new_[7514]_ ;
  assign \new_[7523]_  = ~A169 & A170;
  assign \new_[7527]_  = ~A166 & A167;
  assign \new_[7528]_  = ~A168 & \new_[7527]_ ;
  assign \new_[7529]_  = \new_[7528]_  & \new_[7523]_ ;
  assign \new_[7533]_  = ~A298 & A200;
  assign \new_[7534]_  = A199 & \new_[7533]_ ;
  assign \new_[7538]_  = A301 & A300;
  assign \new_[7539]_  = A299 & \new_[7538]_ ;
  assign \new_[7540]_  = \new_[7539]_  & \new_[7534]_ ;
  assign \new_[7543]_  = ~A169 & A170;
  assign \new_[7547]_  = ~A166 & A167;
  assign \new_[7548]_  = ~A168 & \new_[7547]_ ;
  assign \new_[7549]_  = \new_[7548]_  & \new_[7543]_ ;
  assign \new_[7553]_  = ~A298 & A200;
  assign \new_[7554]_  = A199 & \new_[7553]_ ;
  assign \new_[7558]_  = A302 & A300;
  assign \new_[7559]_  = A299 & \new_[7558]_ ;
  assign \new_[7560]_  = \new_[7559]_  & \new_[7554]_ ;
  assign \new_[7563]_  = ~A169 & A170;
  assign \new_[7567]_  = ~A166 & A167;
  assign \new_[7568]_  = ~A168 & \new_[7567]_ ;
  assign \new_[7569]_  = \new_[7568]_  & \new_[7563]_ ;
  assign \new_[7573]_  = A298 & ~A200;
  assign \new_[7574]_  = ~A199 & \new_[7573]_ ;
  assign \new_[7578]_  = A301 & A300;
  assign \new_[7579]_  = ~A299 & \new_[7578]_ ;
  assign \new_[7580]_  = \new_[7579]_  & \new_[7574]_ ;
  assign \new_[7583]_  = ~A169 & A170;
  assign \new_[7587]_  = ~A166 & A167;
  assign \new_[7588]_  = ~A168 & \new_[7587]_ ;
  assign \new_[7589]_  = \new_[7588]_  & \new_[7583]_ ;
  assign \new_[7593]_  = A298 & ~A200;
  assign \new_[7594]_  = ~A199 & \new_[7593]_ ;
  assign \new_[7598]_  = A302 & A300;
  assign \new_[7599]_  = ~A299 & \new_[7598]_ ;
  assign \new_[7600]_  = \new_[7599]_  & \new_[7594]_ ;
  assign \new_[7603]_  = ~A169 & A170;
  assign \new_[7607]_  = ~A166 & A167;
  assign \new_[7608]_  = ~A168 & \new_[7607]_ ;
  assign \new_[7609]_  = \new_[7608]_  & \new_[7603]_ ;
  assign \new_[7613]_  = ~A298 & ~A200;
  assign \new_[7614]_  = ~A199 & \new_[7613]_ ;
  assign \new_[7618]_  = A301 & A300;
  assign \new_[7619]_  = A299 & \new_[7618]_ ;
  assign \new_[7620]_  = \new_[7619]_  & \new_[7614]_ ;
  assign \new_[7623]_  = ~A169 & A170;
  assign \new_[7627]_  = ~A166 & A167;
  assign \new_[7628]_  = ~A168 & \new_[7627]_ ;
  assign \new_[7629]_  = \new_[7628]_  & \new_[7623]_ ;
  assign \new_[7633]_  = ~A298 & ~A200;
  assign \new_[7634]_  = ~A199 & \new_[7633]_ ;
  assign \new_[7638]_  = A302 & A300;
  assign \new_[7639]_  = A299 & \new_[7638]_ ;
  assign \new_[7640]_  = \new_[7639]_  & \new_[7634]_ ;
  assign \new_[7643]_  = ~A169 & A170;
  assign \new_[7647]_  = A166 & ~A167;
  assign \new_[7648]_  = ~A168 & \new_[7647]_ ;
  assign \new_[7649]_  = \new_[7648]_  & \new_[7643]_ ;
  assign \new_[7653]_  = A298 & A202;
  assign \new_[7654]_  = ~A201 & \new_[7653]_ ;
  assign \new_[7658]_  = A301 & A300;
  assign \new_[7659]_  = ~A299 & \new_[7658]_ ;
  assign \new_[7660]_  = \new_[7659]_  & \new_[7654]_ ;
  assign \new_[7663]_  = ~A169 & A170;
  assign \new_[7667]_  = A166 & ~A167;
  assign \new_[7668]_  = ~A168 & \new_[7667]_ ;
  assign \new_[7669]_  = \new_[7668]_  & \new_[7663]_ ;
  assign \new_[7673]_  = A298 & A202;
  assign \new_[7674]_  = ~A201 & \new_[7673]_ ;
  assign \new_[7678]_  = A302 & A300;
  assign \new_[7679]_  = ~A299 & \new_[7678]_ ;
  assign \new_[7680]_  = \new_[7679]_  & \new_[7674]_ ;
  assign \new_[7683]_  = ~A169 & A170;
  assign \new_[7687]_  = A166 & ~A167;
  assign \new_[7688]_  = ~A168 & \new_[7687]_ ;
  assign \new_[7689]_  = \new_[7688]_  & \new_[7683]_ ;
  assign \new_[7693]_  = ~A298 & A202;
  assign \new_[7694]_  = ~A201 & \new_[7693]_ ;
  assign \new_[7698]_  = A301 & A300;
  assign \new_[7699]_  = A299 & \new_[7698]_ ;
  assign \new_[7700]_  = \new_[7699]_  & \new_[7694]_ ;
  assign \new_[7703]_  = ~A169 & A170;
  assign \new_[7707]_  = A166 & ~A167;
  assign \new_[7708]_  = ~A168 & \new_[7707]_ ;
  assign \new_[7709]_  = \new_[7708]_  & \new_[7703]_ ;
  assign \new_[7713]_  = ~A298 & A202;
  assign \new_[7714]_  = ~A201 & \new_[7713]_ ;
  assign \new_[7718]_  = A302 & A300;
  assign \new_[7719]_  = A299 & \new_[7718]_ ;
  assign \new_[7720]_  = \new_[7719]_  & \new_[7714]_ ;
  assign \new_[7723]_  = ~A169 & A170;
  assign \new_[7727]_  = A166 & ~A167;
  assign \new_[7728]_  = ~A168 & \new_[7727]_ ;
  assign \new_[7729]_  = \new_[7728]_  & \new_[7723]_ ;
  assign \new_[7733]_  = A298 & A203;
  assign \new_[7734]_  = ~A201 & \new_[7733]_ ;
  assign \new_[7738]_  = A301 & A300;
  assign \new_[7739]_  = ~A299 & \new_[7738]_ ;
  assign \new_[7740]_  = \new_[7739]_  & \new_[7734]_ ;
  assign \new_[7743]_  = ~A169 & A170;
  assign \new_[7747]_  = A166 & ~A167;
  assign \new_[7748]_  = ~A168 & \new_[7747]_ ;
  assign \new_[7749]_  = \new_[7748]_  & \new_[7743]_ ;
  assign \new_[7753]_  = A298 & A203;
  assign \new_[7754]_  = ~A201 & \new_[7753]_ ;
  assign \new_[7758]_  = A302 & A300;
  assign \new_[7759]_  = ~A299 & \new_[7758]_ ;
  assign \new_[7760]_  = \new_[7759]_  & \new_[7754]_ ;
  assign \new_[7763]_  = ~A169 & A170;
  assign \new_[7767]_  = A166 & ~A167;
  assign \new_[7768]_  = ~A168 & \new_[7767]_ ;
  assign \new_[7769]_  = \new_[7768]_  & \new_[7763]_ ;
  assign \new_[7773]_  = ~A298 & A203;
  assign \new_[7774]_  = ~A201 & \new_[7773]_ ;
  assign \new_[7778]_  = A301 & A300;
  assign \new_[7779]_  = A299 & \new_[7778]_ ;
  assign \new_[7780]_  = \new_[7779]_  & \new_[7774]_ ;
  assign \new_[7783]_  = ~A169 & A170;
  assign \new_[7787]_  = A166 & ~A167;
  assign \new_[7788]_  = ~A168 & \new_[7787]_ ;
  assign \new_[7789]_  = \new_[7788]_  & \new_[7783]_ ;
  assign \new_[7793]_  = ~A298 & A203;
  assign \new_[7794]_  = ~A201 & \new_[7793]_ ;
  assign \new_[7798]_  = A302 & A300;
  assign \new_[7799]_  = A299 & \new_[7798]_ ;
  assign \new_[7800]_  = \new_[7799]_  & \new_[7794]_ ;
  assign \new_[7803]_  = ~A169 & A170;
  assign \new_[7807]_  = A166 & ~A167;
  assign \new_[7808]_  = ~A168 & \new_[7807]_ ;
  assign \new_[7809]_  = \new_[7808]_  & \new_[7803]_ ;
  assign \new_[7813]_  = A298 & A200;
  assign \new_[7814]_  = A199 & \new_[7813]_ ;
  assign \new_[7818]_  = A301 & A300;
  assign \new_[7819]_  = ~A299 & \new_[7818]_ ;
  assign \new_[7820]_  = \new_[7819]_  & \new_[7814]_ ;
  assign \new_[7823]_  = ~A169 & A170;
  assign \new_[7827]_  = A166 & ~A167;
  assign \new_[7828]_  = ~A168 & \new_[7827]_ ;
  assign \new_[7829]_  = \new_[7828]_  & \new_[7823]_ ;
  assign \new_[7833]_  = A298 & A200;
  assign \new_[7834]_  = A199 & \new_[7833]_ ;
  assign \new_[7838]_  = A302 & A300;
  assign \new_[7839]_  = ~A299 & \new_[7838]_ ;
  assign \new_[7840]_  = \new_[7839]_  & \new_[7834]_ ;
  assign \new_[7843]_  = ~A169 & A170;
  assign \new_[7847]_  = A166 & ~A167;
  assign \new_[7848]_  = ~A168 & \new_[7847]_ ;
  assign \new_[7849]_  = \new_[7848]_  & \new_[7843]_ ;
  assign \new_[7853]_  = ~A298 & A200;
  assign \new_[7854]_  = A199 & \new_[7853]_ ;
  assign \new_[7858]_  = A301 & A300;
  assign \new_[7859]_  = A299 & \new_[7858]_ ;
  assign \new_[7860]_  = \new_[7859]_  & \new_[7854]_ ;
  assign \new_[7863]_  = ~A169 & A170;
  assign \new_[7867]_  = A166 & ~A167;
  assign \new_[7868]_  = ~A168 & \new_[7867]_ ;
  assign \new_[7869]_  = \new_[7868]_  & \new_[7863]_ ;
  assign \new_[7873]_  = ~A298 & A200;
  assign \new_[7874]_  = A199 & \new_[7873]_ ;
  assign \new_[7878]_  = A302 & A300;
  assign \new_[7879]_  = A299 & \new_[7878]_ ;
  assign \new_[7880]_  = \new_[7879]_  & \new_[7874]_ ;
  assign \new_[7883]_  = ~A169 & A170;
  assign \new_[7887]_  = A166 & ~A167;
  assign \new_[7888]_  = ~A168 & \new_[7887]_ ;
  assign \new_[7889]_  = \new_[7888]_  & \new_[7883]_ ;
  assign \new_[7893]_  = A298 & ~A200;
  assign \new_[7894]_  = ~A199 & \new_[7893]_ ;
  assign \new_[7898]_  = A301 & A300;
  assign \new_[7899]_  = ~A299 & \new_[7898]_ ;
  assign \new_[7900]_  = \new_[7899]_  & \new_[7894]_ ;
  assign \new_[7903]_  = ~A169 & A170;
  assign \new_[7907]_  = A166 & ~A167;
  assign \new_[7908]_  = ~A168 & \new_[7907]_ ;
  assign \new_[7909]_  = \new_[7908]_  & \new_[7903]_ ;
  assign \new_[7913]_  = A298 & ~A200;
  assign \new_[7914]_  = ~A199 & \new_[7913]_ ;
  assign \new_[7918]_  = A302 & A300;
  assign \new_[7919]_  = ~A299 & \new_[7918]_ ;
  assign \new_[7920]_  = \new_[7919]_  & \new_[7914]_ ;
  assign \new_[7923]_  = ~A169 & A170;
  assign \new_[7927]_  = A166 & ~A167;
  assign \new_[7928]_  = ~A168 & \new_[7927]_ ;
  assign \new_[7929]_  = \new_[7928]_  & \new_[7923]_ ;
  assign \new_[7933]_  = ~A298 & ~A200;
  assign \new_[7934]_  = ~A199 & \new_[7933]_ ;
  assign \new_[7938]_  = A301 & A300;
  assign \new_[7939]_  = A299 & \new_[7938]_ ;
  assign \new_[7940]_  = \new_[7939]_  & \new_[7934]_ ;
  assign \new_[7943]_  = ~A169 & A170;
  assign \new_[7947]_  = A166 & ~A167;
  assign \new_[7948]_  = ~A168 & \new_[7947]_ ;
  assign \new_[7949]_  = \new_[7948]_  & \new_[7943]_ ;
  assign \new_[7953]_  = ~A298 & ~A200;
  assign \new_[7954]_  = ~A199 & \new_[7953]_ ;
  assign \new_[7958]_  = A302 & A300;
  assign \new_[7959]_  = A299 & \new_[7958]_ ;
  assign \new_[7960]_  = \new_[7959]_  & \new_[7954]_ ;
  assign \new_[7964]_  = ~A199 & A166;
  assign \new_[7965]_  = A167 & \new_[7964]_ ;
  assign \new_[7969]_  = ~A202 & ~A201;
  assign \new_[7970]_  = A200 & \new_[7969]_ ;
  assign \new_[7971]_  = \new_[7970]_  & \new_[7965]_ ;
  assign \new_[7975]_  = ~A299 & A298;
  assign \new_[7976]_  = ~A203 & \new_[7975]_ ;
  assign \new_[7980]_  = ~A302 & ~A301;
  assign \new_[7981]_  = ~A300 & \new_[7980]_ ;
  assign \new_[7982]_  = \new_[7981]_  & \new_[7976]_ ;
  assign \new_[7986]_  = ~A199 & A166;
  assign \new_[7987]_  = A167 & \new_[7986]_ ;
  assign \new_[7991]_  = ~A202 & ~A201;
  assign \new_[7992]_  = A200 & \new_[7991]_ ;
  assign \new_[7993]_  = \new_[7992]_  & \new_[7987]_ ;
  assign \new_[7997]_  = A299 & ~A298;
  assign \new_[7998]_  = ~A203 & \new_[7997]_ ;
  assign \new_[8002]_  = ~A302 & ~A301;
  assign \new_[8003]_  = ~A300 & \new_[8002]_ ;
  assign \new_[8004]_  = \new_[8003]_  & \new_[7998]_ ;
  assign \new_[8008]_  = A199 & A166;
  assign \new_[8009]_  = A167 & \new_[8008]_ ;
  assign \new_[8013]_  = ~A202 & ~A201;
  assign \new_[8014]_  = ~A200 & \new_[8013]_ ;
  assign \new_[8015]_  = \new_[8014]_  & \new_[8009]_ ;
  assign \new_[8019]_  = ~A299 & A298;
  assign \new_[8020]_  = ~A203 & \new_[8019]_ ;
  assign \new_[8024]_  = ~A302 & ~A301;
  assign \new_[8025]_  = ~A300 & \new_[8024]_ ;
  assign \new_[8026]_  = \new_[8025]_  & \new_[8020]_ ;
  assign \new_[8030]_  = A199 & A166;
  assign \new_[8031]_  = A167 & \new_[8030]_ ;
  assign \new_[8035]_  = ~A202 & ~A201;
  assign \new_[8036]_  = ~A200 & \new_[8035]_ ;
  assign \new_[8037]_  = \new_[8036]_  & \new_[8031]_ ;
  assign \new_[8041]_  = A299 & ~A298;
  assign \new_[8042]_  = ~A203 & \new_[8041]_ ;
  assign \new_[8046]_  = ~A302 & ~A301;
  assign \new_[8047]_  = ~A300 & \new_[8046]_ ;
  assign \new_[8048]_  = \new_[8047]_  & \new_[8042]_ ;
  assign \new_[8052]_  = ~A199 & ~A166;
  assign \new_[8053]_  = ~A167 & \new_[8052]_ ;
  assign \new_[8057]_  = ~A202 & ~A201;
  assign \new_[8058]_  = A200 & \new_[8057]_ ;
  assign \new_[8059]_  = \new_[8058]_  & \new_[8053]_ ;
  assign \new_[8063]_  = ~A299 & A298;
  assign \new_[8064]_  = ~A203 & \new_[8063]_ ;
  assign \new_[8068]_  = ~A302 & ~A301;
  assign \new_[8069]_  = ~A300 & \new_[8068]_ ;
  assign \new_[8070]_  = \new_[8069]_  & \new_[8064]_ ;
  assign \new_[8074]_  = ~A199 & ~A166;
  assign \new_[8075]_  = ~A167 & \new_[8074]_ ;
  assign \new_[8079]_  = ~A202 & ~A201;
  assign \new_[8080]_  = A200 & \new_[8079]_ ;
  assign \new_[8081]_  = \new_[8080]_  & \new_[8075]_ ;
  assign \new_[8085]_  = A299 & ~A298;
  assign \new_[8086]_  = ~A203 & \new_[8085]_ ;
  assign \new_[8090]_  = ~A302 & ~A301;
  assign \new_[8091]_  = ~A300 & \new_[8090]_ ;
  assign \new_[8092]_  = \new_[8091]_  & \new_[8086]_ ;
  assign \new_[8096]_  = A199 & ~A166;
  assign \new_[8097]_  = ~A167 & \new_[8096]_ ;
  assign \new_[8101]_  = ~A202 & ~A201;
  assign \new_[8102]_  = ~A200 & \new_[8101]_ ;
  assign \new_[8103]_  = \new_[8102]_  & \new_[8097]_ ;
  assign \new_[8107]_  = ~A299 & A298;
  assign \new_[8108]_  = ~A203 & \new_[8107]_ ;
  assign \new_[8112]_  = ~A302 & ~A301;
  assign \new_[8113]_  = ~A300 & \new_[8112]_ ;
  assign \new_[8114]_  = \new_[8113]_  & \new_[8108]_ ;
  assign \new_[8118]_  = A199 & ~A166;
  assign \new_[8119]_  = ~A167 & \new_[8118]_ ;
  assign \new_[8123]_  = ~A202 & ~A201;
  assign \new_[8124]_  = ~A200 & \new_[8123]_ ;
  assign \new_[8125]_  = \new_[8124]_  & \new_[8119]_ ;
  assign \new_[8129]_  = A299 & ~A298;
  assign \new_[8130]_  = ~A203 & \new_[8129]_ ;
  assign \new_[8134]_  = ~A302 & ~A301;
  assign \new_[8135]_  = ~A300 & \new_[8134]_ ;
  assign \new_[8136]_  = \new_[8135]_  & \new_[8130]_ ;
  assign \new_[8140]_  = A167 & A168;
  assign \new_[8141]_  = ~A170 & \new_[8140]_ ;
  assign \new_[8145]_  = ~A202 & A201;
  assign \new_[8146]_  = ~A166 & \new_[8145]_ ;
  assign \new_[8147]_  = \new_[8146]_  & \new_[8141]_ ;
  assign \new_[8151]_  = ~A299 & A298;
  assign \new_[8152]_  = ~A203 & \new_[8151]_ ;
  assign \new_[8156]_  = ~A302 & ~A301;
  assign \new_[8157]_  = ~A300 & \new_[8156]_ ;
  assign \new_[8158]_  = \new_[8157]_  & \new_[8152]_ ;
  assign \new_[8162]_  = A167 & A168;
  assign \new_[8163]_  = ~A170 & \new_[8162]_ ;
  assign \new_[8167]_  = ~A202 & A201;
  assign \new_[8168]_  = ~A166 & \new_[8167]_ ;
  assign \new_[8169]_  = \new_[8168]_  & \new_[8163]_ ;
  assign \new_[8173]_  = A299 & ~A298;
  assign \new_[8174]_  = ~A203 & \new_[8173]_ ;
  assign \new_[8178]_  = ~A302 & ~A301;
  assign \new_[8179]_  = ~A300 & \new_[8178]_ ;
  assign \new_[8180]_  = \new_[8179]_  & \new_[8174]_ ;
  assign \new_[8184]_  = ~A167 & A168;
  assign \new_[8185]_  = ~A170 & \new_[8184]_ ;
  assign \new_[8189]_  = ~A202 & A201;
  assign \new_[8190]_  = A166 & \new_[8189]_ ;
  assign \new_[8191]_  = \new_[8190]_  & \new_[8185]_ ;
  assign \new_[8195]_  = ~A299 & A298;
  assign \new_[8196]_  = ~A203 & \new_[8195]_ ;
  assign \new_[8200]_  = ~A302 & ~A301;
  assign \new_[8201]_  = ~A300 & \new_[8200]_ ;
  assign \new_[8202]_  = \new_[8201]_  & \new_[8196]_ ;
  assign \new_[8206]_  = ~A167 & A168;
  assign \new_[8207]_  = ~A170 & \new_[8206]_ ;
  assign \new_[8211]_  = ~A202 & A201;
  assign \new_[8212]_  = A166 & \new_[8211]_ ;
  assign \new_[8213]_  = \new_[8212]_  & \new_[8207]_ ;
  assign \new_[8217]_  = A299 & ~A298;
  assign \new_[8218]_  = ~A203 & \new_[8217]_ ;
  assign \new_[8222]_  = ~A302 & ~A301;
  assign \new_[8223]_  = ~A300 & \new_[8222]_ ;
  assign \new_[8224]_  = \new_[8223]_  & \new_[8218]_ ;
  assign \new_[8228]_  = ~A199 & ~A168;
  assign \new_[8229]_  = ~A170 & \new_[8228]_ ;
  assign \new_[8233]_  = ~A202 & ~A201;
  assign \new_[8234]_  = A200 & \new_[8233]_ ;
  assign \new_[8235]_  = \new_[8234]_  & \new_[8229]_ ;
  assign \new_[8239]_  = ~A299 & A298;
  assign \new_[8240]_  = ~A203 & \new_[8239]_ ;
  assign \new_[8244]_  = ~A302 & ~A301;
  assign \new_[8245]_  = ~A300 & \new_[8244]_ ;
  assign \new_[8246]_  = \new_[8245]_  & \new_[8240]_ ;
  assign \new_[8250]_  = ~A199 & ~A168;
  assign \new_[8251]_  = ~A170 & \new_[8250]_ ;
  assign \new_[8255]_  = ~A202 & ~A201;
  assign \new_[8256]_  = A200 & \new_[8255]_ ;
  assign \new_[8257]_  = \new_[8256]_  & \new_[8251]_ ;
  assign \new_[8261]_  = A299 & ~A298;
  assign \new_[8262]_  = ~A203 & \new_[8261]_ ;
  assign \new_[8266]_  = ~A302 & ~A301;
  assign \new_[8267]_  = ~A300 & \new_[8266]_ ;
  assign \new_[8268]_  = \new_[8267]_  & \new_[8262]_ ;
  assign \new_[8272]_  = A199 & ~A168;
  assign \new_[8273]_  = ~A170 & \new_[8272]_ ;
  assign \new_[8277]_  = ~A202 & ~A201;
  assign \new_[8278]_  = ~A200 & \new_[8277]_ ;
  assign \new_[8279]_  = \new_[8278]_  & \new_[8273]_ ;
  assign \new_[8283]_  = ~A299 & A298;
  assign \new_[8284]_  = ~A203 & \new_[8283]_ ;
  assign \new_[8288]_  = ~A302 & ~A301;
  assign \new_[8289]_  = ~A300 & \new_[8288]_ ;
  assign \new_[8290]_  = \new_[8289]_  & \new_[8284]_ ;
  assign \new_[8294]_  = A199 & ~A168;
  assign \new_[8295]_  = ~A170 & \new_[8294]_ ;
  assign \new_[8299]_  = ~A202 & ~A201;
  assign \new_[8300]_  = ~A200 & \new_[8299]_ ;
  assign \new_[8301]_  = \new_[8300]_  & \new_[8295]_ ;
  assign \new_[8305]_  = A299 & ~A298;
  assign \new_[8306]_  = ~A203 & \new_[8305]_ ;
  assign \new_[8310]_  = ~A302 & ~A301;
  assign \new_[8311]_  = ~A300 & \new_[8310]_ ;
  assign \new_[8312]_  = \new_[8311]_  & \new_[8306]_ ;
  assign \new_[8316]_  = A167 & A168;
  assign \new_[8317]_  = A169 & \new_[8316]_ ;
  assign \new_[8321]_  = ~A202 & A201;
  assign \new_[8322]_  = ~A166 & \new_[8321]_ ;
  assign \new_[8323]_  = \new_[8322]_  & \new_[8317]_ ;
  assign \new_[8327]_  = ~A299 & A298;
  assign \new_[8328]_  = ~A203 & \new_[8327]_ ;
  assign \new_[8332]_  = ~A302 & ~A301;
  assign \new_[8333]_  = ~A300 & \new_[8332]_ ;
  assign \new_[8334]_  = \new_[8333]_  & \new_[8328]_ ;
  assign \new_[8338]_  = A167 & A168;
  assign \new_[8339]_  = A169 & \new_[8338]_ ;
  assign \new_[8343]_  = ~A202 & A201;
  assign \new_[8344]_  = ~A166 & \new_[8343]_ ;
  assign \new_[8345]_  = \new_[8344]_  & \new_[8339]_ ;
  assign \new_[8349]_  = A299 & ~A298;
  assign \new_[8350]_  = ~A203 & \new_[8349]_ ;
  assign \new_[8354]_  = ~A302 & ~A301;
  assign \new_[8355]_  = ~A300 & \new_[8354]_ ;
  assign \new_[8356]_  = \new_[8355]_  & \new_[8350]_ ;
  assign \new_[8360]_  = ~A167 & A168;
  assign \new_[8361]_  = A169 & \new_[8360]_ ;
  assign \new_[8365]_  = ~A202 & A201;
  assign \new_[8366]_  = A166 & \new_[8365]_ ;
  assign \new_[8367]_  = \new_[8366]_  & \new_[8361]_ ;
  assign \new_[8371]_  = ~A299 & A298;
  assign \new_[8372]_  = ~A203 & \new_[8371]_ ;
  assign \new_[8376]_  = ~A302 & ~A301;
  assign \new_[8377]_  = ~A300 & \new_[8376]_ ;
  assign \new_[8378]_  = \new_[8377]_  & \new_[8372]_ ;
  assign \new_[8382]_  = ~A167 & A168;
  assign \new_[8383]_  = A169 & \new_[8382]_ ;
  assign \new_[8387]_  = ~A202 & A201;
  assign \new_[8388]_  = A166 & \new_[8387]_ ;
  assign \new_[8389]_  = \new_[8388]_  & \new_[8383]_ ;
  assign \new_[8393]_  = A299 & ~A298;
  assign \new_[8394]_  = ~A203 & \new_[8393]_ ;
  assign \new_[8398]_  = ~A302 & ~A301;
  assign \new_[8399]_  = ~A300 & \new_[8398]_ ;
  assign \new_[8400]_  = \new_[8399]_  & \new_[8394]_ ;
  assign \new_[8404]_  = ~A199 & ~A168;
  assign \new_[8405]_  = A169 & \new_[8404]_ ;
  assign \new_[8409]_  = ~A202 & ~A201;
  assign \new_[8410]_  = A200 & \new_[8409]_ ;
  assign \new_[8411]_  = \new_[8410]_  & \new_[8405]_ ;
  assign \new_[8415]_  = ~A299 & A298;
  assign \new_[8416]_  = ~A203 & \new_[8415]_ ;
  assign \new_[8420]_  = ~A302 & ~A301;
  assign \new_[8421]_  = ~A300 & \new_[8420]_ ;
  assign \new_[8422]_  = \new_[8421]_  & \new_[8416]_ ;
  assign \new_[8426]_  = ~A199 & ~A168;
  assign \new_[8427]_  = A169 & \new_[8426]_ ;
  assign \new_[8431]_  = ~A202 & ~A201;
  assign \new_[8432]_  = A200 & \new_[8431]_ ;
  assign \new_[8433]_  = \new_[8432]_  & \new_[8427]_ ;
  assign \new_[8437]_  = A299 & ~A298;
  assign \new_[8438]_  = ~A203 & \new_[8437]_ ;
  assign \new_[8442]_  = ~A302 & ~A301;
  assign \new_[8443]_  = ~A300 & \new_[8442]_ ;
  assign \new_[8444]_  = \new_[8443]_  & \new_[8438]_ ;
  assign \new_[8448]_  = A199 & ~A168;
  assign \new_[8449]_  = A169 & \new_[8448]_ ;
  assign \new_[8453]_  = ~A202 & ~A201;
  assign \new_[8454]_  = ~A200 & \new_[8453]_ ;
  assign \new_[8455]_  = \new_[8454]_  & \new_[8449]_ ;
  assign \new_[8459]_  = ~A299 & A298;
  assign \new_[8460]_  = ~A203 & \new_[8459]_ ;
  assign \new_[8464]_  = ~A302 & ~A301;
  assign \new_[8465]_  = ~A300 & \new_[8464]_ ;
  assign \new_[8466]_  = \new_[8465]_  & \new_[8460]_ ;
  assign \new_[8470]_  = A199 & ~A168;
  assign \new_[8471]_  = A169 & \new_[8470]_ ;
  assign \new_[8475]_  = ~A202 & ~A201;
  assign \new_[8476]_  = ~A200 & \new_[8475]_ ;
  assign \new_[8477]_  = \new_[8476]_  & \new_[8471]_ ;
  assign \new_[8481]_  = A299 & ~A298;
  assign \new_[8482]_  = ~A203 & \new_[8481]_ ;
  assign \new_[8486]_  = ~A302 & ~A301;
  assign \new_[8487]_  = ~A300 & \new_[8486]_ ;
  assign \new_[8488]_  = \new_[8487]_  & \new_[8482]_ ;
  assign \new_[8492]_  = A168 & ~A169;
  assign \new_[8493]_  = A170 & \new_[8492]_ ;
  assign \new_[8497]_  = A201 & A200;
  assign \new_[8498]_  = ~A199 & \new_[8497]_ ;
  assign \new_[8499]_  = \new_[8498]_  & \new_[8493]_ ;
  assign \new_[8503]_  = ~A299 & A298;
  assign \new_[8504]_  = A202 & \new_[8503]_ ;
  assign \new_[8508]_  = ~A302 & ~A301;
  assign \new_[8509]_  = ~A300 & \new_[8508]_ ;
  assign \new_[8510]_  = \new_[8509]_  & \new_[8504]_ ;
  assign \new_[8514]_  = A168 & ~A169;
  assign \new_[8515]_  = A170 & \new_[8514]_ ;
  assign \new_[8519]_  = A201 & A200;
  assign \new_[8520]_  = ~A199 & \new_[8519]_ ;
  assign \new_[8521]_  = \new_[8520]_  & \new_[8515]_ ;
  assign \new_[8525]_  = A299 & ~A298;
  assign \new_[8526]_  = A202 & \new_[8525]_ ;
  assign \new_[8530]_  = ~A302 & ~A301;
  assign \new_[8531]_  = ~A300 & \new_[8530]_ ;
  assign \new_[8532]_  = \new_[8531]_  & \new_[8526]_ ;
  assign \new_[8536]_  = A168 & ~A169;
  assign \new_[8537]_  = A170 & \new_[8536]_ ;
  assign \new_[8541]_  = A201 & A200;
  assign \new_[8542]_  = ~A199 & \new_[8541]_ ;
  assign \new_[8543]_  = \new_[8542]_  & \new_[8537]_ ;
  assign \new_[8547]_  = ~A299 & A298;
  assign \new_[8548]_  = A203 & \new_[8547]_ ;
  assign \new_[8552]_  = ~A302 & ~A301;
  assign \new_[8553]_  = ~A300 & \new_[8552]_ ;
  assign \new_[8554]_  = \new_[8553]_  & \new_[8548]_ ;
  assign \new_[8558]_  = A168 & ~A169;
  assign \new_[8559]_  = A170 & \new_[8558]_ ;
  assign \new_[8563]_  = A201 & A200;
  assign \new_[8564]_  = ~A199 & \new_[8563]_ ;
  assign \new_[8565]_  = \new_[8564]_  & \new_[8559]_ ;
  assign \new_[8569]_  = A299 & ~A298;
  assign \new_[8570]_  = A203 & \new_[8569]_ ;
  assign \new_[8574]_  = ~A302 & ~A301;
  assign \new_[8575]_  = ~A300 & \new_[8574]_ ;
  assign \new_[8576]_  = \new_[8575]_  & \new_[8570]_ ;
  assign \new_[8580]_  = A168 & ~A169;
  assign \new_[8581]_  = A170 & \new_[8580]_ ;
  assign \new_[8585]_  = ~A201 & A200;
  assign \new_[8586]_  = ~A199 & \new_[8585]_ ;
  assign \new_[8587]_  = \new_[8586]_  & \new_[8581]_ ;
  assign \new_[8591]_  = A298 & ~A203;
  assign \new_[8592]_  = ~A202 & \new_[8591]_ ;
  assign \new_[8596]_  = A301 & A300;
  assign \new_[8597]_  = ~A299 & \new_[8596]_ ;
  assign \new_[8598]_  = \new_[8597]_  & \new_[8592]_ ;
  assign \new_[8602]_  = A168 & ~A169;
  assign \new_[8603]_  = A170 & \new_[8602]_ ;
  assign \new_[8607]_  = ~A201 & A200;
  assign \new_[8608]_  = ~A199 & \new_[8607]_ ;
  assign \new_[8609]_  = \new_[8608]_  & \new_[8603]_ ;
  assign \new_[8613]_  = A298 & ~A203;
  assign \new_[8614]_  = ~A202 & \new_[8613]_ ;
  assign \new_[8618]_  = A302 & A300;
  assign \new_[8619]_  = ~A299 & \new_[8618]_ ;
  assign \new_[8620]_  = \new_[8619]_  & \new_[8614]_ ;
  assign \new_[8624]_  = A168 & ~A169;
  assign \new_[8625]_  = A170 & \new_[8624]_ ;
  assign \new_[8629]_  = ~A201 & A200;
  assign \new_[8630]_  = ~A199 & \new_[8629]_ ;
  assign \new_[8631]_  = \new_[8630]_  & \new_[8625]_ ;
  assign \new_[8635]_  = ~A298 & ~A203;
  assign \new_[8636]_  = ~A202 & \new_[8635]_ ;
  assign \new_[8640]_  = A301 & A300;
  assign \new_[8641]_  = A299 & \new_[8640]_ ;
  assign \new_[8642]_  = \new_[8641]_  & \new_[8636]_ ;
  assign \new_[8646]_  = A168 & ~A169;
  assign \new_[8647]_  = A170 & \new_[8646]_ ;
  assign \new_[8651]_  = ~A201 & A200;
  assign \new_[8652]_  = ~A199 & \new_[8651]_ ;
  assign \new_[8653]_  = \new_[8652]_  & \new_[8647]_ ;
  assign \new_[8657]_  = ~A298 & ~A203;
  assign \new_[8658]_  = ~A202 & \new_[8657]_ ;
  assign \new_[8662]_  = A302 & A300;
  assign \new_[8663]_  = A299 & \new_[8662]_ ;
  assign \new_[8664]_  = \new_[8663]_  & \new_[8658]_ ;
  assign \new_[8668]_  = A168 & ~A169;
  assign \new_[8669]_  = A170 & \new_[8668]_ ;
  assign \new_[8673]_  = A201 & ~A200;
  assign \new_[8674]_  = A199 & \new_[8673]_ ;
  assign \new_[8675]_  = \new_[8674]_  & \new_[8669]_ ;
  assign \new_[8679]_  = ~A299 & A298;
  assign \new_[8680]_  = A202 & \new_[8679]_ ;
  assign \new_[8684]_  = ~A302 & ~A301;
  assign \new_[8685]_  = ~A300 & \new_[8684]_ ;
  assign \new_[8686]_  = \new_[8685]_  & \new_[8680]_ ;
  assign \new_[8690]_  = A168 & ~A169;
  assign \new_[8691]_  = A170 & \new_[8690]_ ;
  assign \new_[8695]_  = A201 & ~A200;
  assign \new_[8696]_  = A199 & \new_[8695]_ ;
  assign \new_[8697]_  = \new_[8696]_  & \new_[8691]_ ;
  assign \new_[8701]_  = A299 & ~A298;
  assign \new_[8702]_  = A202 & \new_[8701]_ ;
  assign \new_[8706]_  = ~A302 & ~A301;
  assign \new_[8707]_  = ~A300 & \new_[8706]_ ;
  assign \new_[8708]_  = \new_[8707]_  & \new_[8702]_ ;
  assign \new_[8712]_  = A168 & ~A169;
  assign \new_[8713]_  = A170 & \new_[8712]_ ;
  assign \new_[8717]_  = A201 & ~A200;
  assign \new_[8718]_  = A199 & \new_[8717]_ ;
  assign \new_[8719]_  = \new_[8718]_  & \new_[8713]_ ;
  assign \new_[8723]_  = ~A299 & A298;
  assign \new_[8724]_  = A203 & \new_[8723]_ ;
  assign \new_[8728]_  = ~A302 & ~A301;
  assign \new_[8729]_  = ~A300 & \new_[8728]_ ;
  assign \new_[8730]_  = \new_[8729]_  & \new_[8724]_ ;
  assign \new_[8734]_  = A168 & ~A169;
  assign \new_[8735]_  = A170 & \new_[8734]_ ;
  assign \new_[8739]_  = A201 & ~A200;
  assign \new_[8740]_  = A199 & \new_[8739]_ ;
  assign \new_[8741]_  = \new_[8740]_  & \new_[8735]_ ;
  assign \new_[8745]_  = A299 & ~A298;
  assign \new_[8746]_  = A203 & \new_[8745]_ ;
  assign \new_[8750]_  = ~A302 & ~A301;
  assign \new_[8751]_  = ~A300 & \new_[8750]_ ;
  assign \new_[8752]_  = \new_[8751]_  & \new_[8746]_ ;
  assign \new_[8756]_  = A168 & ~A169;
  assign \new_[8757]_  = A170 & \new_[8756]_ ;
  assign \new_[8761]_  = ~A201 & ~A200;
  assign \new_[8762]_  = A199 & \new_[8761]_ ;
  assign \new_[8763]_  = \new_[8762]_  & \new_[8757]_ ;
  assign \new_[8767]_  = A298 & ~A203;
  assign \new_[8768]_  = ~A202 & \new_[8767]_ ;
  assign \new_[8772]_  = A301 & A300;
  assign \new_[8773]_  = ~A299 & \new_[8772]_ ;
  assign \new_[8774]_  = \new_[8773]_  & \new_[8768]_ ;
  assign \new_[8778]_  = A168 & ~A169;
  assign \new_[8779]_  = A170 & \new_[8778]_ ;
  assign \new_[8783]_  = ~A201 & ~A200;
  assign \new_[8784]_  = A199 & \new_[8783]_ ;
  assign \new_[8785]_  = \new_[8784]_  & \new_[8779]_ ;
  assign \new_[8789]_  = A298 & ~A203;
  assign \new_[8790]_  = ~A202 & \new_[8789]_ ;
  assign \new_[8794]_  = A302 & A300;
  assign \new_[8795]_  = ~A299 & \new_[8794]_ ;
  assign \new_[8796]_  = \new_[8795]_  & \new_[8790]_ ;
  assign \new_[8800]_  = A168 & ~A169;
  assign \new_[8801]_  = A170 & \new_[8800]_ ;
  assign \new_[8805]_  = ~A201 & ~A200;
  assign \new_[8806]_  = A199 & \new_[8805]_ ;
  assign \new_[8807]_  = \new_[8806]_  & \new_[8801]_ ;
  assign \new_[8811]_  = ~A298 & ~A203;
  assign \new_[8812]_  = ~A202 & \new_[8811]_ ;
  assign \new_[8816]_  = A301 & A300;
  assign \new_[8817]_  = A299 & \new_[8816]_ ;
  assign \new_[8818]_  = \new_[8817]_  & \new_[8812]_ ;
  assign \new_[8822]_  = A168 & ~A169;
  assign \new_[8823]_  = A170 & \new_[8822]_ ;
  assign \new_[8827]_  = ~A201 & ~A200;
  assign \new_[8828]_  = A199 & \new_[8827]_ ;
  assign \new_[8829]_  = \new_[8828]_  & \new_[8823]_ ;
  assign \new_[8833]_  = ~A298 & ~A203;
  assign \new_[8834]_  = ~A202 & \new_[8833]_ ;
  assign \new_[8838]_  = A302 & A300;
  assign \new_[8839]_  = A299 & \new_[8838]_ ;
  assign \new_[8840]_  = \new_[8839]_  & \new_[8834]_ ;
  assign \new_[8844]_  = ~A168 & ~A169;
  assign \new_[8845]_  = A170 & \new_[8844]_ ;
  assign \new_[8849]_  = A201 & ~A166;
  assign \new_[8850]_  = A167 & \new_[8849]_ ;
  assign \new_[8851]_  = \new_[8850]_  & \new_[8845]_ ;
  assign \new_[8855]_  = A298 & ~A203;
  assign \new_[8856]_  = ~A202 & \new_[8855]_ ;
  assign \new_[8860]_  = A301 & A300;
  assign \new_[8861]_  = ~A299 & \new_[8860]_ ;
  assign \new_[8862]_  = \new_[8861]_  & \new_[8856]_ ;
  assign \new_[8866]_  = ~A168 & ~A169;
  assign \new_[8867]_  = A170 & \new_[8866]_ ;
  assign \new_[8871]_  = A201 & ~A166;
  assign \new_[8872]_  = A167 & \new_[8871]_ ;
  assign \new_[8873]_  = \new_[8872]_  & \new_[8867]_ ;
  assign \new_[8877]_  = A298 & ~A203;
  assign \new_[8878]_  = ~A202 & \new_[8877]_ ;
  assign \new_[8882]_  = A302 & A300;
  assign \new_[8883]_  = ~A299 & \new_[8882]_ ;
  assign \new_[8884]_  = \new_[8883]_  & \new_[8878]_ ;
  assign \new_[8888]_  = ~A168 & ~A169;
  assign \new_[8889]_  = A170 & \new_[8888]_ ;
  assign \new_[8893]_  = A201 & ~A166;
  assign \new_[8894]_  = A167 & \new_[8893]_ ;
  assign \new_[8895]_  = \new_[8894]_  & \new_[8889]_ ;
  assign \new_[8899]_  = ~A298 & ~A203;
  assign \new_[8900]_  = ~A202 & \new_[8899]_ ;
  assign \new_[8904]_  = A301 & A300;
  assign \new_[8905]_  = A299 & \new_[8904]_ ;
  assign \new_[8906]_  = \new_[8905]_  & \new_[8900]_ ;
  assign \new_[8910]_  = ~A168 & ~A169;
  assign \new_[8911]_  = A170 & \new_[8910]_ ;
  assign \new_[8915]_  = A201 & ~A166;
  assign \new_[8916]_  = A167 & \new_[8915]_ ;
  assign \new_[8917]_  = \new_[8916]_  & \new_[8911]_ ;
  assign \new_[8921]_  = ~A298 & ~A203;
  assign \new_[8922]_  = ~A202 & \new_[8921]_ ;
  assign \new_[8926]_  = A302 & A300;
  assign \new_[8927]_  = A299 & \new_[8926]_ ;
  assign \new_[8928]_  = \new_[8927]_  & \new_[8922]_ ;
  assign \new_[8932]_  = ~A168 & ~A169;
  assign \new_[8933]_  = A170 & \new_[8932]_ ;
  assign \new_[8937]_  = ~A201 & ~A166;
  assign \new_[8938]_  = A167 & \new_[8937]_ ;
  assign \new_[8939]_  = \new_[8938]_  & \new_[8933]_ ;
  assign \new_[8943]_  = ~A299 & A298;
  assign \new_[8944]_  = A202 & \new_[8943]_ ;
  assign \new_[8948]_  = ~A302 & ~A301;
  assign \new_[8949]_  = ~A300 & \new_[8948]_ ;
  assign \new_[8950]_  = \new_[8949]_  & \new_[8944]_ ;
  assign \new_[8954]_  = ~A168 & ~A169;
  assign \new_[8955]_  = A170 & \new_[8954]_ ;
  assign \new_[8959]_  = ~A201 & ~A166;
  assign \new_[8960]_  = A167 & \new_[8959]_ ;
  assign \new_[8961]_  = \new_[8960]_  & \new_[8955]_ ;
  assign \new_[8965]_  = A299 & ~A298;
  assign \new_[8966]_  = A202 & \new_[8965]_ ;
  assign \new_[8970]_  = ~A302 & ~A301;
  assign \new_[8971]_  = ~A300 & \new_[8970]_ ;
  assign \new_[8972]_  = \new_[8971]_  & \new_[8966]_ ;
  assign \new_[8976]_  = ~A168 & ~A169;
  assign \new_[8977]_  = A170 & \new_[8976]_ ;
  assign \new_[8981]_  = ~A201 & ~A166;
  assign \new_[8982]_  = A167 & \new_[8981]_ ;
  assign \new_[8983]_  = \new_[8982]_  & \new_[8977]_ ;
  assign \new_[8987]_  = ~A299 & A298;
  assign \new_[8988]_  = A203 & \new_[8987]_ ;
  assign \new_[8992]_  = ~A302 & ~A301;
  assign \new_[8993]_  = ~A300 & \new_[8992]_ ;
  assign \new_[8994]_  = \new_[8993]_  & \new_[8988]_ ;
  assign \new_[8998]_  = ~A168 & ~A169;
  assign \new_[8999]_  = A170 & \new_[8998]_ ;
  assign \new_[9003]_  = ~A201 & ~A166;
  assign \new_[9004]_  = A167 & \new_[9003]_ ;
  assign \new_[9005]_  = \new_[9004]_  & \new_[8999]_ ;
  assign \new_[9009]_  = A299 & ~A298;
  assign \new_[9010]_  = A203 & \new_[9009]_ ;
  assign \new_[9014]_  = ~A302 & ~A301;
  assign \new_[9015]_  = ~A300 & \new_[9014]_ ;
  assign \new_[9016]_  = \new_[9015]_  & \new_[9010]_ ;
  assign \new_[9020]_  = ~A168 & ~A169;
  assign \new_[9021]_  = A170 & \new_[9020]_ ;
  assign \new_[9025]_  = A199 & ~A166;
  assign \new_[9026]_  = A167 & \new_[9025]_ ;
  assign \new_[9027]_  = \new_[9026]_  & \new_[9021]_ ;
  assign \new_[9031]_  = ~A299 & A298;
  assign \new_[9032]_  = A200 & \new_[9031]_ ;
  assign \new_[9036]_  = ~A302 & ~A301;
  assign \new_[9037]_  = ~A300 & \new_[9036]_ ;
  assign \new_[9038]_  = \new_[9037]_  & \new_[9032]_ ;
  assign \new_[9042]_  = ~A168 & ~A169;
  assign \new_[9043]_  = A170 & \new_[9042]_ ;
  assign \new_[9047]_  = A199 & ~A166;
  assign \new_[9048]_  = A167 & \new_[9047]_ ;
  assign \new_[9049]_  = \new_[9048]_  & \new_[9043]_ ;
  assign \new_[9053]_  = A299 & ~A298;
  assign \new_[9054]_  = A200 & \new_[9053]_ ;
  assign \new_[9058]_  = ~A302 & ~A301;
  assign \new_[9059]_  = ~A300 & \new_[9058]_ ;
  assign \new_[9060]_  = \new_[9059]_  & \new_[9054]_ ;
  assign \new_[9064]_  = ~A168 & ~A169;
  assign \new_[9065]_  = A170 & \new_[9064]_ ;
  assign \new_[9069]_  = ~A199 & ~A166;
  assign \new_[9070]_  = A167 & \new_[9069]_ ;
  assign \new_[9071]_  = \new_[9070]_  & \new_[9065]_ ;
  assign \new_[9075]_  = ~A299 & A298;
  assign \new_[9076]_  = ~A200 & \new_[9075]_ ;
  assign \new_[9080]_  = ~A302 & ~A301;
  assign \new_[9081]_  = ~A300 & \new_[9080]_ ;
  assign \new_[9082]_  = \new_[9081]_  & \new_[9076]_ ;
  assign \new_[9086]_  = ~A168 & ~A169;
  assign \new_[9087]_  = A170 & \new_[9086]_ ;
  assign \new_[9091]_  = ~A199 & ~A166;
  assign \new_[9092]_  = A167 & \new_[9091]_ ;
  assign \new_[9093]_  = \new_[9092]_  & \new_[9087]_ ;
  assign \new_[9097]_  = A299 & ~A298;
  assign \new_[9098]_  = ~A200 & \new_[9097]_ ;
  assign \new_[9102]_  = ~A302 & ~A301;
  assign \new_[9103]_  = ~A300 & \new_[9102]_ ;
  assign \new_[9104]_  = \new_[9103]_  & \new_[9098]_ ;
  assign \new_[9108]_  = ~A168 & ~A169;
  assign \new_[9109]_  = A170 & \new_[9108]_ ;
  assign \new_[9113]_  = A201 & A166;
  assign \new_[9114]_  = ~A167 & \new_[9113]_ ;
  assign \new_[9115]_  = \new_[9114]_  & \new_[9109]_ ;
  assign \new_[9119]_  = A298 & ~A203;
  assign \new_[9120]_  = ~A202 & \new_[9119]_ ;
  assign \new_[9124]_  = A301 & A300;
  assign \new_[9125]_  = ~A299 & \new_[9124]_ ;
  assign \new_[9126]_  = \new_[9125]_  & \new_[9120]_ ;
  assign \new_[9130]_  = ~A168 & ~A169;
  assign \new_[9131]_  = A170 & \new_[9130]_ ;
  assign \new_[9135]_  = A201 & A166;
  assign \new_[9136]_  = ~A167 & \new_[9135]_ ;
  assign \new_[9137]_  = \new_[9136]_  & \new_[9131]_ ;
  assign \new_[9141]_  = A298 & ~A203;
  assign \new_[9142]_  = ~A202 & \new_[9141]_ ;
  assign \new_[9146]_  = A302 & A300;
  assign \new_[9147]_  = ~A299 & \new_[9146]_ ;
  assign \new_[9148]_  = \new_[9147]_  & \new_[9142]_ ;
  assign \new_[9152]_  = ~A168 & ~A169;
  assign \new_[9153]_  = A170 & \new_[9152]_ ;
  assign \new_[9157]_  = A201 & A166;
  assign \new_[9158]_  = ~A167 & \new_[9157]_ ;
  assign \new_[9159]_  = \new_[9158]_  & \new_[9153]_ ;
  assign \new_[9163]_  = ~A298 & ~A203;
  assign \new_[9164]_  = ~A202 & \new_[9163]_ ;
  assign \new_[9168]_  = A301 & A300;
  assign \new_[9169]_  = A299 & \new_[9168]_ ;
  assign \new_[9170]_  = \new_[9169]_  & \new_[9164]_ ;
  assign \new_[9174]_  = ~A168 & ~A169;
  assign \new_[9175]_  = A170 & \new_[9174]_ ;
  assign \new_[9179]_  = A201 & A166;
  assign \new_[9180]_  = ~A167 & \new_[9179]_ ;
  assign \new_[9181]_  = \new_[9180]_  & \new_[9175]_ ;
  assign \new_[9185]_  = ~A298 & ~A203;
  assign \new_[9186]_  = ~A202 & \new_[9185]_ ;
  assign \new_[9190]_  = A302 & A300;
  assign \new_[9191]_  = A299 & \new_[9190]_ ;
  assign \new_[9192]_  = \new_[9191]_  & \new_[9186]_ ;
  assign \new_[9196]_  = ~A168 & ~A169;
  assign \new_[9197]_  = A170 & \new_[9196]_ ;
  assign \new_[9201]_  = ~A201 & A166;
  assign \new_[9202]_  = ~A167 & \new_[9201]_ ;
  assign \new_[9203]_  = \new_[9202]_  & \new_[9197]_ ;
  assign \new_[9207]_  = ~A299 & A298;
  assign \new_[9208]_  = A202 & \new_[9207]_ ;
  assign \new_[9212]_  = ~A302 & ~A301;
  assign \new_[9213]_  = ~A300 & \new_[9212]_ ;
  assign \new_[9214]_  = \new_[9213]_  & \new_[9208]_ ;
  assign \new_[9218]_  = ~A168 & ~A169;
  assign \new_[9219]_  = A170 & \new_[9218]_ ;
  assign \new_[9223]_  = ~A201 & A166;
  assign \new_[9224]_  = ~A167 & \new_[9223]_ ;
  assign \new_[9225]_  = \new_[9224]_  & \new_[9219]_ ;
  assign \new_[9229]_  = A299 & ~A298;
  assign \new_[9230]_  = A202 & \new_[9229]_ ;
  assign \new_[9234]_  = ~A302 & ~A301;
  assign \new_[9235]_  = ~A300 & \new_[9234]_ ;
  assign \new_[9236]_  = \new_[9235]_  & \new_[9230]_ ;
  assign \new_[9240]_  = ~A168 & ~A169;
  assign \new_[9241]_  = A170 & \new_[9240]_ ;
  assign \new_[9245]_  = ~A201 & A166;
  assign \new_[9246]_  = ~A167 & \new_[9245]_ ;
  assign \new_[9247]_  = \new_[9246]_  & \new_[9241]_ ;
  assign \new_[9251]_  = ~A299 & A298;
  assign \new_[9252]_  = A203 & \new_[9251]_ ;
  assign \new_[9256]_  = ~A302 & ~A301;
  assign \new_[9257]_  = ~A300 & \new_[9256]_ ;
  assign \new_[9258]_  = \new_[9257]_  & \new_[9252]_ ;
  assign \new_[9262]_  = ~A168 & ~A169;
  assign \new_[9263]_  = A170 & \new_[9262]_ ;
  assign \new_[9267]_  = ~A201 & A166;
  assign \new_[9268]_  = ~A167 & \new_[9267]_ ;
  assign \new_[9269]_  = \new_[9268]_  & \new_[9263]_ ;
  assign \new_[9273]_  = A299 & ~A298;
  assign \new_[9274]_  = A203 & \new_[9273]_ ;
  assign \new_[9278]_  = ~A302 & ~A301;
  assign \new_[9279]_  = ~A300 & \new_[9278]_ ;
  assign \new_[9280]_  = \new_[9279]_  & \new_[9274]_ ;
  assign \new_[9284]_  = ~A168 & ~A169;
  assign \new_[9285]_  = A170 & \new_[9284]_ ;
  assign \new_[9289]_  = A199 & A166;
  assign \new_[9290]_  = ~A167 & \new_[9289]_ ;
  assign \new_[9291]_  = \new_[9290]_  & \new_[9285]_ ;
  assign \new_[9295]_  = ~A299 & A298;
  assign \new_[9296]_  = A200 & \new_[9295]_ ;
  assign \new_[9300]_  = ~A302 & ~A301;
  assign \new_[9301]_  = ~A300 & \new_[9300]_ ;
  assign \new_[9302]_  = \new_[9301]_  & \new_[9296]_ ;
  assign \new_[9306]_  = ~A168 & ~A169;
  assign \new_[9307]_  = A170 & \new_[9306]_ ;
  assign \new_[9311]_  = A199 & A166;
  assign \new_[9312]_  = ~A167 & \new_[9311]_ ;
  assign \new_[9313]_  = \new_[9312]_  & \new_[9307]_ ;
  assign \new_[9317]_  = A299 & ~A298;
  assign \new_[9318]_  = A200 & \new_[9317]_ ;
  assign \new_[9322]_  = ~A302 & ~A301;
  assign \new_[9323]_  = ~A300 & \new_[9322]_ ;
  assign \new_[9324]_  = \new_[9323]_  & \new_[9318]_ ;
  assign \new_[9328]_  = ~A168 & ~A169;
  assign \new_[9329]_  = A170 & \new_[9328]_ ;
  assign \new_[9333]_  = ~A199 & A166;
  assign \new_[9334]_  = ~A167 & \new_[9333]_ ;
  assign \new_[9335]_  = \new_[9334]_  & \new_[9329]_ ;
  assign \new_[9339]_  = ~A299 & A298;
  assign \new_[9340]_  = ~A200 & \new_[9339]_ ;
  assign \new_[9344]_  = ~A302 & ~A301;
  assign \new_[9345]_  = ~A300 & \new_[9344]_ ;
  assign \new_[9346]_  = \new_[9345]_  & \new_[9340]_ ;
  assign \new_[9350]_  = ~A168 & ~A169;
  assign \new_[9351]_  = A170 & \new_[9350]_ ;
  assign \new_[9355]_  = ~A199 & A166;
  assign \new_[9356]_  = ~A167 & \new_[9355]_ ;
  assign \new_[9357]_  = \new_[9356]_  & \new_[9351]_ ;
  assign \new_[9361]_  = A299 & ~A298;
  assign \new_[9362]_  = ~A200 & \new_[9361]_ ;
  assign \new_[9366]_  = ~A302 & ~A301;
  assign \new_[9367]_  = ~A300 & \new_[9366]_ ;
  assign \new_[9368]_  = \new_[9367]_  & \new_[9362]_ ;
  assign \new_[9372]_  = A168 & ~A169;
  assign \new_[9373]_  = A170 & \new_[9372]_ ;
  assign \new_[9377]_  = ~A201 & A200;
  assign \new_[9378]_  = ~A199 & \new_[9377]_ ;
  assign \new_[9379]_  = \new_[9378]_  & \new_[9373]_ ;
  assign \new_[9383]_  = A298 & ~A203;
  assign \new_[9384]_  = ~A202 & \new_[9383]_ ;
  assign \new_[9387]_  = ~A300 & ~A299;
  assign \new_[9390]_  = ~A302 & ~A301;
  assign \new_[9391]_  = \new_[9390]_  & \new_[9387]_ ;
  assign \new_[9392]_  = \new_[9391]_  & \new_[9384]_ ;
  assign \new_[9396]_  = A168 & ~A169;
  assign \new_[9397]_  = A170 & \new_[9396]_ ;
  assign \new_[9401]_  = ~A201 & A200;
  assign \new_[9402]_  = ~A199 & \new_[9401]_ ;
  assign \new_[9403]_  = \new_[9402]_  & \new_[9397]_ ;
  assign \new_[9407]_  = ~A298 & ~A203;
  assign \new_[9408]_  = ~A202 & \new_[9407]_ ;
  assign \new_[9411]_  = ~A300 & A299;
  assign \new_[9414]_  = ~A302 & ~A301;
  assign \new_[9415]_  = \new_[9414]_  & \new_[9411]_ ;
  assign \new_[9416]_  = \new_[9415]_  & \new_[9408]_ ;
  assign \new_[9420]_  = A168 & ~A169;
  assign \new_[9421]_  = A170 & \new_[9420]_ ;
  assign \new_[9425]_  = ~A201 & ~A200;
  assign \new_[9426]_  = A199 & \new_[9425]_ ;
  assign \new_[9427]_  = \new_[9426]_  & \new_[9421]_ ;
  assign \new_[9431]_  = A298 & ~A203;
  assign \new_[9432]_  = ~A202 & \new_[9431]_ ;
  assign \new_[9435]_  = ~A300 & ~A299;
  assign \new_[9438]_  = ~A302 & ~A301;
  assign \new_[9439]_  = \new_[9438]_  & \new_[9435]_ ;
  assign \new_[9440]_  = \new_[9439]_  & \new_[9432]_ ;
  assign \new_[9444]_  = A168 & ~A169;
  assign \new_[9445]_  = A170 & \new_[9444]_ ;
  assign \new_[9449]_  = ~A201 & ~A200;
  assign \new_[9450]_  = A199 & \new_[9449]_ ;
  assign \new_[9451]_  = \new_[9450]_  & \new_[9445]_ ;
  assign \new_[9455]_  = ~A298 & ~A203;
  assign \new_[9456]_  = ~A202 & \new_[9455]_ ;
  assign \new_[9459]_  = ~A300 & A299;
  assign \new_[9462]_  = ~A302 & ~A301;
  assign \new_[9463]_  = \new_[9462]_  & \new_[9459]_ ;
  assign \new_[9464]_  = \new_[9463]_  & \new_[9456]_ ;
  assign \new_[9468]_  = ~A168 & ~A169;
  assign \new_[9469]_  = A170 & \new_[9468]_ ;
  assign \new_[9473]_  = A201 & ~A166;
  assign \new_[9474]_  = A167 & \new_[9473]_ ;
  assign \new_[9475]_  = \new_[9474]_  & \new_[9469]_ ;
  assign \new_[9479]_  = A298 & ~A203;
  assign \new_[9480]_  = ~A202 & \new_[9479]_ ;
  assign \new_[9483]_  = ~A300 & ~A299;
  assign \new_[9486]_  = ~A302 & ~A301;
  assign \new_[9487]_  = \new_[9486]_  & \new_[9483]_ ;
  assign \new_[9488]_  = \new_[9487]_  & \new_[9480]_ ;
  assign \new_[9492]_  = ~A168 & ~A169;
  assign \new_[9493]_  = A170 & \new_[9492]_ ;
  assign \new_[9497]_  = A201 & ~A166;
  assign \new_[9498]_  = A167 & \new_[9497]_ ;
  assign \new_[9499]_  = \new_[9498]_  & \new_[9493]_ ;
  assign \new_[9503]_  = ~A298 & ~A203;
  assign \new_[9504]_  = ~A202 & \new_[9503]_ ;
  assign \new_[9507]_  = ~A300 & A299;
  assign \new_[9510]_  = ~A302 & ~A301;
  assign \new_[9511]_  = \new_[9510]_  & \new_[9507]_ ;
  assign \new_[9512]_  = \new_[9511]_  & \new_[9504]_ ;
  assign \new_[9516]_  = ~A168 & ~A169;
  assign \new_[9517]_  = A170 & \new_[9516]_ ;
  assign \new_[9521]_  = A201 & A166;
  assign \new_[9522]_  = ~A167 & \new_[9521]_ ;
  assign \new_[9523]_  = \new_[9522]_  & \new_[9517]_ ;
  assign \new_[9527]_  = A298 & ~A203;
  assign \new_[9528]_  = ~A202 & \new_[9527]_ ;
  assign \new_[9531]_  = ~A300 & ~A299;
  assign \new_[9534]_  = ~A302 & ~A301;
  assign \new_[9535]_  = \new_[9534]_  & \new_[9531]_ ;
  assign \new_[9536]_  = \new_[9535]_  & \new_[9528]_ ;
  assign \new_[9540]_  = ~A168 & ~A169;
  assign \new_[9541]_  = A170 & \new_[9540]_ ;
  assign \new_[9545]_  = A201 & A166;
  assign \new_[9546]_  = ~A167 & \new_[9545]_ ;
  assign \new_[9547]_  = \new_[9546]_  & \new_[9541]_ ;
  assign \new_[9551]_  = ~A298 & ~A203;
  assign \new_[9552]_  = ~A202 & \new_[9551]_ ;
  assign \new_[9555]_  = ~A300 & A299;
  assign \new_[9558]_  = ~A302 & ~A301;
  assign \new_[9559]_  = \new_[9558]_  & \new_[9555]_ ;
  assign \new_[9560]_  = \new_[9559]_  & \new_[9552]_ ;
endmodule


