// Benchmark "top" written by ABC on Thu Oct  8 22:52:01 2020

module top ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_;
  assign new_n137_ = ~\A[125]  & \A[127] ;
  assign new_n138_ = \A[126]  & \A[127] ;
  assign new_n139_ = \A[126]  & ~new_n138_;
  assign new_n140_ = \A[125]  & ~new_n139_;
  assign new_n141_ = ~new_n137_ & ~new_n140_;
  assign new_n142_ = ~\A[123]  & ~new_n141_;
  assign new_n143_ = ~\A[124]  & ~new_n139_;
  assign new_n144_ = \A[124]  & ~new_n141_;
  assign new_n145_ = ~new_n143_ & ~new_n144_;
  assign new_n146_ = \A[123]  & ~new_n145_;
  assign new_n147_ = ~new_n142_ & ~new_n146_;
  assign new_n148_ = ~\A[121]  & ~new_n147_;
  assign new_n149_ = ~\A[122]  & ~new_n145_;
  assign new_n150_ = \A[122]  & ~new_n147_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = \A[121]  & ~new_n151_;
  assign new_n153_ = ~new_n148_ & ~new_n152_;
  assign new_n154_ = ~\A[119]  & ~new_n153_;
  assign new_n155_ = ~\A[120]  & ~new_n151_;
  assign new_n156_ = \A[120]  & ~new_n153_;
  assign new_n157_ = ~new_n155_ & ~new_n156_;
  assign new_n158_ = \A[119]  & ~new_n157_;
  assign new_n159_ = ~new_n154_ & ~new_n158_;
  assign new_n160_ = ~\A[117]  & ~new_n159_;
  assign new_n161_ = ~\A[118]  & ~new_n157_;
  assign new_n162_ = \A[118]  & ~new_n159_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = \A[117]  & ~new_n163_;
  assign new_n165_ = ~new_n160_ & ~new_n164_;
  assign new_n166_ = ~\A[115]  & ~new_n165_;
  assign new_n167_ = ~\A[116]  & ~new_n163_;
  assign new_n168_ = \A[116]  & ~new_n165_;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = \A[115]  & ~new_n169_;
  assign new_n171_ = ~new_n166_ & ~new_n170_;
  assign new_n172_ = ~\A[113]  & ~new_n171_;
  assign new_n173_ = ~\A[114]  & ~new_n169_;
  assign new_n174_ = \A[114]  & ~new_n171_;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = \A[113]  & ~new_n175_;
  assign new_n177_ = ~new_n172_ & ~new_n176_;
  assign new_n178_ = ~\A[111]  & ~new_n177_;
  assign new_n179_ = ~\A[112]  & ~new_n175_;
  assign new_n180_ = \A[112]  & ~new_n177_;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign new_n182_ = \A[111]  & ~new_n181_;
  assign new_n183_ = ~new_n178_ & ~new_n182_;
  assign new_n184_ = ~\A[109]  & ~new_n183_;
  assign new_n185_ = ~\A[110]  & ~new_n181_;
  assign new_n186_ = \A[110]  & ~new_n183_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = \A[109]  & ~new_n187_;
  assign new_n189_ = ~new_n184_ & ~new_n188_;
  assign new_n190_ = ~\A[107]  & ~new_n189_;
  assign new_n191_ = ~\A[108]  & ~new_n187_;
  assign new_n192_ = \A[108]  & ~new_n189_;
  assign new_n193_ = ~new_n191_ & ~new_n192_;
  assign new_n194_ = \A[107]  & ~new_n193_;
  assign new_n195_ = ~new_n190_ & ~new_n194_;
  assign new_n196_ = ~\A[105]  & ~new_n195_;
  assign new_n197_ = ~\A[106]  & ~new_n193_;
  assign new_n198_ = \A[106]  & ~new_n195_;
  assign new_n199_ = ~new_n197_ & ~new_n198_;
  assign new_n200_ = \A[105]  & ~new_n199_;
  assign new_n201_ = ~new_n196_ & ~new_n200_;
  assign new_n202_ = ~\A[103]  & ~new_n201_;
  assign new_n203_ = ~\A[104]  & ~new_n199_;
  assign new_n204_ = \A[104]  & ~new_n201_;
  assign new_n205_ = ~new_n203_ & ~new_n204_;
  assign new_n206_ = \A[103]  & ~new_n205_;
  assign new_n207_ = ~new_n202_ & ~new_n206_;
  assign new_n208_ = ~\A[101]  & ~new_n207_;
  assign new_n209_ = ~\A[102]  & ~new_n205_;
  assign new_n210_ = \A[102]  & ~new_n207_;
  assign new_n211_ = ~new_n209_ & ~new_n210_;
  assign new_n212_ = \A[101]  & ~new_n211_;
  assign new_n213_ = ~new_n208_ & ~new_n212_;
  assign new_n214_ = ~\A[99]  & ~new_n213_;
  assign new_n215_ = ~\A[100]  & ~new_n211_;
  assign new_n216_ = \A[100]  & ~new_n213_;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = \A[99]  & ~new_n217_;
  assign new_n219_ = ~new_n214_ & ~new_n218_;
  assign new_n220_ = ~\A[97]  & ~new_n219_;
  assign new_n221_ = ~\A[98]  & ~new_n217_;
  assign new_n222_ = \A[98]  & ~new_n219_;
  assign new_n223_ = ~new_n221_ & ~new_n222_;
  assign new_n224_ = \A[97]  & ~new_n223_;
  assign new_n225_ = ~new_n220_ & ~new_n224_;
  assign new_n226_ = ~\A[95]  & ~new_n225_;
  assign new_n227_ = ~\A[96]  & ~new_n223_;
  assign new_n228_ = \A[96]  & ~new_n225_;
  assign new_n229_ = ~new_n227_ & ~new_n228_;
  assign new_n230_ = \A[95]  & ~new_n229_;
  assign new_n231_ = ~new_n226_ & ~new_n230_;
  assign new_n232_ = ~\A[93]  & ~new_n231_;
  assign new_n233_ = ~\A[94]  & ~new_n229_;
  assign new_n234_ = \A[94]  & ~new_n231_;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = \A[93]  & ~new_n235_;
  assign new_n237_ = ~new_n232_ & ~new_n236_;
  assign new_n238_ = ~\A[91]  & ~new_n237_;
  assign new_n239_ = ~\A[92]  & ~new_n235_;
  assign new_n240_ = \A[92]  & ~new_n237_;
  assign new_n241_ = ~new_n239_ & ~new_n240_;
  assign new_n242_ = \A[91]  & ~new_n241_;
  assign new_n243_ = ~new_n238_ & ~new_n242_;
  assign new_n244_ = ~\A[89]  & ~new_n243_;
  assign new_n245_ = ~\A[90]  & ~new_n241_;
  assign new_n246_ = \A[90]  & ~new_n243_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = \A[89]  & ~new_n247_;
  assign new_n249_ = ~new_n244_ & ~new_n248_;
  assign new_n250_ = ~\A[87]  & ~new_n249_;
  assign new_n251_ = ~\A[88]  & ~new_n247_;
  assign new_n252_ = \A[88]  & ~new_n249_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = \A[87]  & ~new_n253_;
  assign new_n255_ = ~new_n250_ & ~new_n254_;
  assign new_n256_ = ~\A[85]  & ~new_n255_;
  assign new_n257_ = ~\A[86]  & ~new_n253_;
  assign new_n258_ = \A[86]  & ~new_n255_;
  assign new_n259_ = ~new_n257_ & ~new_n258_;
  assign new_n260_ = \A[85]  & ~new_n259_;
  assign new_n261_ = ~new_n256_ & ~new_n260_;
  assign new_n262_ = ~\A[83]  & ~new_n261_;
  assign new_n263_ = ~\A[84]  & ~new_n259_;
  assign new_n264_ = \A[84]  & ~new_n261_;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = \A[83]  & ~new_n265_;
  assign new_n267_ = ~new_n262_ & ~new_n266_;
  assign new_n268_ = ~\A[81]  & ~new_n267_;
  assign new_n269_ = ~\A[82]  & ~new_n265_;
  assign new_n270_ = \A[82]  & ~new_n267_;
  assign new_n271_ = ~new_n269_ & ~new_n270_;
  assign new_n272_ = \A[81]  & ~new_n271_;
  assign new_n273_ = ~new_n268_ & ~new_n272_;
  assign new_n274_ = ~\A[79]  & ~new_n273_;
  assign new_n275_ = ~\A[80]  & ~new_n271_;
  assign new_n276_ = \A[80]  & ~new_n273_;
  assign new_n277_ = ~new_n275_ & ~new_n276_;
  assign new_n278_ = \A[79]  & ~new_n277_;
  assign new_n279_ = ~new_n274_ & ~new_n278_;
  assign new_n280_ = ~\A[77]  & ~new_n279_;
  assign new_n281_ = ~\A[78]  & ~new_n277_;
  assign new_n282_ = \A[78]  & ~new_n279_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = \A[77]  & ~new_n283_;
  assign new_n285_ = ~new_n280_ & ~new_n284_;
  assign new_n286_ = ~\A[75]  & ~new_n285_;
  assign new_n287_ = ~\A[76]  & ~new_n283_;
  assign new_n288_ = \A[76]  & ~new_n285_;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign new_n290_ = \A[75]  & ~new_n289_;
  assign new_n291_ = ~new_n286_ & ~new_n290_;
  assign new_n292_ = ~\A[73]  & ~new_n291_;
  assign new_n293_ = ~\A[74]  & ~new_n289_;
  assign new_n294_ = \A[74]  & ~new_n291_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = \A[73]  & ~new_n295_;
  assign new_n297_ = ~new_n292_ & ~new_n296_;
  assign new_n298_ = ~\A[71]  & ~new_n297_;
  assign new_n299_ = ~\A[72]  & ~new_n295_;
  assign new_n300_ = \A[72]  & ~new_n297_;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = \A[71]  & ~new_n301_;
  assign new_n303_ = ~new_n298_ & ~new_n302_;
  assign new_n304_ = ~\A[69]  & ~new_n303_;
  assign new_n305_ = ~\A[70]  & ~new_n301_;
  assign new_n306_ = \A[70]  & ~new_n303_;
  assign new_n307_ = ~new_n305_ & ~new_n306_;
  assign new_n308_ = \A[69]  & ~new_n307_;
  assign new_n309_ = ~new_n304_ & ~new_n308_;
  assign new_n310_ = ~\A[67]  & ~new_n309_;
  assign new_n311_ = ~\A[68]  & ~new_n307_;
  assign new_n312_ = \A[68]  & ~new_n309_;
  assign new_n313_ = ~new_n311_ & ~new_n312_;
  assign new_n314_ = \A[67]  & ~new_n313_;
  assign new_n315_ = ~new_n310_ & ~new_n314_;
  assign new_n316_ = ~\A[65]  & ~new_n315_;
  assign new_n317_ = ~\A[66]  & ~new_n313_;
  assign new_n318_ = \A[66]  & ~new_n315_;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = \A[65]  & ~new_n319_;
  assign new_n321_ = ~new_n316_ & ~new_n320_;
  assign new_n322_ = ~\A[63]  & ~new_n321_;
  assign new_n323_ = ~\A[64]  & ~new_n319_;
  assign new_n324_ = \A[64]  & ~new_n321_;
  assign new_n325_ = ~new_n323_ & ~new_n324_;
  assign new_n326_ = \A[63]  & ~new_n325_;
  assign new_n327_ = ~new_n322_ & ~new_n326_;
  assign new_n328_ = ~\A[61]  & ~new_n327_;
  assign new_n329_ = ~\A[62]  & ~new_n325_;
  assign new_n330_ = \A[62]  & ~new_n327_;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = \A[61]  & ~new_n331_;
  assign new_n333_ = ~new_n328_ & ~new_n332_;
  assign new_n334_ = ~\A[59]  & ~new_n333_;
  assign new_n335_ = ~\A[60]  & ~new_n331_;
  assign new_n336_ = \A[60]  & ~new_n333_;
  assign new_n337_ = ~new_n335_ & ~new_n336_;
  assign new_n338_ = \A[59]  & ~new_n337_;
  assign new_n339_ = ~new_n334_ & ~new_n338_;
  assign new_n340_ = ~\A[57]  & ~new_n339_;
  assign new_n341_ = ~\A[58]  & ~new_n337_;
  assign new_n342_ = \A[58]  & ~new_n339_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = \A[57]  & ~new_n343_;
  assign new_n345_ = ~new_n340_ & ~new_n344_;
  assign new_n346_ = ~\A[55]  & ~new_n345_;
  assign new_n347_ = ~\A[56]  & ~new_n343_;
  assign new_n348_ = \A[56]  & ~new_n345_;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_ = \A[55]  & ~new_n349_;
  assign new_n351_ = ~new_n346_ & ~new_n350_;
  assign new_n352_ = ~\A[53]  & ~new_n351_;
  assign new_n353_ = ~\A[54]  & ~new_n349_;
  assign new_n354_ = \A[54]  & ~new_n351_;
  assign new_n355_ = ~new_n353_ & ~new_n354_;
  assign new_n356_ = \A[53]  & ~new_n355_;
  assign new_n357_ = ~new_n352_ & ~new_n356_;
  assign new_n358_ = ~\A[51]  & ~new_n357_;
  assign new_n359_ = ~\A[52]  & ~new_n355_;
  assign new_n360_ = \A[52]  & ~new_n357_;
  assign new_n361_ = ~new_n359_ & ~new_n360_;
  assign new_n362_ = \A[51]  & ~new_n361_;
  assign new_n363_ = ~new_n358_ & ~new_n362_;
  assign new_n364_ = ~\A[49]  & ~new_n363_;
  assign new_n365_ = ~\A[50]  & ~new_n361_;
  assign new_n366_ = \A[50]  & ~new_n363_;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = \A[49]  & ~new_n367_;
  assign new_n369_ = ~new_n364_ & ~new_n368_;
  assign new_n370_ = ~\A[47]  & ~new_n369_;
  assign new_n371_ = ~\A[48]  & ~new_n367_;
  assign new_n372_ = \A[48]  & ~new_n369_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = \A[47]  & ~new_n373_;
  assign new_n375_ = ~new_n370_ & ~new_n374_;
  assign new_n376_ = ~\A[45]  & ~new_n375_;
  assign new_n377_ = ~\A[46]  & ~new_n373_;
  assign new_n378_ = \A[46]  & ~new_n375_;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_ = \A[45]  & ~new_n379_;
  assign new_n381_ = ~new_n376_ & ~new_n380_;
  assign new_n382_ = ~\A[43]  & ~new_n381_;
  assign new_n383_ = ~\A[44]  & ~new_n379_;
  assign new_n384_ = \A[44]  & ~new_n381_;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = \A[43]  & ~new_n385_;
  assign new_n387_ = ~new_n382_ & ~new_n386_;
  assign new_n388_ = ~\A[41]  & ~new_n387_;
  assign new_n389_ = ~\A[42]  & ~new_n385_;
  assign new_n390_ = \A[42]  & ~new_n387_;
  assign new_n391_ = ~new_n389_ & ~new_n390_;
  assign new_n392_ = \A[41]  & ~new_n391_;
  assign new_n393_ = ~new_n388_ & ~new_n392_;
  assign new_n394_ = ~\A[39]  & ~new_n393_;
  assign new_n395_ = ~\A[40]  & ~new_n391_;
  assign new_n396_ = \A[40]  & ~new_n393_;
  assign new_n397_ = ~new_n395_ & ~new_n396_;
  assign new_n398_ = \A[39]  & ~new_n397_;
  assign new_n399_ = ~new_n394_ & ~new_n398_;
  assign new_n400_ = ~\A[37]  & ~new_n399_;
  assign new_n401_ = ~\A[38]  & ~new_n397_;
  assign new_n402_ = \A[38]  & ~new_n399_;
  assign new_n403_ = ~new_n401_ & ~new_n402_;
  assign new_n404_ = \A[37]  & ~new_n403_;
  assign new_n405_ = ~new_n400_ & ~new_n404_;
  assign new_n406_ = ~\A[35]  & ~new_n405_;
  assign new_n407_ = ~\A[36]  & ~new_n403_;
  assign new_n408_ = \A[36]  & ~new_n405_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = \A[35]  & ~new_n409_;
  assign new_n411_ = ~new_n406_ & ~new_n410_;
  assign new_n412_ = ~\A[33]  & ~new_n411_;
  assign new_n413_ = ~\A[34]  & ~new_n409_;
  assign new_n414_ = \A[34]  & ~new_n411_;
  assign new_n415_ = ~new_n413_ & ~new_n414_;
  assign new_n416_ = \A[33]  & ~new_n415_;
  assign new_n417_ = ~new_n412_ & ~new_n416_;
  assign new_n418_ = ~\A[31]  & ~new_n417_;
  assign new_n419_ = ~\A[32]  & ~new_n415_;
  assign new_n420_ = \A[32]  & ~new_n417_;
  assign new_n421_ = ~new_n419_ & ~new_n420_;
  assign new_n422_ = \A[31]  & ~new_n421_;
  assign new_n423_ = ~new_n418_ & ~new_n422_;
  assign new_n424_ = ~\A[29]  & ~new_n423_;
  assign new_n425_ = ~\A[30]  & ~new_n421_;
  assign new_n426_ = \A[30]  & ~new_n423_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = \A[29]  & ~new_n427_;
  assign new_n429_ = ~new_n424_ & ~new_n428_;
  assign new_n430_ = ~\A[27]  & ~new_n429_;
  assign new_n431_ = ~\A[28]  & ~new_n427_;
  assign new_n432_ = \A[28]  & ~new_n429_;
  assign new_n433_ = ~new_n431_ & ~new_n432_;
  assign new_n434_ = \A[27]  & ~new_n433_;
  assign new_n435_ = ~new_n430_ & ~new_n434_;
  assign new_n436_ = ~\A[25]  & ~new_n435_;
  assign new_n437_ = ~\A[26]  & ~new_n433_;
  assign new_n438_ = \A[26]  & ~new_n435_;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign new_n440_ = \A[25]  & ~new_n439_;
  assign new_n441_ = ~new_n436_ & ~new_n440_;
  assign new_n442_ = ~\A[23]  & ~new_n441_;
  assign new_n443_ = ~\A[24]  & ~new_n439_;
  assign new_n444_ = \A[24]  & ~new_n441_;
  assign new_n445_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = \A[23]  & ~new_n445_;
  assign new_n447_ = ~new_n442_ & ~new_n446_;
  assign new_n448_ = ~\A[21]  & ~new_n447_;
  assign new_n449_ = ~\A[22]  & ~new_n445_;
  assign new_n450_ = \A[22]  & ~new_n447_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = \A[21]  & ~new_n451_;
  assign new_n453_ = ~new_n448_ & ~new_n452_;
  assign new_n454_ = ~\A[19]  & ~new_n453_;
  assign new_n455_ = ~\A[20]  & ~new_n451_;
  assign new_n456_ = \A[20]  & ~new_n453_;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_ = \A[19]  & ~new_n457_;
  assign new_n459_ = ~new_n454_ & ~new_n458_;
  assign new_n460_ = ~\A[17]  & ~new_n459_;
  assign new_n461_ = ~\A[18]  & ~new_n457_;
  assign new_n462_ = \A[18]  & ~new_n459_;
  assign new_n463_ = ~new_n461_ & ~new_n462_;
  assign new_n464_ = \A[17]  & ~new_n463_;
  assign new_n465_ = ~new_n460_ & ~new_n464_;
  assign new_n466_ = ~\A[15]  & ~new_n465_;
  assign new_n467_ = ~\A[16]  & ~new_n463_;
  assign new_n468_ = \A[16]  & ~new_n465_;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_ = \A[15]  & ~new_n469_;
  assign new_n471_ = ~new_n466_ & ~new_n470_;
  assign new_n472_ = ~\A[13]  & ~new_n471_;
  assign new_n473_ = ~\A[14]  & ~new_n469_;
  assign new_n474_ = \A[14]  & ~new_n471_;
  assign new_n475_ = ~new_n473_ & ~new_n474_;
  assign new_n476_ = \A[13]  & ~new_n475_;
  assign new_n477_ = ~new_n472_ & ~new_n476_;
  assign new_n478_ = ~\A[11]  & ~new_n477_;
  assign new_n479_ = ~\A[12]  & ~new_n475_;
  assign new_n480_ = \A[12]  & ~new_n477_;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = \A[11]  & ~new_n481_;
  assign new_n483_ = ~new_n478_ & ~new_n482_;
  assign new_n484_ = ~\A[9]  & ~new_n483_;
  assign new_n485_ = ~\A[10]  & ~new_n481_;
  assign new_n486_ = \A[10]  & ~new_n483_;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = \A[9]  & ~new_n487_;
  assign new_n489_ = ~new_n484_ & ~new_n488_;
  assign new_n490_ = ~\A[7]  & ~new_n489_;
  assign new_n491_ = ~\A[8]  & ~new_n487_;
  assign new_n492_ = \A[8]  & ~new_n489_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = \A[7]  & ~new_n493_;
  assign new_n495_ = ~new_n490_ & ~new_n494_;
  assign new_n496_ = ~\A[5]  & ~new_n495_;
  assign new_n497_ = ~\A[6]  & ~new_n493_;
  assign new_n498_ = \A[6]  & ~new_n495_;
  assign new_n499_ = ~new_n497_ & ~new_n498_;
  assign new_n500_ = \A[5]  & ~new_n499_;
  assign new_n501_ = ~new_n496_ & ~new_n500_;
  assign new_n502_ = ~\A[3]  & ~new_n501_;
  assign new_n503_ = ~\A[4]  & ~new_n499_;
  assign new_n504_ = \A[4]  & ~new_n501_;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = \A[3]  & ~new_n505_;
  assign new_n507_ = ~new_n502_ & ~new_n506_;
  assign new_n508_ = \A[1]  & ~\A[2] ;
  assign new_n509_ = new_n507_ & ~new_n508_;
  assign new_n510_ = new_n505_ & new_n508_;
  assign \P[0]  = ~new_n509_ & ~new_n510_;
  assign new_n512_ = ~\A[126]  & \A[127] ;
  assign new_n513_ = ~\A[126]  & ~new_n512_;
  assign new_n514_ = ~\A[124]  & ~\A[125] ;
  assign new_n515_ = ~\A[122]  & ~\A[123] ;
  assign new_n516_ = \A[121]  & new_n515_;
  assign new_n517_ = new_n514_ & ~new_n516_;
  assign new_n518_ = new_n513_ & ~new_n517_;
  assign new_n519_ = ~\A[120]  & ~new_n518_;
  assign new_n520_ = new_n514_ & ~new_n515_;
  assign new_n521_ = new_n513_ & ~new_n520_;
  assign new_n522_ = \A[120]  & ~new_n521_;
  assign new_n523_ = ~new_n519_ & ~new_n522_;
  assign new_n524_ = ~\A[118]  & ~\A[119] ;
  assign new_n525_ = new_n523_ & ~new_n524_;
  assign new_n526_ = new_n521_ & new_n524_;
  assign new_n527_ = ~new_n525_ & ~new_n526_;
  assign new_n528_ = ~\A[116]  & ~\A[117] ;
  assign new_n529_ = new_n527_ & ~new_n528_;
  assign new_n530_ = ~new_n523_ & new_n528_;
  assign new_n531_ = ~new_n529_ & ~new_n530_;
  assign new_n532_ = ~\A[114]  & ~\A[115] ;
  assign new_n533_ = new_n531_ & ~new_n532_;
  assign new_n534_ = ~new_n527_ & new_n532_;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~\A[112]  & ~\A[113] ;
  assign new_n537_ = new_n535_ & ~new_n536_;
  assign new_n538_ = ~new_n531_ & new_n536_;
  assign new_n539_ = ~new_n537_ & ~new_n538_;
  assign new_n540_ = ~\A[110]  & ~\A[111] ;
  assign new_n541_ = new_n539_ & ~new_n540_;
  assign new_n542_ = ~new_n535_ & new_n540_;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = ~\A[108]  & ~\A[109] ;
  assign new_n545_ = new_n543_ & ~new_n544_;
  assign new_n546_ = ~new_n539_ & new_n544_;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = ~\A[106]  & ~\A[107] ;
  assign new_n549_ = new_n547_ & ~new_n548_;
  assign new_n550_ = ~new_n543_ & new_n548_;
  assign new_n551_ = ~new_n549_ & ~new_n550_;
  assign new_n552_ = ~\A[104]  & ~\A[105] ;
  assign new_n553_ = new_n551_ & ~new_n552_;
  assign new_n554_ = ~new_n547_ & new_n552_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = ~\A[102]  & ~\A[103] ;
  assign new_n557_ = new_n555_ & ~new_n556_;
  assign new_n558_ = ~new_n551_ & new_n556_;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = ~\A[100]  & ~\A[101] ;
  assign new_n561_ = new_n559_ & ~new_n560_;
  assign new_n562_ = ~new_n555_ & new_n560_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = ~\A[98]  & ~\A[99] ;
  assign new_n565_ = new_n563_ & ~new_n564_;
  assign new_n566_ = ~new_n559_ & new_n564_;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = ~\A[96]  & ~\A[97] ;
  assign new_n569_ = new_n567_ & ~new_n568_;
  assign new_n570_ = ~new_n563_ & new_n568_;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign new_n572_ = ~\A[94]  & ~\A[95] ;
  assign new_n573_ = new_n571_ & ~new_n572_;
  assign new_n574_ = ~new_n567_ & new_n572_;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = ~\A[92]  & ~\A[93] ;
  assign new_n577_ = new_n575_ & ~new_n576_;
  assign new_n578_ = ~new_n571_ & new_n576_;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign new_n580_ = ~\A[90]  & ~\A[91] ;
  assign new_n581_ = new_n579_ & ~new_n580_;
  assign new_n582_ = ~new_n575_ & new_n580_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = ~\A[88]  & ~\A[89] ;
  assign new_n585_ = new_n583_ & ~new_n584_;
  assign new_n586_ = ~new_n579_ & new_n584_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~\A[86]  & ~\A[87] ;
  assign new_n589_ = new_n587_ & ~new_n588_;
  assign new_n590_ = ~new_n583_ & new_n588_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~\A[84]  & ~\A[85] ;
  assign new_n593_ = new_n591_ & ~new_n592_;
  assign new_n594_ = ~new_n587_ & new_n592_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~\A[82]  & ~\A[83] ;
  assign new_n597_ = new_n595_ & ~new_n596_;
  assign new_n598_ = ~new_n591_ & new_n596_;
  assign new_n599_ = ~new_n597_ & ~new_n598_;
  assign new_n600_ = ~\A[80]  & ~\A[81] ;
  assign new_n601_ = new_n599_ & ~new_n600_;
  assign new_n602_ = ~new_n595_ & new_n600_;
  assign new_n603_ = ~new_n601_ & ~new_n602_;
  assign new_n604_ = ~\A[78]  & ~\A[79] ;
  assign new_n605_ = new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n599_ & new_n604_;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign new_n608_ = ~\A[76]  & ~\A[77] ;
  assign new_n609_ = new_n607_ & ~new_n608_;
  assign new_n610_ = ~new_n603_ & new_n608_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = ~\A[74]  & ~\A[75] ;
  assign new_n613_ = new_n611_ & ~new_n612_;
  assign new_n614_ = ~new_n607_ & new_n612_;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign new_n616_ = ~\A[72]  & ~\A[73] ;
  assign new_n617_ = new_n615_ & ~new_n616_;
  assign new_n618_ = ~new_n611_ & new_n616_;
  assign new_n619_ = ~new_n617_ & ~new_n618_;
  assign new_n620_ = ~\A[70]  & ~\A[71] ;
  assign new_n621_ = new_n619_ & ~new_n620_;
  assign new_n622_ = ~new_n615_ & new_n620_;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_ = ~\A[68]  & ~\A[69] ;
  assign new_n625_ = new_n623_ & ~new_n624_;
  assign new_n626_ = ~new_n619_ & new_n624_;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign new_n628_ = ~\A[66]  & ~\A[67] ;
  assign new_n629_ = new_n627_ & ~new_n628_;
  assign new_n630_ = ~new_n623_ & new_n628_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = ~\A[64]  & ~\A[65] ;
  assign new_n633_ = new_n631_ & ~new_n632_;
  assign new_n634_ = ~new_n627_ & new_n632_;
  assign new_n635_ = ~new_n633_ & ~new_n634_;
  assign new_n636_ = ~\A[62]  & ~\A[63] ;
  assign new_n637_ = new_n635_ & ~new_n636_;
  assign new_n638_ = ~new_n631_ & new_n636_;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign new_n640_ = ~\A[60]  & ~\A[61] ;
  assign new_n641_ = new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n635_ & new_n640_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = ~\A[58]  & ~\A[59] ;
  assign new_n645_ = new_n643_ & ~new_n644_;
  assign new_n646_ = ~new_n639_ & new_n644_;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = ~\A[56]  & ~\A[57] ;
  assign new_n649_ = new_n647_ & ~new_n648_;
  assign new_n650_ = ~new_n643_ & new_n648_;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = ~\A[54]  & ~\A[55] ;
  assign new_n653_ = new_n651_ & ~new_n652_;
  assign new_n654_ = ~new_n647_ & new_n652_;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign new_n656_ = ~\A[52]  & ~\A[53] ;
  assign new_n657_ = new_n655_ & ~new_n656_;
  assign new_n658_ = ~new_n651_ & new_n656_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~\A[50]  & ~\A[51] ;
  assign new_n661_ = new_n659_ & ~new_n660_;
  assign new_n662_ = ~new_n655_ & new_n660_;
  assign new_n663_ = ~new_n661_ & ~new_n662_;
  assign new_n664_ = ~\A[48]  & ~\A[49] ;
  assign new_n665_ = new_n663_ & ~new_n664_;
  assign new_n666_ = ~new_n659_ & new_n664_;
  assign new_n667_ = ~new_n665_ & ~new_n666_;
  assign new_n668_ = ~\A[46]  & ~\A[47] ;
  assign new_n669_ = new_n667_ & ~new_n668_;
  assign new_n670_ = ~new_n663_ & new_n668_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~\A[44]  & ~\A[45] ;
  assign new_n673_ = new_n671_ & ~new_n672_;
  assign new_n674_ = ~new_n667_ & new_n672_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = ~\A[42]  & ~\A[43] ;
  assign new_n677_ = new_n675_ & ~new_n676_;
  assign new_n678_ = ~new_n671_ & new_n676_;
  assign new_n679_ = ~new_n677_ & ~new_n678_;
  assign new_n680_ = ~\A[40]  & ~\A[41] ;
  assign new_n681_ = new_n679_ & ~new_n680_;
  assign new_n682_ = ~new_n675_ & new_n680_;
  assign new_n683_ = ~new_n681_ & ~new_n682_;
  assign new_n684_ = ~\A[38]  & ~\A[39] ;
  assign new_n685_ = new_n683_ & ~new_n684_;
  assign new_n686_ = ~new_n679_ & new_n684_;
  assign new_n687_ = ~new_n685_ & ~new_n686_;
  assign new_n688_ = ~\A[36]  & ~\A[37] ;
  assign new_n689_ = new_n687_ & ~new_n688_;
  assign new_n690_ = ~new_n683_ & new_n688_;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = ~\A[34]  & ~\A[35] ;
  assign new_n693_ = new_n691_ & ~new_n692_;
  assign new_n694_ = ~new_n687_ & new_n692_;
  assign new_n695_ = ~new_n693_ & ~new_n694_;
  assign new_n696_ = ~\A[32]  & ~\A[33] ;
  assign new_n697_ = new_n695_ & ~new_n696_;
  assign new_n698_ = ~new_n691_ & new_n696_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign new_n700_ = ~\A[30]  & ~\A[31] ;
  assign new_n701_ = new_n699_ & ~new_n700_;
  assign new_n702_ = ~new_n695_ & new_n700_;
  assign new_n703_ = ~new_n701_ & ~new_n702_;
  assign new_n704_ = ~\A[28]  & ~\A[29] ;
  assign new_n705_ = new_n703_ & ~new_n704_;
  assign new_n706_ = ~new_n699_ & new_n704_;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign new_n708_ = ~\A[26]  & ~\A[27] ;
  assign new_n709_ = new_n707_ & ~new_n708_;
  assign new_n710_ = ~new_n703_ & new_n708_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = ~\A[24]  & ~\A[25] ;
  assign new_n713_ = new_n711_ & ~new_n712_;
  assign new_n714_ = ~new_n707_ & new_n712_;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = ~\A[22]  & ~\A[23] ;
  assign new_n717_ = new_n715_ & ~new_n716_;
  assign new_n718_ = ~new_n711_ & new_n716_;
  assign new_n719_ = ~new_n717_ & ~new_n718_;
  assign new_n720_ = ~\A[20]  & ~\A[21] ;
  assign new_n721_ = new_n719_ & ~new_n720_;
  assign new_n722_ = ~new_n715_ & new_n720_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = ~\A[18]  & ~\A[19] ;
  assign new_n725_ = new_n723_ & ~new_n724_;
  assign new_n726_ = ~new_n719_ & new_n724_;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = ~\A[16]  & ~\A[17] ;
  assign new_n729_ = new_n727_ & ~new_n728_;
  assign new_n730_ = ~new_n723_ & new_n728_;
  assign new_n731_ = ~new_n729_ & ~new_n730_;
  assign new_n732_ = ~\A[14]  & ~\A[15] ;
  assign new_n733_ = new_n731_ & ~new_n732_;
  assign new_n734_ = ~new_n727_ & new_n732_;
  assign new_n735_ = ~new_n733_ & ~new_n734_;
  assign new_n736_ = ~\A[12]  & ~\A[13] ;
  assign new_n737_ = new_n735_ & ~new_n736_;
  assign new_n738_ = ~new_n731_ & new_n736_;
  assign new_n739_ = ~new_n737_ & ~new_n738_;
  assign new_n740_ = ~\A[10]  & ~\A[11] ;
  assign new_n741_ = new_n739_ & ~new_n740_;
  assign new_n742_ = ~new_n735_ & new_n740_;
  assign new_n743_ = ~new_n741_ & ~new_n742_;
  assign new_n744_ = ~\A[8]  & ~\A[9] ;
  assign new_n745_ = new_n743_ & ~new_n744_;
  assign new_n746_ = ~new_n739_ & new_n744_;
  assign new_n747_ = ~new_n745_ & ~new_n746_;
  assign new_n748_ = ~\A[6]  & ~\A[7] ;
  assign new_n749_ = new_n747_ & ~new_n748_;
  assign new_n750_ = ~new_n743_ & new_n748_;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign new_n752_ = ~\A[4]  & ~\A[5] ;
  assign new_n753_ = new_n751_ & ~new_n752_;
  assign new_n754_ = ~new_n747_ & new_n752_;
  assign new_n755_ = ~new_n753_ & ~new_n754_;
  assign new_n756_ = ~\A[2]  & ~\A[3] ;
  assign new_n757_ = new_n755_ & ~new_n756_;
  assign new_n758_ = ~new_n751_ & new_n756_;
  assign \P[1]  = ~new_n757_ & ~new_n758_;
  assign new_n760_ = new_n513_ & new_n514_;
  assign new_n761_ = ~\A[120]  & ~\A[121] ;
  assign new_n762_ = new_n515_ & new_n761_;
  assign new_n763_ = ~\A[117]  & new_n524_;
  assign new_n764_ = ~\A[116]  & new_n763_;
  assign new_n765_ = new_n762_ & ~new_n764_;
  assign new_n766_ = new_n760_ & ~new_n765_;
  assign new_n767_ = ~\A[113]  & ~\A[114] ;
  assign new_n768_ = ~\A[112]  & new_n767_;
  assign new_n769_ = new_n766_ & ~new_n768_;
  assign new_n770_ = \A[115]  & new_n764_;
  assign new_n771_ = new_n762_ & ~new_n770_;
  assign new_n772_ = new_n760_ & ~new_n771_;
  assign new_n773_ = new_n768_ & new_n772_;
  assign new_n774_ = ~new_n769_ & ~new_n773_;
  assign new_n775_ = ~\A[109]  & new_n540_;
  assign new_n776_ = ~\A[108]  & new_n775_;
  assign new_n777_ = new_n774_ & ~new_n776_;
  assign new_n778_ = ~new_n766_ & new_n776_;
  assign new_n779_ = ~new_n777_ & ~new_n778_;
  assign new_n780_ = ~\A[105]  & new_n548_;
  assign new_n781_ = ~\A[104]  & new_n780_;
  assign new_n782_ = new_n779_ & ~new_n781_;
  assign new_n783_ = ~new_n774_ & new_n781_;
  assign new_n784_ = ~new_n782_ & ~new_n783_;
  assign new_n785_ = ~\A[101]  & new_n556_;
  assign new_n786_ = ~\A[100]  & new_n785_;
  assign new_n787_ = new_n784_ & ~new_n786_;
  assign new_n788_ = ~new_n779_ & new_n786_;
  assign new_n789_ = ~new_n787_ & ~new_n788_;
  assign new_n790_ = ~\A[97]  & new_n564_;
  assign new_n791_ = ~\A[96]  & new_n790_;
  assign new_n792_ = new_n789_ & ~new_n791_;
  assign new_n793_ = ~new_n784_ & new_n791_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = ~\A[93]  & new_n572_;
  assign new_n796_ = ~\A[92]  & new_n795_;
  assign new_n797_ = new_n794_ & ~new_n796_;
  assign new_n798_ = ~new_n789_ & new_n796_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = ~\A[89]  & new_n580_;
  assign new_n801_ = ~\A[88]  & new_n800_;
  assign new_n802_ = new_n799_ & ~new_n801_;
  assign new_n803_ = ~new_n794_ & new_n801_;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = ~\A[85]  & new_n588_;
  assign new_n806_ = ~\A[84]  & new_n805_;
  assign new_n807_ = new_n804_ & ~new_n806_;
  assign new_n808_ = ~new_n799_ & new_n806_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = ~\A[81]  & new_n596_;
  assign new_n811_ = ~\A[80]  & new_n810_;
  assign new_n812_ = new_n809_ & ~new_n811_;
  assign new_n813_ = ~new_n804_ & new_n811_;
  assign new_n814_ = ~new_n812_ & ~new_n813_;
  assign new_n815_ = ~\A[77]  & new_n604_;
  assign new_n816_ = ~\A[76]  & new_n815_;
  assign new_n817_ = new_n814_ & ~new_n816_;
  assign new_n818_ = ~new_n809_ & new_n816_;
  assign new_n819_ = ~new_n817_ & ~new_n818_;
  assign new_n820_ = ~\A[73]  & new_n612_;
  assign new_n821_ = ~\A[72]  & new_n820_;
  assign new_n822_ = new_n819_ & ~new_n821_;
  assign new_n823_ = ~new_n814_ & new_n821_;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = ~\A[69]  & new_n620_;
  assign new_n826_ = ~\A[68]  & new_n825_;
  assign new_n827_ = new_n824_ & ~new_n826_;
  assign new_n828_ = ~new_n819_ & new_n826_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~\A[65]  & new_n628_;
  assign new_n831_ = ~\A[64]  & new_n830_;
  assign new_n832_ = new_n829_ & ~new_n831_;
  assign new_n833_ = ~new_n824_ & new_n831_;
  assign new_n834_ = ~new_n832_ & ~new_n833_;
  assign new_n835_ = ~\A[61]  & new_n636_;
  assign new_n836_ = ~\A[60]  & new_n835_;
  assign new_n837_ = new_n834_ & ~new_n836_;
  assign new_n838_ = ~new_n829_ & new_n836_;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = ~\A[57]  & new_n644_;
  assign new_n841_ = ~\A[56]  & new_n840_;
  assign new_n842_ = new_n839_ & ~new_n841_;
  assign new_n843_ = ~new_n834_ & new_n841_;
  assign new_n844_ = ~new_n842_ & ~new_n843_;
  assign new_n845_ = ~\A[53]  & new_n652_;
  assign new_n846_ = ~\A[52]  & new_n845_;
  assign new_n847_ = new_n844_ & ~new_n846_;
  assign new_n848_ = ~new_n839_ & new_n846_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = ~\A[49]  & new_n660_;
  assign new_n851_ = ~\A[48]  & new_n850_;
  assign new_n852_ = new_n849_ & ~new_n851_;
  assign new_n853_ = ~new_n844_ & new_n851_;
  assign new_n854_ = ~new_n852_ & ~new_n853_;
  assign new_n855_ = ~\A[45]  & new_n668_;
  assign new_n856_ = ~\A[44]  & new_n855_;
  assign new_n857_ = new_n854_ & ~new_n856_;
  assign new_n858_ = ~new_n849_ & new_n856_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~\A[41]  & new_n676_;
  assign new_n861_ = ~\A[40]  & new_n860_;
  assign new_n862_ = new_n859_ & ~new_n861_;
  assign new_n863_ = ~new_n854_ & new_n861_;
  assign new_n864_ = ~new_n862_ & ~new_n863_;
  assign new_n865_ = ~\A[37]  & new_n684_;
  assign new_n866_ = ~\A[36]  & new_n865_;
  assign new_n867_ = new_n864_ & ~new_n866_;
  assign new_n868_ = ~new_n859_ & new_n866_;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = ~\A[33]  & new_n692_;
  assign new_n871_ = ~\A[32]  & new_n870_;
  assign new_n872_ = new_n869_ & ~new_n871_;
  assign new_n873_ = ~new_n864_ & new_n871_;
  assign new_n874_ = ~new_n872_ & ~new_n873_;
  assign new_n875_ = ~\A[29]  & new_n700_;
  assign new_n876_ = ~\A[28]  & new_n875_;
  assign new_n877_ = new_n874_ & ~new_n876_;
  assign new_n878_ = ~new_n869_ & new_n876_;
  assign new_n879_ = ~new_n877_ & ~new_n878_;
  assign new_n880_ = ~\A[25]  & new_n708_;
  assign new_n881_ = ~\A[24]  & new_n880_;
  assign new_n882_ = new_n879_ & ~new_n881_;
  assign new_n883_ = ~new_n874_ & new_n881_;
  assign new_n884_ = ~new_n882_ & ~new_n883_;
  assign new_n885_ = ~\A[21]  & new_n716_;
  assign new_n886_ = ~\A[20]  & new_n885_;
  assign new_n887_ = new_n884_ & ~new_n886_;
  assign new_n888_ = ~new_n879_ & new_n886_;
  assign new_n889_ = ~new_n887_ & ~new_n888_;
  assign new_n890_ = ~\A[17]  & new_n724_;
  assign new_n891_ = ~\A[16]  & new_n890_;
  assign new_n892_ = new_n889_ & ~new_n891_;
  assign new_n893_ = ~new_n884_ & new_n891_;
  assign new_n894_ = ~new_n892_ & ~new_n893_;
  assign new_n895_ = ~\A[13]  & new_n732_;
  assign new_n896_ = ~\A[12]  & new_n895_;
  assign new_n897_ = new_n894_ & ~new_n896_;
  assign new_n898_ = ~new_n889_ & new_n896_;
  assign new_n899_ = ~new_n897_ & ~new_n898_;
  assign new_n900_ = ~\A[9]  & new_n740_;
  assign new_n901_ = ~\A[8]  & new_n900_;
  assign new_n902_ = new_n899_ & ~new_n901_;
  assign new_n903_ = ~new_n894_ & new_n901_;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = ~\A[5]  & new_n748_;
  assign new_n906_ = ~\A[4]  & new_n905_;
  assign new_n907_ = new_n904_ & ~new_n906_;
  assign new_n908_ = ~new_n899_ & new_n906_;
  assign \P[2]  = new_n907_ | new_n908_;
  assign new_n910_ = new_n760_ & new_n762_;
  assign new_n911_ = ~\A[113]  & new_n532_;
  assign new_n912_ = ~\A[112]  & new_n764_;
  assign new_n913_ = new_n911_ & new_n912_;
  assign new_n914_ = ~\A[107]  & new_n776_;
  assign new_n915_ = ~\A[106]  & new_n914_;
  assign new_n916_ = ~\A[105]  & new_n915_;
  assign new_n917_ = ~\A[104]  & new_n916_;
  assign new_n918_ = new_n913_ & ~new_n917_;
  assign new_n919_ = new_n910_ & ~new_n918_;
  assign new_n920_ = ~\A[101]  & ~\A[102] ;
  assign new_n921_ = ~\A[100]  & new_n920_;
  assign new_n922_ = ~\A[99]  & new_n921_;
  assign new_n923_ = ~\A[98]  & new_n922_;
  assign new_n924_ = ~\A[97]  & new_n923_;
  assign new_n925_ = ~\A[96]  & new_n924_;
  assign new_n926_ = new_n919_ & ~new_n925_;
  assign new_n927_ = \A[103]  & new_n917_;
  assign new_n928_ = new_n913_ & ~new_n927_;
  assign new_n929_ = new_n910_ & ~new_n928_;
  assign new_n930_ = new_n925_ & new_n929_;
  assign new_n931_ = ~new_n926_ & ~new_n930_;
  assign new_n932_ = ~\A[91]  & new_n796_;
  assign new_n933_ = ~\A[90]  & new_n932_;
  assign new_n934_ = ~\A[89]  & new_n933_;
  assign new_n935_ = ~\A[88]  & new_n934_;
  assign new_n936_ = new_n931_ & ~new_n935_;
  assign new_n937_ = ~new_n919_ & new_n935_;
  assign new_n938_ = ~new_n936_ & ~new_n937_;
  assign new_n939_ = ~\A[83]  & new_n806_;
  assign new_n940_ = ~\A[82]  & new_n939_;
  assign new_n941_ = ~\A[81]  & new_n940_;
  assign new_n942_ = ~\A[80]  & new_n941_;
  assign new_n943_ = new_n938_ & ~new_n942_;
  assign new_n944_ = ~new_n931_ & new_n942_;
  assign new_n945_ = ~new_n943_ & ~new_n944_;
  assign new_n946_ = ~\A[75]  & new_n816_;
  assign new_n947_ = ~\A[74]  & new_n946_;
  assign new_n948_ = ~\A[73]  & new_n947_;
  assign new_n949_ = ~\A[72]  & new_n948_;
  assign new_n950_ = new_n945_ & ~new_n949_;
  assign new_n951_ = ~new_n938_ & new_n949_;
  assign new_n952_ = ~new_n950_ & ~new_n951_;
  assign new_n953_ = ~\A[67]  & new_n826_;
  assign new_n954_ = ~\A[66]  & new_n953_;
  assign new_n955_ = ~\A[65]  & new_n954_;
  assign new_n956_ = ~\A[64]  & new_n955_;
  assign new_n957_ = new_n952_ & ~new_n956_;
  assign new_n958_ = ~new_n945_ & new_n956_;
  assign new_n959_ = ~new_n957_ & ~new_n958_;
  assign new_n960_ = ~\A[59]  & new_n836_;
  assign new_n961_ = ~\A[58]  & new_n960_;
  assign new_n962_ = ~\A[57]  & new_n961_;
  assign new_n963_ = ~\A[56]  & new_n962_;
  assign new_n964_ = new_n959_ & ~new_n963_;
  assign new_n965_ = ~new_n952_ & new_n963_;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = ~\A[51]  & new_n846_;
  assign new_n968_ = ~\A[50]  & new_n967_;
  assign new_n969_ = ~\A[49]  & new_n968_;
  assign new_n970_ = ~\A[48]  & new_n969_;
  assign new_n971_ = new_n966_ & ~new_n970_;
  assign new_n972_ = ~new_n959_ & new_n970_;
  assign new_n973_ = ~new_n971_ & ~new_n972_;
  assign new_n974_ = ~\A[43]  & new_n856_;
  assign new_n975_ = ~\A[42]  & new_n974_;
  assign new_n976_ = ~\A[41]  & new_n975_;
  assign new_n977_ = ~\A[40]  & new_n976_;
  assign new_n978_ = new_n973_ & ~new_n977_;
  assign new_n979_ = ~new_n966_ & new_n977_;
  assign new_n980_ = ~new_n978_ & ~new_n979_;
  assign new_n981_ = ~\A[35]  & new_n866_;
  assign new_n982_ = ~\A[34]  & new_n981_;
  assign new_n983_ = ~\A[33]  & new_n982_;
  assign new_n984_ = ~\A[32]  & new_n983_;
  assign new_n985_ = new_n980_ & ~new_n984_;
  assign new_n986_ = ~new_n973_ & new_n984_;
  assign new_n987_ = ~new_n985_ & ~new_n986_;
  assign new_n988_ = ~\A[27]  & new_n876_;
  assign new_n989_ = ~\A[26]  & new_n988_;
  assign new_n990_ = ~\A[25]  & new_n989_;
  assign new_n991_ = ~\A[24]  & new_n990_;
  assign new_n992_ = new_n987_ & ~new_n991_;
  assign new_n993_ = ~new_n980_ & new_n991_;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign new_n995_ = ~\A[19]  & new_n886_;
  assign new_n996_ = ~\A[18]  & new_n995_;
  assign new_n997_ = ~\A[17]  & new_n996_;
  assign new_n998_ = ~\A[16]  & new_n997_;
  assign new_n999_ = new_n994_ & ~new_n998_;
  assign new_n1000_ = ~new_n987_ & new_n998_;
  assign new_n1001_ = ~new_n999_ & ~new_n1000_;
  assign new_n1002_ = ~\A[11]  & new_n896_;
  assign new_n1003_ = ~\A[10]  & new_n1002_;
  assign new_n1004_ = ~\A[9]  & new_n1003_;
  assign new_n1005_ = ~\A[8]  & new_n1004_;
  assign new_n1006_ = new_n1001_ & ~new_n1005_;
  assign new_n1007_ = ~new_n994_ & new_n1005_;
  assign \P[3]  = new_n1006_ | new_n1007_;
  assign new_n1009_ = new_n910_ & new_n913_;
  assign new_n1010_ = ~\A[99]  & new_n786_;
  assign new_n1011_ = ~\A[98]  & new_n917_;
  assign new_n1012_ = ~\A[97]  & new_n1011_;
  assign new_n1013_ = ~\A[96]  & new_n1012_;
  assign new_n1014_ = new_n1010_ & new_n1013_;
  assign new_n1015_ = ~\A[87]  & new_n935_;
  assign new_n1016_ = ~\A[86]  & new_n1015_;
  assign new_n1017_ = ~\A[85]  & new_n1016_;
  assign new_n1018_ = ~\A[84]  & new_n1017_;
  assign new_n1019_ = ~\A[83]  & new_n1018_;
  assign new_n1020_ = ~\A[82]  & new_n1019_;
  assign new_n1021_ = ~\A[81]  & new_n1020_;
  assign new_n1022_ = ~\A[80]  & new_n1021_;
  assign new_n1023_ = new_n1014_ & ~new_n1022_;
  assign new_n1024_ = new_n1009_ & ~new_n1023_;
  assign new_n1025_ = ~\A[77]  & ~\A[78] ;
  assign new_n1026_ = ~\A[76]  & new_n1025_;
  assign new_n1027_ = ~\A[75]  & new_n1026_;
  assign new_n1028_ = ~\A[74]  & new_n1027_;
  assign new_n1029_ = ~\A[73]  & new_n1028_;
  assign new_n1030_ = ~\A[72]  & new_n1029_;
  assign new_n1031_ = ~\A[71]  & new_n1030_;
  assign new_n1032_ = ~\A[70]  & new_n1031_;
  assign new_n1033_ = ~\A[69]  & new_n1032_;
  assign new_n1034_ = ~\A[68]  & new_n1033_;
  assign new_n1035_ = ~\A[67]  & new_n1034_;
  assign new_n1036_ = ~\A[66]  & new_n1035_;
  assign new_n1037_ = ~\A[65]  & new_n1036_;
  assign new_n1038_ = ~\A[64]  & new_n1037_;
  assign new_n1039_ = new_n1024_ & ~new_n1038_;
  assign new_n1040_ = \A[79]  & new_n1022_;
  assign new_n1041_ = new_n1014_ & ~new_n1040_;
  assign new_n1042_ = new_n1009_ & ~new_n1041_;
  assign new_n1043_ = new_n1038_ & new_n1042_;
  assign new_n1044_ = ~new_n1039_ & ~new_n1043_;
  assign new_n1045_ = ~\A[55]  & new_n963_;
  assign new_n1046_ = ~\A[54]  & new_n1045_;
  assign new_n1047_ = ~\A[53]  & new_n1046_;
  assign new_n1048_ = ~\A[52]  & new_n1047_;
  assign new_n1049_ = ~\A[51]  & new_n1048_;
  assign new_n1050_ = ~\A[50]  & new_n1049_;
  assign new_n1051_ = ~\A[49]  & new_n1050_;
  assign new_n1052_ = ~\A[48]  & new_n1051_;
  assign new_n1053_ = new_n1044_ & ~new_n1052_;
  assign new_n1054_ = ~new_n1024_ & new_n1052_;
  assign new_n1055_ = ~new_n1053_ & ~new_n1054_;
  assign new_n1056_ = ~\A[39]  & new_n977_;
  assign new_n1057_ = ~\A[38]  & new_n1056_;
  assign new_n1058_ = ~\A[37]  & new_n1057_;
  assign new_n1059_ = ~\A[36]  & new_n1058_;
  assign new_n1060_ = ~\A[35]  & new_n1059_;
  assign new_n1061_ = ~\A[34]  & new_n1060_;
  assign new_n1062_ = ~\A[33]  & new_n1061_;
  assign new_n1063_ = ~\A[32]  & new_n1062_;
  assign new_n1064_ = new_n1055_ & ~new_n1063_;
  assign new_n1065_ = ~new_n1044_ & new_n1063_;
  assign new_n1066_ = ~new_n1064_ & ~new_n1065_;
  assign new_n1067_ = ~\A[23]  & new_n991_;
  assign new_n1068_ = ~\A[22]  & new_n1067_;
  assign new_n1069_ = ~\A[21]  & new_n1068_;
  assign new_n1070_ = ~\A[20]  & new_n1069_;
  assign new_n1071_ = ~\A[19]  & new_n1070_;
  assign new_n1072_ = ~\A[18]  & new_n1071_;
  assign new_n1073_ = ~\A[17]  & new_n1072_;
  assign new_n1074_ = ~\A[16]  & new_n1073_;
  assign new_n1075_ = new_n1066_ & ~new_n1074_;
  assign new_n1076_ = ~new_n1055_ & new_n1074_;
  assign \P[4]  = new_n1075_ | new_n1076_;
  assign new_n1078_ = new_n1009_ & new_n1014_;
  assign new_n1079_ = ~\A[71]  & new_n949_;
  assign new_n1080_ = ~\A[70]  & new_n1022_;
  assign new_n1081_ = ~\A[69]  & new_n1080_;
  assign new_n1082_ = ~\A[68]  & new_n1081_;
  assign new_n1083_ = ~\A[67]  & new_n1082_;
  assign new_n1084_ = ~\A[66]  & new_n1083_;
  assign new_n1085_ = ~\A[65]  & new_n1084_;
  assign new_n1086_ = ~\A[64]  & new_n1085_;
  assign new_n1087_ = new_n1079_ & new_n1086_;
  assign new_n1088_ = ~\A[47]  & new_n1052_;
  assign new_n1089_ = ~\A[46]  & new_n1088_;
  assign new_n1090_ = ~\A[45]  & new_n1089_;
  assign new_n1091_ = ~\A[44]  & new_n1090_;
  assign new_n1092_ = ~\A[43]  & new_n1091_;
  assign new_n1093_ = ~\A[42]  & new_n1092_;
  assign new_n1094_ = ~\A[41]  & new_n1093_;
  assign new_n1095_ = ~\A[40]  & new_n1094_;
  assign new_n1096_ = ~\A[39]  & new_n1095_;
  assign new_n1097_ = ~\A[38]  & new_n1096_;
  assign new_n1098_ = ~\A[37]  & new_n1097_;
  assign new_n1099_ = ~\A[36]  & new_n1098_;
  assign new_n1100_ = ~\A[35]  & new_n1099_;
  assign new_n1101_ = ~\A[34]  & new_n1100_;
  assign new_n1102_ = ~\A[33]  & new_n1101_;
  assign new_n1103_ = ~\A[32]  & new_n1102_;
  assign new_n1104_ = new_n1087_ & ~new_n1103_;
  assign \P[5]  = ~new_n1078_ | new_n1104_;
  assign \P[6]  = ~new_n1078_ | ~new_n1087_;
  assign new_n1107_ = ~\A[0]  & ~\P[6] ;
  assign new_n1108_ = new_n1005_ & new_n1107_;
  assign new_n1109_ = ~\A[3]  & new_n1108_;
  assign new_n1110_ = ~\A[2]  & new_n1109_;
  assign new_n1111_ = new_n1074_ & new_n1103_;
  assign new_n1112_ = new_n906_ & new_n1111_;
  assign new_n1113_ = ~\A[1]  & new_n1112_;
  assign F = ~new_n1110_ | ~new_n1113_;
endmodule


