module top ( 
    pv28_20_, pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv120_16_, pv120_29_,
    pv168_9_, pv180_10_, pv28_10_, pv56_13_, pv56_22_, pv88_7_, pv88_29_,
    pv120_15_, pv180_4_, pv56_14_, pv56_25_, pv88_8_, pv88_17_, pv88_28_,
    pv120_18_, pv180_5_, pv180_12_, pv192_0_, pv56_15_, pv56_24_, pv88_9_,
    pv88_18_, pv88_27_, pv120_17_, pv168_8_, pv180_6_, pv88_2_, pv88_15_,
    pv88_26_, pv120_12_, pv88_3_, pv88_16_, pv88_25_, pv120_11_, pv180_0_,
    pv56_10_, pv56_21_, pv88_4_, pv88_13_, pv88_24_, pv120_14_, pv126_5_,
    pv180_1_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_, pv120_13_,
    pv180_2_, pv28_8_, pv56_5_, pv88_11_, pv88_22_, pv120_5_, pv132_0_,
    pv156_6_, pv168_1_, pv189_0_, pv28_9_, pv56_4_, pv88_12_, pv88_21_,
    pv120_6_, pv156_5_, pv156_10_, pv168_2_, pv189_1_, pv28_6_, pv56_7_,
    pv88_20_, pv120_3_, pv120_10_, pv156_8_, pv189_2_, pv28_7_, pv56_6_,
    pv88_10_, pv120_4_, pv168_0_, pv28_4_, pv56_9_, pv120_1_, pv168_5_,
    pv28_5_, pv56_8_, pv120_2_, pv156_9_, pv156_14_, pv168_6_, pv28_2_,
    pv156_13_, pv28_3_, pv120_0_, pv156_12_, pv168_4_, pv28_0_, pv186_1_,
    pv28_1_, pv144_4_, pv186_2_, pv144_5_, pv156_0_, pv132_5_, pv144_6_,
    pv56_1_, pv120_9_, pv120_30_, pv132_4_, pv156_2_, pv56_0_, pv88_30_,
    pv132_3_, pv144_8_, pv156_1_, pv28_19_, pv56_3_, pv88_31_, pv120_7_,
    pv132_2_, pv144_9_, pv156_4_, pv56_2_, pv120_8_, pv120_20_, pv132_1_,
    pv186_0_, pv28_17_, pv120_21_, pv126_3_, pv144_10_, pv168_12_,
    pv183_2_, pv28_18_, pv28_27_, pv120_22_, pv126_4_, pv28_15_, pv28_26_,
    pv88_0_, pv120_23_, pv126_1_, pv144_12_, pv168_14_, pv28_16_, pv28_25_,
    pv88_1_, pv120_24_, pv120_31_, pv126_2_, pv168_13_, pv28_13_, pv28_24_,
    pv56_16_, pv56_27_, pv120_25_, pv144_14_, pv180_14_, pv192_2_,
    pv28_14_, pv28_23_, pv56_17_, pv56_26_, pv120_19_, pv120_26_, pv126_0_,
    pv144_0_, pv144_13_, pv180_8_, pv180_13_, pv192_1_, pv28_11_, pv28_22_,
    pv56_18_, pv120_27_, pv144_1_, pv168_10_, pv180_9_, pv183_0_, pv28_12_,
    pv28_21_, pv56_19_, pv120_28_, pv144_2_, pv183_1_,
    pv198_3_, pv198_0_, pv198_2_, pv198_1_, pv194_0_, pv194_1_  );
  input  pv28_20_, pv56_12_, pv56_23_, pv88_6_, pv88_19_, pv120_16_,
    pv120_29_, pv168_9_, pv180_10_, pv28_10_, pv56_13_, pv56_22_, pv88_7_,
    pv88_29_, pv120_15_, pv180_4_, pv56_14_, pv56_25_, pv88_8_, pv88_17_,
    pv88_28_, pv120_18_, pv180_5_, pv180_12_, pv192_0_, pv56_15_, pv56_24_,
    pv88_9_, pv88_18_, pv88_27_, pv120_17_, pv168_8_, pv180_6_, pv88_2_,
    pv88_15_, pv88_26_, pv120_12_, pv88_3_, pv88_16_, pv88_25_, pv120_11_,
    pv180_0_, pv56_10_, pv56_21_, pv88_4_, pv88_13_, pv88_24_, pv120_14_,
    pv126_5_, pv180_1_, pv56_11_, pv56_20_, pv88_5_, pv88_14_, pv88_23_,
    pv120_13_, pv180_2_, pv28_8_, pv56_5_, pv88_11_, pv88_22_, pv120_5_,
    pv132_0_, pv156_6_, pv168_1_, pv189_0_, pv28_9_, pv56_4_, pv88_12_,
    pv88_21_, pv120_6_, pv156_5_, pv156_10_, pv168_2_, pv189_1_, pv28_6_,
    pv56_7_, pv88_20_, pv120_3_, pv120_10_, pv156_8_, pv189_2_, pv28_7_,
    pv56_6_, pv88_10_, pv120_4_, pv168_0_, pv28_4_, pv56_9_, pv120_1_,
    pv168_5_, pv28_5_, pv56_8_, pv120_2_, pv156_9_, pv156_14_, pv168_6_,
    pv28_2_, pv156_13_, pv28_3_, pv120_0_, pv156_12_, pv168_4_, pv28_0_,
    pv186_1_, pv28_1_, pv144_4_, pv186_2_, pv144_5_, pv156_0_, pv132_5_,
    pv144_6_, pv56_1_, pv120_9_, pv120_30_, pv132_4_, pv156_2_, pv56_0_,
    pv88_30_, pv132_3_, pv144_8_, pv156_1_, pv28_19_, pv56_3_, pv88_31_,
    pv120_7_, pv132_2_, pv144_9_, pv156_4_, pv56_2_, pv120_8_, pv120_20_,
    pv132_1_, pv186_0_, pv28_17_, pv120_21_, pv126_3_, pv144_10_,
    pv168_12_, pv183_2_, pv28_18_, pv28_27_, pv120_22_, pv126_4_, pv28_15_,
    pv28_26_, pv88_0_, pv120_23_, pv126_1_, pv144_12_, pv168_14_, pv28_16_,
    pv28_25_, pv88_1_, pv120_24_, pv120_31_, pv126_2_, pv168_13_, pv28_13_,
    pv28_24_, pv56_16_, pv56_27_, pv120_25_, pv144_14_, pv180_14_,
    pv192_2_, pv28_14_, pv28_23_, pv56_17_, pv56_26_, pv120_19_, pv120_26_,
    pv126_0_, pv144_0_, pv144_13_, pv180_8_, pv180_13_, pv192_1_, pv28_11_,
    pv28_22_, pv56_18_, pv120_27_, pv144_1_, pv168_10_, pv180_9_, pv183_0_,
    pv28_12_, pv28_21_, pv56_19_, pv120_28_, pv144_2_, pv183_1_;
  output pv198_3_, pv198_0_, pv198_2_, pv198_1_, pv194_0_, pv194_1_;
  wire new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_;
  assign new_n199_ = pv88_22_ & pv120_22_;
  assign new_n200_ = pv180_0_ & pv120_24_;
  assign new_n201_ = pv88_24_ & new_n200_;
  assign new_n202_ = pv180_1_ & new_n201_;
  assign new_n203_ = pv180_1_ & pv120_25_;
  assign new_n204_ = pv180_0_ & new_n203_;
  assign new_n205_ = pv88_25_ & new_n204_;
  assign new_n206_ = pv180_2_ & new_n205_;
  assign new_n207_ = pv88_23_ & pv120_23_;
  assign new_n208_ = pv180_0_ & new_n207_;
  assign new_n209_ = pv132_1_ & pv180_9_;
  assign new_n210_ = pv180_8_ & new_n209_;
  assign new_n211_ = pv126_1_ & new_n210_;
  assign new_n212_ = pv180_10_ & new_n211_;
  assign new_n213_ = pv120_30_ & pv88_30_;
  assign new_n214_ = pv88_31_ & pv120_31_;
  assign new_n215_ = pv180_8_ & new_n214_;
  assign new_n216_ = pv132_0_ & pv180_8_;
  assign new_n217_ = pv126_0_ & new_n216_;
  assign new_n218_ = pv180_9_ & new_n217_;
  assign new_n219_ = ~new_n215_ & ~new_n218_;
  assign new_n220_ = ~new_n212_ & ~new_n213_;
  assign new_n221_ = new_n219_ & new_n220_;
  assign new_n222_ = pv192_0_ & ~new_n221_;
  assign new_n223_ = pv192_1_ & new_n222_;
  assign new_n224_ = pv120_29_ & pv180_5_;
  assign new_n225_ = pv180_4_ & new_n224_;
  assign new_n226_ = pv88_29_ & new_n225_;
  assign new_n227_ = pv180_6_ & new_n226_;
  assign new_n228_ = pv88_26_ & pv120_26_;
  assign new_n229_ = pv88_27_ & pv120_27_;
  assign new_n230_ = pv180_4_ & new_n229_;
  assign new_n231_ = pv180_4_ & pv120_28_;
  assign new_n232_ = pv88_28_ & new_n231_;
  assign new_n233_ = pv180_5_ & new_n232_;
  assign new_n234_ = ~new_n230_ & ~new_n233_;
  assign new_n235_ = ~new_n227_ & ~new_n228_;
  assign new_n236_ = new_n234_ & new_n235_;
  assign new_n237_ = pv192_0_ & ~new_n236_;
  assign new_n238_ = pv132_5_ & pv180_13_;
  assign new_n239_ = pv180_12_ & new_n238_;
  assign new_n240_ = pv126_5_ & new_n239_;
  assign new_n241_ = pv180_14_ & new_n240_;
  assign new_n242_ = pv132_2_ & pv126_2_;
  assign new_n243_ = pv132_3_ & pv126_3_;
  assign new_n244_ = pv180_12_ & new_n243_;
  assign new_n245_ = pv180_12_ & pv132_4_;
  assign new_n246_ = pv126_4_ & new_n245_;
  assign new_n247_ = pv180_13_ & new_n246_;
  assign new_n248_ = ~new_n244_ & ~new_n247_;
  assign new_n249_ = ~new_n241_ & ~new_n242_;
  assign new_n250_ = new_n248_ & new_n249_;
  assign new_n251_ = pv192_0_ & pv192_1_;
  assign new_n252_ = ~new_n250_ & new_n251_;
  assign new_n253_ = pv192_2_ & new_n252_;
  assign new_n254_ = ~new_n223_ & ~new_n237_;
  assign new_n255_ = ~new_n253_ & new_n254_;
  assign new_n256_ = ~new_n206_ & ~new_n208_;
  assign new_n257_ = ~new_n199_ & ~new_n202_;
  assign new_n258_ = new_n256_ & new_n257_;
  assign pv198_3_ = ~new_n255_ | ~new_n258_;
  assign new_n260_ = pv28_2_ & pv56_2_;
  assign new_n261_ = pv56_4_ & pv144_0_;
  assign new_n262_ = pv28_4_ & new_n261_;
  assign new_n263_ = pv144_1_ & new_n262_;
  assign new_n264_ = pv56_5_ & pv144_1_;
  assign new_n265_ = pv144_0_ & new_n264_;
  assign new_n266_ = pv28_5_ & new_n265_;
  assign new_n267_ = pv144_2_ & new_n266_;
  assign new_n268_ = pv28_3_ & pv56_3_;
  assign new_n269_ = pv144_0_ & new_n268_;
  assign new_n270_ = pv56_13_ & pv144_9_;
  assign new_n271_ = pv144_8_ & new_n270_;
  assign new_n272_ = pv28_13_ & new_n271_;
  assign new_n273_ = pv144_10_ & new_n272_;
  assign new_n274_ = pv28_10_ & pv56_10_;
  assign new_n275_ = pv56_11_ & pv28_11_;
  assign new_n276_ = pv144_8_ & new_n275_;
  assign new_n277_ = pv56_12_ & pv144_8_;
  assign new_n278_ = pv28_12_ & new_n277_;
  assign new_n279_ = pv144_9_ & new_n278_;
  assign new_n280_ = ~new_n276_ & ~new_n279_;
  assign new_n281_ = ~new_n273_ & ~new_n274_;
  assign new_n282_ = new_n280_ & new_n281_;
  assign new_n283_ = pv183_0_ & ~new_n282_;
  assign new_n284_ = pv183_1_ & new_n283_;
  assign new_n285_ = pv56_9_ & pv144_5_;
  assign new_n286_ = pv144_4_ & new_n285_;
  assign new_n287_ = pv28_9_ & new_n286_;
  assign new_n288_ = pv144_6_ & new_n287_;
  assign new_n289_ = pv28_6_ & pv56_6_;
  assign new_n290_ = pv56_7_ & pv28_7_;
  assign new_n291_ = pv144_4_ & new_n290_;
  assign new_n292_ = pv56_8_ & pv144_4_;
  assign new_n293_ = pv28_8_ & new_n292_;
  assign new_n294_ = pv144_5_ & new_n293_;
  assign new_n295_ = ~new_n291_ & ~new_n294_;
  assign new_n296_ = ~new_n288_ & ~new_n289_;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = pv183_0_ & ~new_n297_;
  assign new_n299_ = pv56_17_ & pv144_13_;
  assign new_n300_ = pv144_12_ & new_n299_;
  assign new_n301_ = pv28_17_ & new_n300_;
  assign new_n302_ = pv144_14_ & new_n301_;
  assign new_n303_ = pv56_14_ & pv28_14_;
  assign new_n304_ = pv56_15_ & pv28_15_;
  assign new_n305_ = pv144_12_ & new_n304_;
  assign new_n306_ = pv144_12_ & pv56_16_;
  assign new_n307_ = pv28_16_ & new_n306_;
  assign new_n308_ = pv144_13_ & new_n307_;
  assign new_n309_ = ~new_n305_ & ~new_n308_;
  assign new_n310_ = ~new_n302_ & ~new_n303_;
  assign new_n311_ = new_n309_ & new_n310_;
  assign new_n312_ = pv183_0_ & pv183_1_;
  assign new_n313_ = ~new_n311_ & new_n312_;
  assign new_n314_ = pv183_2_ & new_n313_;
  assign new_n315_ = ~new_n284_ & ~new_n298_;
  assign new_n316_ = ~new_n314_ & new_n315_;
  assign new_n317_ = ~new_n267_ & ~new_n269_;
  assign new_n318_ = ~new_n260_ & ~new_n263_;
  assign new_n319_ = new_n317_ & new_n318_;
  assign pv198_0_ = ~new_n316_ | ~new_n319_;
  assign new_n321_ = pv88_6_ & pv120_6_;
  assign new_n322_ = pv168_0_ & pv120_8_;
  assign new_n323_ = pv88_8_ & new_n322_;
  assign new_n324_ = pv168_1_ & new_n323_;
  assign new_n325_ = pv168_1_ & pv120_9_;
  assign new_n326_ = pv168_0_ & new_n325_;
  assign new_n327_ = pv88_9_ & new_n326_;
  assign new_n328_ = pv168_2_ & new_n327_;
  assign new_n329_ = pv88_7_ & pv120_7_;
  assign new_n330_ = pv168_0_ & new_n329_;
  assign new_n331_ = pv168_9_ & pv120_17_;
  assign new_n332_ = pv168_8_ & new_n331_;
  assign new_n333_ = pv88_17_ & new_n332_;
  assign new_n334_ = pv168_10_ & new_n333_;
  assign new_n335_ = pv120_14_ & pv88_14_;
  assign new_n336_ = pv120_15_ & pv88_15_;
  assign new_n337_ = pv168_8_ & new_n336_;
  assign new_n338_ = pv120_16_ & pv168_8_;
  assign new_n339_ = pv88_16_ & new_n338_;
  assign new_n340_ = pv168_9_ & new_n339_;
  assign new_n341_ = ~new_n337_ & ~new_n340_;
  assign new_n342_ = ~new_n334_ & ~new_n335_;
  assign new_n343_ = new_n341_ & new_n342_;
  assign new_n344_ = pv189_0_ & ~new_n343_;
  assign new_n345_ = pv189_1_ & new_n344_;
  assign new_n346_ = pv120_13_ & pv168_5_;
  assign new_n347_ = pv168_4_ & new_n346_;
  assign new_n348_ = pv88_13_ & new_n347_;
  assign new_n349_ = pv168_6_ & new_n348_;
  assign new_n350_ = pv120_10_ & pv88_10_;
  assign new_n351_ = pv120_11_ & pv88_11_;
  assign new_n352_ = pv168_4_ & new_n351_;
  assign new_n353_ = pv120_12_ & pv168_4_;
  assign new_n354_ = pv88_12_ & new_n353_;
  assign new_n355_ = pv168_5_ & new_n354_;
  assign new_n356_ = ~new_n352_ & ~new_n355_;
  assign new_n357_ = ~new_n349_ & ~new_n350_;
  assign new_n358_ = new_n356_ & new_n357_;
  assign new_n359_ = pv189_0_ & ~new_n358_;
  assign new_n360_ = pv120_21_ & pv168_13_;
  assign new_n361_ = pv168_12_ & new_n360_;
  assign new_n362_ = pv88_21_ & new_n361_;
  assign new_n363_ = pv168_14_ & new_n362_;
  assign new_n364_ = pv120_18_ & pv88_18_;
  assign new_n365_ = pv88_19_ & pv120_19_;
  assign new_n366_ = pv168_12_ & new_n365_;
  assign new_n367_ = pv120_20_ & pv168_12_;
  assign new_n368_ = pv88_20_ & new_n367_;
  assign new_n369_ = pv168_13_ & new_n368_;
  assign new_n370_ = ~new_n366_ & ~new_n369_;
  assign new_n371_ = ~new_n363_ & ~new_n364_;
  assign new_n372_ = new_n370_ & new_n371_;
  assign new_n373_ = pv189_0_ & pv189_1_;
  assign new_n374_ = ~new_n372_ & new_n373_;
  assign new_n375_ = pv189_2_ & new_n374_;
  assign new_n376_ = ~new_n345_ & ~new_n359_;
  assign new_n377_ = ~new_n375_ & new_n376_;
  assign new_n378_ = ~new_n328_ & ~new_n330_;
  assign new_n379_ = ~new_n321_ & ~new_n324_;
  assign new_n380_ = new_n378_ & new_n379_;
  assign pv198_2_ = ~new_n377_ | ~new_n380_;
  assign new_n382_ = pv28_18_ & pv56_18_;
  assign new_n383_ = pv56_20_ & pv156_0_;
  assign new_n384_ = pv28_20_ & new_n383_;
  assign new_n385_ = pv156_1_ & new_n384_;
  assign new_n386_ = pv56_21_ & pv156_1_;
  assign new_n387_ = pv156_0_ & new_n386_;
  assign new_n388_ = pv28_21_ & new_n387_;
  assign new_n389_ = pv156_2_ & new_n388_;
  assign new_n390_ = pv28_19_ & pv56_19_;
  assign new_n391_ = pv156_0_ & new_n390_;
  assign new_n392_ = pv120_1_ & pv156_9_;
  assign new_n393_ = pv156_8_ & new_n392_;
  assign new_n394_ = pv88_1_ & new_n393_;
  assign new_n395_ = pv156_10_ & new_n394_;
  assign new_n396_ = pv28_26_ & pv56_26_;
  assign new_n397_ = pv28_27_ & pv56_27_;
  assign new_n398_ = pv156_8_ & new_n397_;
  assign new_n399_ = pv156_8_ & pv120_0_;
  assign new_n400_ = pv88_0_ & new_n399_;
  assign new_n401_ = pv156_9_ & new_n400_;
  assign new_n402_ = ~new_n398_ & ~new_n401_;
  assign new_n403_ = ~new_n395_ & ~new_n396_;
  assign new_n404_ = new_n402_ & new_n403_;
  assign new_n405_ = pv186_0_ & ~new_n404_;
  assign new_n406_ = pv186_1_ & new_n405_;
  assign new_n407_ = pv56_25_ & pv156_5_;
  assign new_n408_ = pv156_4_ & new_n407_;
  assign new_n409_ = pv28_25_ & new_n408_;
  assign new_n410_ = pv156_6_ & new_n409_;
  assign new_n411_ = pv56_22_ & pv28_22_;
  assign new_n412_ = pv56_23_ & pv28_23_;
  assign new_n413_ = pv156_4_ & new_n412_;
  assign new_n414_ = pv56_24_ & pv156_4_;
  assign new_n415_ = pv28_24_ & new_n414_;
  assign new_n416_ = pv156_5_ & new_n415_;
  assign new_n417_ = ~new_n413_ & ~new_n416_;
  assign new_n418_ = ~new_n410_ & ~new_n411_;
  assign new_n419_ = new_n417_ & new_n418_;
  assign new_n420_ = pv186_0_ & ~new_n419_;
  assign new_n421_ = pv120_5_ & pv156_13_;
  assign new_n422_ = pv156_12_ & new_n421_;
  assign new_n423_ = pv88_5_ & new_n422_;
  assign new_n424_ = pv156_14_ & new_n423_;
  assign new_n425_ = pv88_2_ & pv120_2_;
  assign new_n426_ = pv88_3_ & pv120_3_;
  assign new_n427_ = pv156_12_ & new_n426_;
  assign new_n428_ = pv120_4_ & pv156_12_;
  assign new_n429_ = pv88_4_ & new_n428_;
  assign new_n430_ = pv156_13_ & new_n429_;
  assign new_n431_ = ~new_n427_ & ~new_n430_;
  assign new_n432_ = ~new_n424_ & ~new_n425_;
  assign new_n433_ = new_n431_ & new_n432_;
  assign new_n434_ = pv186_1_ & pv186_0_;
  assign new_n435_ = ~new_n433_ & new_n434_;
  assign new_n436_ = pv186_2_ & new_n435_;
  assign new_n437_ = ~new_n406_ & ~new_n420_;
  assign new_n438_ = ~new_n436_ & new_n437_;
  assign new_n439_ = ~new_n389_ & ~new_n391_;
  assign new_n440_ = ~new_n382_ & ~new_n385_;
  assign new_n441_ = new_n439_ & new_n440_;
  assign pv198_1_ = ~new_n438_ | ~new_n441_;
  assign pv194_0_ = pv28_0_ & pv56_0_;
  assign pv194_1_ = pv28_1_ & pv56_1_;
endmodule

