module i6 ( 
    \V138(0) , \V138(2) , \V32(27) , \V32(26) , \V32(25) , \V32(24) ,
    \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) ,
    \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) ,
    \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) ,
    \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V64(27) , \V64(26) ,
    \V64(25) , \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) ,
    \V64(19) , \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) ,
    \V64(13) , \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) ,
    \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) ,
    \V64(0) , \V96(27) , \V138(4) , \V96(26) , \V96(25) , \V96(24) ,
    \V96(23) , \V96(22) , \V96(21) , \V96(20) , \V96(19) , \V96(18) ,
    \V96(17) , \V96(16) , \V96(15) , \V96(14) , \V96(13) , \V96(12) ,
    \V96(11) , \V96(10) , \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) ,
    \V96(4) , \V96(3) , \V96(2) , \V96(1) , \V96(0) , \V32(31) , \V32(30) ,
    \V32(29) , \V32(28) , \V131(27) , \V131(26) , \V131(25) , \V131(24) ,
    \V131(23) , \V131(22) , \V131(21) , \V131(20) , \V131(19) , \V131(18) ,
    \V131(17) , \V131(16) , \V131(15) , \V131(14) , \V131(13) , \V131(12) ,
    \V131(11) , \V131(10) , \V131(9) , \V131(8) , \V131(7) , \V131(6) ,
    \V131(5) , \V131(4) , \V131(3) , \V131(2) , \V131(1) , \V131(0) ,
    \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V99(0) , \V138(3) ,
    \V98(0) , \V97(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) ,
    \V134(0) , \V133(1) , \V133(0) , \V131(31) , \V131(30) , \V131(29) ,
    \V131(28) ,
    \V166(27) , \V166(26) , \V166(25) , \V166(24) , \V166(23) , \V166(22) ,
    \V166(21) , \V166(20) , \V166(19) , \V166(18) , \V166(17) , \V166(16) ,
    \V166(15) , \V166(14) , \V166(13) , \V166(12) , \V166(11) , \V166(10) ,
    \V166(9) , \V166(8) , \V166(7) , \V166(6) , \V166(5) , \V166(4) ,
    \V166(3) , \V166(2) , \V166(1) , \V166(0) , \V198(31) , \V198(30) ,
    \V198(29) , \V198(28) , \V198(27) , \V198(26) , \V198(25) , \V198(24) ,
    \V198(23) , \V198(22) , \V198(21) , \V198(20) , \V198(19) , \V198(18) ,
    \V198(17) , \V198(16) , \V198(15) , \V198(14) , \V198(13) , \V198(12) ,
    \V198(11) , \V198(10) , \V198(9) , \V198(8) , \V198(7) , \V198(6) ,
    \V198(5) , \V198(4) , \V198(3) , \V198(2) , \V198(1) , \V198(0) ,
    \V205(6) , \V205(5) , \V205(4) , \V205(3) , \V205(2) , \V205(1) ,
    \V205(0)   );
  input  \V138(0) , \V138(2) , \V32(27) , \V32(26) , \V32(25) ,
    \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) ,
    \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) ,
    \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) ,
    \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) ,
    \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) , \V64(22) ,
    \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) , \V64(16) ,
    \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) , \V64(10) ,
    \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) ,
    \V64(2) , \V64(1) , \V64(0) , \V96(27) , \V138(4) , \V96(26) ,
    \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) ,
    \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) ,
    \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) ,
    \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) ,
    \V96(0) , \V32(31) , \V32(30) , \V32(29) , \V32(28) , \V131(27) ,
    \V131(26) , \V131(25) , \V131(24) , \V131(23) , \V131(22) , \V131(21) ,
    \V131(20) , \V131(19) , \V131(18) , \V131(17) , \V131(16) , \V131(15) ,
    \V131(14) , \V131(13) , \V131(12) , \V131(11) , \V131(10) , \V131(9) ,
    \V131(8) , \V131(7) , \V131(6) , \V131(5) , \V131(4) , \V131(3) ,
    \V131(2) , \V131(1) , \V131(0) , \V64(31) , \V64(30) , \V64(29) ,
    \V64(28) , \V99(0) , \V138(3) , \V98(0) , \V97(0) , \V96(31) ,
    \V96(30) , \V96(29) , \V96(28) , \V134(0) , \V133(1) , \V133(0) ,
    \V131(31) , \V131(30) , \V131(29) , \V131(28) ;
  output \V166(27) , \V166(26) , \V166(25) , \V166(24) , \V166(23) ,
    \V166(22) , \V166(21) , \V166(20) , \V166(19) , \V166(18) , \V166(17) ,
    \V166(16) , \V166(15) , \V166(14) , \V166(13) , \V166(12) , \V166(11) ,
    \V166(10) , \V166(9) , \V166(8) , \V166(7) , \V166(6) , \V166(5) ,
    \V166(4) , \V166(3) , \V166(2) , \V166(1) , \V166(0) , \V198(31) ,
    \V198(30) , \V198(29) , \V198(28) , \V198(27) , \V198(26) , \V198(25) ,
    \V198(24) , \V198(23) , \V198(22) , \V198(21) , \V198(20) , \V198(19) ,
    \V198(18) , \V198(17) , \V198(16) , \V198(15) , \V198(14) , \V198(13) ,
    \V198(12) , \V198(11) , \V198(10) , \V198(9) , \V198(8) , \V198(7) ,
    \V198(6) , \V198(5) , \V198(4) , \V198(3) , \V198(2) , \V198(1) ,
    \V198(0) , \V205(6) , \V205(5) , \V205(4) , \V205(3) , \V205(2) ,
    \V205(1) , \V205(0) ;
  wire new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_;
  assign new_n206_ = ~\V138(2)  & \V32(27) ;
  assign new_n207_ = ~\V138(0)  & new_n206_;
  assign new_n208_ = ~\V138(2)  & \V64(27) ;
  assign new_n209_ = \V138(0)  & new_n208_;
  assign new_n210_ = \V138(2)  & ~\V64(27) ;
  assign new_n211_ = \V138(0)  & new_n210_;
  assign new_n212_ = ~new_n207_ & ~new_n209_;
  assign \V166(27)  = new_n211_ | ~new_n212_;
  assign new_n214_ = ~\V138(2)  & \V32(26) ;
  assign new_n215_ = ~\V138(0)  & new_n214_;
  assign new_n216_ = ~\V138(2)  & \V64(26) ;
  assign new_n217_ = \V138(0)  & new_n216_;
  assign new_n218_ = \V138(2)  & ~\V64(26) ;
  assign new_n219_ = \V138(0)  & new_n218_;
  assign new_n220_ = ~new_n215_ & ~new_n217_;
  assign \V166(26)  = new_n219_ | ~new_n220_;
  assign new_n222_ = ~\V138(2)  & \V32(25) ;
  assign new_n223_ = ~\V138(0)  & new_n222_;
  assign new_n224_ = ~\V138(2)  & \V64(25) ;
  assign new_n225_ = \V138(0)  & new_n224_;
  assign new_n226_ = \V138(2)  & ~\V64(25) ;
  assign new_n227_ = \V138(0)  & new_n226_;
  assign new_n228_ = ~new_n223_ & ~new_n225_;
  assign \V166(25)  = new_n227_ | ~new_n228_;
  assign new_n230_ = ~\V138(2)  & \V32(24) ;
  assign new_n231_ = ~\V138(0)  & new_n230_;
  assign new_n232_ = ~\V138(2)  & \V64(24) ;
  assign new_n233_ = \V138(0)  & new_n232_;
  assign new_n234_ = \V138(2)  & ~\V64(24) ;
  assign new_n235_ = \V138(0)  & new_n234_;
  assign new_n236_ = ~new_n231_ & ~new_n233_;
  assign \V166(24)  = new_n235_ | ~new_n236_;
  assign new_n238_ = ~\V138(2)  & \V32(23) ;
  assign new_n239_ = ~\V138(0)  & new_n238_;
  assign new_n240_ = ~\V138(2)  & \V64(23) ;
  assign new_n241_ = \V138(0)  & new_n240_;
  assign new_n242_ = \V138(2)  & ~\V64(23) ;
  assign new_n243_ = \V138(0)  & new_n242_;
  assign new_n244_ = ~new_n239_ & ~new_n241_;
  assign \V166(23)  = new_n243_ | ~new_n244_;
  assign new_n246_ = ~\V138(2)  & \V32(22) ;
  assign new_n247_ = ~\V138(0)  & new_n246_;
  assign new_n248_ = ~\V138(2)  & \V64(22) ;
  assign new_n249_ = \V138(0)  & new_n248_;
  assign new_n250_ = \V138(2)  & ~\V64(22) ;
  assign new_n251_ = \V138(0)  & new_n250_;
  assign new_n252_ = ~new_n247_ & ~new_n249_;
  assign \V166(22)  = new_n251_ | ~new_n252_;
  assign new_n254_ = ~\V138(2)  & \V32(21) ;
  assign new_n255_ = ~\V138(0)  & new_n254_;
  assign new_n256_ = ~\V138(2)  & \V64(21) ;
  assign new_n257_ = \V138(0)  & new_n256_;
  assign new_n258_ = \V138(2)  & ~\V64(21) ;
  assign new_n259_ = \V138(0)  & new_n258_;
  assign new_n260_ = ~new_n255_ & ~new_n257_;
  assign \V166(21)  = new_n259_ | ~new_n260_;
  assign new_n262_ = ~\V138(2)  & \V32(20) ;
  assign new_n263_ = ~\V138(0)  & new_n262_;
  assign new_n264_ = ~\V138(2)  & \V64(20) ;
  assign new_n265_ = \V138(0)  & new_n264_;
  assign new_n266_ = \V138(2)  & ~\V64(20) ;
  assign new_n267_ = \V138(0)  & new_n266_;
  assign new_n268_ = ~new_n263_ & ~new_n265_;
  assign \V166(20)  = new_n267_ | ~new_n268_;
  assign new_n270_ = ~\V138(2)  & \V32(19) ;
  assign new_n271_ = ~\V138(0)  & new_n270_;
  assign new_n272_ = ~\V138(2)  & \V64(19) ;
  assign new_n273_ = \V138(0)  & new_n272_;
  assign new_n274_ = \V138(2)  & ~\V64(19) ;
  assign new_n275_ = \V138(0)  & new_n274_;
  assign new_n276_ = ~new_n271_ & ~new_n273_;
  assign \V166(19)  = new_n275_ | ~new_n276_;
  assign new_n278_ = ~\V138(2)  & \V32(18) ;
  assign new_n279_ = ~\V138(0)  & new_n278_;
  assign new_n280_ = ~\V138(2)  & \V64(18) ;
  assign new_n281_ = \V138(0)  & new_n280_;
  assign new_n282_ = \V138(2)  & ~\V64(18) ;
  assign new_n283_ = \V138(0)  & new_n282_;
  assign new_n284_ = ~new_n279_ & ~new_n281_;
  assign \V166(18)  = new_n283_ | ~new_n284_;
  assign new_n286_ = ~\V138(2)  & \V32(17) ;
  assign new_n287_ = ~\V138(0)  & new_n286_;
  assign new_n288_ = ~\V138(2)  & \V64(17) ;
  assign new_n289_ = \V138(0)  & new_n288_;
  assign new_n290_ = \V138(2)  & ~\V64(17) ;
  assign new_n291_ = \V138(0)  & new_n290_;
  assign new_n292_ = ~new_n287_ & ~new_n289_;
  assign \V166(17)  = new_n291_ | ~new_n292_;
  assign new_n294_ = ~\V138(2)  & \V32(16) ;
  assign new_n295_ = ~\V138(0)  & new_n294_;
  assign new_n296_ = ~\V138(2)  & \V64(16) ;
  assign new_n297_ = \V138(0)  & new_n296_;
  assign new_n298_ = \V138(2)  & ~\V64(16) ;
  assign new_n299_ = \V138(0)  & new_n298_;
  assign new_n300_ = ~new_n295_ & ~new_n297_;
  assign \V166(16)  = new_n299_ | ~new_n300_;
  assign new_n302_ = ~\V138(2)  & \V32(15) ;
  assign new_n303_ = ~\V138(0)  & new_n302_;
  assign new_n304_ = ~\V138(2)  & \V64(15) ;
  assign new_n305_ = \V138(0)  & new_n304_;
  assign new_n306_ = \V138(2)  & ~\V64(15) ;
  assign new_n307_ = \V138(0)  & new_n306_;
  assign new_n308_ = ~new_n303_ & ~new_n305_;
  assign \V166(15)  = new_n307_ | ~new_n308_;
  assign new_n310_ = ~\V138(2)  & \V32(14) ;
  assign new_n311_ = ~\V138(0)  & new_n310_;
  assign new_n312_ = ~\V138(2)  & \V64(14) ;
  assign new_n313_ = \V138(0)  & new_n312_;
  assign new_n314_ = \V138(2)  & ~\V64(14) ;
  assign new_n315_ = \V138(0)  & new_n314_;
  assign new_n316_ = ~new_n311_ & ~new_n313_;
  assign \V166(14)  = new_n315_ | ~new_n316_;
  assign new_n318_ = ~\V138(2)  & \V32(13) ;
  assign new_n319_ = ~\V138(0)  & new_n318_;
  assign new_n320_ = ~\V138(2)  & \V64(13) ;
  assign new_n321_ = \V138(0)  & new_n320_;
  assign new_n322_ = \V138(2)  & ~\V64(13) ;
  assign new_n323_ = \V138(0)  & new_n322_;
  assign new_n324_ = ~new_n319_ & ~new_n321_;
  assign \V166(13)  = new_n323_ | ~new_n324_;
  assign new_n326_ = ~\V138(2)  & \V32(12) ;
  assign new_n327_ = ~\V138(0)  & new_n326_;
  assign new_n328_ = ~\V138(2)  & \V64(12) ;
  assign new_n329_ = \V138(0)  & new_n328_;
  assign new_n330_ = \V138(2)  & ~\V64(12) ;
  assign new_n331_ = \V138(0)  & new_n330_;
  assign new_n332_ = ~new_n327_ & ~new_n329_;
  assign \V166(12)  = new_n331_ | ~new_n332_;
  assign new_n334_ = ~\V138(2)  & \V32(11) ;
  assign new_n335_ = ~\V138(0)  & new_n334_;
  assign new_n336_ = ~\V138(2)  & \V64(11) ;
  assign new_n337_ = \V138(0)  & new_n336_;
  assign new_n338_ = \V138(2)  & ~\V64(11) ;
  assign new_n339_ = \V138(0)  & new_n338_;
  assign new_n340_ = ~new_n335_ & ~new_n337_;
  assign \V166(11)  = new_n339_ | ~new_n340_;
  assign new_n342_ = ~\V138(2)  & \V32(10) ;
  assign new_n343_ = ~\V138(0)  & new_n342_;
  assign new_n344_ = ~\V138(2)  & \V64(10) ;
  assign new_n345_ = \V138(0)  & new_n344_;
  assign new_n346_ = \V138(2)  & ~\V64(10) ;
  assign new_n347_ = \V138(0)  & new_n346_;
  assign new_n348_ = ~new_n343_ & ~new_n345_;
  assign \V166(10)  = new_n347_ | ~new_n348_;
  assign new_n350_ = ~\V138(2)  & \V32(9) ;
  assign new_n351_ = ~\V138(0)  & new_n350_;
  assign new_n352_ = ~\V138(2)  & \V64(9) ;
  assign new_n353_ = \V138(0)  & new_n352_;
  assign new_n354_ = \V138(2)  & ~\V64(9) ;
  assign new_n355_ = \V138(0)  & new_n354_;
  assign new_n356_ = ~new_n351_ & ~new_n353_;
  assign \V166(9)  = new_n355_ | ~new_n356_;
  assign new_n358_ = ~\V138(2)  & \V32(8) ;
  assign new_n359_ = ~\V138(0)  & new_n358_;
  assign new_n360_ = ~\V138(2)  & \V64(8) ;
  assign new_n361_ = \V138(0)  & new_n360_;
  assign new_n362_ = \V138(2)  & ~\V64(8) ;
  assign new_n363_ = \V138(0)  & new_n362_;
  assign new_n364_ = ~new_n359_ & ~new_n361_;
  assign \V166(8)  = new_n363_ | ~new_n364_;
  assign new_n366_ = ~\V138(2)  & \V32(7) ;
  assign new_n367_ = ~\V138(0)  & new_n366_;
  assign new_n368_ = ~\V138(2)  & \V64(7) ;
  assign new_n369_ = \V138(0)  & new_n368_;
  assign new_n370_ = \V138(2)  & ~\V64(7) ;
  assign new_n371_ = \V138(0)  & new_n370_;
  assign new_n372_ = ~new_n367_ & ~new_n369_;
  assign \V166(7)  = new_n371_ | ~new_n372_;
  assign new_n374_ = ~\V138(2)  & \V32(6) ;
  assign new_n375_ = ~\V138(0)  & new_n374_;
  assign new_n376_ = ~\V138(2)  & \V64(6) ;
  assign new_n377_ = \V138(0)  & new_n376_;
  assign new_n378_ = \V138(2)  & ~\V64(6) ;
  assign new_n379_ = \V138(0)  & new_n378_;
  assign new_n380_ = ~new_n375_ & ~new_n377_;
  assign \V166(6)  = new_n379_ | ~new_n380_;
  assign new_n382_ = ~\V138(2)  & \V32(5) ;
  assign new_n383_ = ~\V138(0)  & new_n382_;
  assign new_n384_ = ~\V138(2)  & \V64(5) ;
  assign new_n385_ = \V138(0)  & new_n384_;
  assign new_n386_ = \V138(2)  & ~\V64(5) ;
  assign new_n387_ = \V138(0)  & new_n386_;
  assign new_n388_ = ~new_n383_ & ~new_n385_;
  assign \V166(5)  = new_n387_ | ~new_n388_;
  assign new_n390_ = ~\V138(2)  & \V32(4) ;
  assign new_n391_ = ~\V138(0)  & new_n390_;
  assign new_n392_ = ~\V138(2)  & \V64(4) ;
  assign new_n393_ = \V138(0)  & new_n392_;
  assign new_n394_ = \V138(2)  & ~\V64(4) ;
  assign new_n395_ = \V138(0)  & new_n394_;
  assign new_n396_ = ~new_n391_ & ~new_n393_;
  assign \V166(4)  = new_n395_ | ~new_n396_;
  assign new_n398_ = ~\V138(2)  & \V32(3) ;
  assign new_n399_ = ~\V138(0)  & new_n398_;
  assign new_n400_ = ~\V138(2)  & \V64(3) ;
  assign new_n401_ = \V138(0)  & new_n400_;
  assign new_n402_ = \V138(2)  & ~\V64(3) ;
  assign new_n403_ = \V138(0)  & new_n402_;
  assign new_n404_ = ~new_n399_ & ~new_n401_;
  assign \V166(3)  = new_n403_ | ~new_n404_;
  assign new_n406_ = ~\V138(2)  & \V32(2) ;
  assign new_n407_ = ~\V138(0)  & new_n406_;
  assign new_n408_ = ~\V138(2)  & \V64(2) ;
  assign new_n409_ = \V138(0)  & new_n408_;
  assign new_n410_ = \V138(2)  & ~\V64(2) ;
  assign new_n411_ = \V138(0)  & new_n410_;
  assign new_n412_ = ~new_n407_ & ~new_n409_;
  assign \V166(2)  = new_n411_ | ~new_n412_;
  assign new_n414_ = ~\V138(2)  & \V32(1) ;
  assign new_n415_ = ~\V138(0)  & new_n414_;
  assign new_n416_ = ~\V138(2)  & \V64(1) ;
  assign new_n417_ = \V138(0)  & new_n416_;
  assign new_n418_ = \V138(2)  & ~\V64(1) ;
  assign new_n419_ = \V138(0)  & new_n418_;
  assign new_n420_ = ~new_n415_ & ~new_n417_;
  assign \V166(1)  = new_n419_ | ~new_n420_;
  assign new_n422_ = ~\V138(2)  & \V32(0) ;
  assign new_n423_ = ~\V138(0)  & new_n422_;
  assign new_n424_ = ~\V138(2)  & \V64(0) ;
  assign new_n425_ = \V138(0)  & new_n424_;
  assign new_n426_ = \V138(2)  & ~\V64(0) ;
  assign new_n427_ = \V138(0)  & new_n426_;
  assign new_n428_ = ~new_n423_ & ~new_n425_;
  assign \V166(0)  = new_n427_ | ~new_n428_;
  assign new_n430_ = ~\V138(0)  & \V96(27) ;
  assign new_n431_ = ~\V138(2)  & new_n430_;
  assign new_n432_ = \V138(4)  & new_n431_;
  assign new_n433_ = \V138(0)  & \V131(27) ;
  assign new_n434_ = ~\V138(2)  & new_n433_;
  assign new_n435_ = \V138(4)  & new_n434_;
  assign new_n436_ = \V138(0)  & ~\V131(27) ;
  assign new_n437_ = \V138(2)  & new_n436_;
  assign new_n438_ = \V138(4)  & new_n437_;
  assign new_n439_ = \V138(2)  & ~\V138(4) ;
  assign new_n440_ = ~new_n432_ & ~new_n435_;
  assign new_n441_ = ~new_n438_ & ~new_n439_;
  assign \V198(31)  = ~new_n440_ | ~new_n441_;
  assign new_n443_ = ~\V138(0)  & \V96(26) ;
  assign new_n444_ = ~\V138(2)  & new_n443_;
  assign new_n445_ = \V138(4)  & new_n444_;
  assign new_n446_ = \V138(0)  & \V131(26) ;
  assign new_n447_ = ~\V138(2)  & new_n446_;
  assign new_n448_ = \V138(4)  & new_n447_;
  assign new_n449_ = \V138(0)  & ~\V131(26) ;
  assign new_n450_ = \V138(2)  & new_n449_;
  assign new_n451_ = \V138(4)  & new_n450_;
  assign new_n452_ = ~new_n445_ & ~new_n448_;
  assign new_n453_ = ~new_n439_ & ~new_n451_;
  assign \V198(30)  = ~new_n452_ | ~new_n453_;
  assign new_n455_ = ~\V138(0)  & \V96(25) ;
  assign new_n456_ = ~\V138(2)  & new_n455_;
  assign new_n457_ = \V138(4)  & new_n456_;
  assign new_n458_ = \V138(0)  & \V131(25) ;
  assign new_n459_ = ~\V138(2)  & new_n458_;
  assign new_n460_ = \V138(4)  & new_n459_;
  assign new_n461_ = \V138(0)  & ~\V131(25) ;
  assign new_n462_ = \V138(2)  & new_n461_;
  assign new_n463_ = \V138(4)  & new_n462_;
  assign new_n464_ = ~new_n457_ & ~new_n460_;
  assign new_n465_ = ~new_n439_ & ~new_n463_;
  assign \V198(29)  = ~new_n464_ | ~new_n465_;
  assign new_n467_ = ~\V138(0)  & \V96(24) ;
  assign new_n468_ = ~\V138(2)  & new_n467_;
  assign new_n469_ = \V138(4)  & new_n468_;
  assign new_n470_ = \V138(0)  & \V131(24) ;
  assign new_n471_ = ~\V138(2)  & new_n470_;
  assign new_n472_ = \V138(4)  & new_n471_;
  assign new_n473_ = \V138(0)  & ~\V131(24) ;
  assign new_n474_ = \V138(2)  & new_n473_;
  assign new_n475_ = \V138(4)  & new_n474_;
  assign new_n476_ = ~new_n469_ & ~new_n472_;
  assign new_n477_ = ~new_n439_ & ~new_n475_;
  assign \V198(28)  = ~new_n476_ | ~new_n477_;
  assign new_n479_ = ~\V138(0)  & \V96(23) ;
  assign new_n480_ = ~\V138(2)  & new_n479_;
  assign new_n481_ = \V138(4)  & new_n480_;
  assign new_n482_ = \V138(0)  & \V131(23) ;
  assign new_n483_ = ~\V138(2)  & new_n482_;
  assign new_n484_ = \V138(4)  & new_n483_;
  assign new_n485_ = \V138(0)  & ~\V131(23) ;
  assign new_n486_ = \V138(2)  & new_n485_;
  assign new_n487_ = \V138(4)  & new_n486_;
  assign new_n488_ = ~new_n481_ & ~new_n484_;
  assign new_n489_ = ~new_n439_ & ~new_n487_;
  assign \V198(27)  = ~new_n488_ | ~new_n489_;
  assign new_n491_ = ~\V138(0)  & \V96(22) ;
  assign new_n492_ = ~\V138(2)  & new_n491_;
  assign new_n493_ = \V138(4)  & new_n492_;
  assign new_n494_ = \V138(0)  & \V131(22) ;
  assign new_n495_ = ~\V138(2)  & new_n494_;
  assign new_n496_ = \V138(4)  & new_n495_;
  assign new_n497_ = \V138(0)  & ~\V131(22) ;
  assign new_n498_ = \V138(2)  & new_n497_;
  assign new_n499_ = \V138(4)  & new_n498_;
  assign new_n500_ = ~new_n493_ & ~new_n496_;
  assign new_n501_ = ~new_n439_ & ~new_n499_;
  assign \V198(26)  = ~new_n500_ | ~new_n501_;
  assign new_n503_ = ~\V138(0)  & \V96(21) ;
  assign new_n504_ = ~\V138(2)  & new_n503_;
  assign new_n505_ = \V138(4)  & new_n504_;
  assign new_n506_ = \V138(0)  & \V131(21) ;
  assign new_n507_ = ~\V138(2)  & new_n506_;
  assign new_n508_ = \V138(4)  & new_n507_;
  assign new_n509_ = \V138(0)  & ~\V131(21) ;
  assign new_n510_ = \V138(2)  & new_n509_;
  assign new_n511_ = \V138(4)  & new_n510_;
  assign new_n512_ = ~new_n505_ & ~new_n508_;
  assign new_n513_ = ~new_n439_ & ~new_n511_;
  assign \V198(25)  = ~new_n512_ | ~new_n513_;
  assign new_n515_ = ~\V138(0)  & \V96(20) ;
  assign new_n516_ = ~\V138(2)  & new_n515_;
  assign new_n517_ = \V138(4)  & new_n516_;
  assign new_n518_ = \V138(0)  & \V131(20) ;
  assign new_n519_ = ~\V138(2)  & new_n518_;
  assign new_n520_ = \V138(4)  & new_n519_;
  assign new_n521_ = \V138(0)  & ~\V131(20) ;
  assign new_n522_ = \V138(2)  & new_n521_;
  assign new_n523_ = \V138(4)  & new_n522_;
  assign new_n524_ = ~new_n517_ & ~new_n520_;
  assign new_n525_ = ~new_n439_ & ~new_n523_;
  assign \V198(24)  = ~new_n524_ | ~new_n525_;
  assign new_n527_ = ~\V138(0)  & \V96(19) ;
  assign new_n528_ = ~\V138(2)  & new_n527_;
  assign new_n529_ = \V138(4)  & new_n528_;
  assign new_n530_ = \V138(0)  & \V131(19) ;
  assign new_n531_ = ~\V138(2)  & new_n530_;
  assign new_n532_ = \V138(4)  & new_n531_;
  assign new_n533_ = \V138(0)  & ~\V131(19) ;
  assign new_n534_ = \V138(2)  & new_n533_;
  assign new_n535_ = \V138(4)  & new_n534_;
  assign new_n536_ = ~new_n529_ & ~new_n532_;
  assign new_n537_ = ~new_n439_ & ~new_n535_;
  assign \V198(23)  = ~new_n536_ | ~new_n537_;
  assign new_n539_ = ~\V138(0)  & \V96(18) ;
  assign new_n540_ = ~\V138(2)  & new_n539_;
  assign new_n541_ = \V138(4)  & new_n540_;
  assign new_n542_ = \V138(0)  & \V131(18) ;
  assign new_n543_ = ~\V138(2)  & new_n542_;
  assign new_n544_ = \V138(4)  & new_n543_;
  assign new_n545_ = \V138(0)  & ~\V131(18) ;
  assign new_n546_ = \V138(2)  & new_n545_;
  assign new_n547_ = \V138(4)  & new_n546_;
  assign new_n548_ = ~new_n541_ & ~new_n544_;
  assign new_n549_ = ~new_n439_ & ~new_n547_;
  assign \V198(22)  = ~new_n548_ | ~new_n549_;
  assign new_n551_ = ~\V138(0)  & \V96(17) ;
  assign new_n552_ = ~\V138(2)  & new_n551_;
  assign new_n553_ = \V138(4)  & new_n552_;
  assign new_n554_ = \V138(0)  & \V131(17) ;
  assign new_n555_ = ~\V138(2)  & new_n554_;
  assign new_n556_ = \V138(4)  & new_n555_;
  assign new_n557_ = \V138(0)  & ~\V131(17) ;
  assign new_n558_ = \V138(2)  & new_n557_;
  assign new_n559_ = \V138(4)  & new_n558_;
  assign new_n560_ = ~new_n553_ & ~new_n556_;
  assign new_n561_ = ~new_n439_ & ~new_n559_;
  assign \V198(21)  = ~new_n560_ | ~new_n561_;
  assign new_n563_ = ~\V138(0)  & \V96(16) ;
  assign new_n564_ = ~\V138(2)  & new_n563_;
  assign new_n565_ = \V138(4)  & new_n564_;
  assign new_n566_ = \V138(0)  & \V131(16) ;
  assign new_n567_ = ~\V138(2)  & new_n566_;
  assign new_n568_ = \V138(4)  & new_n567_;
  assign new_n569_ = \V138(0)  & ~\V131(16) ;
  assign new_n570_ = \V138(2)  & new_n569_;
  assign new_n571_ = \V138(4)  & new_n570_;
  assign new_n572_ = ~new_n565_ & ~new_n568_;
  assign new_n573_ = ~new_n439_ & ~new_n571_;
  assign \V198(20)  = ~new_n572_ | ~new_n573_;
  assign new_n575_ = ~\V138(0)  & \V96(15) ;
  assign new_n576_ = ~\V138(2)  & new_n575_;
  assign new_n577_ = \V138(4)  & new_n576_;
  assign new_n578_ = \V138(0)  & \V131(15) ;
  assign new_n579_ = ~\V138(2)  & new_n578_;
  assign new_n580_ = \V138(4)  & new_n579_;
  assign new_n581_ = \V138(0)  & ~\V131(15) ;
  assign new_n582_ = \V138(2)  & new_n581_;
  assign new_n583_ = \V138(4)  & new_n582_;
  assign new_n584_ = ~new_n577_ & ~new_n580_;
  assign new_n585_ = ~new_n439_ & ~new_n583_;
  assign \V198(19)  = ~new_n584_ | ~new_n585_;
  assign new_n587_ = ~\V138(0)  & \V96(14) ;
  assign new_n588_ = ~\V138(2)  & new_n587_;
  assign new_n589_ = \V138(4)  & new_n588_;
  assign new_n590_ = \V138(0)  & \V131(14) ;
  assign new_n591_ = ~\V138(2)  & new_n590_;
  assign new_n592_ = \V138(4)  & new_n591_;
  assign new_n593_ = \V138(0)  & ~\V131(14) ;
  assign new_n594_ = \V138(2)  & new_n593_;
  assign new_n595_ = \V138(4)  & new_n594_;
  assign new_n596_ = ~new_n589_ & ~new_n592_;
  assign new_n597_ = ~new_n439_ & ~new_n595_;
  assign \V198(18)  = ~new_n596_ | ~new_n597_;
  assign new_n599_ = ~\V138(0)  & \V96(13) ;
  assign new_n600_ = ~\V138(2)  & new_n599_;
  assign new_n601_ = \V138(4)  & new_n600_;
  assign new_n602_ = \V138(0)  & \V131(13) ;
  assign new_n603_ = ~\V138(2)  & new_n602_;
  assign new_n604_ = \V138(4)  & new_n603_;
  assign new_n605_ = \V138(0)  & ~\V131(13) ;
  assign new_n606_ = \V138(2)  & new_n605_;
  assign new_n607_ = \V138(4)  & new_n606_;
  assign new_n608_ = ~new_n601_ & ~new_n604_;
  assign new_n609_ = ~new_n439_ & ~new_n607_;
  assign \V198(17)  = ~new_n608_ | ~new_n609_;
  assign new_n611_ = ~\V138(0)  & \V96(12) ;
  assign new_n612_ = ~\V138(2)  & new_n611_;
  assign new_n613_ = \V138(4)  & new_n612_;
  assign new_n614_ = \V138(0)  & \V131(12) ;
  assign new_n615_ = ~\V138(2)  & new_n614_;
  assign new_n616_ = \V138(4)  & new_n615_;
  assign new_n617_ = \V138(0)  & ~\V131(12) ;
  assign new_n618_ = \V138(2)  & new_n617_;
  assign new_n619_ = \V138(4)  & new_n618_;
  assign new_n620_ = ~new_n613_ & ~new_n616_;
  assign new_n621_ = ~new_n439_ & ~new_n619_;
  assign \V198(16)  = ~new_n620_ | ~new_n621_;
  assign new_n623_ = ~\V138(0)  & \V96(11) ;
  assign new_n624_ = ~\V138(2)  & new_n623_;
  assign new_n625_ = \V138(4)  & new_n624_;
  assign new_n626_ = \V138(0)  & \V131(11) ;
  assign new_n627_ = ~\V138(2)  & new_n626_;
  assign new_n628_ = \V138(4)  & new_n627_;
  assign new_n629_ = \V138(0)  & ~\V131(11) ;
  assign new_n630_ = \V138(2)  & new_n629_;
  assign new_n631_ = \V138(4)  & new_n630_;
  assign new_n632_ = ~new_n625_ & ~new_n628_;
  assign new_n633_ = ~new_n439_ & ~new_n631_;
  assign \V198(15)  = ~new_n632_ | ~new_n633_;
  assign new_n635_ = ~\V138(0)  & \V96(10) ;
  assign new_n636_ = ~\V138(2)  & new_n635_;
  assign new_n637_ = \V138(4)  & new_n636_;
  assign new_n638_ = \V138(0)  & \V131(10) ;
  assign new_n639_ = ~\V138(2)  & new_n638_;
  assign new_n640_ = \V138(4)  & new_n639_;
  assign new_n641_ = \V138(0)  & ~\V131(10) ;
  assign new_n642_ = \V138(2)  & new_n641_;
  assign new_n643_ = \V138(4)  & new_n642_;
  assign new_n644_ = ~new_n637_ & ~new_n640_;
  assign new_n645_ = ~new_n439_ & ~new_n643_;
  assign \V198(14)  = ~new_n644_ | ~new_n645_;
  assign new_n647_ = ~\V138(0)  & \V96(9) ;
  assign new_n648_ = ~\V138(2)  & new_n647_;
  assign new_n649_ = \V138(4)  & new_n648_;
  assign new_n650_ = \V138(0)  & \V131(9) ;
  assign new_n651_ = ~\V138(2)  & new_n650_;
  assign new_n652_ = \V138(4)  & new_n651_;
  assign new_n653_ = \V138(0)  & ~\V131(9) ;
  assign new_n654_ = \V138(2)  & new_n653_;
  assign new_n655_ = \V138(4)  & new_n654_;
  assign new_n656_ = ~new_n649_ & ~new_n652_;
  assign new_n657_ = ~new_n439_ & ~new_n655_;
  assign \V198(13)  = ~new_n656_ | ~new_n657_;
  assign new_n659_ = ~\V138(0)  & \V96(8) ;
  assign new_n660_ = ~\V138(2)  & new_n659_;
  assign new_n661_ = \V138(4)  & new_n660_;
  assign new_n662_ = \V138(0)  & \V131(8) ;
  assign new_n663_ = ~\V138(2)  & new_n662_;
  assign new_n664_ = \V138(4)  & new_n663_;
  assign new_n665_ = \V138(0)  & ~\V131(8) ;
  assign new_n666_ = \V138(2)  & new_n665_;
  assign new_n667_ = \V138(4)  & new_n666_;
  assign new_n668_ = ~new_n661_ & ~new_n664_;
  assign new_n669_ = ~new_n439_ & ~new_n667_;
  assign \V198(12)  = ~new_n668_ | ~new_n669_;
  assign new_n671_ = ~\V138(0)  & \V96(7) ;
  assign new_n672_ = ~\V138(2)  & new_n671_;
  assign new_n673_ = \V138(4)  & new_n672_;
  assign new_n674_ = \V138(0)  & \V131(7) ;
  assign new_n675_ = ~\V138(2)  & new_n674_;
  assign new_n676_ = \V138(4)  & new_n675_;
  assign new_n677_ = \V138(0)  & ~\V131(7) ;
  assign new_n678_ = \V138(2)  & new_n677_;
  assign new_n679_ = \V138(4)  & new_n678_;
  assign new_n680_ = ~new_n673_ & ~new_n676_;
  assign new_n681_ = ~new_n439_ & ~new_n679_;
  assign \V198(11)  = ~new_n680_ | ~new_n681_;
  assign new_n683_ = ~\V138(0)  & \V96(6) ;
  assign new_n684_ = ~\V138(2)  & new_n683_;
  assign new_n685_ = \V138(4)  & new_n684_;
  assign new_n686_ = \V138(0)  & \V131(6) ;
  assign new_n687_ = ~\V138(2)  & new_n686_;
  assign new_n688_ = \V138(4)  & new_n687_;
  assign new_n689_ = \V138(0)  & ~\V131(6) ;
  assign new_n690_ = \V138(2)  & new_n689_;
  assign new_n691_ = \V138(4)  & new_n690_;
  assign new_n692_ = ~new_n685_ & ~new_n688_;
  assign new_n693_ = ~new_n439_ & ~new_n691_;
  assign \V198(10)  = ~new_n692_ | ~new_n693_;
  assign new_n695_ = ~\V138(0)  & \V96(5) ;
  assign new_n696_ = ~\V138(2)  & new_n695_;
  assign new_n697_ = \V138(4)  & new_n696_;
  assign new_n698_ = \V138(0)  & \V131(5) ;
  assign new_n699_ = ~\V138(2)  & new_n698_;
  assign new_n700_ = \V138(4)  & new_n699_;
  assign new_n701_ = \V138(0)  & ~\V131(5) ;
  assign new_n702_ = \V138(2)  & new_n701_;
  assign new_n703_ = \V138(4)  & new_n702_;
  assign new_n704_ = ~new_n697_ & ~new_n700_;
  assign new_n705_ = ~new_n439_ & ~new_n703_;
  assign \V198(9)  = ~new_n704_ | ~new_n705_;
  assign new_n707_ = ~\V138(0)  & \V96(4) ;
  assign new_n708_ = ~\V138(2)  & new_n707_;
  assign new_n709_ = \V138(4)  & new_n708_;
  assign new_n710_ = \V138(0)  & \V131(4) ;
  assign new_n711_ = ~\V138(2)  & new_n710_;
  assign new_n712_ = \V138(4)  & new_n711_;
  assign new_n713_ = \V138(0)  & ~\V131(4) ;
  assign new_n714_ = \V138(2)  & new_n713_;
  assign new_n715_ = \V138(4)  & new_n714_;
  assign new_n716_ = ~new_n709_ & ~new_n712_;
  assign new_n717_ = ~new_n439_ & ~new_n715_;
  assign \V198(8)  = ~new_n716_ | ~new_n717_;
  assign new_n719_ = ~\V138(0)  & \V96(3) ;
  assign new_n720_ = ~\V138(2)  & new_n719_;
  assign new_n721_ = \V138(4)  & new_n720_;
  assign new_n722_ = \V138(0)  & \V131(3) ;
  assign new_n723_ = ~\V138(2)  & new_n722_;
  assign new_n724_ = \V138(4)  & new_n723_;
  assign new_n725_ = \V138(0)  & ~\V131(3) ;
  assign new_n726_ = \V138(2)  & new_n725_;
  assign new_n727_ = \V138(4)  & new_n726_;
  assign new_n728_ = ~new_n721_ & ~new_n724_;
  assign new_n729_ = ~new_n439_ & ~new_n727_;
  assign \V198(7)  = ~new_n728_ | ~new_n729_;
  assign new_n731_ = ~\V138(0)  & \V96(2) ;
  assign new_n732_ = ~\V138(2)  & new_n731_;
  assign new_n733_ = \V138(4)  & new_n732_;
  assign new_n734_ = \V138(0)  & \V131(2) ;
  assign new_n735_ = ~\V138(2)  & new_n734_;
  assign new_n736_ = \V138(4)  & new_n735_;
  assign new_n737_ = \V138(0)  & ~\V131(2) ;
  assign new_n738_ = \V138(2)  & new_n737_;
  assign new_n739_ = \V138(4)  & new_n738_;
  assign new_n740_ = ~new_n733_ & ~new_n736_;
  assign new_n741_ = ~new_n439_ & ~new_n739_;
  assign \V198(6)  = ~new_n740_ | ~new_n741_;
  assign new_n743_ = ~\V138(0)  & \V96(1) ;
  assign new_n744_ = ~\V138(2)  & new_n743_;
  assign new_n745_ = \V138(4)  & new_n744_;
  assign new_n746_ = \V138(0)  & \V131(1) ;
  assign new_n747_ = ~\V138(2)  & new_n746_;
  assign new_n748_ = \V138(4)  & new_n747_;
  assign new_n749_ = \V138(0)  & ~\V131(1) ;
  assign new_n750_ = \V138(2)  & new_n749_;
  assign new_n751_ = \V138(4)  & new_n750_;
  assign new_n752_ = ~new_n745_ & ~new_n748_;
  assign new_n753_ = ~new_n439_ & ~new_n751_;
  assign \V198(5)  = ~new_n752_ | ~new_n753_;
  assign new_n755_ = ~\V138(0)  & \V96(0) ;
  assign new_n756_ = ~\V138(2)  & new_n755_;
  assign new_n757_ = \V138(4)  & new_n756_;
  assign new_n758_ = \V138(0)  & \V131(0) ;
  assign new_n759_ = ~\V138(2)  & new_n758_;
  assign new_n760_ = \V138(4)  & new_n759_;
  assign new_n761_ = \V138(0)  & ~\V131(0) ;
  assign new_n762_ = \V138(2)  & new_n761_;
  assign new_n763_ = \V138(4)  & new_n762_;
  assign new_n764_ = ~new_n757_ & ~new_n760_;
  assign new_n765_ = ~new_n439_ & ~new_n763_;
  assign \V198(4)  = ~new_n764_ | ~new_n765_;
  assign new_n767_ = ~\V138(0)  & \V32(31) ;
  assign new_n768_ = ~\V138(2)  & new_n767_;
  assign new_n769_ = \V138(4)  & new_n768_;
  assign new_n770_ = \V138(0)  & \V64(31) ;
  assign new_n771_ = ~\V138(2)  & new_n770_;
  assign new_n772_ = \V138(4)  & new_n771_;
  assign new_n773_ = \V138(0)  & ~\V64(31) ;
  assign new_n774_ = \V138(2)  & new_n773_;
  assign new_n775_ = \V138(4)  & new_n774_;
  assign new_n776_ = ~new_n769_ & ~new_n772_;
  assign new_n777_ = ~new_n439_ & ~new_n775_;
  assign \V198(3)  = ~new_n776_ | ~new_n777_;
  assign new_n779_ = ~\V138(0)  & \V32(30) ;
  assign new_n780_ = ~\V138(2)  & new_n779_;
  assign new_n781_ = \V138(4)  & new_n780_;
  assign new_n782_ = \V138(0)  & \V64(30) ;
  assign new_n783_ = ~\V138(2)  & new_n782_;
  assign new_n784_ = \V138(4)  & new_n783_;
  assign new_n785_ = \V138(0)  & ~\V64(30) ;
  assign new_n786_ = \V138(2)  & new_n785_;
  assign new_n787_ = \V138(4)  & new_n786_;
  assign new_n788_ = ~new_n781_ & ~new_n784_;
  assign new_n789_ = ~new_n439_ & ~new_n787_;
  assign \V198(2)  = ~new_n788_ | ~new_n789_;
  assign new_n791_ = ~\V138(0)  & \V32(29) ;
  assign new_n792_ = ~\V138(2)  & new_n791_;
  assign new_n793_ = \V138(4)  & new_n792_;
  assign new_n794_ = \V138(0)  & \V64(29) ;
  assign new_n795_ = ~\V138(2)  & new_n794_;
  assign new_n796_ = \V138(4)  & new_n795_;
  assign new_n797_ = \V138(0)  & ~\V64(29) ;
  assign new_n798_ = \V138(2)  & new_n797_;
  assign new_n799_ = \V138(4)  & new_n798_;
  assign new_n800_ = ~new_n793_ & ~new_n796_;
  assign new_n801_ = ~new_n439_ & ~new_n799_;
  assign \V198(1)  = ~new_n800_ | ~new_n801_;
  assign new_n803_ = ~\V138(0)  & \V32(28) ;
  assign new_n804_ = ~\V138(2)  & new_n803_;
  assign new_n805_ = \V138(4)  & new_n804_;
  assign new_n806_ = \V138(0)  & \V64(28) ;
  assign new_n807_ = ~\V138(2)  & new_n806_;
  assign new_n808_ = \V138(4)  & new_n807_;
  assign new_n809_ = \V138(0)  & ~\V64(28) ;
  assign new_n810_ = \V138(2)  & new_n809_;
  assign new_n811_ = \V138(4)  & new_n810_;
  assign new_n812_ = ~new_n805_ & ~new_n808_;
  assign new_n813_ = ~new_n439_ & ~new_n811_;
  assign \V198(0)  = ~new_n812_ | ~new_n813_;
  assign new_n815_ = ~\V138(0)  & \V99(0) ;
  assign new_n816_ = ~\V138(2)  & new_n815_;
  assign new_n817_ = \V138(3)  & new_n816_;
  assign new_n818_ = \V138(0)  & \V134(0) ;
  assign new_n819_ = ~\V138(2)  & new_n818_;
  assign new_n820_ = \V138(3)  & new_n819_;
  assign new_n821_ = \V138(2)  & new_n818_;
  assign new_n822_ = \V138(3)  & new_n821_;
  assign new_n823_ = ~new_n817_ & ~new_n820_;
  assign \V205(6)  = new_n822_ | ~new_n823_;
  assign new_n825_ = ~\V138(0)  & \V98(0) ;
  assign new_n826_ = ~\V138(2)  & new_n825_;
  assign new_n827_ = \V138(3)  & new_n826_;
  assign new_n828_ = \V138(0)  & \V133(1) ;
  assign new_n829_ = ~\V138(2)  & new_n828_;
  assign new_n830_ = \V138(3)  & new_n829_;
  assign new_n831_ = \V138(0)  & ~\V133(1) ;
  assign new_n832_ = \V138(2)  & new_n831_;
  assign new_n833_ = \V138(3)  & new_n832_;
  assign new_n834_ = \V138(2)  & ~\V138(3) ;
  assign new_n835_ = ~new_n827_ & ~new_n830_;
  assign new_n836_ = ~new_n833_ & ~new_n834_;
  assign \V205(5)  = ~new_n835_ | ~new_n836_;
  assign new_n838_ = ~\V138(0)  & \V97(0) ;
  assign new_n839_ = ~\V138(2)  & new_n838_;
  assign new_n840_ = \V138(3)  & new_n839_;
  assign new_n841_ = \V138(0)  & \V133(0) ;
  assign new_n842_ = ~\V138(2)  & new_n841_;
  assign new_n843_ = \V138(3)  & new_n842_;
  assign new_n844_ = \V138(0)  & ~\V133(0) ;
  assign new_n845_ = \V138(2)  & new_n844_;
  assign new_n846_ = \V138(3)  & new_n845_;
  assign new_n847_ = ~new_n840_ & ~new_n843_;
  assign new_n848_ = ~new_n834_ & ~new_n846_;
  assign \V205(4)  = ~new_n847_ | ~new_n848_;
  assign new_n850_ = ~\V138(0)  & \V96(31) ;
  assign new_n851_ = ~\V138(2)  & new_n850_;
  assign new_n852_ = \V138(3)  & new_n851_;
  assign new_n853_ = \V138(0)  & \V131(31) ;
  assign new_n854_ = ~\V138(2)  & new_n853_;
  assign new_n855_ = \V138(3)  & new_n854_;
  assign new_n856_ = \V138(0)  & ~\V131(31) ;
  assign new_n857_ = \V138(2)  & new_n856_;
  assign new_n858_ = \V138(3)  & new_n857_;
  assign new_n859_ = ~new_n852_ & ~new_n855_;
  assign new_n860_ = ~new_n834_ & ~new_n858_;
  assign \V205(3)  = ~new_n859_ | ~new_n860_;
  assign new_n862_ = ~\V138(0)  & \V96(30) ;
  assign new_n863_ = ~\V138(2)  & new_n862_;
  assign new_n864_ = \V138(3)  & new_n863_;
  assign new_n865_ = \V138(0)  & \V131(30) ;
  assign new_n866_ = ~\V138(2)  & new_n865_;
  assign new_n867_ = \V138(3)  & new_n866_;
  assign new_n868_ = \V138(0)  & ~\V131(30) ;
  assign new_n869_ = \V138(2)  & new_n868_;
  assign new_n870_ = \V138(3)  & new_n869_;
  assign new_n871_ = ~new_n864_ & ~new_n867_;
  assign new_n872_ = ~new_n834_ & ~new_n870_;
  assign \V205(2)  = ~new_n871_ | ~new_n872_;
  assign new_n874_ = ~\V138(0)  & \V96(29) ;
  assign new_n875_ = ~\V138(2)  & new_n874_;
  assign new_n876_ = \V138(3)  & new_n875_;
  assign new_n877_ = \V138(0)  & \V131(29) ;
  assign new_n878_ = ~\V138(2)  & new_n877_;
  assign new_n879_ = \V138(3)  & new_n878_;
  assign new_n880_ = \V138(0)  & ~\V131(29) ;
  assign new_n881_ = \V138(2)  & new_n880_;
  assign new_n882_ = \V138(3)  & new_n881_;
  assign new_n883_ = ~new_n876_ & ~new_n879_;
  assign new_n884_ = ~new_n834_ & ~new_n882_;
  assign \V205(1)  = ~new_n883_ | ~new_n884_;
  assign new_n886_ = ~\V138(0)  & \V96(28) ;
  assign new_n887_ = ~\V138(2)  & new_n886_;
  assign new_n888_ = \V138(3)  & new_n887_;
  assign new_n889_ = \V138(0)  & \V131(28) ;
  assign new_n890_ = ~\V138(2)  & new_n889_;
  assign new_n891_ = \V138(3)  & new_n890_;
  assign new_n892_ = \V138(0)  & ~\V131(28) ;
  assign new_n893_ = \V138(2)  & new_n892_;
  assign new_n894_ = \V138(3)  & new_n893_;
  assign new_n895_ = ~new_n888_ & ~new_n891_;
  assign new_n896_ = ~new_n834_ & ~new_n894_;
  assign \V205(0)  = ~new_n895_ | ~new_n896_;
endmodule

