module top ( 
    p_193_130_, p_257_171_, p_2435_225_, p_79_60_, p_135_106_, p_142_113_,
    p_192_129_, p_209_146_, p_2096_218_, p_2454_230_, p_4_3_, p_51_36_,
    p_52_37_, p_112_87_, p_126_99_, p_179_118_, p_189_126_, p_21_14_,
    p_25_18_, p_90_69_, p_206_143_, p_253_167_, p_277_187_, p_60_43_,
    p_61_44_, p_66_49_, p_202_139_, p_22_15_, p_24_17_, p_119_94_,
    p_132_105_, p_203_140_, p_250_164_, p_267_177_, p_270_180_, p_559_193_,
    p_2443_227_, p_3_2_, p_53_38_, p_54_39_, p_102_79_, p_182_121_,
    p_212_149_, p_1961_204_, p_1986_209_, p_2090_217_, p_2430_224_,
    p_23_16_, p_169_114_, p_213_150_, p_242_156_, p_28_21_, p_29_22_,
    p_93_72_, p_94_73_, p_95_74_, p_96_75_, p_128_101_, p_651_195_,
    p_661_196_, p_14_9_, p_32_23_, p_34_25_, p_36_27_, p_67_50_, p_69_52_,
    p_104_81_, p_106_83_, p_252_166_, p_269_179_, p_276_186_, p_2_1_,
    p_72_53_, p_99_76_, p_100_77_, p_113_88_, p_125_98_, p_2451_229_,
    p_35_26_, p_116_91_, p_136_107_, p_240_154_, p_273_183_, p_62_45_,
    p_63_46_, p_64_47_, p_65_48_, p_183_122_, p_199_136_, p_1981_208_,
    p_1996_211_, p_11_8_, p_26_19_, p_140_111_, p_207_144_, p_214_151_,
    p_243_157_, p_263_173_, p_1_0_, p_186_125_, p_196_133_, p_247_161_,
    p_33_24_, p_68_51_, p_204_141_, p_266_176_, p_279_189_, p_2678_232_,
    p_19_12_, p_85_64_, p_86_65_, p_87_66_, p_88_67_, p_89_68_, p_120_95_,
    p_181_120_, p_200_137_, p_2100_219_, p_130_103_, p_180_119_,
    p_241_155_, p_265_175_, p_272_182_, p_567_194_, p_8_7_, p_15_10_,
    p_16_11_, p_80_61_, p_81_62_, p_127_100_, p_174_115_, p_184_123_,
    p_198_135_, p_210_147_, p_56_41_, p_103_80_, p_107_84_, p_244_158_,
    p_268_178_, p_1976_207_, p_195_132_, p_248_162_, p_2066_212_,
    p_2106_222_, p_2474_231_, p_43_30_, p_57_42_, p_117_92_, p_137_108_,
    p_278_188_, p_483_191_, p_1384_202_, p_1971_206_, p_7_6_, p_73_54_,
    p_74_55_, p_123_96_, p_177_116_, p_256_170_, p_1083_199_, p_1341_200_,
    p_1991_210_, p_2067_213_, p_2078_215_, p_2105_221_, p_37_28_, p_44_31_,
    p_191_128_, p_208_145_, p_255_169_, p_262_172_, p_275_185_, p_868_198_,
    p_27_20_, p_91_70_, p_92_71_, p_178_117_, p_185_124_, p_197_134_,
    p_211_148_, p_239_153_, p_246_160_, p_2084_216_, p_2104_220_,
    p_108_85_, p_205_142_, p_245_159_, p_2446_228_, p_6_5_, p_40_29_,
    p_75_56_, p_76_57_, p_194_131_, p_201_138_, p_249_163_, p_452_190_,
    p_47_32_, p_131_104_, p_141_112_, p_215_152_, p_264_174_, p_2427_223_,
    p_1966_205_, p_2438_226_, p_20_13_, p_48_33_, p_55_40_, p_115_90_,
    p_190_127_, p_254_168_, p_274_184_, p_543_192_, p_1956_203_, p_5_4_,
    p_50_35_, p_77_58_, p_78_59_, p_82_63_, p_101_78_, p_111_86_,
    p_114_89_, p_124_97_, p_129_102_, p_139_110_, p_860_197_, p_1348_201_,
    p_49_34_, p_105_82_, p_118_93_, p_138_109_, p_251_165_, p_271_181_,
    p_2072_214_,
    p_284_847_, p_171_621_, p_145_1358_, p_150_1277_, p_188_761_,
    p_221_305_, p_311_1278_, p_158_349_, p_235_307_, p_259_414_,
    p_299_692_, p_160_609_, p_367_288_, p_288_700_, p_301_694_, p_384_262_,
    p_218_311_, p_261_506_, p_236_303_, p_319_656_, p_321_848_, p_350_301_,
    p_397_1406_, p_148_851_, p_220_306_, p_369_289_, p_164_607_,
    p_411_264_, p_231_1422_, p_297_849_, p_168_623_, p_156_1046_,
    p_337_263_, p_153_671_, p_223_413_, p_303_698_, p_331_1401_,
    p_391_379_, p_395_1392_, p_282_922_, p_173_389_, p_217_423_,
    p_229_1180_, p_280_850_, p_335_299_, p_162_612_, p_227_1179_,
    p_237_309_, p_176_803_, p_305_702_, p_290_704_, p_329_1414_,
    p_286_696_, p_295_1400_, p_401_1276_, p_238_304_, p_323_923_,
    p_325_507_, p_219_302_, p_166_625_, p_409_298_, p_234_376_,
    p_308_1425_, p_225_1424_  );
  input  p_193_130_, p_257_171_, p_2435_225_, p_79_60_, p_135_106_,
    p_142_113_, p_192_129_, p_209_146_, p_2096_218_, p_2454_230_, p_4_3_,
    p_51_36_, p_52_37_, p_112_87_, p_126_99_, p_179_118_, p_189_126_,
    p_21_14_, p_25_18_, p_90_69_, p_206_143_, p_253_167_, p_277_187_,
    p_60_43_, p_61_44_, p_66_49_, p_202_139_, p_22_15_, p_24_17_,
    p_119_94_, p_132_105_, p_203_140_, p_250_164_, p_267_177_, p_270_180_,
    p_559_193_, p_2443_227_, p_3_2_, p_53_38_, p_54_39_, p_102_79_,
    p_182_121_, p_212_149_, p_1961_204_, p_1986_209_, p_2090_217_,
    p_2430_224_, p_23_16_, p_169_114_, p_213_150_, p_242_156_, p_28_21_,
    p_29_22_, p_93_72_, p_94_73_, p_95_74_, p_96_75_, p_128_101_,
    p_651_195_, p_661_196_, p_14_9_, p_32_23_, p_34_25_, p_36_27_,
    p_67_50_, p_69_52_, p_104_81_, p_106_83_, p_252_166_, p_269_179_,
    p_276_186_, p_2_1_, p_72_53_, p_99_76_, p_100_77_, p_113_88_,
    p_125_98_, p_2451_229_, p_35_26_, p_116_91_, p_136_107_, p_240_154_,
    p_273_183_, p_62_45_, p_63_46_, p_64_47_, p_65_48_, p_183_122_,
    p_199_136_, p_1981_208_, p_1996_211_, p_11_8_, p_26_19_, p_140_111_,
    p_207_144_, p_214_151_, p_243_157_, p_263_173_, p_1_0_, p_186_125_,
    p_196_133_, p_247_161_, p_33_24_, p_68_51_, p_204_141_, p_266_176_,
    p_279_189_, p_2678_232_, p_19_12_, p_85_64_, p_86_65_, p_87_66_,
    p_88_67_, p_89_68_, p_120_95_, p_181_120_, p_200_137_, p_2100_219_,
    p_130_103_, p_180_119_, p_241_155_, p_265_175_, p_272_182_, p_567_194_,
    p_8_7_, p_15_10_, p_16_11_, p_80_61_, p_81_62_, p_127_100_, p_174_115_,
    p_184_123_, p_198_135_, p_210_147_, p_56_41_, p_103_80_, p_107_84_,
    p_244_158_, p_268_178_, p_1976_207_, p_195_132_, p_248_162_,
    p_2066_212_, p_2106_222_, p_2474_231_, p_43_30_, p_57_42_, p_117_92_,
    p_137_108_, p_278_188_, p_483_191_, p_1384_202_, p_1971_206_, p_7_6_,
    p_73_54_, p_74_55_, p_123_96_, p_177_116_, p_256_170_, p_1083_199_,
    p_1341_200_, p_1991_210_, p_2067_213_, p_2078_215_, p_2105_221_,
    p_37_28_, p_44_31_, p_191_128_, p_208_145_, p_255_169_, p_262_172_,
    p_275_185_, p_868_198_, p_27_20_, p_91_70_, p_92_71_, p_178_117_,
    p_185_124_, p_197_134_, p_211_148_, p_239_153_, p_246_160_,
    p_2084_216_, p_2104_220_, p_108_85_, p_205_142_, p_245_159_,
    p_2446_228_, p_6_5_, p_40_29_, p_75_56_, p_76_57_, p_194_131_,
    p_201_138_, p_249_163_, p_452_190_, p_47_32_, p_131_104_, p_141_112_,
    p_215_152_, p_264_174_, p_2427_223_, p_1966_205_, p_2438_226_,
    p_20_13_, p_48_33_, p_55_40_, p_115_90_, p_190_127_, p_254_168_,
    p_274_184_, p_543_192_, p_1956_203_, p_5_4_, p_50_35_, p_77_58_,
    p_78_59_, p_82_63_, p_101_78_, p_111_86_, p_114_89_, p_124_97_,
    p_129_102_, p_139_110_, p_860_197_, p_1348_201_, p_49_34_, p_105_82_,
    p_118_93_, p_138_109_, p_251_165_, p_271_181_, p_2072_214_;
  output p_284_847_, p_171_621_, p_145_1358_, p_150_1277_, p_188_761_,
    p_221_305_, p_311_1278_, p_158_349_, p_235_307_, p_259_414_,
    p_299_692_, p_160_609_, p_367_288_, p_288_700_, p_301_694_, p_384_262_,
    p_218_311_, p_261_506_, p_236_303_, p_319_656_, p_321_848_, p_350_301_,
    p_397_1406_, p_148_851_, p_220_306_, p_369_289_, p_164_607_,
    p_411_264_, p_231_1422_, p_297_849_, p_168_623_, p_156_1046_,
    p_337_263_, p_153_671_, p_223_413_, p_303_698_, p_331_1401_,
    p_391_379_, p_395_1392_, p_282_922_, p_173_389_, p_217_423_,
    p_229_1180_, p_280_850_, p_335_299_, p_162_612_, p_227_1179_,
    p_237_309_, p_176_803_, p_305_702_, p_290_704_, p_329_1414_,
    p_286_696_, p_295_1400_, p_401_1276_, p_238_304_, p_323_923_,
    p_325_507_, p_219_302_, p_166_625_, p_409_298_, p_234_376_,
    p_308_1425_, p_225_1424_;
  wire new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n577_, new_n578_, new_n580_, new_n581_, new_n583_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n940_, new_n941_, new_n942_, new_n943_;
  assign new_n299_ = p_651_195_ & p_543_192_;
  assign new_n300_ = p_77_58_ & new_n299_;
  assign new_n301_ = ~p_651_195_ & p_543_192_;
  assign new_n302_ = p_52_37_ & new_n301_;
  assign new_n303_ = p_651_195_ & ~p_543_192_;
  assign new_n304_ = p_64_47_ & new_n303_;
  assign new_n305_ = ~p_651_195_ & ~p_543_192_;
  assign new_n306_ = p_90_69_ & new_n305_;
  assign new_n307_ = ~new_n300_ & ~new_n302_;
  assign new_n308_ = ~new_n304_ & new_n307_;
  assign p_171_621_ = ~new_n306_ & new_n308_;
  assign new_n310_ = p_868_198_ & ~p_171_621_;
  assign new_n311_ = p_79_60_ & new_n299_;
  assign new_n312_ = p_54_39_ & new_n301_;
  assign new_n313_ = p_66_49_ & new_n303_;
  assign new_n314_ = p_92_71_ & new_n305_;
  assign new_n315_ = ~new_n311_ & ~new_n312_;
  assign new_n316_ = ~new_n313_ & new_n315_;
  assign new_n317_ = ~new_n314_ & new_n316_;
  assign new_n318_ = ~p_868_198_ & ~new_n317_;
  assign p_284_847_ = new_n310_ | new_n318_;
  assign new_n320_ = p_80_61_ & new_n299_;
  assign new_n321_ = p_55_40_ & new_n301_;
  assign new_n322_ = p_67_50_ & new_n303_;
  assign new_n323_ = p_93_72_ & new_n305_;
  assign new_n324_ = ~new_n320_ & ~new_n321_;
  assign new_n325_ = ~new_n322_ & new_n324_;
  assign new_n326_ = ~new_n323_ & new_n325_;
  assign new_n327_ = p_860_197_ & ~new_n326_;
  assign new_n328_ = p_68_51_ & new_n299_;
  assign new_n329_ = p_43_30_ & new_n301_;
  assign new_n330_ = p_56_41_ & new_n303_;
  assign new_n331_ = p_81_62_ & new_n305_;
  assign new_n332_ = ~new_n328_ & ~new_n329_;
  assign new_n333_ = ~new_n330_ & new_n332_;
  assign new_n334_ = ~new_n331_ & new_n333_;
  assign new_n335_ = ~new_n317_ & new_n334_;
  assign new_n336_ = new_n317_ & ~new_n334_;
  assign new_n337_ = ~new_n335_ & ~new_n336_;
  assign new_n338_ = ~p_559_193_ & new_n317_;
  assign new_n339_ = new_n337_ & new_n338_;
  assign new_n340_ = ~new_n337_ & ~new_n338_;
  assign new_n341_ = ~new_n339_ & ~new_n340_;
  assign new_n342_ = ~new_n326_ & new_n341_;
  assign new_n343_ = new_n326_ & ~new_n341_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = ~p_860_197_ & ~new_n344_;
  assign p_145_1358_ = new_n327_ | new_n345_;
  assign new_n347_ = p_2105_221_ & p_2104_220_;
  assign new_n348_ = p_116_91_ & new_n347_;
  assign new_n349_ = ~p_2105_221_ & p_2104_220_;
  assign new_n350_ = p_104_81_ & new_n349_;
  assign new_n351_ = p_2105_221_ & ~p_2104_220_;
  assign new_n352_ = p_128_101_ & new_n351_;
  assign new_n353_ = ~p_2105_221_ & ~p_2104_220_;
  assign new_n354_ = p_140_111_ & new_n353_;
  assign new_n355_ = ~new_n348_ & ~new_n350_;
  assign new_n356_ = ~new_n352_ & new_n355_;
  assign new_n357_ = ~new_n354_ & new_n356_;
  assign new_n358_ = p_29_22_ & ~new_n357_;
  assign new_n359_ = ~p_29_22_ & p_26_19_;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~p_2067_213_ & new_n360_;
  assign new_n362_ = p_2067_213_ & ~new_n360_;
  assign new_n363_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = p_117_92_ & new_n347_;
  assign new_n365_ = p_105_82_ & new_n349_;
  assign new_n366_ = p_129_102_ & new_n351_;
  assign new_n367_ = p_141_112_ & new_n353_;
  assign new_n368_ = ~new_n364_ & ~new_n365_;
  assign new_n369_ = ~new_n366_ & new_n368_;
  assign new_n370_ = ~new_n367_ & new_n369_;
  assign new_n371_ = p_29_22_ & ~new_n370_;
  assign new_n372_ = ~p_29_22_ & p_32_23_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = ~p_1996_211_ & new_n373_;
  assign new_n375_ = p_1996_211_ & ~new_n373_;
  assign new_n376_ = ~new_n374_ & ~new_n375_;
  assign new_n377_ = p_114_89_ & new_n347_;
  assign new_n378_ = p_102_79_ & new_n349_;
  assign new_n379_ = p_126_99_ & new_n351_;
  assign new_n380_ = p_138_109_ & new_n353_;
  assign new_n381_ = ~new_n377_ & ~new_n378_;
  assign new_n382_ = ~new_n379_ & new_n381_;
  assign p_164_607_ = ~new_n380_ & new_n382_;
  assign new_n384_ = p_29_22_ & ~p_164_607_;
  assign new_n385_ = ~p_29_22_ & p_27_20_;
  assign new_n386_ = ~new_n384_ & ~new_n385_;
  assign new_n387_ = ~p_2078_215_ & new_n386_;
  assign new_n388_ = p_2078_215_ & ~new_n386_;
  assign new_n389_ = ~new_n387_ & ~new_n388_;
  assign new_n390_ = p_115_90_ & new_n347_;
  assign new_n391_ = p_103_80_ & new_n349_;
  assign new_n392_ = p_127_100_ & new_n351_;
  assign new_n393_ = p_139_110_ & new_n353_;
  assign new_n394_ = ~new_n390_ & ~new_n391_;
  assign new_n395_ = ~new_n392_ & new_n394_;
  assign new_n396_ = ~new_n393_ & new_n395_;
  assign new_n397_ = p_29_22_ & ~new_n396_;
  assign new_n398_ = ~p_29_22_ & p_33_24_;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = ~p_2072_214_ & new_n399_;
  assign new_n401_ = p_2072_214_ & ~new_n399_;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign new_n403_ = p_113_88_ & new_n347_;
  assign new_n404_ = p_101_78_ & new_n349_;
  assign new_n405_ = p_125_98_ & new_n351_;
  assign new_n406_ = p_137_108_ & new_n353_;
  assign new_n407_ = ~new_n403_ & ~new_n404_;
  assign new_n408_ = ~new_n405_ & new_n407_;
  assign p_160_609_ = ~new_n406_ & new_n408_;
  assign new_n410_ = p_29_22_ & ~p_160_609_;
  assign new_n411_ = ~p_29_22_ & p_34_25_;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = ~p_2084_216_ & new_n412_;
  assign new_n414_ = p_2084_216_ & ~new_n412_;
  assign new_n415_ = ~new_n413_ & ~new_n414_;
  assign new_n416_ = new_n363_ & new_n376_;
  assign new_n417_ = new_n389_ & new_n416_;
  assign new_n418_ = new_n402_ & new_n417_;
  assign new_n419_ = new_n415_ & new_n418_;
  assign new_n420_ = p_112_87_ & new_n347_;
  assign new_n421_ = p_100_77_ & new_n349_;
  assign new_n422_ = p_124_97_ & new_n351_;
  assign new_n423_ = p_136_107_ & new_n353_;
  assign new_n424_ = ~new_n420_ & ~new_n421_;
  assign new_n425_ = ~new_n422_ & new_n424_;
  assign p_162_612_ = ~new_n423_ & new_n425_;
  assign new_n427_ = p_29_22_ & ~p_162_612_;
  assign new_n428_ = ~p_29_22_ & p_35_26_;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = ~p_2090_217_ & new_n429_;
  assign new_n431_ = p_2090_217_ & ~new_n429_;
  assign new_n432_ = ~new_n430_ & ~new_n431_;
  assign new_n433_ = p_111_86_ & new_n347_;
  assign new_n434_ = p_99_76_ & new_n349_;
  assign new_n435_ = p_123_96_ & new_n351_;
  assign new_n436_ = p_135_106_ & new_n353_;
  assign new_n437_ = ~new_n433_ & ~new_n434_;
  assign new_n438_ = ~new_n435_ & new_n437_;
  assign new_n439_ = ~new_n436_ & new_n438_;
  assign new_n440_ = p_29_22_ & ~new_n439_;
  assign new_n441_ = p_28_21_ & ~p_29_22_;
  assign new_n442_ = ~new_n440_ & ~new_n441_;
  assign new_n443_ = new_n432_ & ~new_n442_;
  assign new_n444_ = new_n419_ & new_n443_;
  assign new_n445_ = p_11_8_ & p_868_198_;
  assign new_n446_ = p_11_8_ & ~p_868_198_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = p_16_11_ & ~new_n317_;
  assign new_n449_ = p_4_3_ & ~p_16_11_;
  assign new_n450_ = ~new_n448_ & ~new_n449_;
  assign new_n451_ = ~p_1348_201_ & new_n450_;
  assign new_n452_ = p_1348_201_ & ~new_n450_;
  assign new_n453_ = ~new_n451_ & ~new_n452_;
  assign new_n454_ = p_16_11_ & ~new_n334_;
  assign new_n455_ = p_19_12_ & ~p_16_11_;
  assign new_n456_ = ~new_n454_ & ~new_n455_;
  assign new_n457_ = ~p_1341_200_ & new_n456_;
  assign new_n458_ = p_1341_200_ & ~new_n456_;
  assign new_n459_ = ~new_n457_ & ~new_n458_;
  assign new_n460_ = p_16_11_ & ~p_171_621_;
  assign new_n461_ = ~p_16_11_ & p_5_4_;
  assign new_n462_ = ~new_n460_ & ~new_n461_;
  assign new_n463_ = ~p_1961_204_ & new_n462_;
  assign new_n464_ = p_1961_204_ & ~new_n462_;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign new_n466_ = p_78_59_ & new_n299_;
  assign new_n467_ = p_53_38_ & new_n301_;
  assign new_n468_ = p_65_48_ & new_n303_;
  assign new_n469_ = p_91_70_ & new_n305_;
  assign new_n470_ = ~new_n466_ & ~new_n467_;
  assign new_n471_ = ~new_n468_ & new_n470_;
  assign p_299_692_ = new_n469_ | ~new_n471_;
  assign new_n473_ = p_16_11_ & p_299_692_;
  assign new_n474_ = ~p_16_11_ & p_20_13_;
  assign new_n475_ = ~new_n473_ & ~new_n474_;
  assign new_n476_ = ~p_1956_203_ & new_n475_;
  assign new_n477_ = p_1956_203_ & ~new_n475_;
  assign new_n478_ = ~new_n476_ & ~new_n477_;
  assign new_n479_ = p_76_57_ & new_n299_;
  assign new_n480_ = p_51_36_ & new_n301_;
  assign new_n481_ = p_63_46_ & new_n303_;
  assign new_n482_ = p_89_68_ & new_n305_;
  assign new_n483_ = ~new_n479_ & ~new_n480_;
  assign new_n484_ = ~new_n481_ & new_n483_;
  assign p_168_623_ = ~new_n482_ & new_n484_;
  assign new_n486_ = p_16_11_ & ~p_168_623_;
  assign new_n487_ = p_21_14_ & ~p_16_11_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = ~p_1966_205_ & new_n488_;
  assign new_n490_ = p_1966_205_ & ~new_n488_;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = new_n453_ & new_n459_;
  assign new_n493_ = new_n465_ & new_n492_;
  assign new_n494_ = new_n478_ & new_n493_;
  assign new_n495_ = new_n491_ & new_n494_;
  assign new_n496_ = p_74_55_ & new_n299_;
  assign new_n497_ = p_49_34_ & new_n301_;
  assign new_n498_ = p_87_66_ & new_n305_;
  assign new_n499_ = ~new_n496_ & ~new_n497_;
  assign new_n500_ = ~new_n303_ & new_n499_;
  assign p_288_700_ = new_n498_ | ~new_n500_;
  assign new_n502_ = p_16_11_ & p_288_700_;
  assign new_n503_ = p_23_16_ & ~p_16_11_;
  assign new_n504_ = ~new_n502_ & ~new_n503_;
  assign new_n505_ = ~p_1976_207_ & new_n504_;
  assign new_n506_ = p_1976_207_ & ~new_n504_;
  assign new_n507_ = ~new_n505_ & ~new_n506_;
  assign new_n508_ = p_75_56_ & new_n299_;
  assign new_n509_ = p_50_35_ & new_n301_;
  assign new_n510_ = p_62_45_ & new_n303_;
  assign new_n511_ = p_88_67_ & new_n305_;
  assign new_n512_ = ~new_n508_ & ~new_n509_;
  assign new_n513_ = ~new_n510_ & new_n512_;
  assign p_166_625_ = ~new_n511_ & new_n513_;
  assign new_n515_ = p_16_11_ & ~p_166_625_;
  assign new_n516_ = p_22_15_ & ~p_16_11_;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_ = ~p_1971_206_ & new_n517_;
  assign new_n519_ = p_1971_206_ & ~new_n517_;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = p_72_53_ & new_n299_;
  assign new_n522_ = p_47_32_ & new_n301_;
  assign new_n523_ = p_60_43_ & new_n303_;
  assign new_n524_ = p_85_64_ & new_n305_;
  assign new_n525_ = ~new_n521_ & ~new_n522_;
  assign new_n526_ = ~new_n523_ & new_n525_;
  assign p_290_704_ = new_n524_ | ~new_n526_;
  assign new_n528_ = p_16_11_ & p_290_704_;
  assign new_n529_ = p_24_17_ & ~p_16_11_;
  assign new_n530_ = ~new_n528_ & ~new_n529_;
  assign new_n531_ = ~p_1986_209_ & new_n530_;
  assign new_n532_ = p_1986_209_ & ~new_n530_;
  assign new_n533_ = ~new_n531_ & ~new_n532_;
  assign new_n534_ = p_73_54_ & new_n299_;
  assign new_n535_ = p_48_33_ & new_n301_;
  assign new_n536_ = p_61_44_ & new_n303_;
  assign new_n537_ = p_86_65_ & new_n305_;
  assign new_n538_ = ~new_n534_ & ~new_n535_;
  assign new_n539_ = ~new_n536_ & new_n538_;
  assign p_305_702_ = new_n537_ | ~new_n539_;
  assign new_n541_ = p_16_11_ & p_305_702_;
  assign new_n542_ = ~p_16_11_ & p_6_5_;
  assign new_n543_ = ~new_n541_ & ~new_n542_;
  assign new_n544_ = ~p_1981_208_ & new_n543_;
  assign new_n545_ = p_1981_208_ & ~new_n543_;
  assign new_n546_ = ~new_n544_ & ~new_n545_;
  assign new_n547_ = p_107_84_ & new_n347_;
  assign new_n548_ = p_95_74_ & new_n349_;
  assign new_n549_ = p_119_94_ & new_n351_;
  assign new_n550_ = p_131_104_ & new_n353_;
  assign new_n551_ = ~new_n547_ & ~new_n548_;
  assign new_n552_ = ~new_n549_ & new_n551_;
  assign new_n553_ = ~new_n550_ & new_n552_;
  assign new_n554_ = p_29_22_ & ~new_n553_;
  assign new_n555_ = p_25_18_ & ~p_29_22_;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = ~p_1991_210_ & new_n556_;
  assign new_n558_ = p_1991_210_ & ~new_n556_;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = new_n507_ & new_n520_;
  assign new_n561_ = new_n533_ & new_n560_;
  assign new_n562_ = new_n546_ & new_n561_;
  assign new_n563_ = new_n559_ & new_n562_;
  assign new_n564_ = new_n495_ & new_n563_;
  assign new_n565_ = new_n444_ & ~new_n447_;
  assign p_311_1278_ = new_n564_ & new_n565_;
  assign new_n567_ = p_3_2_ & p_1_0_;
  assign new_n568_ = p_69_52_ & p_57_42_;
  assign new_n569_ = p_108_85_ & new_n568_;
  assign new_n570_ = p_120_95_ & new_n569_;
  assign new_n571_ = p_567_194_ & ~new_n570_;
  assign new_n572_ = p_44_31_ & p_82_63_;
  assign new_n573_ = p_96_75_ & new_n572_;
  assign new_n574_ = p_132_105_ & new_n573_;
  assign new_n575_ = p_2106_222_ & ~new_n574_;
  assign p_319_656_ = ~new_n571_ & ~new_n575_;
  assign new_n577_ = p_483_191_ & ~new_n567_;
  assign new_n578_ = p_319_656_ & new_n577_;
  assign p_188_761_ = ~p_661_196_ | ~new_n578_;
  assign new_n580_ = p_2084_216_ & p_2072_214_;
  assign new_n581_ = p_2078_215_ & new_n580_;
  assign p_158_349_ = ~p_2090_217_ | ~new_n581_;
  assign new_n583_ = p_661_196_ & p_15_10_;
  assign p_259_414_ = ~p_2_1_ | ~new_n583_;
  assign p_325_507_ = new_n570_ & new_n574_;
  assign new_n586_ = ~p_288_700_ & ~p_166_625_;
  assign new_n587_ = p_288_700_ & p_166_625_;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = ~p_290_704_ & p_305_702_;
  assign new_n590_ = p_290_704_ & ~p_305_702_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = new_n588_ & ~new_n591_;
  assign new_n593_ = ~new_n588_ & new_n591_;
  assign new_n594_ = ~new_n592_ & ~new_n593_;
  assign new_n595_ = ~new_n326_ & new_n334_;
  assign new_n596_ = new_n326_ & ~new_n334_;
  assign new_n597_ = ~new_n595_ & ~new_n596_;
  assign new_n598_ = ~p_171_621_ & p_168_623_;
  assign new_n599_ = p_171_621_ & ~p_168_623_;
  assign new_n600_ = ~new_n598_ & ~new_n599_;
  assign new_n601_ = ~new_n317_ & ~p_299_692_;
  assign new_n602_ = new_n317_ & p_299_692_;
  assign new_n603_ = ~new_n601_ & ~new_n602_;
  assign new_n604_ = ~new_n597_ & ~new_n600_;
  assign new_n605_ = ~new_n603_ & new_n604_;
  assign new_n606_ = new_n600_ & ~new_n603_;
  assign new_n607_ = new_n597_ & new_n606_;
  assign new_n608_ = ~new_n605_ & ~new_n607_;
  assign new_n609_ = new_n597_ & ~new_n600_;
  assign new_n610_ = new_n603_ & new_n609_;
  assign new_n611_ = new_n600_ & new_n603_;
  assign new_n612_ = ~new_n597_ & new_n611_;
  assign new_n613_ = ~new_n610_ & ~new_n612_;
  assign new_n614_ = new_n608_ & new_n613_;
  assign new_n615_ = new_n594_ & ~new_n614_;
  assign new_n616_ = ~new_n594_ & new_n614_;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign p_397_1406_ = ~p_37_28_ & new_n617_;
  assign new_n619_ = p_860_197_ & ~new_n317_;
  assign new_n620_ = ~p_860_197_ & ~new_n338_;
  assign p_148_851_ = new_n619_ | new_n620_;
  assign new_n622_ = ~p_1384_202_ & ~p_164_607_;
  assign new_n623_ = p_40_29_ & new_n622_;
  assign new_n624_ = p_160_609_ & new_n623_;
  assign new_n625_ = ~p_1348_201_ & ~new_n624_;
  assign new_n626_ = ~p_2067_213_ & new_n624_;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign new_n628_ = new_n317_ & ~new_n627_;
  assign new_n629_ = ~p_1956_203_ & ~new_n624_;
  assign new_n630_ = ~p_2072_214_ & new_n624_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = p_299_692_ & ~new_n631_;
  assign new_n633_ = ~p_299_692_ & new_n631_;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = new_n628_ & ~new_n634_;
  assign new_n636_ = ~p_1341_200_ & ~new_n624_;
  assign new_n637_ = ~p_1996_211_ & new_n624_;
  assign new_n638_ = ~new_n636_ & ~new_n637_;
  assign new_n639_ = new_n334_ & ~new_n638_;
  assign new_n640_ = ~new_n317_ & ~new_n627_;
  assign new_n641_ = new_n317_ & new_n627_;
  assign new_n642_ = ~new_n640_ & ~new_n641_;
  assign new_n643_ = ~new_n634_ & new_n639_;
  assign new_n644_ = ~new_n642_ & new_n643_;
  assign new_n645_ = ~p_299_692_ & ~new_n631_;
  assign new_n646_ = ~new_n635_ & ~new_n644_;
  assign new_n647_ = ~new_n645_ & new_n646_;
  assign new_n648_ = p_305_702_ & ~new_n624_;
  assign new_n649_ = p_8_7_ & new_n648_;
  assign new_n650_ = ~p_1981_208_ & ~new_n624_;
  assign new_n651_ = p_8_7_ & new_n650_;
  assign new_n652_ = new_n649_ & new_n651_;
  assign new_n653_ = ~new_n649_ & ~new_n651_;
  assign new_n654_ = ~new_n652_ & ~new_n653_;
  assign new_n655_ = ~p_168_623_ & new_n624_;
  assign new_n656_ = ~p_168_623_ & ~new_n624_;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = p_8_7_ & ~new_n657_;
  assign new_n659_ = ~p_1966_205_ & ~new_n624_;
  assign new_n660_ = ~p_2084_216_ & new_n624_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = p_8_7_ & ~new_n661_;
  assign new_n663_ = new_n658_ & new_n662_;
  assign new_n664_ = ~new_n658_ & ~new_n662_;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = ~p_1961_204_ & ~new_n624_;
  assign new_n667_ = ~p_2078_215_ & new_n624_;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = ~p_171_621_ & ~new_n668_;
  assign new_n670_ = p_171_621_ & new_n668_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~p_166_625_ & new_n624_;
  assign new_n673_ = ~p_166_625_ & ~new_n624_;
  assign new_n674_ = ~new_n672_ & ~new_n673_;
  assign new_n675_ = p_8_7_ & ~new_n674_;
  assign new_n676_ = ~p_1971_206_ & ~new_n624_;
  assign new_n677_ = ~p_2090_217_ & new_n624_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = p_8_7_ & ~new_n678_;
  assign new_n680_ = new_n675_ & new_n679_;
  assign new_n681_ = ~new_n675_ & ~new_n679_;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = p_288_700_ & ~new_n624_;
  assign new_n684_ = p_8_7_ & new_n683_;
  assign new_n685_ = ~p_1976_207_ & ~new_n624_;
  assign new_n686_ = p_8_7_ & new_n685_;
  assign new_n687_ = new_n684_ & new_n686_;
  assign new_n688_ = ~new_n684_ & ~new_n686_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = ~new_n654_ & ~new_n665_;
  assign new_n691_ = ~new_n671_ & new_n690_;
  assign new_n692_ = ~new_n682_ & new_n691_;
  assign new_n693_ = ~new_n689_ & new_n692_;
  assign new_n694_ = ~new_n647_ & new_n693_;
  assign new_n695_ = ~new_n658_ & new_n662_;
  assign new_n696_ = ~new_n654_ & ~new_n689_;
  assign new_n697_ = new_n695_ & new_n696_;
  assign new_n698_ = ~new_n682_ & new_n697_;
  assign new_n699_ = p_171_621_ & ~new_n668_;
  assign new_n700_ = ~new_n689_ & new_n699_;
  assign new_n701_ = ~new_n682_ & new_n700_;
  assign new_n702_ = ~new_n654_ & new_n701_;
  assign new_n703_ = ~new_n665_ & new_n702_;
  assign new_n704_ = ~new_n684_ & new_n686_;
  assign new_n705_ = ~new_n654_ & new_n704_;
  assign new_n706_ = ~new_n675_ & new_n679_;
  assign new_n707_ = ~new_n654_ & new_n706_;
  assign new_n708_ = ~new_n689_ & new_n707_;
  assign new_n709_ = ~new_n649_ & new_n651_;
  assign new_n710_ = ~new_n698_ & ~new_n703_;
  assign new_n711_ = ~new_n705_ & new_n710_;
  assign new_n712_ = ~new_n708_ & new_n711_;
  assign new_n713_ = ~new_n709_ & new_n712_;
  assign new_n714_ = ~new_n694_ & new_n713_;
  assign new_n715_ = p_160_609_ & ~new_n622_;
  assign new_n716_ = p_40_29_ & new_n715_;
  assign new_n717_ = ~new_n357_ & ~new_n624_;
  assign new_n718_ = new_n716_ & new_n717_;
  assign new_n719_ = ~p_2067_213_ & ~new_n624_;
  assign new_n720_ = new_n716_ & new_n719_;
  assign new_n721_ = new_n718_ & new_n720_;
  assign new_n722_ = ~new_n718_ & ~new_n720_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = p_290_704_ & ~new_n624_;
  assign new_n725_ = new_n716_ & new_n724_;
  assign new_n726_ = ~p_1986_209_ & ~new_n624_;
  assign new_n727_ = new_n716_ & new_n726_;
  assign new_n728_ = new_n725_ & new_n727_;
  assign new_n729_ = ~new_n725_ & ~new_n727_;
  assign new_n730_ = ~new_n728_ & ~new_n729_;
  assign new_n731_ = ~new_n553_ & ~new_n624_;
  assign new_n732_ = new_n716_ & new_n731_;
  assign new_n733_ = ~p_1991_210_ & ~new_n624_;
  assign new_n734_ = new_n716_ & new_n733_;
  assign new_n735_ = new_n732_ & new_n734_;
  assign new_n736_ = ~new_n732_ & ~new_n734_;
  assign new_n737_ = ~new_n735_ & ~new_n736_;
  assign new_n738_ = ~new_n370_ & ~new_n624_;
  assign new_n739_ = new_n716_ & new_n738_;
  assign new_n740_ = ~p_1996_211_ & ~new_n624_;
  assign new_n741_ = new_n716_ & new_n740_;
  assign new_n742_ = new_n739_ & new_n741_;
  assign new_n743_ = ~new_n739_ & ~new_n741_;
  assign new_n744_ = ~new_n742_ & ~new_n743_;
  assign new_n745_ = ~new_n723_ & ~new_n730_;
  assign new_n746_ = ~new_n737_ & new_n745_;
  assign new_n747_ = ~new_n744_ & new_n746_;
  assign new_n748_ = ~new_n725_ & new_n727_;
  assign new_n749_ = ~new_n723_ & ~new_n744_;
  assign new_n750_ = new_n748_ & new_n749_;
  assign new_n751_ = ~new_n737_ & new_n750_;
  assign new_n752_ = ~new_n739_ & new_n741_;
  assign new_n753_ = ~new_n723_ & new_n752_;
  assign new_n754_ = ~new_n732_ & new_n734_;
  assign new_n755_ = ~new_n723_ & new_n754_;
  assign new_n756_ = ~new_n744_ & new_n755_;
  assign new_n757_ = ~new_n718_ & new_n720_;
  assign new_n758_ = ~new_n751_ & ~new_n753_;
  assign new_n759_ = ~new_n756_ & new_n758_;
  assign new_n760_ = ~new_n757_ & new_n759_;
  assign new_n761_ = ~new_n747_ & new_n760_;
  assign new_n762_ = ~new_n714_ & ~new_n761_;
  assign new_n763_ = new_n714_ & ~new_n760_;
  assign p_329_1414_ = new_n762_ | new_n763_;
  assign new_n765_ = p_868_198_ & ~p_168_623_;
  assign new_n766_ = ~p_868_198_ & p_299_692_;
  assign p_297_849_ = new_n765_ | new_n766_;
  assign new_n768_ = ~p_2096_218_ & ~new_n439_;
  assign new_n769_ = ~new_n439_ & ~new_n768_;
  assign new_n770_ = ~p_2096_218_ & ~new_n768_;
  assign new_n771_ = ~new_n769_ & ~new_n770_;
  assign new_n772_ = ~new_n347_ & ~new_n349_;
  assign new_n773_ = ~new_n351_ & new_n772_;
  assign new_n774_ = ~new_n353_ & new_n773_;
  assign new_n775_ = ~p_2100_219_ & ~new_n774_;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign new_n777_ = ~p_2100_219_ & ~new_n775_;
  assign new_n778_ = ~new_n776_ & ~new_n777_;
  assign p_156_1046_ = ~new_n771_ | ~new_n778_;
  assign new_n780_ = p_860_197_ & ~new_n334_;
  assign p_153_671_ = ~p_860_197_ | new_n780_;
  assign p_223_413_ = ~p_661_196_ | ~p_7_6_;
  assign new_n783_ = ~new_n338_ & ~new_n603_;
  assign new_n784_ = ~new_n597_ & new_n783_;
  assign new_n785_ = ~new_n597_ & new_n603_;
  assign new_n786_ = new_n338_ & new_n785_;
  assign new_n787_ = ~new_n784_ & ~new_n786_;
  assign new_n788_ = new_n338_ & ~new_n603_;
  assign new_n789_ = new_n597_ & new_n788_;
  assign new_n790_ = new_n597_ & new_n603_;
  assign new_n791_ = ~new_n338_ & new_n790_;
  assign new_n792_ = ~new_n789_ & ~new_n791_;
  assign new_n793_ = new_n787_ & new_n792_;
  assign new_n794_ = new_n594_ & ~new_n793_;
  assign new_n795_ = ~new_n594_ & new_n793_;
  assign new_n796_ = ~new_n794_ & ~new_n795_;
  assign new_n797_ = p_868_198_ & ~new_n796_;
  assign new_n798_ = ~p_868_198_ & ~new_n326_;
  assign p_331_1401_ = new_n797_ | new_n798_;
  assign new_n800_ = p_160_609_ & ~p_162_612_;
  assign new_n801_ = ~p_160_609_ & p_162_612_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = new_n439_ & ~new_n774_;
  assign new_n804_ = ~new_n439_ & new_n774_;
  assign new_n805_ = ~new_n803_ & ~new_n804_;
  assign new_n806_ = new_n802_ & ~new_n805_;
  assign new_n807_ = ~new_n802_ & new_n805_;
  assign new_n808_ = ~new_n806_ & ~new_n807_;
  assign new_n809_ = p_118_93_ & new_n347_;
  assign new_n810_ = p_106_83_ & new_n349_;
  assign new_n811_ = p_130_103_ & new_n351_;
  assign new_n812_ = p_142_113_ & new_n353_;
  assign new_n813_ = ~new_n809_ & ~new_n810_;
  assign new_n814_ = ~new_n811_ & new_n813_;
  assign new_n815_ = ~new_n812_ & new_n814_;
  assign new_n816_ = ~new_n553_ & new_n815_;
  assign new_n817_ = new_n553_ & ~new_n815_;
  assign new_n818_ = ~new_n816_ & ~new_n817_;
  assign new_n819_ = ~p_164_607_ & new_n396_;
  assign new_n820_ = p_164_607_ & ~new_n396_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign new_n822_ = ~new_n357_ & new_n370_;
  assign new_n823_ = new_n357_ & ~new_n370_;
  assign new_n824_ = ~new_n822_ & ~new_n823_;
  assign new_n825_ = ~new_n818_ & ~new_n821_;
  assign new_n826_ = ~new_n824_ & new_n825_;
  assign new_n827_ = new_n821_ & ~new_n824_;
  assign new_n828_ = new_n818_ & new_n827_;
  assign new_n829_ = ~new_n826_ & ~new_n828_;
  assign new_n830_ = new_n818_ & ~new_n821_;
  assign new_n831_ = new_n824_ & new_n830_;
  assign new_n832_ = new_n821_ & new_n824_;
  assign new_n833_ = ~new_n818_ & new_n832_;
  assign new_n834_ = ~new_n831_ & ~new_n833_;
  assign new_n835_ = new_n829_ & new_n834_;
  assign new_n836_ = new_n808_ & ~new_n835_;
  assign new_n837_ = ~new_n808_ & new_n835_;
  assign new_n838_ = ~new_n836_ & ~new_n837_;
  assign p_395_1392_ = ~p_37_28_ & new_n838_;
  assign new_n840_ = p_868_198_ & ~new_n338_;
  assign new_n841_ = ~p_868_198_ & ~new_n334_;
  assign p_282_922_ = new_n840_ | new_n841_;
  assign p_173_389_ = p_94_73_ & p_452_190_;
  assign p_217_423_ = ~p_2106_222_ | p_223_413_;
  assign new_n845_ = p_1986_209_ & ~p_1981_208_;
  assign new_n846_ = ~p_1986_209_ & p_1981_208_;
  assign new_n847_ = ~new_n845_ & ~new_n846_;
  assign new_n848_ = p_1996_211_ & ~p_1991_210_;
  assign new_n849_ = ~p_1996_211_ & p_1991_210_;
  assign new_n850_ = ~new_n848_ & ~new_n849_;
  assign new_n851_ = new_n847_ & ~new_n850_;
  assign new_n852_ = ~new_n847_ & new_n850_;
  assign new_n853_ = ~new_n851_ & ~new_n852_;
  assign new_n854_ = ~p_2474_231_ & p_1956_203_;
  assign new_n855_ = p_2474_231_ & ~p_1956_203_;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = p_1976_207_ & ~p_1971_206_;
  assign new_n858_ = ~p_1976_207_ & p_1971_206_;
  assign new_n859_ = ~new_n857_ & ~new_n858_;
  assign new_n860_ = ~p_1961_204_ & p_1966_205_;
  assign new_n861_ = p_1961_204_ & ~p_1966_205_;
  assign new_n862_ = ~new_n860_ & ~new_n861_;
  assign new_n863_ = ~new_n856_ & ~new_n859_;
  assign new_n864_ = ~new_n862_ & new_n863_;
  assign new_n865_ = new_n859_ & ~new_n862_;
  assign new_n866_ = new_n856_ & new_n865_;
  assign new_n867_ = ~new_n864_ & ~new_n866_;
  assign new_n868_ = new_n856_ & ~new_n859_;
  assign new_n869_ = new_n862_ & new_n868_;
  assign new_n870_ = new_n859_ & new_n862_;
  assign new_n871_ = ~new_n856_ & new_n870_;
  assign new_n872_ = ~new_n869_ & ~new_n871_;
  assign new_n873_ = new_n867_ & new_n872_;
  assign new_n874_ = new_n853_ & ~new_n873_;
  assign new_n875_ = ~new_n853_ & new_n873_;
  assign p_229_1180_ = ~new_n874_ & ~new_n875_;
  assign new_n877_ = ~p_2096_218_ & p_2100_219_;
  assign new_n878_ = p_2096_218_ & ~p_2100_219_;
  assign new_n879_ = ~new_n877_ & ~new_n878_;
  assign new_n880_ = ~p_2678_232_ & p_2067_213_;
  assign new_n881_ = p_2678_232_ & ~p_2067_213_;
  assign new_n882_ = ~new_n880_ & ~new_n881_;
  assign new_n883_ = p_2090_217_ & ~p_2084_216_;
  assign new_n884_ = ~p_2090_217_ & p_2084_216_;
  assign new_n885_ = ~new_n883_ & ~new_n884_;
  assign new_n886_ = p_2078_215_ & ~p_2072_214_;
  assign new_n887_ = ~p_2078_215_ & p_2072_214_;
  assign new_n888_ = ~new_n886_ & ~new_n887_;
  assign new_n889_ = ~new_n882_ & ~new_n885_;
  assign new_n890_ = ~new_n888_ & new_n889_;
  assign new_n891_ = new_n885_ & ~new_n888_;
  assign new_n892_ = new_n882_ & new_n891_;
  assign new_n893_ = ~new_n890_ & ~new_n892_;
  assign new_n894_ = new_n882_ & ~new_n885_;
  assign new_n895_ = new_n888_ & new_n894_;
  assign new_n896_ = new_n885_ & new_n888_;
  assign new_n897_ = ~new_n882_ & new_n896_;
  assign new_n898_ = ~new_n895_ & ~new_n897_;
  assign new_n899_ = new_n893_ & new_n898_;
  assign new_n900_ = new_n879_ & ~new_n899_;
  assign new_n901_ = ~new_n879_ & new_n899_;
  assign p_227_1179_ = ~new_n900_ & ~new_n901_;
  assign new_n903_ = p_483_191_ & p_319_656_;
  assign new_n904_ = p_36_27_ & new_n903_;
  assign p_176_803_ = ~p_661_196_ | ~new_n904_;
  assign new_n906_ = ~p_2454_230_ & p_2451_229_;
  assign new_n907_ = p_2454_230_ & ~p_2451_229_;
  assign new_n908_ = ~new_n906_ & ~new_n907_;
  assign new_n909_ = ~p_1341_200_ & p_1348_201_;
  assign new_n910_ = p_1341_200_ & ~p_1348_201_;
  assign new_n911_ = ~new_n909_ & ~new_n910_;
  assign new_n912_ = new_n908_ & ~new_n911_;
  assign new_n913_ = ~new_n908_ & new_n911_;
  assign new_n914_ = ~new_n912_ & ~new_n913_;
  assign new_n915_ = ~p_2430_224_ & p_2427_223_;
  assign new_n916_ = p_2430_224_ & ~p_2427_223_;
  assign new_n917_ = ~new_n915_ & ~new_n916_;
  assign new_n918_ = p_2443_227_ & ~p_2446_228_;
  assign new_n919_ = ~p_2443_227_ & p_2446_228_;
  assign new_n920_ = ~new_n918_ & ~new_n919_;
  assign new_n921_ = p_2435_225_ & ~p_2438_226_;
  assign new_n922_ = ~p_2435_225_ & p_2438_226_;
  assign new_n923_ = ~new_n921_ & ~new_n922_;
  assign new_n924_ = ~new_n917_ & ~new_n920_;
  assign new_n925_ = ~new_n923_ & new_n924_;
  assign new_n926_ = new_n920_ & ~new_n923_;
  assign new_n927_ = new_n917_ & new_n926_;
  assign new_n928_ = ~new_n925_ & ~new_n927_;
  assign new_n929_ = new_n917_ & ~new_n920_;
  assign new_n930_ = new_n923_ & new_n929_;
  assign new_n931_ = new_n920_ & new_n923_;
  assign new_n932_ = ~new_n917_ & new_n931_;
  assign new_n933_ = ~new_n930_ & ~new_n932_;
  assign new_n934_ = new_n928_ & new_n933_;
  assign new_n935_ = new_n914_ & ~new_n934_;
  assign new_n936_ = ~new_n914_ & new_n934_;
  assign new_n937_ = ~new_n935_ & ~new_n936_;
  assign p_401_1276_ = p_14_9_ & new_n937_;
  assign p_234_376_ = ~p_567_194_ | p_223_413_;
  assign new_n940_ = ~p_229_1180_ & ~p_401_1276_;
  assign new_n941_ = ~p_397_1406_ & ~p_227_1179_;
  assign new_n942_ = ~p_395_1392_ & new_n941_;
  assign new_n943_ = p_319_656_ & new_n940_;
  assign p_308_1425_ = new_n942_ & new_n943_;
  assign p_231_1422_ = 1'b0;
  assign p_150_1277_ = ~p_311_1278_;
  assign p_221_305_ = ~p_96_75_;
  assign p_235_307_ = ~p_69_52_;
  assign p_301_694_ = ~p_171_621_;
  assign p_218_311_ = ~p_44_31_;
  assign p_261_506_ = ~p_325_507_;
  assign p_236_303_ = ~p_120_95_;
  assign p_220_306_ = ~p_82_63_;
  assign p_303_698_ = ~p_166_625_;
  assign p_237_309_ = ~p_57_42_;
  assign p_286_696_ = ~p_168_623_;
  assign p_238_304_ = ~p_108_85_;
  assign p_219_302_ = ~p_132_105_;
  assign p_225_1424_ = ~p_308_1425_;
  assign p_367_288_ = p_1083_199_;
  assign p_384_262_ = p_2066_212_;
  assign p_321_848_ = p_284_847_;
  assign p_350_301_ = p_452_190_;
  assign p_369_289_ = p_1083_199_;
  assign p_411_264_ = p_2066_212_;
  assign p_337_263_ = p_2066_212_;
  assign p_391_379_ = p_452_190_;
  assign p_280_850_ = p_297_849_;
  assign p_335_299_ = p_452_190_;
  assign p_295_1400_ = p_331_1401_;
  assign p_323_923_ = p_282_922_;
  assign p_409_298_ = p_452_190_;
endmodule

